magic
tech sky130A
timestamp 1756781249
use icellwrapdummy  icell_dummy_left
timestamp 1756780365
transform 1 0 0 0 1 0
box 0 -27 393 243
use icellwrapdummy  icell_dummy_right
timestamp 1756780365
transform 1 0 6681 0 1 0
box 0 -27 393 243
use icellwrap  XIC
array 0 14 393 0 0 232
timestamp 1756690244
transform 1 0 393 0 1 0
box 0 -27 393 243
use icellwrapfinal  XIC_15
timestamp 1756777818
transform 1 0 6288 0 1 0
box 0 -27 393 243
<< end >>
