magic
tech sky130A
magscale 1 2
timestamp 1757605323
<< metal1 >>
rect 1618 38806 1684 38812
rect 1618 38752 1624 38806
rect 1678 38802 1684 38806
rect 1678 38756 14718 38802
rect 1678 38752 1684 38756
rect 1618 38746 1684 38752
rect 1718 38706 1784 38712
rect 1718 38652 1724 38706
rect 1778 38702 1784 38706
rect 1778 38656 14108 38702
rect 1778 38652 1784 38656
rect 1718 38646 1784 38652
rect 1818 38606 1884 38612
rect 1818 38552 1824 38606
rect 1878 38602 1884 38606
rect 1878 38556 12542 38602
rect 1878 38552 1884 38556
rect 1818 38546 1884 38552
rect 1918 38506 1984 38512
rect 1918 38452 1924 38506
rect 1978 38502 1984 38506
rect 1978 38456 12460 38502
rect 1978 38452 1984 38456
rect 1918 38446 1984 38452
rect 2704 38290 2770 38296
rect 2704 38236 2710 38290
rect 2764 38286 2770 38290
rect 2764 38240 4502 38286
rect 2764 38236 2770 38240
rect 2704 38230 2770 38236
rect 2604 38190 2670 38196
rect 2604 38136 2610 38190
rect 2664 38186 2670 38190
rect 2664 38140 4162 38186
rect 2664 38136 2670 38140
rect 2604 38130 2670 38136
rect 2504 38090 2570 38096
rect 2504 38036 2510 38090
rect 2564 38086 2570 38090
rect 2564 38040 3562 38086
rect 2564 38036 2570 38040
rect 2504 38030 2570 38036
rect 3518 37808 3562 38040
rect 4116 37808 4162 38140
rect 4456 37808 4502 38240
rect 12420 37812 12460 38456
rect 12502 37812 12542 38556
rect 14068 37812 14108 38656
rect 14678 37812 14718 38756
rect 1518 30712 1584 30718
rect 1518 30658 1524 30712
rect 1578 30704 1584 30712
rect 1578 30658 2840 30704
rect 1518 30652 1584 30658
rect 1418 30626 1484 30632
rect 1418 30572 1424 30626
rect 1478 30622 1484 30626
rect 1478 30576 2840 30622
rect 1478 30572 1484 30576
rect 1418 30566 1484 30572
rect 1318 29060 1384 29066
rect 1318 29006 1324 29060
rect 1378 29056 1384 29060
rect 1378 29010 2840 29056
rect 1378 29006 1384 29010
rect 1318 29000 1384 29006
rect 1218 28450 1284 28456
rect 1218 28396 1224 28450
rect 1278 28446 1284 28450
rect 1278 28400 2840 28446
rect 1278 28396 1284 28400
rect 1218 28390 1284 28396
rect 1618 26092 1684 26098
rect 1618 26038 1624 26092
rect 1678 26088 1684 26092
rect 1678 26042 14718 26088
rect 1678 26038 1684 26042
rect 1618 26032 1684 26038
rect 1718 25992 1784 25998
rect 1718 25938 1724 25992
rect 1778 25988 1784 25992
rect 1778 25942 14108 25988
rect 1778 25938 1784 25942
rect 1718 25932 1784 25938
rect 1818 25892 1884 25898
rect 1818 25838 1824 25892
rect 1878 25888 1884 25892
rect 1878 25842 12542 25888
rect 1878 25838 1884 25842
rect 1818 25832 1884 25838
rect 1918 25792 1984 25798
rect 1918 25738 1924 25792
rect 1978 25788 1984 25792
rect 1978 25742 12460 25788
rect 1978 25738 1984 25742
rect 1918 25732 1984 25738
rect 2364 25576 2430 25582
rect 2364 25522 2370 25576
rect 2424 25572 2430 25576
rect 2424 25526 4502 25572
rect 2424 25522 2430 25526
rect 2364 25516 2430 25522
rect 2264 25476 2330 25482
rect 2264 25422 2270 25476
rect 2324 25472 2330 25476
rect 2324 25426 4162 25472
rect 2324 25422 2330 25426
rect 2264 25416 2330 25422
rect 2164 25376 2230 25382
rect 2164 25322 2170 25376
rect 2224 25372 2230 25376
rect 2224 25326 3562 25372
rect 2224 25322 2230 25326
rect 2164 25316 2230 25322
rect 3518 25094 3562 25326
rect 4116 25094 4162 25426
rect 4456 25094 4502 25526
rect 12420 25098 12460 25742
rect 12502 25098 12542 25842
rect 14068 25098 14108 25942
rect 14678 25098 14718 26042
rect 1518 17998 1584 18004
rect 1518 17944 1524 17998
rect 1578 17990 1584 17998
rect 1578 17944 2840 17990
rect 1518 17938 1584 17944
rect 1418 17912 1484 17918
rect 1418 17858 1424 17912
rect 1478 17908 1484 17912
rect 1478 17862 2840 17908
rect 1478 17858 1484 17862
rect 1418 17852 1484 17858
rect 1318 16346 1384 16352
rect 1318 16292 1324 16346
rect 1378 16342 1384 16346
rect 1378 16296 2840 16342
rect 1378 16292 1384 16296
rect 1318 16286 1384 16292
rect 1218 15736 1284 15742
rect 1218 15682 1224 15736
rect 1278 15732 1284 15736
rect 1278 15686 2840 15732
rect 1278 15682 1284 15686
rect 1218 15676 1284 15682
rect 1618 13378 1684 13384
rect 1618 13324 1624 13378
rect 1678 13374 1684 13378
rect 1678 13328 14718 13374
rect 1678 13324 1684 13328
rect 1618 13318 1684 13324
rect 1718 13278 1784 13284
rect 1718 13224 1724 13278
rect 1778 13274 1784 13278
rect 1778 13228 14108 13274
rect 1778 13224 1784 13228
rect 1718 13218 1784 13224
rect 1818 13178 1884 13184
rect 1818 13124 1824 13178
rect 1878 13174 1884 13178
rect 1878 13128 12542 13174
rect 1878 13124 1884 13128
rect 1818 13118 1884 13124
rect 1918 13078 1984 13084
rect 1918 13024 1924 13078
rect 1978 13074 1984 13078
rect 1978 13028 12460 13074
rect 1978 13024 1984 13028
rect 1918 13018 1984 13024
rect 2364 12862 2430 12868
rect 2364 12808 2370 12862
rect 2424 12858 2430 12862
rect 2424 12812 4502 12858
rect 2424 12808 2430 12812
rect 2364 12802 2430 12808
rect 2264 12762 2330 12768
rect 2264 12708 2270 12762
rect 2324 12758 2330 12762
rect 2324 12712 4162 12758
rect 2324 12708 2330 12712
rect 2264 12702 2330 12708
rect 2164 12662 2230 12668
rect 2164 12608 2170 12662
rect 2224 12658 2230 12662
rect 2224 12612 3562 12658
rect 2224 12608 2230 12612
rect 2164 12602 2230 12608
rect 3518 12380 3562 12612
rect 4116 12380 4162 12712
rect 4456 12380 4502 12812
rect 12420 12384 12460 13028
rect 12502 12384 12542 13128
rect 14068 12384 14108 13228
rect 14678 12384 14718 13328
rect 1518 5284 1584 5290
rect 1518 5230 1524 5284
rect 1578 5276 1584 5284
rect 1578 5230 2840 5276
rect 1518 5224 1584 5230
rect 1418 5198 1484 5204
rect 1418 5144 1424 5198
rect 1478 5194 1484 5198
rect 1478 5148 2840 5194
rect 1478 5144 1484 5148
rect 1418 5138 1484 5144
rect 1318 3632 1384 3638
rect 1318 3578 1324 3632
rect 1378 3628 1384 3632
rect 1378 3582 2840 3628
rect 1378 3578 1384 3582
rect 1318 3572 1384 3578
rect 1218 3022 1284 3028
rect 1218 2968 1224 3022
rect 1278 3018 1284 3022
rect 1278 2972 2840 3018
rect 1278 2968 1284 2972
rect 1218 2962 1284 2968
<< via1 >>
rect 1624 38752 1678 38806
rect 1724 38652 1778 38706
rect 1824 38552 1878 38606
rect 1924 38452 1978 38506
rect 2710 38236 2764 38290
rect 2610 38136 2664 38190
rect 2510 38036 2564 38090
rect 1524 30658 1578 30712
rect 1424 30572 1478 30626
rect 1324 29006 1378 29060
rect 1224 28396 1278 28450
rect 1624 26038 1678 26092
rect 1724 25938 1778 25992
rect 1824 25838 1878 25892
rect 1924 25738 1978 25792
rect 2370 25522 2424 25576
rect 2270 25422 2324 25476
rect 2170 25322 2224 25376
rect 1524 17944 1578 17998
rect 1424 17858 1478 17912
rect 1324 16292 1378 16346
rect 1224 15682 1278 15736
rect 1624 13324 1678 13378
rect 1724 13224 1778 13278
rect 1824 13124 1878 13178
rect 1924 13024 1978 13078
rect 2370 12808 2424 12862
rect 2270 12708 2324 12762
rect 2170 12608 2224 12662
rect 1524 5230 1578 5284
rect 1424 5144 1478 5198
rect 1324 3578 1378 3632
rect 1224 2968 1278 3022
<< metal2 >>
rect 23788 43616 23868 43626
rect 23788 43610 23798 43616
rect 1228 43564 23798 43610
rect 1228 28456 1274 43564
rect 23788 43558 23798 43564
rect 23858 43610 23868 43616
rect 23858 43564 29618 43610
rect 23858 43558 23868 43564
rect 23788 43548 23868 43558
rect 24340 43516 24420 43526
rect 24340 43510 24350 43516
rect 1328 43464 24350 43510
rect 1328 29066 1374 43464
rect 24340 43458 24350 43464
rect 24410 43510 24420 43516
rect 24410 43464 29618 43510
rect 24410 43458 24420 43464
rect 24340 43448 24420 43458
rect 24892 43418 24972 43428
rect 24892 43410 24902 43418
rect 1428 43364 24902 43410
rect 1428 30632 1474 43364
rect 24892 43360 24902 43364
rect 24962 43410 24972 43418
rect 24962 43364 29618 43410
rect 24962 43360 24972 43364
rect 24892 43350 24972 43360
rect 25444 43314 25524 43324
rect 25444 43310 25454 43314
rect 1528 43264 25454 43310
rect 1528 30718 1574 43264
rect 25444 43256 25454 43264
rect 25514 43310 25524 43314
rect 25514 43264 29618 43310
rect 25514 43256 25524 43264
rect 25444 43246 25524 43256
rect 25996 43216 26076 43226
rect 25996 43210 26006 43216
rect 1628 43164 26006 43210
rect 1628 38812 1674 43164
rect 25996 43158 26006 43164
rect 26066 43210 26076 43216
rect 26066 43164 29618 43210
rect 26066 43158 26076 43164
rect 25996 43148 26076 43158
rect 26548 43116 26628 43126
rect 26548 43110 26558 43116
rect 1728 43064 26558 43110
rect 1618 38806 1684 38812
rect 1618 38752 1624 38806
rect 1678 38752 1684 38806
rect 1618 38746 1684 38752
rect 1518 30712 1584 30718
rect 1518 30658 1524 30712
rect 1578 30658 1584 30712
rect 1518 30652 1584 30658
rect 1418 30626 1484 30632
rect 1418 30572 1424 30626
rect 1478 30572 1484 30626
rect 1418 30566 1484 30572
rect 1318 29060 1384 29066
rect 1318 29006 1324 29060
rect 1378 29006 1384 29060
rect 1318 29000 1384 29006
rect 1218 28450 1284 28456
rect 1218 28396 1224 28450
rect 1278 28396 1284 28450
rect 1218 28390 1284 28396
rect 1228 15742 1274 28390
rect 1328 16352 1374 29000
rect 1428 17918 1474 30566
rect 1528 18004 1574 30652
rect 1628 26098 1674 38746
rect 1728 38712 1774 43064
rect 26548 43058 26558 43064
rect 26618 43110 26628 43116
rect 26618 43064 29618 43110
rect 26618 43058 26628 43064
rect 26548 43048 26628 43058
rect 27100 43016 27180 43026
rect 27100 43010 27110 43016
rect 1828 42964 27110 43010
rect 1718 38706 1784 38712
rect 1718 38652 1724 38706
rect 1778 38652 1784 38706
rect 1718 38646 1784 38652
rect 1618 26092 1684 26098
rect 1618 26038 1624 26092
rect 1678 26038 1684 26092
rect 1618 26032 1684 26038
rect 1518 17998 1584 18004
rect 1518 17944 1524 17998
rect 1578 17944 1584 17998
rect 1518 17938 1584 17944
rect 1418 17912 1484 17918
rect 1418 17858 1424 17912
rect 1478 17858 1484 17912
rect 1418 17852 1484 17858
rect 1318 16346 1384 16352
rect 1318 16292 1324 16346
rect 1378 16292 1384 16346
rect 1318 16286 1384 16292
rect 1218 15736 1284 15742
rect 1218 15682 1224 15736
rect 1278 15682 1284 15736
rect 1218 15676 1284 15682
rect 1228 3028 1274 15676
rect 1328 3638 1374 16286
rect 1428 5204 1474 17852
rect 1528 5290 1574 17938
rect 1628 13384 1674 26032
rect 1728 25998 1774 38646
rect 1828 38612 1874 42964
rect 27100 42958 27110 42964
rect 27170 43010 27180 43016
rect 27170 42964 29618 43010
rect 27170 42958 27180 42964
rect 27100 42948 27180 42958
rect 27652 42916 27732 42926
rect 27652 42910 27662 42916
rect 1928 42864 27662 42910
rect 1818 38606 1884 38612
rect 1818 38552 1824 38606
rect 1878 38552 1884 38606
rect 1818 38546 1884 38552
rect 1718 25992 1784 25998
rect 1718 25938 1724 25992
rect 1778 25938 1784 25992
rect 1718 25932 1784 25938
rect 1618 13378 1684 13384
rect 1618 13324 1624 13378
rect 1678 13324 1684 13378
rect 1618 13318 1684 13324
rect 1518 5284 1584 5290
rect 1518 5230 1524 5284
rect 1578 5230 1584 5284
rect 1518 5224 1584 5230
rect 1418 5198 1484 5204
rect 1418 5144 1424 5198
rect 1478 5144 1484 5198
rect 1418 5138 1484 5144
rect 1318 3632 1384 3638
rect 1318 3578 1324 3632
rect 1378 3578 1384 3632
rect 1318 3572 1384 3578
rect 1218 3022 1284 3028
rect 1218 2968 1224 3022
rect 1278 2968 1284 3022
rect 1328 2972 1374 3572
rect 1428 2972 1474 5138
rect 1528 2972 1574 5224
rect 1628 2972 1674 13318
rect 1728 13284 1774 25932
rect 1828 25898 1874 38546
rect 1928 38512 1974 42864
rect 27652 42858 27662 42864
rect 27722 42910 27732 42916
rect 27722 42864 29618 42910
rect 27722 42858 27732 42864
rect 27652 42848 27732 42858
rect 20476 42642 20556 42652
rect 20476 42636 20486 42642
rect 2174 42590 20486 42636
rect 1918 38506 1984 38512
rect 1918 38452 1924 38506
rect 1978 38452 1984 38506
rect 1918 38446 1984 38452
rect 1818 25892 1884 25898
rect 1818 25838 1824 25892
rect 1878 25838 1884 25892
rect 1818 25832 1884 25838
rect 1718 13278 1784 13284
rect 1718 13224 1724 13278
rect 1778 13224 1784 13278
rect 1718 13218 1784 13224
rect 1728 2972 1774 13218
rect 1828 13184 1874 25832
rect 1928 25798 1974 38446
rect 1918 25792 1984 25798
rect 1918 25738 1924 25792
rect 1978 25738 1984 25792
rect 1918 25732 1984 25738
rect 1818 13178 1884 13184
rect 1818 13124 1824 13178
rect 1878 13124 1884 13178
rect 1818 13118 1884 13124
rect 1828 2972 1874 13118
rect 1928 13084 1974 25732
rect 2174 25382 2220 42590
rect 20476 42584 20486 42590
rect 20546 42636 20556 42642
rect 20546 42590 23644 42636
rect 20546 42584 20556 42590
rect 20476 42574 20556 42584
rect 21028 42542 21108 42552
rect 21028 42536 21038 42542
rect 2274 42490 21038 42536
rect 2274 25482 2320 42490
rect 21028 42484 21038 42490
rect 21098 42536 21108 42542
rect 21098 42490 23644 42536
rect 21098 42484 21108 42490
rect 21028 42474 21108 42484
rect 21580 42442 21660 42452
rect 21580 42436 21590 42442
rect 2374 42390 21590 42436
rect 2374 25582 2420 42390
rect 21580 42384 21590 42390
rect 21650 42436 21660 42442
rect 21650 42390 23644 42436
rect 21650 42384 21660 42390
rect 21580 42374 21660 42384
rect 22132 42302 22212 42312
rect 22132 42296 22142 42302
rect 2514 42250 22142 42296
rect 2514 38096 2560 42250
rect 22132 42244 22142 42250
rect 22202 42296 22212 42302
rect 22202 42250 23644 42296
rect 22202 42244 22212 42250
rect 22132 42234 22212 42244
rect 22684 42202 22764 42212
rect 22684 42196 22694 42202
rect 2614 42150 22694 42196
rect 2614 38196 2660 42150
rect 22684 42144 22694 42150
rect 22754 42196 22764 42202
rect 22754 42150 23644 42196
rect 22754 42144 22764 42150
rect 22684 42134 22764 42144
rect 23236 42102 23316 42112
rect 23236 42096 23246 42102
rect 2714 42050 23246 42096
rect 2714 38296 2760 42050
rect 23236 42044 23246 42050
rect 23306 42096 23316 42102
rect 23306 42050 23644 42096
rect 23306 42044 23316 42050
rect 23236 42034 23316 42044
rect 2704 38290 2770 38296
rect 2704 38236 2710 38290
rect 2764 38236 2770 38290
rect 2704 38230 2770 38236
rect 2604 38190 2670 38196
rect 2604 38136 2610 38190
rect 2664 38136 2670 38190
rect 2604 38130 2670 38136
rect 2504 38090 2570 38096
rect 2504 38036 2510 38090
rect 2564 38036 2570 38090
rect 2614 38040 2660 38130
rect 2714 38040 2760 38230
rect 2504 38030 2570 38036
rect 19008 35722 19102 35734
rect 19008 35720 19906 35722
rect 19008 35664 19028 35720
rect 19084 35664 19906 35720
rect 19008 35662 19906 35664
rect 19962 35662 19971 35722
rect 19008 35658 19102 35662
rect 19028 35655 19084 35658
rect 2364 25576 2430 25582
rect 2364 25522 2370 25576
rect 2424 25522 2430 25576
rect 2364 25516 2430 25522
rect 2264 25476 2330 25482
rect 2264 25422 2270 25476
rect 2324 25422 2330 25476
rect 2264 25416 2330 25422
rect 2164 25376 2230 25382
rect 2164 25322 2170 25376
rect 2224 25322 2230 25376
rect 2164 25316 2230 25322
rect 1918 13078 1984 13084
rect 1918 13024 1924 13078
rect 1978 13024 1984 13078
rect 1918 13018 1984 13024
rect 1928 2972 1974 13018
rect 2174 12668 2220 25316
rect 2274 12768 2320 25416
rect 2374 12868 2420 25516
rect 2364 12862 2430 12868
rect 2364 12808 2370 12862
rect 2424 12808 2430 12862
rect 2364 12802 2430 12808
rect 2264 12762 2330 12768
rect 2264 12708 2270 12762
rect 2324 12708 2330 12762
rect 2264 12702 2330 12708
rect 2164 12662 2230 12668
rect 2164 12608 2170 12662
rect 2224 12608 2230 12662
rect 2274 12612 2320 12702
rect 2374 12612 2420 12802
rect 2164 12602 2230 12608
rect 1218 2962 1284 2968
<< via2 >>
rect 23798 43558 23858 43616
rect 24350 43458 24410 43516
rect 24902 43360 24962 43418
rect 25454 43256 25514 43314
rect 26006 43158 26066 43216
rect 26558 43058 26618 43116
rect 27110 42958 27170 43016
rect 27662 42858 27722 42916
rect 20486 42584 20546 42642
rect 21038 42484 21098 42542
rect 21590 42384 21650 42442
rect 22142 42244 22202 42302
rect 22694 42144 22754 42202
rect 23246 42044 23306 42102
rect 19028 35664 19084 35720
rect 19906 35662 19962 35722
<< metal3 >>
rect 20482 44866 20550 44872
rect 20482 44798 20484 44866
rect 20548 44798 20550 44866
rect 20482 44792 20550 44798
rect 21034 44866 21102 44872
rect 21034 44798 21036 44866
rect 21100 44798 21102 44866
rect 21034 44792 21102 44798
rect 21586 44866 21654 44872
rect 21586 44798 21588 44866
rect 21652 44798 21654 44866
rect 21586 44792 21654 44798
rect 22138 44866 22206 44872
rect 22138 44798 22140 44866
rect 22204 44798 22206 44866
rect 22138 44792 22206 44798
rect 22690 44866 22758 44872
rect 22690 44798 22692 44866
rect 22756 44798 22758 44866
rect 22690 44792 22758 44798
rect 23242 44866 23310 44872
rect 23242 44798 23244 44866
rect 23308 44798 23310 44866
rect 23242 44792 23310 44798
rect 23794 44866 23862 44872
rect 23794 44798 23796 44866
rect 23860 44798 23862 44866
rect 23794 44792 23862 44798
rect 24346 44866 24414 44872
rect 24346 44798 24348 44866
rect 24412 44798 24414 44866
rect 24346 44792 24414 44798
rect 24898 44866 24966 44872
rect 24898 44798 24900 44866
rect 24964 44798 24966 44866
rect 24898 44792 24966 44798
rect 25450 44866 25518 44872
rect 25450 44798 25452 44866
rect 25516 44798 25518 44866
rect 25450 44792 25518 44798
rect 26002 44866 26070 44872
rect 26002 44798 26004 44866
rect 26068 44798 26070 44866
rect 26002 44792 26070 44798
rect 26554 44866 26622 44872
rect 26554 44798 26556 44866
rect 26620 44798 26622 44866
rect 26554 44792 26622 44798
rect 27106 44866 27174 44872
rect 27106 44798 27108 44866
rect 27172 44798 27174 44866
rect 27106 44792 27174 44798
rect 27658 44866 27726 44872
rect 27658 44798 27660 44866
rect 27724 44798 27726 44866
rect 27658 44792 27726 44798
rect 20486 42652 20546 44792
rect 20476 42642 20556 42652
rect 20476 42584 20486 42642
rect 20546 42584 20556 42642
rect 20476 42574 20556 42584
rect 20486 42224 20546 42574
rect 21038 42552 21098 44792
rect 21028 42542 21108 42552
rect 21028 42484 21038 42542
rect 21098 42484 21108 42542
rect 21028 42474 21108 42484
rect 21038 42224 21098 42474
rect 21590 42452 21650 44792
rect 21580 42442 21660 42452
rect 21580 42384 21590 42442
rect 21650 42384 21660 42442
rect 21580 42374 21660 42384
rect 21590 42224 21650 42374
rect 22142 42312 22202 44792
rect 22132 42302 22212 42312
rect 22132 42244 22142 42302
rect 22202 42244 22212 42302
rect 22132 42234 22212 42244
rect 22142 41884 22202 42234
rect 22694 42212 22754 44792
rect 22684 42202 22764 42212
rect 22684 42144 22694 42202
rect 22754 42144 22764 42202
rect 22684 42134 22764 42144
rect 22694 41884 22754 42134
rect 23246 42112 23306 44792
rect 23798 43626 23858 44792
rect 23788 43616 23868 43626
rect 23788 43558 23798 43616
rect 23858 43558 23868 43616
rect 23788 43548 23868 43558
rect 23798 42560 23858 43548
rect 24350 43526 24410 44792
rect 24340 43516 24420 43526
rect 24340 43458 24350 43516
rect 24410 43458 24420 43516
rect 24340 43448 24420 43458
rect 24350 42560 24410 43448
rect 24902 43428 24962 44792
rect 24892 43418 24972 43428
rect 24892 43360 24902 43418
rect 24962 43360 24972 43418
rect 24892 43350 24972 43360
rect 24902 42560 24962 43350
rect 25454 43324 25514 44792
rect 25444 43314 25524 43324
rect 25444 43256 25454 43314
rect 25514 43256 25524 43314
rect 25444 43246 25524 43256
rect 25454 42560 25514 43246
rect 26006 43226 26066 44792
rect 25996 43216 26076 43226
rect 25996 43158 26006 43216
rect 26066 43158 26076 43216
rect 25996 43148 26076 43158
rect 26006 42560 26066 43148
rect 26558 43126 26618 44792
rect 26548 43116 26628 43126
rect 26548 43058 26558 43116
rect 26618 43058 26628 43116
rect 26548 43048 26628 43058
rect 26558 42560 26618 43048
rect 27110 43026 27170 44792
rect 27100 43016 27180 43026
rect 27100 42958 27110 43016
rect 27170 42958 27180 43016
rect 27100 42948 27180 42958
rect 27110 42560 27170 42948
rect 27662 42926 27722 44792
rect 27652 42916 27732 42926
rect 27652 42858 27662 42916
rect 27722 42858 27732 42916
rect 27652 42848 27732 42858
rect 27662 42560 27722 42848
rect 23236 42102 23316 42112
rect 23236 42044 23246 42102
rect 23306 42044 23316 42102
rect 23236 42034 23316 42044
rect 23246 41884 23306 42034
rect 200 37748 3138 37754
rect 200 37280 206 37748
rect 594 37280 2904 37748
rect 3132 37280 3138 37748
rect 200 37274 3138 37280
rect 800 37148 3438 37154
rect 800 36680 806 37148
rect 1194 36680 3204 37148
rect 3432 36680 3438 37148
rect 800 36674 3438 36680
rect 19000 35724 19118 35740
rect 19000 35660 19024 35724
rect 19088 35660 19118 35724
rect 19000 35658 19118 35660
rect 19901 35722 19967 35727
rect 19901 35662 19906 35722
rect 19962 35662 19967 35722
rect 19901 35657 19967 35662
rect 200 25034 3138 25040
rect 200 24566 206 25034
rect 594 24566 2904 25034
rect 3132 24566 3138 25034
rect 200 24560 3138 24566
rect 800 24434 3438 24440
rect 800 23966 806 24434
rect 1194 23966 3204 24434
rect 3432 23966 3438 24434
rect 800 23960 3438 23966
rect 200 12320 3138 12326
rect 200 11852 206 12320
rect 594 11852 2904 12320
rect 3132 11852 3138 12320
rect 200 11846 3138 11852
rect 800 11720 3438 11726
rect 800 11252 806 11720
rect 1194 11252 3204 11720
rect 3432 11252 3438 11720
rect 800 11246 3438 11252
rect 19904 590 19964 35657
rect 19896 526 19902 590
rect 19966 526 19972 590
<< via3 >>
rect 20484 44798 20548 44866
rect 21036 44798 21100 44866
rect 21588 44798 21652 44866
rect 22140 44798 22204 44866
rect 22692 44798 22756 44866
rect 23244 44798 23308 44866
rect 23796 44798 23860 44866
rect 24348 44798 24412 44866
rect 24900 44798 24964 44866
rect 25452 44798 25516 44866
rect 26004 44798 26068 44866
rect 26556 44798 26620 44866
rect 27108 44798 27172 44866
rect 27660 44798 27724 44866
rect 206 37280 594 37748
rect 2904 37280 3132 37748
rect 806 36680 1194 37148
rect 3204 36680 3432 37148
rect 19024 35720 19088 35724
rect 19024 35664 19028 35720
rect 19028 35664 19084 35720
rect 19084 35664 19088 35720
rect 19024 35660 19088 35664
rect 206 24566 594 25034
rect 2904 24566 3132 25034
rect 806 23966 1194 24434
rect 3204 23966 3432 24434
rect 206 11852 594 12320
rect 2904 11852 3132 12320
rect 806 11252 1194 11720
rect 3204 11252 3432 11720
rect 19902 526 19966 590
<< metal4 >>
rect 6134 44804 6194 45152
rect 6686 44804 6746 45152
rect 7238 44804 7298 45152
rect 7790 44804 7850 45152
rect 8342 44804 8402 45152
rect 8894 44804 8954 45152
rect 9446 44804 9506 45152
rect 9998 44804 10058 45152
rect 10550 44804 10610 45152
rect 11102 44804 11162 45152
rect 11654 44804 11714 45152
rect 12206 44804 12266 45152
rect 12758 44804 12818 45152
rect 13310 44804 13370 45152
rect 13862 44804 13922 45152
rect 14414 44804 14474 45152
rect 14966 44804 15026 45152
rect 15518 44804 15578 45152
rect 16070 44804 16130 45152
rect 16622 44804 16682 45152
rect 17174 44804 17234 45152
rect 17726 44804 17786 45152
rect 18278 44804 18338 45152
rect 18830 44804 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44872 20546 45152
rect 21038 44872 21098 45152
rect 21590 44872 21650 45152
rect 22142 44872 22202 45152
rect 22694 44872 22754 45152
rect 23246 44872 23306 45152
rect 23798 44872 23858 45152
rect 24350 44872 24410 45152
rect 24902 44872 24962 45152
rect 25454 44872 25514 45152
rect 26006 44872 26066 45152
rect 26558 44872 26618 45152
rect 27110 44872 27170 45152
rect 27662 44872 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 20482 44866 20550 44872
rect 800 44404 18994 44804
rect 20482 44798 20484 44866
rect 20548 44798 20550 44866
rect 20482 44792 20550 44798
rect 21034 44866 21102 44872
rect 21034 44798 21036 44866
rect 21100 44798 21102 44866
rect 21034 44792 21102 44798
rect 21586 44866 21654 44872
rect 21586 44798 21588 44866
rect 21652 44798 21654 44866
rect 21586 44792 21654 44798
rect 22138 44866 22206 44872
rect 22138 44798 22140 44866
rect 22204 44798 22206 44866
rect 22138 44792 22206 44798
rect 22690 44866 22758 44872
rect 22690 44798 22692 44866
rect 22756 44798 22758 44866
rect 22690 44792 22758 44798
rect 23242 44866 23310 44872
rect 23242 44798 23244 44866
rect 23308 44798 23310 44866
rect 23242 44792 23310 44798
rect 23794 44866 23862 44872
rect 23794 44798 23796 44866
rect 23860 44798 23862 44866
rect 23794 44792 23862 44798
rect 24346 44866 24414 44872
rect 24346 44798 24348 44866
rect 24412 44798 24414 44866
rect 24346 44792 24414 44798
rect 24898 44866 24966 44872
rect 24898 44798 24900 44866
rect 24964 44798 24966 44866
rect 24898 44792 24966 44798
rect 25450 44866 25518 44872
rect 25450 44798 25452 44866
rect 25516 44798 25518 44866
rect 25450 44792 25518 44798
rect 26002 44866 26070 44872
rect 26002 44798 26004 44866
rect 26068 44798 26070 44866
rect 26002 44792 26070 44798
rect 26554 44866 26622 44872
rect 26554 44798 26556 44866
rect 26620 44798 26622 44866
rect 26554 44792 26622 44798
rect 27106 44866 27174 44872
rect 27106 44798 27108 44866
rect 27172 44798 27174 44866
rect 27106 44792 27174 44798
rect 27658 44866 27726 44872
rect 27658 44798 27660 44866
rect 27724 44798 27726 44866
rect 27658 44792 27726 44798
rect 200 37748 600 44152
rect 200 37280 206 37748
rect 594 37280 600 37748
rect 200 25034 600 37280
rect 200 24566 206 25034
rect 594 24566 600 25034
rect 200 12320 600 24566
rect 200 11852 206 12320
rect 594 11852 600 12320
rect 200 1000 600 11852
rect 800 37148 1200 44404
rect 2898 37748 3138 37754
rect 2898 37280 2904 37748
rect 3132 37280 3138 37748
rect 2898 37274 3138 37280
rect 800 36680 806 37148
rect 1194 36680 1200 37148
rect 800 24434 1200 36680
rect 3198 37148 3438 37154
rect 3198 36680 3204 37148
rect 3432 36680 3438 37148
rect 3198 36674 3438 36680
rect 19008 35724 19102 35734
rect 19008 35660 19024 35724
rect 19088 35660 19102 35724
rect 19008 35658 19102 35660
rect 19026 35596 19086 35658
rect 19026 35536 19138 35596
rect 17952 26428 30592 26828
rect 2898 25034 3138 25040
rect 2898 24566 2904 25034
rect 3132 24566 3138 25034
rect 2898 24560 3138 24566
rect 800 23966 806 24434
rect 1194 23966 1200 24434
rect 800 11720 1200 23966
rect 3198 24434 3438 24440
rect 3198 23966 3204 24434
rect 3432 23966 3438 24434
rect 3198 23960 3438 23966
rect 17952 13714 26746 14114
rect 2898 12320 3138 12326
rect 2898 11852 2904 12320
rect 3132 11852 3138 12320
rect 2898 11846 3138 11852
rect 800 11252 806 11720
rect 1194 11252 1200 11720
rect 800 1000 1200 11252
rect 3198 11720 3438 11726
rect 3198 11252 3204 11720
rect 3432 11252 3438 11720
rect 3198 11246 3438 11252
rect 17952 1000 22922 1400
rect 26346 1000 26746 13714
rect 30192 1028 30592 26428
rect 19901 590 19967 591
rect 19901 588 19902 590
rect 18834 528 19902 588
rect 18834 200 18894 528
rect 19901 526 19902 528
rect 19966 526 19967 590
rect 19901 525 19967 526
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 1000
rect 26498 0 26678 1000
rect 30362 0 30542 1028
use csdac255  dac_blue
timestamp 1757605323
transform 1 0 4930 0 1 1000
box -2130 0 14808 11424
use csdac255  dac_green
timestamp 1757605323
transform 1 0 4930 0 1 13714
box -2130 0 14808 11424
use csdac255  dac_red
timestamp 1757605323
transform 1 0 4930 0 1 26428
box -2130 0 14808 11424
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
