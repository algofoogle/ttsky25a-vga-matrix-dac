magic
tech sky130A
timestamp 1757512958
<< metal2 >>
rect 173 3651 217 3669
rect -28 3436 0 3450
rect -28 3204 -14 3218
rect -28 2972 -14 2986
rect -28 2740 -14 2754
rect -28 2508 -14 2522
rect -28 2276 -14 2290
rect -28 2044 -14 2058
rect -28 1812 -14 1826
rect -28 1580 -14 1594
rect -28 1348 -14 1362
rect -28 1116 -14 1130
rect -28 884 -14 898
rect -28 652 -14 666
rect -28 420 -14 434
rect -28 188 -14 202
rect 0 -44 39 77
<< metal3 >>
rect 722 4066 760 4069
rect 722 4034 725 4066
rect 757 4034 760 4066
rect 722 4031 760 4034
rect 1115 4066 1153 4069
rect 1115 4034 1118 4066
rect 1150 4034 1153 4066
rect 1115 4031 1153 4034
rect 1508 4066 1546 4069
rect 1508 4034 1511 4066
rect 1543 4034 1546 4066
rect 1508 4031 1546 4034
rect 1901 4066 1939 4069
rect 1901 4034 1904 4066
rect 1936 4034 1939 4066
rect 1901 4031 1939 4034
rect 2294 4066 2332 4069
rect 2294 4034 2297 4066
rect 2329 4034 2332 4066
rect 2294 4031 2332 4034
rect 2687 4066 2725 4069
rect 2687 4034 2690 4066
rect 2722 4034 2725 4066
rect 2687 4031 2725 4034
rect 3080 4066 3118 4069
rect 3080 4034 3083 4066
rect 3115 4034 3118 4066
rect 3080 4031 3118 4034
rect 3473 4066 3511 4069
rect 3473 4034 3476 4066
rect 3508 4034 3511 4066
rect 3473 4031 3511 4034
rect 3866 4066 3904 4069
rect 3866 4034 3869 4066
rect 3901 4034 3904 4066
rect 3866 4031 3904 4034
rect 4259 4066 4297 4069
rect 4259 4034 4262 4066
rect 4294 4034 4297 4066
rect 4259 4031 4297 4034
rect 4652 4066 4690 4069
rect 4652 4034 4655 4066
rect 4687 4034 4690 4066
rect 4652 4031 4690 4034
rect 5045 4066 5083 4069
rect 5045 4034 5048 4066
rect 5080 4034 5083 4066
rect 5045 4031 5083 4034
rect 5438 4066 5476 4069
rect 5438 4034 5441 4066
rect 5473 4034 5476 4066
rect 5438 4031 5476 4034
rect 5831 4066 5869 4069
rect 5831 4034 5834 4066
rect 5866 4034 5869 4066
rect 5831 4031 5869 4034
rect 6224 4066 6262 4069
rect 6224 4034 6227 4066
rect 6259 4034 6262 4066
rect 6224 4031 6262 4034
rect 6617 4066 6655 4069
rect 6617 4034 6620 4066
rect 6652 4034 6655 4066
rect 6617 4031 6655 4034
rect 173 3998 217 4001
rect 173 3884 176 3998
rect 214 3884 217 3998
rect 0 3848 38 3851
rect 0 3734 3 3848
rect 35 3734 38 3848
rect 0 3731 38 3734
rect 0 3700 30 3731
rect 173 3700 217 3884
rect 566 3998 610 4001
rect 566 3884 569 3998
rect 607 3884 610 3998
rect 393 3848 431 3851
rect 393 3734 396 3848
rect 428 3734 431 3848
rect 393 3731 431 3734
rect 393 3700 423 3731
rect 462 3700 492 3753
rect 566 3700 610 3884
rect 726 3700 756 4031
rect 959 3998 1003 4001
rect 959 3884 962 3998
rect 1000 3884 1003 3998
rect 786 3848 824 3851
rect 786 3734 789 3848
rect 821 3734 824 3848
rect 786 3731 824 3734
rect 786 3700 816 3731
rect 855 3700 885 3753
rect 959 3700 1003 3884
rect 1119 3700 1149 4031
rect 1352 3998 1396 4001
rect 1352 3884 1355 3998
rect 1393 3884 1396 3998
rect 1179 3848 1217 3851
rect 1179 3734 1182 3848
rect 1214 3734 1217 3848
rect 1179 3731 1217 3734
rect 1179 3700 1209 3731
rect 1248 3700 1278 3753
rect 1352 3700 1396 3884
rect 1512 3700 1542 4031
rect 1745 3998 1789 4001
rect 1745 3884 1748 3998
rect 1786 3884 1789 3998
rect 1572 3848 1610 3851
rect 1572 3734 1575 3848
rect 1607 3734 1610 3848
rect 1572 3731 1610 3734
rect 1572 3700 1602 3731
rect 1641 3700 1671 3753
rect 1745 3700 1789 3884
rect 1905 3700 1935 4031
rect 2138 3998 2182 4001
rect 2138 3884 2141 3998
rect 2179 3884 2182 3998
rect 1965 3848 2003 3851
rect 1965 3734 1968 3848
rect 2000 3734 2003 3848
rect 1965 3731 2003 3734
rect 1965 3700 1995 3731
rect 2034 3700 2064 3753
rect 2138 3700 2182 3884
rect 2298 3700 2328 4031
rect 2531 3998 2575 4001
rect 2531 3884 2534 3998
rect 2572 3884 2575 3998
rect 2358 3848 2396 3851
rect 2358 3734 2361 3848
rect 2393 3734 2396 3848
rect 2358 3731 2396 3734
rect 2358 3700 2388 3731
rect 2427 3700 2457 3753
rect 2531 3700 2575 3884
rect 2691 3700 2721 4031
rect 2924 3998 2968 4001
rect 2924 3884 2927 3998
rect 2965 3884 2968 3998
rect 2751 3848 2789 3851
rect 2751 3734 2754 3848
rect 2786 3734 2789 3848
rect 2751 3731 2789 3734
rect 2751 3700 2781 3731
rect 2820 3700 2850 3753
rect 2924 3700 2968 3884
rect 3084 3700 3114 4031
rect 3317 3998 3361 4001
rect 3317 3884 3320 3998
rect 3358 3884 3361 3998
rect 3144 3848 3182 3851
rect 3144 3734 3147 3848
rect 3179 3734 3182 3848
rect 3144 3731 3182 3734
rect 3144 3700 3174 3731
rect 3213 3700 3243 3753
rect 3317 3700 3361 3884
rect 3477 3700 3507 4031
rect 3710 3998 3754 4001
rect 3710 3884 3713 3998
rect 3751 3884 3754 3998
rect 3537 3848 3575 3851
rect 3537 3734 3540 3848
rect 3572 3734 3575 3848
rect 3537 3731 3575 3734
rect 3537 3700 3567 3731
rect 3606 3700 3636 3753
rect 3710 3700 3754 3884
rect 3870 3700 3900 4031
rect 4103 3998 4147 4001
rect 4103 3884 4106 3998
rect 4144 3884 4147 3998
rect 3930 3848 3968 3851
rect 3930 3734 3933 3848
rect 3965 3734 3968 3848
rect 3930 3731 3968 3734
rect 3930 3700 3960 3731
rect 3999 3700 4029 3753
rect 4103 3700 4147 3884
rect 4263 3700 4293 4031
rect 4496 3998 4540 4001
rect 4496 3884 4499 3998
rect 4537 3884 4540 3998
rect 4323 3848 4361 3851
rect 4323 3734 4326 3848
rect 4358 3734 4361 3848
rect 4323 3731 4361 3734
rect 4323 3700 4353 3731
rect 4392 3700 4422 3753
rect 4496 3700 4540 3884
rect 4656 3700 4686 4031
rect 4889 3998 4933 4001
rect 4889 3884 4892 3998
rect 4930 3884 4933 3998
rect 4716 3848 4754 3851
rect 4716 3734 4719 3848
rect 4751 3734 4754 3848
rect 4716 3731 4754 3734
rect 4716 3700 4746 3731
rect 4785 3700 4815 3753
rect 4889 3700 4933 3884
rect 5049 3700 5079 4031
rect 5282 3998 5326 4001
rect 5282 3884 5285 3998
rect 5323 3884 5326 3998
rect 5109 3848 5147 3851
rect 5109 3734 5112 3848
rect 5144 3734 5147 3848
rect 5109 3731 5147 3734
rect 5109 3700 5139 3731
rect 5178 3700 5208 3753
rect 5282 3700 5326 3884
rect 5442 3700 5472 4031
rect 5675 3998 5719 4001
rect 5675 3884 5678 3998
rect 5716 3884 5719 3998
rect 5502 3848 5540 3851
rect 5502 3734 5505 3848
rect 5537 3734 5540 3848
rect 5502 3731 5540 3734
rect 5502 3700 5532 3731
rect 5571 3700 5601 3753
rect 5675 3700 5719 3884
rect 5835 3700 5865 4031
rect 6068 3998 6112 4001
rect 6068 3884 6071 3998
rect 6109 3884 6112 3998
rect 5895 3848 5933 3851
rect 5895 3734 5898 3848
rect 5930 3734 5933 3848
rect 5895 3731 5933 3734
rect 5895 3700 5925 3731
rect 5964 3700 5994 3753
rect 6068 3700 6112 3884
rect 6228 3700 6258 4031
rect 6461 3998 6505 4001
rect 6461 3884 6464 3998
rect 6502 3884 6505 3998
rect 6288 3848 6326 3851
rect 6288 3734 6291 3848
rect 6323 3734 6326 3848
rect 6288 3731 6326 3734
rect 6288 3700 6318 3731
rect 6461 3700 6505 3884
rect 6621 3700 6651 4031
rect 6854 3998 6898 4001
rect 6854 3884 6857 3998
rect 6895 3884 6898 3998
rect 6681 3848 6719 3851
rect 6681 3734 6684 3848
rect 6716 3734 6719 3848
rect 6681 3731 6719 3734
rect 6681 3700 6711 3731
rect 6854 3700 6898 3884
rect 0 -23 30 8
rect 0 -26 38 -23
rect 0 -140 3 -26
rect 35 -140 38 -26
rect 0 -143 38 -140
rect 173 -176 217 8
rect 393 -23 423 8
rect 393 -26 431 -23
rect 393 -140 396 -26
rect 428 -140 431 -26
rect 393 -143 431 -140
rect 173 -290 176 -176
rect 214 -290 217 -176
rect 173 -293 217 -290
rect 566 -176 610 8
rect 566 -290 569 -176
rect 607 -290 610 -176
rect 566 -293 610 -290
rect 653 -323 683 4
rect 786 -23 816 8
rect 786 -26 824 -23
rect 786 -140 789 -26
rect 821 -140 824 -26
rect 786 -143 824 -140
rect 959 -176 1003 8
rect 959 -290 962 -176
rect 1000 -290 1003 -176
rect 959 -293 1003 -290
rect 1046 -323 1076 4
rect 1179 -23 1209 8
rect 1179 -26 1217 -23
rect 1179 -140 1182 -26
rect 1214 -140 1217 -26
rect 1179 -143 1217 -140
rect 1352 -176 1396 8
rect 1352 -290 1355 -176
rect 1393 -290 1396 -176
rect 1352 -293 1396 -290
rect 1439 -323 1469 4
rect 1572 -23 1602 8
rect 1572 -26 1610 -23
rect 1572 -140 1575 -26
rect 1607 -140 1610 -26
rect 1572 -143 1610 -140
rect 1745 -176 1789 8
rect 1745 -290 1748 -176
rect 1786 -290 1789 -176
rect 1745 -293 1789 -290
rect 1832 -323 1862 4
rect 1965 -23 1995 8
rect 1965 -26 2003 -23
rect 1965 -140 1968 -26
rect 2000 -140 2003 -26
rect 1965 -143 2003 -140
rect 2138 -176 2182 8
rect 2138 -290 2141 -176
rect 2179 -290 2182 -176
rect 2138 -293 2182 -290
rect 2225 -323 2255 4
rect 2358 -23 2388 8
rect 2358 -26 2396 -23
rect 2358 -140 2361 -26
rect 2393 -140 2396 -26
rect 2358 -143 2396 -140
rect 2531 -176 2575 8
rect 2531 -290 2534 -176
rect 2572 -290 2575 -176
rect 2531 -293 2575 -290
rect 2618 -323 2648 4
rect 2751 -23 2781 8
rect 2751 -26 2789 -23
rect 2751 -140 2754 -26
rect 2786 -140 2789 -26
rect 2751 -143 2789 -140
rect 2924 -176 2968 8
rect 2924 -290 2927 -176
rect 2965 -290 2968 -176
rect 2924 -293 2968 -290
rect 3011 -323 3041 4
rect 3144 -23 3174 8
rect 3144 -26 3182 -23
rect 3144 -140 3147 -26
rect 3179 -140 3182 -26
rect 3144 -143 3182 -140
rect 3317 -176 3361 8
rect 3317 -290 3320 -176
rect 3358 -290 3361 -176
rect 3317 -293 3361 -290
rect 3404 -323 3434 4
rect 3537 -23 3567 8
rect 3537 -26 3575 -23
rect 3537 -140 3540 -26
rect 3572 -140 3575 -26
rect 3537 -143 3575 -140
rect 3710 -176 3754 8
rect 3710 -290 3713 -176
rect 3751 -290 3754 -176
rect 3710 -293 3754 -290
rect 3797 -323 3827 4
rect 3930 -23 3960 8
rect 3930 -26 3968 -23
rect 3930 -140 3933 -26
rect 3965 -140 3968 -26
rect 3930 -143 3968 -140
rect 4103 -176 4147 8
rect 4103 -290 4106 -176
rect 4144 -290 4147 -176
rect 4103 -293 4147 -290
rect 4190 -323 4220 4
rect 4323 -23 4353 8
rect 4323 -26 4361 -23
rect 4323 -140 4326 -26
rect 4358 -140 4361 -26
rect 4323 -143 4361 -140
rect 4496 -176 4540 8
rect 4496 -290 4499 -176
rect 4537 -290 4540 -176
rect 4496 -293 4540 -290
rect 4583 -323 4613 4
rect 4716 -23 4746 8
rect 4716 -26 4754 -23
rect 4716 -140 4719 -26
rect 4751 -140 4754 -26
rect 4716 -143 4754 -140
rect 4889 -176 4933 8
rect 4889 -290 4892 -176
rect 4930 -290 4933 -176
rect 4889 -293 4933 -290
rect 4976 -323 5006 4
rect 5109 -23 5139 8
rect 5109 -26 5147 -23
rect 5109 -140 5112 -26
rect 5144 -140 5147 -26
rect 5109 -143 5147 -140
rect 5282 -176 5326 8
rect 5282 -290 5285 -176
rect 5323 -290 5326 -176
rect 5282 -293 5326 -290
rect 5369 -323 5399 4
rect 5502 -23 5532 8
rect 5502 -26 5540 -23
rect 5502 -140 5505 -26
rect 5537 -140 5540 -26
rect 5502 -143 5540 -140
rect 5675 -176 5719 8
rect 5675 -290 5678 -176
rect 5716 -290 5719 -176
rect 5675 -293 5719 -290
rect 5762 -323 5792 4
rect 5895 -23 5925 8
rect 5895 -26 5933 -23
rect 5895 -140 5898 -26
rect 5930 -140 5933 -26
rect 5895 -143 5933 -140
rect 6068 -176 6112 8
rect 6068 -290 6071 -176
rect 6109 -290 6112 -176
rect 6068 -293 6112 -290
rect 6155 -323 6185 4
rect 6288 -23 6318 8
rect 6288 -26 6326 -23
rect 6288 -140 6291 -26
rect 6323 -140 6326 -26
rect 6288 -143 6326 -140
rect 6461 -176 6505 8
rect 6461 -290 6464 -176
rect 6502 -290 6505 -176
rect 6461 -293 6505 -290
rect 6548 -323 6578 4
rect 6681 -23 6711 8
rect 6681 -26 6719 -23
rect 6681 -140 6684 -26
rect 6716 -140 6719 -26
rect 6681 -143 6719 -140
rect 6854 -176 6898 8
rect 6854 -290 6857 -176
rect 6895 -290 6898 -176
rect 6854 -293 6898 -290
rect 653 -326 691 -323
rect 653 -520 656 -326
rect 688 -520 691 -326
rect 653 -523 691 -520
rect 1046 -326 1084 -323
rect 1046 -520 1049 -326
rect 1081 -520 1084 -326
rect 1046 -523 1084 -520
rect 1439 -326 1477 -323
rect 1439 -520 1442 -326
rect 1474 -520 1477 -326
rect 1439 -523 1477 -520
rect 1832 -326 1870 -323
rect 1832 -520 1835 -326
rect 1867 -520 1870 -326
rect 1832 -523 1870 -520
rect 2225 -326 2263 -323
rect 2225 -520 2228 -326
rect 2260 -520 2263 -326
rect 2225 -523 2263 -520
rect 2618 -326 2656 -323
rect 2618 -520 2621 -326
rect 2653 -520 2656 -326
rect 2618 -523 2656 -520
rect 3011 -326 3049 -323
rect 3011 -520 3014 -326
rect 3046 -520 3049 -326
rect 3011 -523 3049 -520
rect 3404 -326 3442 -323
rect 3404 -520 3407 -326
rect 3439 -520 3442 -326
rect 3404 -523 3442 -520
rect 3797 -326 3835 -323
rect 3797 -520 3800 -326
rect 3832 -520 3835 -326
rect 3797 -523 3835 -520
rect 4190 -326 4228 -323
rect 4190 -520 4193 -326
rect 4225 -520 4228 -326
rect 4190 -523 4228 -520
rect 4583 -326 4621 -323
rect 4583 -520 4586 -326
rect 4618 -520 4621 -326
rect 4583 -523 4621 -520
rect 4976 -326 5014 -323
rect 4976 -520 4979 -326
rect 5011 -520 5014 -326
rect 4976 -523 5014 -520
rect 5369 -326 5407 -323
rect 5369 -520 5372 -326
rect 5404 -520 5407 -326
rect 5369 -523 5407 -520
rect 5762 -326 5800 -323
rect 5762 -520 5765 -326
rect 5797 -520 5800 -326
rect 5762 -523 5800 -520
rect 6155 -326 6193 -323
rect 6155 -520 6158 -326
rect 6190 -520 6193 -326
rect 6155 -523 6193 -520
rect 6548 -326 6586 -323
rect 6548 -520 6551 -326
rect 6583 -520 6586 -326
rect 6548 -523 6586 -520
<< via3 >>
rect 725 4034 757 4066
rect 1118 4034 1150 4066
rect 1511 4034 1543 4066
rect 1904 4034 1936 4066
rect 2297 4034 2329 4066
rect 2690 4034 2722 4066
rect 3083 4034 3115 4066
rect 3476 4034 3508 4066
rect 3869 4034 3901 4066
rect 4262 4034 4294 4066
rect 4655 4034 4687 4066
rect 5048 4034 5080 4066
rect 5441 4034 5473 4066
rect 5834 4034 5866 4066
rect 6227 4034 6259 4066
rect 6620 4034 6652 4066
rect 176 3884 214 3998
rect 3 3734 35 3848
rect 569 3884 607 3998
rect 396 3734 428 3848
rect 962 3884 1000 3998
rect 789 3734 821 3848
rect 1355 3884 1393 3998
rect 1182 3734 1214 3848
rect 1748 3884 1786 3998
rect 1575 3734 1607 3848
rect 2141 3884 2179 3998
rect 1968 3734 2000 3848
rect 2534 3884 2572 3998
rect 2361 3734 2393 3848
rect 2927 3884 2965 3998
rect 2754 3734 2786 3848
rect 3320 3884 3358 3998
rect 3147 3734 3179 3848
rect 3713 3884 3751 3998
rect 3540 3734 3572 3848
rect 4106 3884 4144 3998
rect 3933 3734 3965 3848
rect 4499 3884 4537 3998
rect 4326 3734 4358 3848
rect 4892 3884 4930 3998
rect 4719 3734 4751 3848
rect 5285 3884 5323 3998
rect 5112 3734 5144 3848
rect 5678 3884 5716 3998
rect 5505 3734 5537 3848
rect 6071 3884 6109 3998
rect 5898 3734 5930 3848
rect 6464 3884 6502 3998
rect 6291 3734 6323 3848
rect 6857 3884 6895 3998
rect 6684 3734 6716 3848
rect 3 -140 35 -26
rect 396 -140 428 -26
rect 176 -290 214 -176
rect 569 -290 607 -176
rect 789 -140 821 -26
rect 962 -290 1000 -176
rect 1182 -140 1214 -26
rect 1355 -290 1393 -176
rect 1575 -140 1607 -26
rect 1748 -290 1786 -176
rect 1968 -140 2000 -26
rect 2141 -290 2179 -176
rect 2361 -140 2393 -26
rect 2534 -290 2572 -176
rect 2754 -140 2786 -26
rect 2927 -290 2965 -176
rect 3147 -140 3179 -26
rect 3320 -290 3358 -176
rect 3540 -140 3572 -26
rect 3713 -290 3751 -176
rect 3933 -140 3965 -26
rect 4106 -290 4144 -176
rect 4326 -140 4358 -26
rect 4499 -290 4537 -176
rect 4719 -140 4751 -26
rect 4892 -290 4930 -176
rect 5112 -140 5144 -26
rect 5285 -290 5323 -176
rect 5505 -140 5537 -26
rect 5678 -290 5716 -176
rect 5898 -140 5930 -26
rect 6071 -290 6109 -176
rect 6291 -140 6323 -26
rect 6464 -290 6502 -176
rect 6684 -140 6716 -26
rect 6857 -290 6895 -176
rect 656 -520 688 -326
rect 1049 -520 1081 -326
rect 1442 -520 1474 -326
rect 1835 -520 1867 -326
rect 2228 -520 2260 -326
rect 2621 -520 2653 -326
rect 3014 -520 3046 -326
rect 3407 -520 3439 -326
rect 3800 -520 3832 -326
rect 4193 -520 4225 -326
rect 4586 -520 4618 -326
rect 4979 -520 5011 -326
rect 5372 -520 5404 -326
rect 5765 -520 5797 -326
rect 6158 -520 6190 -326
rect 6551 -520 6583 -326
<< metal4 >>
rect 722 4066 760 4069
rect 722 4061 725 4066
rect -30 4034 725 4061
rect 757 4061 760 4066
rect 1115 4066 1153 4069
rect 1115 4061 1118 4066
rect 757 4034 1118 4061
rect 1150 4061 1153 4066
rect 1508 4066 1546 4069
rect 1508 4061 1511 4066
rect 1150 4034 1511 4061
rect 1543 4061 1546 4066
rect 1901 4066 1939 4069
rect 1901 4061 1904 4066
rect 1543 4034 1904 4061
rect 1936 4061 1939 4066
rect 2294 4066 2332 4069
rect 2294 4061 2297 4066
rect 1936 4034 2297 4061
rect 2329 4061 2332 4066
rect 2687 4066 2725 4069
rect 2687 4061 2690 4066
rect 2329 4034 2690 4061
rect 2722 4061 2725 4066
rect 3080 4066 3118 4069
rect 3080 4061 3083 4066
rect 2722 4034 3083 4061
rect 3115 4061 3118 4066
rect 3473 4066 3511 4069
rect 3473 4061 3476 4066
rect 3115 4034 3476 4061
rect 3508 4061 3511 4066
rect 3866 4066 3904 4069
rect 3866 4061 3869 4066
rect 3508 4034 3869 4061
rect 3901 4061 3904 4066
rect 4259 4066 4297 4069
rect 4259 4061 4262 4066
rect 3901 4034 4262 4061
rect 4294 4061 4297 4066
rect 4652 4066 4690 4069
rect 4652 4061 4655 4066
rect 4294 4034 4655 4061
rect 4687 4061 4690 4066
rect 5045 4066 5083 4069
rect 5045 4061 5048 4066
rect 4687 4034 5048 4061
rect 5080 4061 5083 4066
rect 5438 4066 5476 4069
rect 5438 4061 5441 4066
rect 5080 4034 5441 4061
rect 5473 4061 5476 4066
rect 5831 4066 5869 4069
rect 5831 4061 5834 4066
rect 5473 4034 5834 4061
rect 5866 4061 5869 4066
rect 6224 4066 6262 4069
rect 6224 4061 6227 4066
rect 5866 4034 6227 4061
rect 6259 4061 6262 4066
rect 6617 4066 6655 4069
rect 6617 4061 6620 4066
rect 6259 4034 6620 4061
rect 6652 4061 6655 4066
rect 6652 4034 7074 4061
rect -30 4031 7074 4034
rect -30 3998 7374 4001
rect -30 3884 176 3998
rect 214 3884 569 3998
rect 607 3884 962 3998
rect 1000 3884 1355 3998
rect 1393 3884 1748 3998
rect 1786 3884 2141 3998
rect 2179 3884 2534 3998
rect 2572 3884 2927 3998
rect 2965 3884 3320 3998
rect 3358 3884 3713 3998
rect 3751 3884 4106 3998
rect 4144 3884 4499 3998
rect 4537 3884 4892 3998
rect 4930 3884 5285 3998
rect 5323 3884 5678 3998
rect 5716 3884 6071 3998
rect 6109 3884 6464 3998
rect 6502 3884 6857 3998
rect 6895 3884 7374 3998
rect -30 3881 7374 3884
rect -30 3848 7224 3851
rect -30 3734 3 3848
rect 35 3734 396 3848
rect 428 3734 789 3848
rect 821 3734 1182 3848
rect 1214 3734 1575 3848
rect 1607 3734 1968 3848
rect 2000 3734 2361 3848
rect 2393 3734 2754 3848
rect 2786 3734 3147 3848
rect 3179 3734 3540 3848
rect 3572 3734 3933 3848
rect 3965 3734 4326 3848
rect 4358 3734 4719 3848
rect 4751 3734 5112 3848
rect 5144 3734 5505 3848
rect 5537 3734 5898 3848
rect 5930 3734 6291 3848
rect 6323 3734 6684 3848
rect 6716 3734 7224 3848
rect -30 3731 7224 3734
rect 7104 -23 7224 3731
rect -30 -26 7224 -23
rect -30 -140 3 -26
rect 35 -140 396 -26
rect 428 -140 789 -26
rect 821 -140 1182 -26
rect 1214 -140 1575 -26
rect 1607 -140 1968 -26
rect 2000 -140 2361 -26
rect 2393 -140 2754 -26
rect 2786 -140 3147 -26
rect 3179 -140 3540 -26
rect 3572 -140 3933 -26
rect 3965 -140 4326 -26
rect 4358 -140 4719 -26
rect 4751 -140 5112 -26
rect 5144 -140 5505 -26
rect 5537 -140 5898 -26
rect 5930 -140 6291 -26
rect 6323 -140 6684 -26
rect 6716 -140 7224 -26
rect -30 -143 7224 -140
rect 7254 -173 7374 3881
rect -30 -176 7374 -173
rect -30 -290 176 -176
rect 214 -290 569 -176
rect 607 -290 962 -176
rect 1000 -290 1355 -176
rect 1393 -290 1748 -176
rect 1786 -290 2141 -176
rect 2179 -290 2534 -176
rect 2572 -290 2927 -176
rect 2965 -290 3320 -176
rect 3358 -290 3713 -176
rect 3751 -290 4106 -176
rect 4144 -290 4499 -176
rect 4537 -290 4892 -176
rect 4930 -290 5285 -176
rect 5323 -290 5678 -176
rect 5716 -290 6071 -176
rect 6109 -290 6464 -176
rect 6502 -290 6857 -176
rect 6895 -290 7374 -176
rect -30 -293 7374 -290
rect 393 -326 6681 -323
rect 393 -520 656 -326
rect 688 -520 1049 -326
rect 1081 -520 1442 -326
rect 1474 -520 1835 -326
rect 1867 -520 2228 -326
rect 2260 -520 2621 -326
rect 2653 -520 3014 -326
rect 3046 -520 3407 -326
rect 3439 -520 3800 -326
rect 3832 -520 4193 -326
rect 4225 -520 4586 -326
rect 4618 -520 4979 -326
rect 5011 -520 5372 -326
rect 5404 -520 5765 -326
rect 5797 -520 6158 -326
rect 6190 -520 6551 -326
rect 6583 -520 6681 -326
rect 393 -523 6681 -520
use row15x  XIR
array 1 1 7074 15 0 232
timestamp 1757512958
transform 1 0 0 0 1 0
box -28 -55 7074 243
<< labels >>
flabel metal2 -28 3436 -14 3450 0 FreeSans 40 0 0 0 Rn[0]
port 0 nsew
flabel metal2 -28 3204 -14 3218 0 FreeSans 40 0 0 0 Rn[1]
port 1 nsew
flabel metal2 -28 2972 -14 2986 0 FreeSans 40 0 0 0 Rn[2]
port 2 nsew
flabel metal2 -28 2740 -14 2754 0 FreeSans 40 0 0 0 Rn[3]
port 3 nsew
flabel metal2 -28 2508 -14 2522 0 FreeSans 40 0 0 0 Rn[4]
port 4 nsew
flabel metal2 -28 2276 -14 2290 0 FreeSans 40 0 0 0 Rn[5]
port 5 nsew
flabel metal2 -28 2044 -14 2058 0 FreeSans 40 0 0 0 Rn[6]
port 6 nsew
flabel metal2 -28 1812 -14 1826 0 FreeSans 40 0 0 0 Rn[7]
port 7 nsew
flabel metal2 -28 1580 -14 1594 0 FreeSans 40 0 0 0 Rn[8]
port 8 nsew
flabel metal2 -28 1348 -14 1362 0 FreeSans 40 0 0 0 Rn[9]
port 9 nsew
flabel metal2 -28 1116 -14 1130 0 FreeSans 40 0 0 0 Rn[10]
port 10 nsew
flabel metal2 -28 884 -14 898 0 FreeSans 40 0 0 0 Rn[11]
port 11 nsew
flabel metal2 -28 652 -14 666 0 FreeSans 40 0 0 0 Rn[12]
port 12 nsew
flabel metal2 -28 420 -14 434 0 FreeSans 40 0 0 0 Rn[13]
port 13 nsew
flabel metal2 -28 188 -14 202 0 FreeSans 40 0 0 0 Rn[14]
port 14 nsew
flabel metal3 462 3738 492 3753 0 FreeSans 40 0 0 0 Cn[0]
port 100 nsew
flabel metal3 855 3738 885 3753 0 FreeSans 40 0 0 0 Cn[1]
port 101 nsew
flabel metal3 1248 3738 1278 3753 0 FreeSans 40 0 0 0 Cn[2]
port 102 nsew
flabel metal3 1641 3738 1671 3753 0 FreeSans 40 0 0 0 Cn[3]
port 103 nsew
flabel metal3 2034 3738 2064 3753 0 FreeSans 40 0 0 0 Cn[4]
port 104 nsew
flabel metal3 2427 3738 2457 3753 0 FreeSans 40 0 0 0 Cn[5]
port 105 nsew
flabel metal3 2820 3738 2850 3753 0 FreeSans 40 0 0 0 Cn[6]
port 106 nsew
flabel metal3 3213 3738 3243 3753 0 FreeSans 40 0 0 0 Cn[7]
port 107 nsew
flabel metal3 3606 3738 3636 3753 0 FreeSans 40 0 0 0 Cn[8]
port 108 nsew
flabel metal3 3999 3738 4029 3753 0 FreeSans 40 0 0 0 Cn[9]
port 109 nsew
flabel metal3 4392 3738 4422 3753 0 FreeSans 40 0 0 0 Cn[10]
port 110 nsew
flabel metal3 4785 3738 4815 3753 0 FreeSans 40 0 0 0 Cn[11]
port 111 nsew
flabel metal3 5178 3738 5208 3753 0 FreeSans 40 0 0 0 Cn[12]
port 112 nsew
flabel metal3 5571 3738 5601 3753 0 FreeSans 40 0 0 0 Cn[13]
port 113 nsew
flabel metal3 5964 3738 5994 3753 0 FreeSans 40 0 0 0 Cn[14]
port 114 nsew
flabel metal4 -30 3731 0 3851 0 FreeSans 80 90 0 0 VPWR
port 201 nsew
flabel metal4 -30 4031 0 4061 0 FreeSans 80 90 0 0 Vbias
port 202 nsew
flabel metal4 6581 -523 6681 -423 0 FreeSans 80 0 0 0 Iout
port 203 nsew
flabel metal4 -30 3881 0 4001 0 FreeSans 80 90 0 0 VGND
port 200 nsew
<< end >>
