magic
tech sky130A
magscale 1 2
timestamp 1757605323
<< metal1 >>
rect -1412 10662 -1368 11424
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect -1330 10662 -1192 10750
rect -814 10662 -768 11424
rect -474 10662 -428 11424
rect 7490 11384 7530 11424
rect 7572 11384 7612 11424
rect 9138 11384 9178 11424
rect 9748 11384 9788 11424
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect 684 10662 1268 10796
rect -2130 4230 -2090 4270
rect -2130 4148 -2090 4188
rect -2130 2582 -2090 2622
rect -2130 1972 -2090 2012
<< via1 >>
rect -1320 10750 -1202 11316
rect 694 10796 1258 11016
<< metal2 >>
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect 684 10786 1268 10796
rect -1330 10740 -1192 10750
rect 808 9650 886 9734
rect 788 9640 906 9650
rect 788 9118 798 9640
rect 896 9118 906 9640
rect 3182 9630 3238 9639
rect 3436 9632 3492 9639
rect 3182 9565 3238 9574
rect 3434 9630 3680 9632
rect 3434 9574 3436 9630
rect 3492 9574 3680 9630
rect 3434 9572 3680 9574
rect 3436 9565 3492 9572
rect 3620 9490 3680 9572
rect 4233 9568 4242 9624
rect 4298 9568 4307 9624
rect 4862 9238 4922 9610
rect 8524 9506 8580 9515
rect 3342 9236 4922 9238
rect 3335 9180 3344 9236
rect 3400 9180 4922 9236
rect 3342 9178 4922 9180
rect 5654 9136 5714 9414
rect 4128 9134 5714 9136
rect 788 9108 906 9118
rect 4121 9078 4130 9134
rect 4186 9078 5714 9134
rect 4128 9076 5714 9078
rect 6120 9018 6180 9426
rect 4914 9016 6180 9018
rect 4907 8960 4916 9016
rect 4972 8960 6180 9016
rect 4914 8958 6180 8960
rect 5702 8912 5758 8919
rect 6582 8912 6642 9396
rect 5700 8910 6642 8912
rect 5700 8854 5702 8910
rect 5758 8854 6642 8910
rect 5700 8852 6642 8854
rect 5702 8845 5758 8852
rect 6526 8802 6582 8809
rect 7044 8802 7104 9506
rect 7424 9492 7480 9501
rect 7424 9427 7480 9436
rect 8198 9462 8254 9471
rect 9604 9500 9660 9509
rect 8524 9441 8580 9450
rect 9245 9414 9254 9470
rect 9310 9414 9319 9470
rect 9604 9435 9660 9444
rect 10332 9470 10388 9479
rect 8198 9397 8254 9406
rect 10332 9405 10388 9414
rect 11346 9396 11402 9403
rect 10702 9394 11404 9396
rect 10702 9338 11346 9394
rect 11402 9338 11404 9394
rect 10702 9336 11404 9338
rect 11346 9329 11402 9336
rect 6524 8800 7104 8802
rect 6524 8744 6526 8800
rect 6582 8744 7104 8800
rect 6524 8742 7104 8744
rect 6526 8735 6582 8742
rect -44 7912 16 7952
rect -44 7448 16 7488
rect -44 6984 16 7024
rect -44 6520 16 6560
rect -44 6056 16 6096
rect -44 5592 16 5632
rect -44 5128 16 5168
rect -44 4664 16 4704
rect -44 4200 16 4240
rect -44 3736 16 3776
rect -44 3272 16 3312
rect -44 2808 16 2848
rect -44 2344 16 2384
rect -44 1880 16 1920
rect -44 1416 16 1456
<< via2 >>
rect -1320 10750 -1202 11316
rect 694 10796 1258 11016
rect 798 9118 896 9640
rect 3182 9574 3238 9630
rect 3436 9574 3492 9630
rect 4242 9568 4298 9624
rect 3344 9180 3400 9236
rect 4130 9078 4186 9134
rect 4916 8960 4972 9016
rect 5702 8854 5758 8910
rect 7424 9436 7480 9492
rect 8198 9406 8254 9462
rect 8524 9450 8580 9506
rect 9254 9414 9310 9470
rect 9604 9444 9660 9500
rect 10332 9414 10388 9470
rect 11346 9338 11402 9394
rect 6526 8744 6582 8800
<< metal3 >>
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect 14268 11320 14508 11326
rect 14268 11092 14274 11320
rect 14502 11092 14508 11320
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect 684 10786 1268 10796
rect -1330 10740 -1192 10750
rect 788 9640 906 9650
rect 788 9118 798 9640
rect 896 9118 906 9640
rect 3177 9632 3243 9635
rect 788 9108 906 9118
rect 984 9630 3243 9632
rect 984 9574 3182 9630
rect 3238 9574 3243 9630
rect 984 9572 3243 9574
rect 984 8492 1044 9572
rect 3177 9569 3243 9572
rect 3431 9630 3497 9635
rect 3431 9574 3436 9630
rect 3492 9574 3497 9630
rect 3431 9569 3497 9574
rect 4237 9624 4303 9629
rect 3434 9496 3494 9569
rect 4237 9568 4242 9624
rect 4298 9568 4303 9624
rect 4237 9563 4303 9568
rect 1770 9436 3494 9496
rect 1770 8492 1830 9436
rect 4240 9368 4300 9563
rect 8519 9508 8585 9511
rect 8519 9506 8904 9508
rect 7419 9494 7485 9497
rect 2556 9308 4300 9368
rect 7272 9492 7485 9494
rect 7272 9436 7424 9492
rect 7480 9436 7485 9492
rect 8193 9464 8259 9467
rect 7272 9434 7485 9436
rect 2556 8492 2616 9308
rect 3339 9236 3405 9241
rect 3339 9180 3344 9236
rect 3400 9180 3405 9236
rect 3339 9175 3405 9180
rect 3342 8492 3402 9175
rect 4125 9134 4191 9139
rect 4125 9078 4130 9134
rect 4186 9078 4191 9134
rect 4125 9073 4191 9078
rect 4128 8492 4188 9073
rect 4911 9016 4977 9021
rect 4911 8960 4916 9016
rect 4972 8960 4977 9016
rect 4911 8955 4977 8960
rect 4914 8492 4974 8955
rect 5697 8910 5763 8915
rect 5697 8854 5702 8910
rect 5758 8854 5763 8910
rect 5697 8849 5763 8854
rect 5700 8492 5760 8849
rect 6521 8802 6587 8805
rect 6486 8800 6587 8802
rect 6486 8744 6526 8800
rect 6582 8744 6587 8800
rect 6486 8739 6587 8744
rect 6486 8492 6546 8739
rect 7272 8492 7332 9434
rect 7419 9431 7485 9434
rect 8058 9462 8259 9464
rect 8058 9406 8198 9462
rect 8254 9406 8259 9462
rect 8519 9450 8524 9506
rect 8580 9450 8904 9506
rect 9599 9502 9665 9505
rect 9599 9500 9994 9502
rect 8519 9448 8904 9450
rect 8519 9445 8585 9448
rect 8058 9404 8259 9406
rect 8058 8492 8118 9404
rect 8193 9401 8259 9404
rect 8844 8492 8904 9448
rect 9249 9470 9315 9475
rect 9249 9414 9254 9470
rect 9310 9414 9315 9470
rect 9599 9444 9604 9500
rect 9660 9444 9994 9500
rect 9599 9442 9994 9444
rect 9599 9439 9665 9442
rect 9249 9409 9315 9414
rect 9252 9320 9312 9409
rect 9934 9322 9994 9442
rect 10327 9472 10393 9475
rect 10327 9470 11262 9472
rect 10327 9414 10332 9470
rect 10388 9414 11262 9470
rect 10327 9412 11262 9414
rect 10327 9409 10393 9412
rect 9252 9260 9690 9320
rect 9934 9262 10476 9322
rect 9630 8492 9690 9260
rect 10416 8492 10476 9262
rect 11202 8492 11262 9412
rect 11341 9396 11407 9399
rect 11341 9394 12048 9396
rect 11341 9338 11346 9394
rect 11402 9338 12048 9394
rect 11341 9336 12048 9338
rect 11341 9333 11407 9336
rect 11988 8492 12048 9336
rect 14268 8742 14508 11092
rect 14268 8514 14274 8742
rect 14502 8514 14508 8742
rect 14268 8508 14508 8514
rect -1385 1050 -1147 1055
rect -2038 810 -2032 1050
rect -1794 1049 -1146 1050
rect -1794 811 -1385 1049
rect -1147 811 -1146 1049
rect -1794 810 -1146 811
rect -1385 805 -1147 810
<< via3 >>
rect -1320 11096 -1202 11316
rect 14274 11092 14502 11320
rect 694 10796 1258 11016
rect 798 9118 896 9640
rect 14274 8514 14502 8742
rect -2032 810 -1794 1050
rect -1385 811 -1147 1049
<< metal4 >>
rect -2032 11316 3228 11326
rect -2032 11096 -1320 11316
rect -1202 11096 3228 11316
rect -2032 11086 3228 11096
rect 10900 11320 14508 11326
rect 10900 11092 14274 11320
rect 14502 11092 14508 11320
rect 10900 11086 14508 11092
rect -2032 8680 -1792 11086
rect -1732 11016 3212 11026
rect -1732 10796 694 11016
rect 1258 10796 3212 11016
rect -1732 10786 3212 10796
rect 10810 10786 14808 11026
rect -1732 8680 -1492 10786
rect 788 9640 906 9650
rect 788 9118 798 9640
rect 896 9118 906 9640
rect 788 9108 906 9118
rect 14066 9108 14208 9168
rect 14568 8694 14808 10786
rect -2033 1050 -1793 1051
rect -2033 810 -2032 1050
rect -1794 810 -1793 1050
rect -1386 1049 -518 1050
rect -2033 809 -1793 810
rect -1732 700 -1492 950
rect -1386 811 -1385 1049
rect -1147 1000 -518 1049
rect -1147 811 370 1000
rect -1386 810 370 811
rect -758 760 370 810
rect -1732 460 202 700
rect 13022 0 13422 400
use array255x  XA
timestamp 1757605323
transform 1 0 60 0 1 1046
box -60 -1046 14748 8138
use thermo15  XThC
timestamp 1757605323
transform 0 -1 3524 -1 0 10408
box -1016 -7616 1090 640
use thermo15  XThR
timestamp 1757605323
transform 1 0 -1114 0 1 8236
box -1016 -7616 1090 640
use vbias  XVB
timestamp 1757605323
transform 1 0 -1412 0 1 9690
box 0 0 2716 1016
<< labels >>
flabel metal4 13022 0 13422 400 0 FreeSans 1600 0 0 0 Iout
port 0 nsew
flabel metal4 -2032 11086 3228 11326 0 FreeSans 1600 0 0 0 VPWR
port 1 nsew
flabel metal4 -1732 10786 3212 11026 0 FreeSans 1600 0 0 0 VGND
port 2 nsew
flabel metal4 14066 9108 14208 9168 0 FreeSans 160 0 0 0 Vbias
port 3 nsew
flabel metal1 -1412 11380 -1368 11424 0 FreeSans 80 0 0 0 bias[2]
port 5 nsew
flabel metal1 -814 11380 -768 11424 0 FreeSans 80 0 0 0 bias[1]
port 6 nsew
flabel metal1 -474 11380 -428 11424 0 FreeSans 80 0 0 0 bias[0]
port 7 nsew
flabel metal1 -2130 1972 -2090 2012 0 FreeSans 80 0 0 0 data[7]
port 1807 nsew
flabel metal1 -2130 2582 -2090 2622 0 FreeSans 80 0 0 0 data[6]
port 1806 nsew
flabel metal1 -2130 4148 -2090 4188 0 FreeSans 80 0 0 0 data[5]
port 1805 nsew
flabel metal1 -2130 4230 -2090 4270 0 FreeSans 80 0 0 0 data[4]
port 1804 nsew
flabel metal1 9748 11384 9788 11424 0 FreeSans 80 0 0 0 data[3]
port 1803 nsew
flabel metal1 9138 11384 9178 11424 0 FreeSans 80 0 0 0 data[2]
port 1802 nsew
flabel metal1 7572 11384 7612 11424 0 FreeSans 80 0 0 0 data[1]
port 1801 nsew
flabel metal1 7490 11384 7530 11424 0 FreeSans 80 0 0 0 data[0]
port 1800 nsew
<< end >>
