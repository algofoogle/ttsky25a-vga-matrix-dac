* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias bias[2] bias[1] bias[0] data[0] data[1]
+ data[2] data[3] data[4] data[5] data[6] data[7]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1753 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t781 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t780 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t103 VGND.t775 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1793 VPWR.t1795 VPWR.t1794 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t1737 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t1736 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t2489 XThR.TBN.t4 a_n997_2667# VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t351 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t311 VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t11 XThC.TBN.t4 VGND.t2057 VGND.t2056 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t2347 VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t2119 VGND.t2118 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t2058 XThC.TBN.t5 XThC.Tn[5].t11 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t378 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t236 VGND.t2483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t2413 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t2412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t176 VGND.t1408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t149 VGND.t1290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t11 XThC.TB5 VPWR.t1271 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t2349 VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t147 VGND.t1288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t1150 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.TBN.t6 XThC.Tn[0].t4 VPWR.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1791 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1792 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t197 VGND.t1723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.TB4.t2 VPWR.t1340 VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.TBN.t7 XThC.Tn[5].t7 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1926 VGND.t1928 VGND.t1927 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t1733 VGND.t1732 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t7 XThR.TBN.t5 a_n1049_5611# VPWR.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t11 XThC.TB5 VGND.t2098 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t2059 XThC.TBN.t8 XThC.Tn[2].t11 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.TB2 XThR.TA2 VPWR.t32 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t175 VGND.t1407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t2069 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t2068 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t1790 VPWR.t1788 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1789 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t2351 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t1022 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1021 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t672 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t816 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t471 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t2353 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t1115 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t1114 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t697 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1785 VPWR.t1787 VPWR.t1786 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.TB1.t3 XThC.Tn[8].t7 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t674 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t1286 VPWR.t1285 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.TB6 XThC.Tn[13].t3 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t1930 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t1929 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.TB5 XThC.TAN VGND.t756 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t7 XThC.TBN.t9 VPWR.t1242 VPWR.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t2121 VGND.t2120 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t1318 XThR.TB7 XThR.Tn[6].t3 VGND.t1317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t210 VPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t1829 XThR.TBN.t6 XThR.Tn[9].t3 VPWR.t1828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.TB7 XThR.TA3 VGND.t2674 VGND.t2673 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1024 VPWR.t1023 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t1026 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t2106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t779 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t778 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t353 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t1784 VPWR.t1782 XA.XIR[2].XIC_15.icell.PUM VPWR.t1783 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.TB7 VPWR.t658 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t1735 VGND.t1734 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t7 XThR.TBN.t7 VPWR.t1831 VPWR.t1830 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t810 VGND.t809 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.TBN.t10 VGND.t1353 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t676 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t643 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t143 VGND.t1284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t94 VGND.t746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t2355 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t2354 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t2491 XThR.TBN.t8 XThR.Tn[5].t11 VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t678 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t680 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t1988 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t1987 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t2415 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t2414 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t1321 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t212 VPWR.t211 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t1141 XThR.TB6 a_n1049_5611# VPWR.t800 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t513 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t682 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t2071 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t2070 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t954 VPWR.t953 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t2356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 a_n1049_7787# XThR.TB2 VPWR.t1908 VPWR.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 VGND.t483 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X96 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X97 VGND.t684 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X98 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X99 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t973 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X100 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1780 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1781 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 VGND.t686 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X102 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t812 VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X103 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1249 VPWR.t1248 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X104 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t638 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X105 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t640 VGND.t639 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t603 VPWR.t602 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X107 VGND.t2046 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2045 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X108 VPWR.t951 XThC.TB3.t3 a_4067_9615# VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X109 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X110 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 VPWR.t822 data[4].t0 a_n1335_4229# VPWR.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X112 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t777 VPWR.t776 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X113 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t128 VGND.t1158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X114 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t2122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X115 VGND.t132 XThR.TBN.t9 XThR.Tn[7].t3 VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X116 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t2076 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X117 a_n1319_5317# XThR.TA3 VPWR.t1917 VPWR.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X118 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t641 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X119 VPWR.t1 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X120 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X121 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X122 XThC.Tn[9].t7 XThC.TB2 VPWR.t404 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 XA.XIR[15].XIC[4].icell.Ien VPWR.t1777 VPWR.t1779 VPWR.t1778 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X124 VGND.t688 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X125 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t109 VGND.t849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X126 VGND.t690 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X127 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1774 VPWR.t1776 VPWR.t1775 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X128 XThC.Tn[5].t10 XThC.TBN.t11 VGND.t1354 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X130 VGND.t930 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X131 VGND.t932 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t931 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t645 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X133 VPWR.t512 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t511 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X134 VPWR.t62 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VGND.t1925 VGND.t1923 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X136 XThR.Tn[9].t7 XThR.TB2 a_n997_3755# VGND.t1784 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X137 XThC.Tn[0].t3 XThC.TBN.t12 a_2979_9615# VPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t2358 VGND.t2357 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X139 XThC.Tn[5].t6 XThC.TBN.t13 a_5949_9615# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X140 VGND.t2097 XThC.TB5 XThC.Tn[4].t10 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X141 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t817 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X142 VGND.t934 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t933 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X143 a_9827_9569# XThC.TB5 XThC.Tn[12].t7 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X144 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X145 XThC.Tn[7].t3 XThC.TBN.t14 VGND.t1356 VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X146 XThC.Tn[2].t10 XThC.TBN.t15 VGND.t1357 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 VGND.t1739 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t1738 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X148 a_n997_1579# XThR.TBN.t10 VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X149 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t347 VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X150 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t349 VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1772 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t8 VGND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X153 VGND.t1637 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t1636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X154 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t870 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X155 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t1178 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X156 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t416 VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t108 VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X159 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X160 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t872 VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t117 VGND.t1009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X162 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t53 VGND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X164 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1229 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X166 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t25 VGND.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X167 XA.XIR[15].XIC[0].icell.Ien VPWR.t1769 VPWR.t1771 VPWR.t1770 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X168 VGND.t936 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t935 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X169 VGND.t1181 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t1180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X170 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1766 VPWR.t1768 VPWR.t1767 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X171 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X172 VGND.t1208 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t1207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X173 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t313 VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X174 VGND.t1358 XThC.TBN.t16 XThC.Tn[1].t11 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VGND.t938 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t937 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X176 VPWR.t66 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X177 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X178 XA.XIR[2].XIC_15.icell.PUM VPWR.t1764 XA.XIR[2].XIC_15.icell.Ien VPWR.t1765 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t1697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X180 VPWR.t1300 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t1299 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X181 VPWR.t638 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t637 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VGND.t940 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X183 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t2360 VGND.t2359 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X184 VPWR.t1763 VPWR.t1761 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X185 VPWR.t832 XThC.TBN.t17 XThC.Tn[10].t9 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VGND.t136 XThR.TBN.t11 XThR.Tn[3].t11 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t1696 VGND.t1695 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X188 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t355 VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X189 XThR.Tn[0].t7 XThR.TBN.t12 a_n1049_8581# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X191 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t96 VGND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X192 VPWR.t1097 VGND.t2689 XA.XIR[0].XIC[8].icell.PUM VPWR.t1096 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X193 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X194 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XThC.Tn[12].t10 XThC.TB5 VPWR.t1270 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X196 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X197 XThR.Tn[11].t11 XThR.TBN.t13 VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t596 VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X199 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t1694 VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X200 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t874 VGND.t873 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X203 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X204 VGND.t2417 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t2416 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XThR.Tn[2].t0 XThR.TBN.t14 VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VGND.t2419 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t2418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X208 VGND.t1922 VGND.t1920 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1921 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X209 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t68 VPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X210 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1247 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X211 VPWR.t85 XThR.TBN.t15 XThR.Tn[12].t11 VPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X212 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X213 XThC.TA3 data[0].t0 VPWR.t717 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 VPWR.t1302 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t1301 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X215 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t375 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X216 VGND.t942 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X217 XA.XIR[0].XIC[13].icell.PDM VGND.t1917 VGND.t1919 VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X218 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 VGND.t2362 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t2073 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t2072 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t944 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X222 XThC.Tn[9].t3 XThC.TB2 a_7875_9569# VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 VGND.t419 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X224 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t442 VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X225 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t2364 VGND.t2363 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X226 VGND.t2075 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t2074 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t473 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t2366 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 a_n1319_5611# XThR.TA2 VPWR.t30 VPWR.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X230 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X231 VGND.t139 XThR.TBN.t16 a_n997_3979# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X232 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t144 VGND.t1285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X233 VPWR.t833 XThC.TBN.t18 XThC.Tn[14].t11 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 VGND.t946 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t945 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X235 VPWR.t70 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X236 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X237 VGND.t948 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t947 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X238 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t398 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X239 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t598 VPWR.t597 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X241 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t1692 VGND.t1691 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X242 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t357 VPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X243 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X244 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t216 VGND.t2067 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X245 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t60 VPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X246 VGND.t950 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X247 VGND.t1966 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t1965 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X248 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t353 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 VPWR.t1401 XThR.TB4 a_n1049_6699# VPWR.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X250 VGND.t2368 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t2367 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X251 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t121 VGND.t1142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X252 VPWR.t1095 VGND.t2690 XA.XIR[0].XIC[3].icell.PUM VPWR.t1094 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X253 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X254 VPWR.t395 XThC.TB6 a_5949_9615# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VPWR.t1064 XThR.TB1.t3 a_n1049_8581# VPWR.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X256 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X257 VPWR.t956 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t955 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X258 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t600 VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X259 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X260 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t89 VGND.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X261 VGND.t952 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X262 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t1342 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X263 VGND.t647 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t2302 XThR.TAN a_n1335_8107# VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VPWR.t466 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X266 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X267 VPWR.t1760 VPWR.t1758 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1759 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X268 VGND.t649 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X269 VGND.t954 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X270 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t468 VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X271 XThC.TB4.t1 XThC.TAN VPWR.t562 VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X272 VGND.t1916 VGND.t1914 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X273 VGND.t1990 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X274 VPWR.t1757 VPWR.t1755 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1756 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X275 XThR.Tn[2].t1 XThR.TB3.t3 VGND.t217 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X276 VGND.t141 XThR.TBN.t17 a_n997_2891# VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 VPWR.t1304 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t1303 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X278 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t138 VGND.t1203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X279 VPWR.t972 XThR.TB5 XThR.Tn[12].t7 VPWR.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t1038 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X281 VGND.t1755 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t1754 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t692 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X283 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X284 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t54 VGND.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X285 VGND.t143 XThR.TBN.t18 XThR.Tn[6].t11 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1614 VGND.t1613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X287 VPWR.t87 XThR.TBN.t19 XThR.Tn[9].t2 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t78 VGND.t597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X289 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X290 VGND.t1913 VGND.t1911 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X291 XA.XIR[14].XIC_15.icell.PUM VPWR.t1753 XA.XIR[14].XIC_15.icell.Ien VPWR.t1754 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X292 a_n997_715# XThR.TBN.t20 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X293 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X294 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XThC.Tn[1].t10 XThC.TBN.t19 VGND.t1359 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 VPWR.t858 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t857 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X297 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t975 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X298 XThR.Tn[14].t7 XThR.TB7 VPWR.t815 VPWR.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t1230 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X300 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t73 VGND.t555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X301 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t228 VGND.t2285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t2370 VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X303 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t33 VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X304 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X305 VGND.t694 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X306 VGND.t696 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t695 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X308 VPWR.t470 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X309 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X310 VPWR.t970 XThR.TB5 a_n1049_6405# VPWR.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X311 VPWR.t860 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t859 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X312 XThR.TAN data[6].t0 VPWR.t628 VPWR.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X313 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t705 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X314 VPWR.t1341 XThC.TB4.t3 a_4861_9615# VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t152 VGND.t1295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X316 VGND.t698 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X317 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t640 VPWR.t639 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X318 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1750 VPWR.t1752 VPWR.t1751 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 VGND.t2607 XThR.TB2 XThR.Tn[1].t11 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t814 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X321 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t1427 VGND.t1426 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X322 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t206 VGND.t1973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X323 XThR.TA3 data[4].t1 a_n1331_2891# VGND.t1327 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t67 VGND.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X325 VGND.t700 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X326 XA.XIR[15].XIC[13].icell.Ien VPWR.t1747 VPWR.t1749 VPWR.t1748 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X327 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t190 VGND.t1655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X328 VPWR.t238 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t237 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X329 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t2371 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X330 VPWR.t642 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t641 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X331 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X332 a_n1049_7787# XThR.TBN.t21 XThR.Tn[1].t3 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X333 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t43 VGND.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X334 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t1028 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X335 VGND.t1360 XThC.TBN.t20 XThC.Tn[4].t7 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X336 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X337 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t29 VGND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X338 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t225 VGND.t2278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1745 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1746 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X340 VGND.t1910 VGND.t1908 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X341 XThC.TA1 data[1].t0 a_7331_10587# VPWR.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X342 VGND.t230 data[1].t1 a_8739_10571# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 XA.XIR[0].XIC[1].icell.PDM VGND.t1905 VGND.t1907 VGND.t1906 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X344 VPWR.t1907 XThR.TB2 XThR.Tn[9].t11 VPWR.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND.t147 XThR.TBN.t22 XThR.Tn[7].t2 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VGND.t1968 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t1967 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X347 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t65 VGND.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X348 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X349 XThR.Tn[13].t11 XThR.TBN.t23 VPWR.t90 VPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X350 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t560 VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X351 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t98 VGND.t759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X352 VGND.t702 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X353 VGND.t1904 VGND.t1902 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t644 VPWR.t643 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X355 VPWR.t775 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X356 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1742 VPWR.t1744 VPWR.t1743 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X357 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t72 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 VPWR.t359 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X359 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t376 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X360 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1739 VPWR.t1741 VPWR.t1740 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X361 VPWR.t240 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X362 VGND.t1323 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X363 VGND.t1957 XThR.TB6 XThR.Tn[5].t3 VGND.t1628 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X365 XThR.Tn[9].t6 XThR.TB2 a_n997_3755# VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 VGND.t704 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X367 XThR.TB6 XThR.TA2 VGND.t61 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X368 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t2374 VGND.t2373 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X369 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t6 VGND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X370 a_n997_1579# XThR.TBN.t24 VGND.t149 VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 VGND.t2570 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t2569 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X372 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t142 VGND.t1281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X373 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t827 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X374 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t828 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 VPWR.t315 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X376 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1737 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1738 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X377 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t2488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X378 VPWR.t9 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X379 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X380 XA.XIR[15].XIC[6].icell.Ien VPWR.t1734 VPWR.t1736 VPWR.t1735 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X381 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t2376 VGND.t2375 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X382 VGND.t706 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X383 VPWR.t1202 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t1201 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X384 VPWR.t566 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t2377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X386 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t605 VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X387 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t562 VGND.t561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X388 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t380 VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t2379 VGND.t2378 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 VPWR.t997 XThR.TAN2 XThR.TBN.t3 VPWR.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X392 VPWR.t242 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X393 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t2078 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X394 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t976 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X395 VPWR.t317 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X396 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t11 VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X397 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X398 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t977 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1732 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1733 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 a_3523_10575# XThC.TAN VGND.t755 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X401 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t2080 VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X402 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t2082 VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t1152 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t168 VGND.t1394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X405 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t698 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X406 VPWR.t834 XThC.TBN.t21 XThC.Tn[13].t11 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X408 VGND.t708 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X409 VGND.t1639 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t1638 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X410 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X411 XThC.Tn[5].t3 XThC.TB6 VGND.t504 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 XThC.Tn[4].t9 XThC.TB5 VGND.t2096 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X414 VGND.t2381 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t2380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X415 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t829 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X416 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X417 VPWR.t321 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X418 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X419 a_n997_1579# XThR.TB6 XThR.Tn[13].t7 VGND.t1627 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 VPWR.t325 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X421 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t2012 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X422 VPWR.t1306 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t1305 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X423 XA.XIR[15].XIC[1].icell.Ien VPWR.t1729 VPWR.t1731 VPWR.t1730 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X424 VGND.t710 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t709 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X425 VGND.t712 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1726 VPWR.t1728 VPWR.t1727 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X427 VGND.t1185 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t1184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X428 VGND.t1210 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t1209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 a_7875_9569# XThC.TB2 XThC.Tn[9].t2 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 XThC.Tn[4].t6 XThC.TBN.t22 VGND.t1361 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VPWR.t176 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X432 a_n1049_5317# XThR.TB7 VPWR.t813 VPWR.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t327 VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X434 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t164 VGND.t1390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X435 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t382 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X436 VGND.t714 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VGND.t1901 VGND.t1899 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VPWR.t568 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t567 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X439 VPWR.t168 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 XThC.TB6 XThC.TAN VGND.t754 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VPWR.t1725 VPWR.t1723 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1724 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X442 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t2382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X443 VPWR.t472 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X444 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X445 a_6243_9615# XThC.TBN.t23 XThC.Tn[6].t7 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t1632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X447 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X448 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t10 VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X450 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X451 XThC.Tn[13].t7 XThC.TB6 VPWR.t394 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X452 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t13 VGND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X453 VGND.t1362 XThC.TBN.t24 XThC.Tn[0].t8 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 XThR.Tn[3].t7 XThR.TBN.t25 a_n1049_6699# VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X456 VGND.t1325 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t1324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X457 VGND.t2283 XThR.TB4 XThR.Tn[3].t3 VGND.t1037 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t830 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X459 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t308 VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X460 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X462 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t1231 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X463 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t227 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t74 VGND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X465 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t2385 VGND.t2384 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X466 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t76 VGND.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X467 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t2125 VGND.t2124 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X468 VGND.t716 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X469 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t1206 VPWR.t1205 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X470 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t1153 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X471 VGND.t956 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t955 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X472 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t3 VGND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X473 XThR.Tn[11].t7 XThR.TB4 VPWR.t1400 VPWR.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X474 VGND.t1212 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X475 VGND.t1187 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t1186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 XThC.Tn[14].t3 XThC.TB7 a_10915_9569# VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 VPWR.t178 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X478 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t323 VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X479 VGND.t2048 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t2047 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X480 VPWR.t170 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X481 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t2013 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X482 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X483 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t2386 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X484 VPWR.t1722 VPWR.t1720 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1721 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X485 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t1179 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X486 VGND.t2173 XThC.TB4.t4 XThC.Tn[3].t11 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VPWR.t403 XThC.TB2 XThC.Tn[9].t6 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X488 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t244 VPWR.t243 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X489 VGND.t475 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X490 VGND.t958 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t957 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X491 VGND.t2388 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X492 VPWR.t968 XThR.TB5 XThR.Tn[12].t6 VPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VGND.t2572 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t2571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X494 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t75 VGND.t574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X495 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t889 VPWR.t888 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X496 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t570 VPWR.t569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X498 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X499 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t2583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 VPWR.t811 XThR.TB7 XThR.Tn[14].t6 VPWR.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X502 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t388 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X503 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t1882 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X504 XThR.Tn[8].t3 XThR.TB1.t4 a_n997_3979# VGND.t1784 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t1029 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X506 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 VGND.t2421 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t2420 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t2390 VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 VPWR.t474 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X510 VPWR.t1284 data[2].t0 XThC.TAN VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X511 VGND.t1898 VGND.t1896 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X512 VPWR.t444 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X513 VGND.t1741 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t1740 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X514 XThC.Tn[13].t2 XThC.TB6 a_10051_9569# VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X515 XThR.Tn[4].t7 XThR.TBN.t26 a_n1049_6405# VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 XThR.TB5 XThR.TAN a_n1319_6405# VPWR.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X517 VGND.t960 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t959 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X518 XThC.Tn[8].t3 XThC.TBN.t25 VPWR.t836 VPWR.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X519 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t390 VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X520 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t1827 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t1541 VGND.t1540 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 a_n1335_4229# data[5].t0 XThR.TA1 VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X523 VGND.t1160 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X524 VGND.t962 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t961 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X525 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t1888 VPWR.t1887 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X526 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t246 VPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t2015 VGND.t2014 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X528 VGND.t1992 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t1991 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t964 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t963 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X530 VGND.t966 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t965 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 XThC.Tn[8].t6 XThC.TB1.t4 a_7651_9569# VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 XThC.Tn[13].t10 XThC.TBN.t26 VPWR.t34 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X533 VGND.t477 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X534 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t891 VPWR.t890 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X535 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t57 VGND.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X536 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t58 VGND.t421 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 VPWR.t1093 VGND.t2691 XA.XIR[0].XIC[9].icell.PUM VPWR.t1092 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X538 VGND.t503 XThC.TB6 XThC.Tn[5].t2 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t819 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X540 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1717 VPWR.t1719 VPWR.t1718 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X541 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t832 VGND.t831 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X542 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t834 VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X544 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X545 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 VGND.t968 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t967 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X548 VGND.t1641 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t1640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X549 a_n1049_5611# XThR.TB6 VPWR.t1140 VPWR.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 XA.XIR[13].XIC_15.icell.PUM VPWR.t1715 XA.XIR[13].XIC_15.icell.Ien VPWR.t1716 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X551 XThR.Tn[10].t4 XThR.TB3.t4 a_n997_2891# VGND.t1319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X552 VGND.t970 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t969 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X553 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X554 VGND.t2175 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t2174 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X555 VGND.t2574 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t2573 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VPWR.t36 XThC.TBN.t27 XThC.Tn[7].t6 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t2584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X558 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 VPWR.t446 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X560 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1713 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1714 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X561 VPWR.t1906 XThR.TB2 XThR.Tn[9].t10 VPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 XThC.Tn[6].t6 XThC.TBN.t28 a_6243_9615# VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X563 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t1344 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X564 VGND.t972 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t971 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X565 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t572 VPWR.t571 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X566 VGND.t1763 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t1762 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X567 VPWR.t607 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X568 VPWR.t838 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X569 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X570 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t862 VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X571 VGND.t974 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X572 VGND.t1994 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t1993 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X573 XA.XIR[15].XIC_15.icell.Ien VPWR.t1710 VPWR.t1712 VPWR.t1711 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X574 VPWR.t448 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X575 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X576 VPWR.t248 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t247 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X577 a_n1049_7493# XThR.TBN.t27 XThR.Tn[2].t11 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X578 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X579 XThC.Tn[0].t7 XThC.TBN.t29 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 VGND.t976 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X581 VPWR.t1709 VPWR.t1707 XA.XIR[9].XIC_15.icell.PUM VPWR.t1708 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X582 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t234 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X583 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t236 VGND.t235 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X584 VGND.t978 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t977 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X585 a_4067_9615# XThC.TBN.t30 XThC.Tn[2].t7 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X586 XThR.Tn[0].t1 XThR.TB1.t5 VGND.t1786 VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X587 VGND.t2678 XThR.TBN.t28 XThR.Tn[5].t10 VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X588 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t184 VGND.t1615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X589 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t250 VPWR.t249 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X590 VGND.t980 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X591 XThR.Tn[14].t3 XThR.TB7 a_n997_715# VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t2017 VGND.t2016 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X593 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t1403 VGND.t1402 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X594 VGND.t877 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X595 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t893 VPWR.t892 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X596 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t2339 VGND.t2338 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X597 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t20 VGND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X598 VGND.t2392 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X599 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t2585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X600 VGND.t2679 XThR.TBN.t29 XThR.Tn[4].t11 VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X601 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t836 VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X602 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X603 VGND.t2394 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t2393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 a_8963_9569# XThC.TB4.t5 XThC.Tn[11].t11 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X605 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t1328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 VGND.t879 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X607 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t178 VGND.t1522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X608 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1705 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1706 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X609 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t1329 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X610 VGND.t881 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X611 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X612 VGND.t1643 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X613 VGND.t1757 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X614 VGND.t883 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X615 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t864 VPWR.t863 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X616 VGND.t2050 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t2049 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X617 VPWR.t609 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t608 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X618 VGND.t885 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t884 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X619 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t1208 VPWR.t1207 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X620 VGND.t69 XThC.TBN.t31 a_8739_9569# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X621 VGND.t2142 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X622 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t2395 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X623 VGND.t887 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t886 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X624 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t172 VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X625 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t574 VPWR.t573 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X626 VGND.t889 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X627 VGND.t1214 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t1213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X628 VGND.t1189 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X629 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t866 VPWR.t865 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X630 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t1405 VGND.t1404 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t237 VGND.t2484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X632 a_9827_9569# XThC.TBN.t32 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X633 VGND.t891 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t890 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X634 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t207 VGND.t1974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X635 VPWR.t223 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X636 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X637 VPWR.t158 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X638 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t2396 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X639 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t140 VGND.t1205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X640 VPWR.t174 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X641 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t1428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X642 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t838 VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X643 VPWR.t1704 VPWR.t1702 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X644 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t2397 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X645 VGND.t1292 XThC.TB1.t5 XThC.Tn[0].t0 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X646 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t219 VGND.t218 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X647 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t133 VGND.t1196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X648 XThR.TA3 data[5].t1 VPWR.t461 VPWR.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X649 VGND.t1743 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t1742 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X650 VPWR.t1210 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t1209 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X651 VGND.t2087 XThC.TAN2 XThC.TBN.t1 VGND.t2086 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X652 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X653 VPWR.t1410 XThR.TAN XThR.TB1.t2 VPWR.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X654 a_n997_1579# XThR.TB6 XThR.Tn[13].t6 VGND.t1626 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t77 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X656 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t611 VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X657 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t46 VGND.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X658 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t2399 VGND.t2398 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1699 VPWR.t1701 VPWR.t1700 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t200 VGND.t1950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X661 VPWR.t225 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X662 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t1047 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X663 XThC.Tn[7].t5 XThC.TBN.t33 VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X664 VGND.t2301 XThR.TAN a_n1335_7243# VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X665 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t1048 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X666 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X667 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X668 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t2401 VGND.t2400 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[12].XIC_15.icell.PUM VPWR.t1697 XA.XIR[12].XIC_15.icell.Ien VPWR.t1698 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t1335 VGND.t1334 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t2018 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X672 VGND.t479 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t706 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X674 VGND.t2576 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t2575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X675 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t174 VGND.t1401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X676 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t773 VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X677 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t185 VGND.t1616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X678 XThC.Tn[11].t0 XThC.TB4.t6 VPWR.t287 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X679 VGND.t2578 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t2577 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X680 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t179 VGND.t1585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1694 VPWR.t1696 VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X682 a_n997_1803# XThR.TBN.t30 VGND.t2680 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X683 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t1417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X684 XThR.Tn[3].t6 XThR.TBN.t31 a_n1049_6699# VPWR.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X685 VPWR.t895 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t894 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X686 VGND.t2681 XThR.TBN.t32 XThR.Tn[3].t10 VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X687 VGND.t893 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t892 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X688 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t1809 VPWR.t1808 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X689 VGND.t2403 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t2402 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X690 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t2405 VGND.t2404 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X691 XThC.Tn[2].t6 XThC.TBN.t34 a_4067_9615# VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X692 VPWR.t160 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X693 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t329 VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X694 VPWR.t613 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X695 VPWR.t1212 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t1211 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X696 XThR.Tn[11].t6 XThR.TB4 VPWR.t1399 VPWR.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X697 VPWR.t1693 VPWR.t1691 XA.XIR[8].XIC_15.icell.PUM VPWR.t1692 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 VPWR.t402 XThC.TB2 a_3773_9615# VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 a_n1049_8581# XThR.TB1.t6 VPWR.t1066 VPWR.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1689 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1690 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X701 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t1699 VGND.t1698 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X702 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t360 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X703 VGND.t895 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X704 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t2341 VGND.t2340 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 VGND.t261 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X706 VGND.t1895 VGND.t1893 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X707 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t329 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t1543 VGND.t1542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t241 VGND.t2597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X710 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t771 VPWR.t770 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X711 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t250 VGND.t2663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X712 VGND.t1040 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X713 VPWR.t716 XThC.TA2 a_5949_10571# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X714 VPWR.t227 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X715 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t1365 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X717 VGND.t1634 XThR.TB3.t5 XThR.Tn[2].t8 VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X718 VPWR.t665 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t664 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X719 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1860 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X720 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t675 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X721 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t700 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X722 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t1337 VGND.t1336 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t120 VGND.t1141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X724 XThC.TBN.t3 XThC.TAN2 VPWR.t1253 VPWR.t1252 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X725 VGND.t897 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t896 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X726 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X727 VGND.t2252 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t2251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X728 VGND.t899 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t898 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X729 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t1811 VPWR.t1810 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X730 XThR.Tn[8].t4 XThR.TB1.t7 a_n997_3979# VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 XA.XIR[6].XIC_15.icell.PUM VPWR.t1687 XA.XIR[6].XIC_15.icell.Ien VPWR.t1688 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X732 VGND.t2546 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t2545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X733 VGND.t901 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X734 VGND.t2254 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t2253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t442 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X736 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t840 VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X737 VGND.t1042 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t1041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 VGND.t2177 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t2176 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X739 VGND.t2144 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X740 VGND.t72 XThC.TBN.t35 a_9827_9569# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X741 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VPWR.t897 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t896 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X743 VPWR.t657 XThC.TB7 XThC.Tn[14].t7 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X744 XThR.Tn[4].t6 XThR.TBN.t33 a_n1049_6405# VPWR.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X745 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X746 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X747 VGND.t444 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X748 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t1813 VPWR.t1812 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X749 VGND.t446 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X750 VPWR.t1398 XThR.TB4 a_n1049_6699# VPWR.t965 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X751 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t252 VPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X752 VGND.t448 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X753 VPWR.t162 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X754 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t667 VPWR.t666 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X755 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t899 VPWR.t898 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X756 VGND.t450 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X757 VPWR.t615 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t614 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X758 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t192 VGND.t1710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X759 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t824 VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X760 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X761 VPWR.t1167 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t1166 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X762 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t2342 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X763 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t1044 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X764 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X765 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t1042 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X766 VGND.t452 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X767 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t36 VGND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X768 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t231 VGND.t2290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X769 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t331 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X770 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t769 VPWR.t768 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X771 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 VGND.t454 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X773 VPWR.t1920 XThR.TBN.t34 XThR.Tn[8].t11 VPWR.t1919 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X774 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t842 VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X775 XThR.Tn[10].t7 XThR.TB3.t6 a_n997_2891# VGND.t2103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X776 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X777 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t1030 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X778 XThC.TB3.t0 XThC.TAN VPWR.t560 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X779 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t243 VGND.t2599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X780 VGND.t456 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X781 VGND.t1892 VGND.t1890 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1891 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X782 VGND.t458 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X783 VPWR.t715 XThC.TA2 XThC.TB2 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X784 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t1419 VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X785 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t1421 VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X786 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t245 VGND.t2601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X787 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t844 VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X788 VGND.t460 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X789 VGND.t1759 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X790 VGND.t1434 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t1433 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X791 XThR.TB3.t1 XThR.TA3 VPWR.t1916 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X792 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t162 VGND.t1352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X793 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t2019 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X794 VGND.t2146 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X795 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t1406 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X796 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t1046 VGND.t1045 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X797 a_n997_715# XThR.TB7 XThR.Tn[14].t2 VGND.t1315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X798 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X799 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X800 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t1255 VPWR.t1254 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X801 VGND.t462 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X802 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t19 VGND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X803 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t166 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 XThR.Tn[0].t11 XThR.TBN.t35 VGND.t2682 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X805 VPWR.t966 XThR.TB5 a_n1049_6405# VPWR.t965 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X806 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 VGND.t464 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X808 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t210 VGND.t2027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X809 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t2343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X810 XThC.Tn[10].t11 XThC.TB3.t4 VPWR.t952 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t1296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X812 VPWR.t1921 XThR.TBN.t36 XThR.Tn[10].t11 VPWR.t1828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t1167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X814 VPWR.t854 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X815 VPWR.t41 XThC.TBN.t36 XThC.Tn[13].t9 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X816 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t1544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X817 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t1338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X818 a_3773_9615# XThC.TB2 VPWR.t401 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XThC.Tn[5].t1 XThC.TB6 VGND.t502 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X820 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t31 VGND.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X821 XThC.Tn[2].t3 XThC.TB3.t5 VGND.t1603 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 VPWR.t1169 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t1168 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X823 VPWR.t767 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t766 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X824 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t2021 VGND.t2020 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X825 VGND.t1745 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t1744 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X826 VPWR.t1890 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t1889 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t37 VGND.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X828 VPWR.t791 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X829 VGND.t2683 XThR.TBN.t37 a_n997_3755# VGND.t1529 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X830 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1345 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X831 VPWR.t785 XThC.TB1.t6 a_2979_9615# VPWR.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t1546 VGND.t1545 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X833 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t1048 VGND.t1047 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X834 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X835 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t1257 VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X836 VGND.t466 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X837 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t2023 VGND.t2022 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X838 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t39 VGND.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X839 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t1423 VGND.t1422 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X840 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t91 VGND.t743 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X841 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X842 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t182 VGND.t1606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X843 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t872 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X844 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t234 VGND.t2429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 VGND.t423 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X846 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t1050 VGND.t1049 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X847 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t186 VGND.t1617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X849 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X850 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t16 VGND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t1547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1854 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X853 a_5155_9615# XThC.TB5 VPWR.t1269 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X854 XA.XIR[5].XIC_15.icell.PUM VPWR.t1685 XA.XIR[5].XIC_15.icell.Ien VPWR.t1686 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X855 VPWR.t856 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t855 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X856 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t2587 VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X857 a_n1049_7493# XThR.TB3.t7 VPWR.t660 VPWR.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X858 VGND.t2548 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t2547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X859 XA.XIR[9].XIC_15.icell.PUM VPWR.t1683 XA.XIR[9].XIC_15.icell.Ien VPWR.t1684 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X860 VGND.t1162 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t1161 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X861 VPWR.t765 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t764 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X862 VPWR.t1892 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t1891 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X863 VGND.t1052 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t1051 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X864 XThC.Tn[8].t11 XThC.TB1.t7 VPWR.t787 VPWR.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X865 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t619 VPWR.t618 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X866 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t1171 VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X867 VGND.t1629 XThR.TB5 XThR.Tn[4].t3 VGND.t1628 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X868 a_5155_9615# XThC.TBN.t37 XThC.Tn[4].t3 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X869 VGND.t1054 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X870 VPWR.t1173 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X871 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t2025 VGND.t2024 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X872 VPWR.t763 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X873 XThR.TB5 XThR.TA1 VGND.t60 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X874 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t1425 VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X875 VPWR.t1894 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t1893 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X876 VPWR.t1259 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t1258 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X877 VPWR.t793 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t792 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X878 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X879 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X880 VPWR.t1682 VPWR.t1680 XA.XIR[1].XIC_15.icell.PUM VPWR.t1681 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X881 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t840 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X882 VPWR.t1679 VPWR.t1677 XA.XIR[5].XIC_15.icell.PUM VPWR.t1678 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X883 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X884 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t2589 VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X885 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t1261 VPWR.t1260 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X886 VGND.t2638 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t2637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X887 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t26 VGND.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X888 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t84 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 VGND.t2640 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t2639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X890 VGND.t1057 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X891 VGND.t2642 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t2641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X892 VGND.t1765 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VPWR.t1676 VPWR.t1674 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X894 XThC.Tn[14].t2 XThC.TB7 a_10915_9569# VGND.t1021 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X895 XThC.TB3.t1 XThC.TA3 a_4387_10575# VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X896 a_n997_1803# XThR.TBN.t38 VGND.t2684 VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X897 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X898 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1175 VPWR.t1174 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X899 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t245 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X900 a_3773_9615# XThC.TBN.t38 XThC.Tn[1].t7 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X901 VGND.t2550 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t203 VGND.t1958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X903 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t247 VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 VGND.t2644 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t2643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X905 VGND.t2148 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 VPWR.t464 XThC.TA1 XThC.TB1.t0 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X907 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t1058 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X908 VGND.t2150 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X909 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t1059 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X910 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t2091 VGND.t2090 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X911 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t1931 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 VGND.t2646 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t2645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X913 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X914 VGND.t2648 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t2647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X915 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1177 VPWR.t1176 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X916 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t2026 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X917 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1672 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X918 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t761 VPWR.t760 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X919 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t252 VGND.t2675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X920 VGND.t1199 XThC.TB3.t6 XThC.Tn[2].t1 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X921 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1346 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X922 a_8739_9569# XThC.TB3.t7 XThC.Tn[10].t6 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t1339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X924 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X925 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t1978 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X926 a_n1319_6405# XThR.TA1 VPWR.t28 VPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X927 VPWR.t182 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X928 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t1932 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X930 VPWR.t1671 VPWR.t1669 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1670 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X931 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t122 VGND.t1143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X932 a_2979_9615# XThC.TB1.t8 VPWR.t789 VPWR.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X933 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t1000 VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X934 VGND.t2650 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t2649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X935 VGND.t2652 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t2651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X936 XThR.Tn[12].t10 XThR.TBN.t39 VPWR.t1922 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X937 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t2028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X938 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1666 VPWR.t1668 VPWR.t1667 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X939 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t80 VGND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X940 XThC.Tn[11].t10 XThC.TBN.t39 VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X941 VGND.t1329 data[4].t2 XThR.TA1 VGND.t1328 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X942 XThR.TBN.t1 XThR.TAN2 VGND.t1708 VGND.t1707 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X943 VGND.t1169 data[3].t0 XThC.TAN2 VGND.t1168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X944 VGND.t2654 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t2653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X945 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t1061 VGND.t1060 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X946 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t1341 VGND.t1340 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X947 a_n997_1803# XThR.TB5 XThR.Tn[12].t3 VGND.t1627 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X948 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X949 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t82 VGND.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X950 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t1063 VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t169 VGND.t1395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X952 a_n997_2667# XThR.TBN.t40 VGND.t2685 VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X953 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1664 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1665 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X954 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t212 VGND.t2063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X955 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X956 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t2093 VGND.t2092 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X957 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t1933 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X958 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X959 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t198 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t522 VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 VPWR.t184 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X962 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t1343 VGND.t1342 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t906 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 VGND.t2580 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t2579 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t227 VGND.t2284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X966 XThC.Tn[4].t2 XThC.TBN.t40 a_5155_9615# VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X967 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t1979 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X968 VGND.t1065 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t1064 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 VPWR.t1214 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t1213 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X970 VPWR.t1924 XThR.TBN.t41 XThR.Tn[8].t10 VPWR.t1923 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X971 VGND.t1191 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t1190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X972 VGND.t1550 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X974 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X975 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1661 VPWR.t1663 VPWR.t1662 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X976 a_7651_9569# XThC.TB1.t9 XThC.Tn[8].t5 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X977 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X978 VGND.t2656 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t2655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X979 VPWR.t1268 XThC.TB5 XThC.Tn[12].t9 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t1066 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X981 VPWR.t1099 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t1098 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X982 VPWR.t1660 VPWR.t1658 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X983 VGND.t2658 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t2657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X984 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t1896 VPWR.t1895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X985 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t795 VPWR.t794 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X986 VGND.t2179 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t2178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X987 VGND.t2686 XThR.TBN.t42 XThR.Tn[1].t7 VGND.t2499 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X988 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t251 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X989 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t1299 VGND.t1298 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X990 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t901 VPWR.t900 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X991 VPWR.t1091 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t1090 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X992 VPWR.t1657 VPWR.t1655 XA.XIR[4].XIC_15.icell.PUM VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X993 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t1002 VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X994 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t1144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X995 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X996 VGND.t2660 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t2659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X997 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X998 XThR.Tn[6].t2 XThR.TB7 VGND.t1314 VGND.t1313 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 a_9827_9569# XThC.TBN.t41 VGND.t73 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1000 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1001 XThR.Tn[9].t1 XThR.TBN.t43 VPWR.t1925 VPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1002 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t2101 VGND.t2100 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1003 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t1301 VGND.t1300 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1004 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t1711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1006 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t204 VGND.t1971 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1007 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t1713 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1008 XThC.Tn[1].t6 XThC.TBN.t42 a_3773_9615# VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1009 VGND.t425 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1010 XThR.Tn[0].t10 XThR.TBN.t44 VGND.t2687 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1011 XThC.Tn[13].t1 XThC.TB6 a_10051_9569# VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1012 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1013 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1014 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t677 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1015 VPWR.t878 XThR.TBN.t45 XThR.Tn[10].t10 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1016 VPWR.t903 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t902 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1017 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1018 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t524 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1652 VPWR.t1654 VPWR.t1653 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1020 XA.XIR[0].XIC[12].icell.PDM VGND.t1887 VGND.t1889 VGND.t1888 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1021 VGND.t2256 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t2255 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 VGND.t2552 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 VGND.t2662 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t2661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1024 VGND.t2512 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t2511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1025 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t1898 VPWR.t1897 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1026 VPWR.t656 XThC.TB7 a_6243_9615# VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t134 VGND.t1197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1028 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t1068 VGND.t1067 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1029 VGND.t2554 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1030 VGND.t2181 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t2180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1031 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t669 VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1032 VGND.t1164 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t1163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VPWR.t1089 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t1088 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1034 VGND.t2538 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t2537 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t2344 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1036 VGND.t1070 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t1069 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 VGND.t1410 XThC.TBN.t43 a_8963_9569# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1038 VGND.t2514 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t2513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1039 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t1366 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1040 VPWR.t1107 XThR.TB1.t8 XThR.Tn[8].t5 VPWR.t1106 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1041 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1650 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1042 VGND.t2516 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t2515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1043 VGND.t2518 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t2517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1044 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t1900 VPWR.t1899 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1045 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t211 VGND.t2060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1046 VGND.t1761 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t1760 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1047 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t1263 VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1048 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t797 VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 VGND.t1436 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t1435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1050 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t1303 VGND.t1302 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1051 XThR.TAN2 data[7].t0 VPWR.t515 VPWR.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1052 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t905 VPWR.t904 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t416 VPWR.t415 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1054 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t132 VGND.t1195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1055 a_6243_10571# XThC.TAN XThC.TB7 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1056 VPWR.t1087 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t1086 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1057 VPWR.t1905 XThR.TB2 a_n1049_7787# VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1058 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t2345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1059 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t2590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1060 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t1004 VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1061 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1062 VPWR.t1101 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1063 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t2102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t41 VGND.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1065 XA.XIR[0].XIC[10].icell.PDM VGND.t1884 VGND.t1886 VGND.t1885 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1066 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t1714 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1067 VGND.t2520 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t2519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1068 a_n1049_7493# XThR.TBN.t46 XThR.Tn[2].t4 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1069 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t66 VGND.t508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1070 VGND.t1767 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1071 XThC.Tn[8].t10 XThC.TB1.t10 VPWR.t1294 VPWR.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1072 VPWR.t122 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1073 VPWR.t1649 VPWR.t1647 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1074 VGND.t1883 VGND.t1881 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1075 VGND.t263 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1076 XThR.Tn[0].t2 XThR.TB1.t9 VGND.t1935 VGND.t1934 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1077 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1078 VGND.t2522 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t2521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1079 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 VPWR.t373 XThR.TB3.t8 XThR.Tn[10].t0 VPWR.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1081 VGND.t1747 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1082 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1083 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t202 VGND.t1953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1085 VPWR.t400 XThC.TB2 a_3773_9615# VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1086 VGND.t1242 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t1241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 VGND.t1524 XThR.TBN.t47 XThR.Tn[4].t10 VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1088 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1645 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1089 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t156 VGND.t1326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1090 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t982 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1092 VPWR.t845 XThC.TBN.t44 XThC.Tn[9].t11 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1093 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t1071 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1094 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1095 VGND.t1411 XThC.TBN.t45 XThC.Tn[5].t9 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1096 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t1981 VGND.t1980 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1097 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t1939 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1098 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t49 VGND.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1099 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t238 VGND.t2485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1100 VGND.t1526 XThR.TBN.t48 a_n997_1579# VGND.t1525 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1101 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1102 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t4 VGND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1103 VGND.t2524 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t2523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1104 VGND.t2526 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t2525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1105 a_2979_9615# XThC.TBN.t46 XThC.Tn[0].t2 VPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1106 VGND.t1684 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t1683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1107 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1108 VGND.t1552 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1109 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1110 VPWR.t1103 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t1102 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1111 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1112 XThC.Tn[12].t6 XThC.TB5 a_9827_9569# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1114 VPWR.t124 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1115 XThR.TA2 data[5].t2 VPWR.t1283 VPWR.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1116 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t232 VGND.t2410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1117 VPWR.t1644 VPWR.t1642 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1118 XThR.Tn[14].t1 XThR.TB7 a_n997_715# VGND.t1312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1119 VPWR.t186 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1120 a_n1049_5317# XThR.TBN.t49 XThR.Tn[6].t7 VPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1121 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1105 VPWR.t1104 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1122 VGND.t2528 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t2527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1123 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t215 VGND.t2066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1124 XA.XIR[15].XIC[12].icell.Ien VPWR.t1639 VPWR.t1641 VPWR.t1640 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1125 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t45 VGND.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1126 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t165 VGND.t1391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1127 VPWR.t217 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1128 VPWR.t1273 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t1272 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1129 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1130 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t1073 VGND.t1072 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1131 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t1716 VGND.t1715 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1132 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t1885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1133 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1134 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t126 VGND.t1156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1135 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t1 VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1136 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t1075 VGND.t1074 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t1032 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t69 VGND.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1139 a_6243_9615# XThC.TB7 VPWR.t655 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1140 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1637 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1638 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1141 VGND.t1880 VGND.t1878 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1142 XThC.Tn[10].t10 XThC.TBN.t47 VPWR.t847 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1143 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1144 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t1983 VGND.t1982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1146 VGND.t1438 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t1437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1147 XA.XIR[1].XIC_15.icell.PUM VPWR.t1635 XA.XIR[1].XIC_15.icell.Ien VPWR.t1636 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1148 XThC.Tn[10].t7 XThC.TB3.t8 a_8739_9569# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1149 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t302 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 VGND.t1020 XThC.TB7 XThC.Tn[6].t3 VGND.t1019 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1151 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t55 VGND.t386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1152 VGND.t1077 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t1076 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1153 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t1079 VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 XThR.Tn[11].t10 XThR.TBN.t50 VPWR.t881 VPWR.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1155 VGND.t2540 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t2539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1156 VPWR.t848 XThC.TBN.t48 XThC.Tn[12].t3 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 VGND.t1081 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t1080 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XA.XIR[15].XIC[10].icell.Ien VPWR.t1632 VPWR.t1634 VPWR.t1633 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1159 VGND.t2530 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t2529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1160 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t1863 VPWR.t1862 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1847 VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1162 VGND.t1083 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t1082 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1163 VPWR.t799 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1164 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t678 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1165 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1629 VPWR.t1631 VPWR.t1630 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VPWR.t1275 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1167 VGND.t2532 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t2531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1168 VGND.t2534 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t2533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1169 VGND.t2183 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1170 VGND.t2536 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t2535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1171 VGND.t1970 XThC.TA3 XThC.TB7 VGND.t1969 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1172 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t767 VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1173 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t759 VPWR.t758 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1174 VPWR.t219 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1175 a_n997_1803# XThR.TB5 XThR.Tn[12].t2 VGND.t1626 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t60 VGND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1177 a_n997_2667# XThR.TBN.t51 VGND.t1528 VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1178 VPWR.t188 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1179 VPWR.t1117 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1180 a_7875_9569# XThC.TBN.t49 VGND.t1412 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1181 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t1718 VGND.t1717 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1182 VGND.t1749 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t1748 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1183 VGND.t1530 XThR.TBN.t52 a_n997_3979# VGND.t1529 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1184 VGND.t545 Vbias.t1 Vbias.t2 VGND.t544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X1185 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t455 VPWR.t454 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1186 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t170 VGND.t1396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1187 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1347 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1188 XThC.Tn[14].t10 XThC.TBN.t50 VPWR.t849 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1189 a_n1049_6699# XThR.TB4 VPWR.t1397 VPWR.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 a_4861_9615# XThC.TBN.t51 XThC.Tn[3].t3 VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1191 VGND.t2611 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t2610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1192 VGND.t265 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1193 VGND.t2613 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t2612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1194 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t1865 VPWR.t1864 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1195 XThC.Tn[2].t2 XThC.TB3.t9 VGND.t1200 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1196 XThC.Tn[9].t10 XThC.TBN.t52 VPWR.t850 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1197 XThC.Tn[5].t8 XThC.TBN.t53 VGND.t1413 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 a_n1335_8107# XThR.TA2 XThR.TB2 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1199 VGND.t2615 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t2614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1200 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t1941 VGND.t1940 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1201 VGND.t2152 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t2151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1202 XA.XIR[15].XIC[5].icell.Ien VPWR.t1626 VPWR.t1628 VPWR.t1627 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1203 VGND.t1877 VGND.t1875 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1204 VPWR.t1296 XThC.TB1.t11 a_2979_9615# VPWR.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1205 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t1084 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1206 XThC.Tn[0].t1 XThC.TBN.t54 a_2979_9615# VPWR.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1207 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t1984 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1208 VPWR.t1277 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t1276 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1209 VPWR.t1119 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1210 XThR.Tn[12].t5 XThR.TB5 VPWR.t964 VPWR.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1211 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t1367 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1212 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t874 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1213 VGND.t2617 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t2616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1214 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1624 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1625 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1215 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t56 VGND.t387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1216 VGND.t1244 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t1243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1217 XThR.Tn[6].t10 XThR.TBN.t53 VGND.t1532 VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1218 a_n1049_5611# XThR.TBN.t54 XThR.Tn[5].t6 VPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1219 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t1331 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 VGND.t1534 XThR.TBN.t55 a_n997_2891# VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 VGND.t2299 XThR.TAN XThR.TB7 VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1222 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t757 VPWR.t756 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1223 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t145 VGND.t1286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1224 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1225 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t1985 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1226 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1227 VPWR.t192 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1228 VGND.t1086 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t1085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1229 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1230 VPWR.t1121 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t1120 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 a_n997_2667# XThR.TB4 XThR.Tn[11].t3 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1232 VPWR.t1623 VPWR.t1621 XA.XIR[12].XIC_15.icell.PUM VPWR.t1622 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1233 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t84 VGND.t614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1234 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t126 VPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1235 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1618 VPWR.t1620 VPWR.t1619 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1236 VGND.t2619 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t2618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1237 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t1294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1238 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t129 VGND.t1192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1239 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t1943 VGND.t1942 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1240 VGND.t2621 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t2620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1241 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1615 VPWR.t1617 VPWR.t1616 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1242 VGND.t1414 XThC.TBN.t55 XThC.Tn[1].t9 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1243 a_n1049_6405# XThR.TB5 VPWR.t962 VPWR.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1244 VGND.t2623 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t2622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1245 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t1867 VPWR.t1866 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1246 VPWR.t576 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1247 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1248 VGND.t1874 VGND.t1872 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1249 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t1087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1250 VGND.t1089 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t1088 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1251 VPWR.t128 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t127 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1252 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1253 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 VPWR.t1109 XThR.TB1.t10 XThR.Tn[8].t6 VPWR.t1108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1255 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t708 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t107 VGND.t846 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1257 VPWR.t883 XThR.TBN.t56 XThR.Tn[7].t6 VPWR.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1613 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1614 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 VGND.t514 XThC.TB2 XThC.Tn[1].t3 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1260 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1611 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1612 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1261 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t99 VGND.t760 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1262 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t1724 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1263 XThC.Tn[12].t2 XThC.TBN.t56 VPWR.t852 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1264 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1265 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1266 VGND.t2606 XThR.TB2 XThR.Tn[1].t10 VGND.t1430 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 XThR.Tn[1].t2 XThR.TBN.t57 a_n1049_7787# VPWR.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1268 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t2052 VGND.t2051 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1269 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t181 VGND.t1605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1270 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1271 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t2558 VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 VGND.t427 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1273 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t137 VGND.t1202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1274 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t578 VPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1275 VGND.t2625 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t2624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1276 VGND.t2627 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t2626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1277 VGND.t1871 VGND.t1869 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1870 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1278 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t130 VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1279 VGND.t1554 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t1553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1280 VGND.t1686 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t1685 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1281 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t196 VPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1282 XThR.Tn[9].t9 XThR.TB2 VPWR.t1904 VPWR.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1283 XThR.Tn[7].t1 XThR.TBN.t58 VGND.t1536 VGND.t1535 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1284 VPWR.t714 data[1].t2 XThC.TA2 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1285 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1856 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1286 VPWR.t580 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t579 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1287 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t1050 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1288 VPWR.t1610 VPWR.t1608 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1609 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1289 VGND.t1415 XThC.TBN.t57 a_7875_9569# VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1290 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1291 VPWR.t886 XThR.TBN.t59 XThR.Tn[13].t10 VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1292 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t221 VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1293 VPWR.t1607 VPWR.t1605 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1606 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1294 VGND.t1166 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t1165 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1295 a_8739_10571# data[0].t1 XThC.TA3 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1296 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t221 VGND.t2105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1297 VGND.t2629 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t2628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1298 VPWR.t1131 XThR.TB3.t9 XThR.Tn[10].t5 VPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1299 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t1279 VPWR.t1278 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1300 VGND.t2582 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t2581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1301 XThC.Tn[3].t2 XThC.TBN.t58 a_4861_9615# VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1303 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1304 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t1849 VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1305 XThR.Tn[5].t2 XThR.TB6 VGND.t1956 VGND.t1624 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1306 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t1548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1307 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t727 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1308 VPWR.t1408 XThR.TAN XThR.TB4 VPWR.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1309 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t2636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1310 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1311 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t2054 VGND.t2053 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1312 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1348 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1313 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t1091 VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t1034 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t2094 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1316 VGND.t2631 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t2630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1317 VGND.t429 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 VPWR.t132 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1319 VGND.t1868 VGND.t1866 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1320 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t582 VPWR.t581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1321 a_n997_715# XThR.TB7 XThR.Tn[14].t0 VGND.t1311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1322 VGND.t2556 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t2555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1323 VGND.t2633 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t2632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1324 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t230 VPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1325 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t2560 VGND.t2559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1326 VGND.t1769 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1327 VGND.t2635 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t2634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1328 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t2507 VGND.t2506 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1329 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t1093 VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 VGND.t853 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1331 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1332 VGND.t2542 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t2541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1333 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t908 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 VGND.t2211 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t2210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1335 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t1281 VPWR.t1280 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1336 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t23 VGND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1337 VPWR.t584 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t583 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1338 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t2592 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1339 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1352 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1340 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1341 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t2594 VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1342 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t2596 VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t1288 VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1344 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t61 VGND.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1345 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1346 VGND.t2213 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t2212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1347 VGND.t2215 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t2214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1348 VGND.t2258 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t2257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1349 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1350 VGND.t1095 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1351 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1352 XThC.Tn[1].t8 XThC.TBN.t59 VGND.t1416 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1353 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1354 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t2055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 VPWR.t1604 VPWR.t1602 XA.XIR[15].XIC_15.icell.PUM VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1356 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1357 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1358 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t1851 VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1359 a_7875_9569# XThC.TB2 XThC.Tn[9].t1 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1360 VPWR.t755 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t754 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1361 VGND.t2217 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t2216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1362 VGND.t1771 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1363 XA.XIR[15].XIC[14].icell.Ien VPWR.t1599 VPWR.t1601 VPWR.t1600 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1364 VGND.t2219 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t2218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1365 VPWR.t134 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t133 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1366 VGND.t267 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1367 VPWR.t291 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t290 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1368 VPWR.t1598 VPWR.t1596 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1597 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 XThR.Tn[13].t5 XThR.TB6 a_n997_1579# VGND.t1623 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1370 a_n1049_8581# XThR.TBN.t60 XThR.Tn[0].t6 VPWR.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1371 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1372 VPWR.t690 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1373 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t2508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1374 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t1726 VGND.t1725 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1375 VGND.t2221 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t2220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1376 VGND.t2223 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t2222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1377 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t105 VGND.t839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1378 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t2510 VGND.t2509 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1379 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t113 VGND.t868 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1380 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1381 VGND.t2225 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t2224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1382 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t692 VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1383 VGND.t2227 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t2226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1384 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t194 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1385 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t368 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1386 VGND.t2114 data[2].t1 XThC.TAN VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1388 VGND.t1537 XThR.TBN.t61 XThR.Tn[2].t5 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1389 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t1728 VGND.t1727 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1390 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t100 VGND.t763 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1391 a_n1049_5317# XThR.TB7 VPWR.t809 VPWR.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1392 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1393 VGND.t2303 XThC.TBN.t60 XThC.Tn[4].t5 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1394 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1395 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t370 VGND.t369 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1396 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t1097 VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1397 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t95 VGND.t747 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1398 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t81 VGND.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1399 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 VGND.t2229 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t2228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1401 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1402 VGND.t2231 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t2230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1403 VGND.t2233 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t2232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t50 VGND.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1405 XThR.Tn[3].t2 XThR.TB4 VGND.t2282 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1406 VGND.t2235 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t2234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1407 VPWR.t753 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t752 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1408 VGND.t1440 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t1439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1409 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t1869 VPWR.t1868 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1410 VPWR.t293 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1411 VPWR.t654 XThC.TB7 a_6243_9615# VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1412 VPWR.t393 XThC.TB6 XThC.Tn[13].t6 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VPWR.t1595 VPWR.t1593 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1594 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1414 VGND.t1253 data[1].t3 XThC.TA1 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1415 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t607 VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1416 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1008 VPWR.t1007 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1417 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t1175 VGND.t1174 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1418 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t1853 VPWR.t1852 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1419 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1590 VPWR.t1592 VPWR.t1591 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 VGND.t1364 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t1363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1421 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t101 VGND.t764 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1422 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t7 VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1423 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1358 VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1424 VPWR.t457 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t456 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1425 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t2246 VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1426 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t1635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1427 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t253 VGND.t2676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1428 VGND.t2305 XThC.TBN.t61 XThC.Tn[7].t2 VGND.t2304 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1429 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1730 VGND.t1729 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1430 VPWR.t1233 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1232 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1431 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1432 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t63 VGND.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1433 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1434 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t609 VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1435 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1436 XThR.Tn[12].t4 XThR.TB5 VPWR.t960 VPWR.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1437 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t372 VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 a_10915_9569# XThC.TBN.t62 VGND.t2307 VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1439 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t180 VGND.t1602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1440 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1036 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1441 XThR.Tn[6].t9 XThR.TBN.t62 VGND.t1539 VGND.t1538 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 VPWR.t1871 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t1870 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1443 XThC.Tn[3].t10 XThC.TB4.t7 VGND.t364 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1444 XThC.Tn[9].t5 XThC.TB2 VPWR.t399 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 VGND.t1751 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1446 a_n997_2667# XThR.TB4 XThR.Tn[11].t2 VGND.t1183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 VGND.t431 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1448 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t652 VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t325 VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1450 VGND.t1366 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t1365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1451 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t1010 VPWR.t1009 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1452 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t233 VGND.t2411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1453 VGND.t1100 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t1099 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1454 VPWR.t1290 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t1289 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1455 VPWR.t459 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t458 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1456 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t586 VPWR.t585 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1457 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1587 VPWR.t1589 VPWR.t1588 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1458 VPWR.t1235 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1234 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1459 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t1101 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1460 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t984 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1461 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t1051 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1462 VGND.t2297 XThR.TAN a_n1335_8331# VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1463 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t1976 VGND.t1975 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1465 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t1177 VGND.t1176 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1466 VGND.t855 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1468 VPWR.t1796 XThC.TBN.t63 XThC.Tn[9].t9 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1469 XA.XIR[15].XIC_15.icell.PUM VPWR.t1585 XA.XIR[15].XIC_15.icell.Ien VPWR.t1586 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t246 VGND.t2602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1471 a_10051_9569# XThC.TBN.t64 VGND.t2308 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1472 VGND.t486 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t485 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1473 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t44 VGND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1474 VPWR.t921 XThR.TBN.t63 XThR.Tn[7].t5 VPWR.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1475 VPWR.t1873 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t1872 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1476 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1368 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1477 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1583 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1584 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1478 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t47 VGND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1479 VPWR.t542 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1480 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1481 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1482 XThC.Tn[11].t1 XThC.TB4.t8 VPWR.t288 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1483 VGND.t1571 XThR.TBN.t64 XThR.Tn[1].t6 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1484 XThR.Tn[1].t1 XThR.TBN.t65 a_n1049_7787# VPWR.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1485 a_7651_9569# XThC.TBN.t65 VGND.t2309 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1486 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1350 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1487 VGND.t1368 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t1367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1488 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1360 VPWR.t1359 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1489 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1490 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t152 VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1491 VGND.t1370 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t1369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1492 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t1103 VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 VPWR.t1875 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t1874 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1494 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t1443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1495 VPWR.t588 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t587 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1496 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t1977 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1497 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1498 XThR.Tn[6].t1 XThR.TB7 VGND.t1310 VGND.t1309 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1499 a_n1049_5611# XThR.TB6 VPWR.t1139 VPWR.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1500 XThR.Tn[9].t8 XThR.TB2 VPWR.t1903 VPWR.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1501 VPWR.t1582 VPWR.t1580 XA.XIR[11].XIC_15.icell.PUM VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1502 VGND.t1372 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t1371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1503 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t2562 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1504 XThC.Tn[4].t4 XThC.TBN.t66 VGND.t2310 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 VGND.t1773 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1506 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t327 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1507 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t654 VGND.t653 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1508 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 VPWR.t924 XThR.TBN.t66 XThR.Tn[13].t9 VPWR.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1510 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t731 VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t751 VPWR.t750 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1512 VGND.t1865 VGND.t1863 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1864 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1513 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t2564 VGND.t2563 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t123 VGND.t1147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1515 VPWR.t1157 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t1156 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1516 VGND.t1105 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t1104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 VPWR.t1237 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1518 VPWR.t544 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1369 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1521 VGND.t1937 XThR.TB1.t11 XThR.Tn[0].t3 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1522 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t2 VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1523 XThR.Tn[5].t9 XThR.TBN.t67 VGND.t1572 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1524 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t709 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1525 XA.XIR[0].XIC[8].icell.PDM VGND.t1860 VGND.t1862 VGND.t1861 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1526 XA.XIR[0].XIC[14].icell.PDM VGND.t1857 VGND.t1859 VGND.t1858 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1527 VGND.t2295 XThR.TAN XThR.TB6 VGND.t2293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1528 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t629 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t985 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t2311 XThC.TBN.t67 XThC.Tn[0].t6 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 VGND.t1374 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t1373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1532 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t590 VPWR.t589 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1533 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t154 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1534 VGND.t1376 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t1375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 VGND.t1645 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1536 VGND.t1107 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t1106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1537 VGND.t1442 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t1441 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1538 VGND.t2312 XThC.TBN.t68 XThC.Tn[3].t7 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 VGND.t1378 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t1377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1540 VGND.t2321 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t2320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t2154 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t2153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1542 VPWR.t546 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1543 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1544 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1545 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1546 XThC.Tn[7].t1 XThC.TBN.t69 VGND.t2314 VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 VPWR.t1797 XThC.TBN.t70 XThC.Tn[12].t1 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 VGND.t1380 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t1379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1549 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t1362 VPWR.t1361 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1550 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t295 VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1551 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1577 VPWR.t1579 VPWR.t1578 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1552 VGND.t1382 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t1381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1553 VGND.t1384 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t1383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1554 VGND.t1556 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1555 VGND.t1688 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t1687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1556 VPWR.t1902 XThR.TB2 a_n1049_7787# VPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1557 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t156 VPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1558 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VGND.t1386 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t1385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1560 VGND.t1388 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t1387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1561 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t223 VGND.t2244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1562 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t694 VPWR.t693 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1563 VGND.t2316 XThC.TBN.t71 a_10915_9569# VGND.t2315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1564 VPWR.t1085 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1565 VPWR.t1012 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t1011 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1566 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t2248 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1567 VPWR.t749 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t748 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t1109 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1569 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t114 VGND.t875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1570 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t114 VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1571 XThC.Tn[11].t2 XThC.TB4.t9 a_8963_9569# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1572 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1573 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t1110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1574 VPWR.t297 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1575 VGND.t365 XThC.TB4.t10 XThC.Tn[3].t9 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1576 VGND.t784 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1577 XThR.Tn[14].t11 XThR.TBN.t68 VPWR.t926 VPWR.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1578 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1579 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1575 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1576 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1580 a_7875_9569# XThC.TBN.t72 VGND.t2317 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1581 VPWR.t1138 XThR.TB6 XThR.Tn[13].t3 VPWR.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1582 VGND.t2158 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t2157 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1584 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1585 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t251 VGND.t2671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1586 XA.XIR[0].XIC[3].icell.PDM VGND.t1854 VGND.t1856 VGND.t1855 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1589 XThC.Tn[11].t3 XThC.TB4.t11 a_8963_9569# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1590 VGND.t786 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t785 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1591 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t592 VPWR.t591 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1592 VGND.t788 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1593 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t299 VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1594 VGND.t1853 VGND.t1851 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1852 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1595 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1573 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1574 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1596 XThC.Tn[0].t9 XThC.TB1.t12 VGND.t2115 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1597 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t159 VGND.t1333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1598 VGND.t2318 XThC.TBN.t73 a_10051_9569# VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1599 VGND.t1246 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t1245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1600 VPWR.t1014 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t1013 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1601 VGND.t181 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1602 XThR.TB1.t0 XThR.TA1 VPWR.t26 VPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1603 VPWR.t1083 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t1082 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1605 XThR.Tn[13].t4 XThR.TB6 a_n997_1579# VGND.t1622 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1606 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1607 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t671 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1608 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t1113 VGND.t1112 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1609 VGND.t2544 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t2543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1610 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 VGND.t2319 XThC.TBN.t74 a_7651_9569# VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1612 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1239 VPWR.t1238 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1613 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t224 VGND.t2277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1614 XThC.TBN.t0 XThC.TAN2 VGND.t2085 VGND.t2084 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1615 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t1016 VPWR.t1015 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1570 VPWR.t1572 VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1617 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t2107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1618 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t24 VGND.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1619 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t2108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1620 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1621 a_n1335_7243# XThR.TA3 XThR.TB3.t2 VGND.t2672 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1622 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t1178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1624 XA.XIR[0].XIC[7].icell.PDM VGND.t1848 VGND.t1850 VGND.t1849 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1625 a_n1049_5317# XThR.TBN.t69 XThR.Tn[6].t6 VPWR.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1626 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t1115 VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_4067_9615# XThC.TB3.t10 VPWR.t702 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1629 VPWR.t1799 XThC.TBN.t75 XThC.Tn[7].t4 VPWR.t1798 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1630 VPWR.t747 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t746 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1631 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t174 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1632 XA.XIR[15].XIC[8].icell.Ien VPWR.t1567 VPWR.t1569 VPWR.t1568 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1633 VPWR.t301 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 VGND.t1573 XThR.TBN.t70 a_n997_1803# VGND.t1525 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1635 VPWR.t232 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1636 XThR.Tn[3].t9 XThR.TBN.t71 VGND.t1575 VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1637 VGND.t2160 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1638 VPWR.t696 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t695 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 VPWR.t932 XThC.TB4.t12 XThC.Tn[11].t4 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1640 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1641 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1642 VGND.t790 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1643 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t2566 VGND.t2565 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1644 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t1292 VPWR.t1291 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1645 VGND.t2276 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t2275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1646 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t176 VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1648 VPWR.t1081 VGND.t2697 Vbias.t4 VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X1649 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1650 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t150 VGND.t1291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1651 VGND.t1117 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t1116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1652 XThC.Tn[0].t5 XThC.TBN.t76 VGND.t815 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1653 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t72 VGND.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1654 VPWR.t1018 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t1017 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1655 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t118 VGND.t1010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 XThC.Tn[3].t6 XThC.TBN.t77 VGND.t816 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1657 VGND.t2005 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t2004 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1658 VGND.t1690 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t1689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1659 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t630 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1661 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t1858 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1663 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[8].XIC_15.icell.PUM VPWR.t1565 XA.XIR[8].XIC_15.icell.Ien VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 a_n1049_8581# XThR.TB1.t12 VPWR.t1111 VPWR.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1666 VGND.t2237 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t2236 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t200 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1668 VPWR.t1564 VPWR.t1562 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1563 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1669 VGND.t792 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1670 VGND.t2323 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1671 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t2109 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1672 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t1877 VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1673 VPWR.t234 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1674 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t978 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1675 VGND.t794 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1676 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 XThC.TB1.t1 XThC.TA1 a_3299_10575# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1678 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t1020 VPWR.t1019 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1679 VPWR.t745 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1680 VGND.t1038 XThR.TB3.t10 XThR.Tn[2].t3 VGND.t1037 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1681 XA.XIR[15].XIC[3].icell.Ien VPWR.t1559 VPWR.t1561 VPWR.t1560 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1682 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t178 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1683 VGND.t796 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1684 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t1364 VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1685 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1686 VPWR.t303 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1687 VPWR.t236 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t235 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1688 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1689 VPWR.t1159 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t1158 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t1731 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1691 VPWR.t478 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 VPWR.t136 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t135 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1693 VGND.t818 XThC.TBN.t78 XThC.Tn[6].t10 VGND.t817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1694 VGND.t798 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1695 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t249 VGND.t2609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1696 XThC.Tn[10].t8 XThC.TB3.t11 VPWR.t703 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1697 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t773 VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1698 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t582 VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1699 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t480 VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1700 VGND.t1847 VGND.t1845 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1846 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1701 VGND.t800 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1702 VGND.t802 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 XThC.Tn[14].t6 XThC.TB7 VPWR.t653 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1704 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t338 VGND.t337 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1705 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t2110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1706 VGND.t1119 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t1118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 VGND.t2116 XThC.TB1.t13 XThC.Tn[0].t10 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1708 VGND.t565 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t564 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t711 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1710 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 VGND.t804 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1713 XThR.Tn[8].t9 XThR.TBN.t72 VPWR.t929 VPWR.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1714 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t172 VGND.t1398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1715 VGND.t806 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1716 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t177 VGND.t1409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t213 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1718 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t547 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1719 VGND.t1248 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t1247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 VGND.t183 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t1879 VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1722 VGND.t185 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 VGND.t808 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t807 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1724 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t282 VPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1725 VGND.t38 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1726 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t1120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1727 a_n1049_5611# XThR.TBN.t73 XThR.Tn[5].t5 VPWR.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1728 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1054 VPWR.t1053 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1729 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t616 VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1730 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t1197 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1731 VGND.t2431 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t2430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1732 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t163 VGND.t1389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1733 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t580 VGND.t579 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1734 XThR.TAN2 data[7].t1 VGND.t319 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1735 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t305 VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1736 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t1774 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1737 XThC.Tn[14].t5 XThC.TB7 VPWR.t652 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1738 VPWR.t434 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1739 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1740 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t1052 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1741 VPWR.t1080 VGND.t2698 XA.XIR[0].XIC[13].icell.PUM VPWR.t1079 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1742 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t1121 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1743 VGND.t777 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1744 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t2249 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 XThC.TB2 XThC.TAN VPWR.t559 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1746 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1334 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1747 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t42 VGND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1748 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t1161 VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1749 XThR.Tn[5].t8 XThR.TBN.t74 VGND.t1577 VGND.t1576 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1750 VGND.t488 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1751 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t659 VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1752 VGND.t2433 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t2432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1753 VGND.t2162 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t2161 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 XThR.Tn[10].t9 XThR.TBN.t75 VPWR.t931 VPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 VPWR.t284 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1756 Vbias.t5 bias[1].t0 VPWR.t1801 VPWR.t1800 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X1757 VGND.t2164 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1758 a_5949_9615# XThC.TB6 VPWR.t392 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1759 VGND.t2435 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t2434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1760 VGND.t2437 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t2436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t219 VGND.t2099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1762 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t661 VGND.t660 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1763 VPWR.t645 XThC.TB3.t12 XThC.Tn[10].t3 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1764 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t549 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1765 VGND.t1844 VGND.t1842 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1766 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t226 VGND.t2279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1767 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t77 VGND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XThC.Tn[13].t8 XThC.TBN.t79 VPWR.t601 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1769 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t1123 VGND.t1122 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1770 a_n997_3755# XThR.TBN.t76 VGND.t1579 VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1771 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t64 VGND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1772 VPWR.t910 XThR.TBN.t77 XThR.Tn[14].t10 VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1773 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t48 VGND.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1774 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t943 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1775 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t202 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t618 VGND.t617 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t1125 VGND.t1124 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 VPWR.t436 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1781 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1782 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t1163 VPWR.t1162 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1783 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t153 VGND.t1304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1784 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t1198 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1785 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t188 VGND.t1631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1786 XThR.Tn[7].t0 XThR.TBN.t78 VGND.t1558 VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1787 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t146 VGND.t1287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1788 VPWR.t1558 VPWR.t1556 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1557 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1789 VGND.t490 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1790 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t519 VPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1791 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1354 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1792 VGND.t1127 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t1126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 XThC.TB4.t0 XThC.TAN VGND.t753 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1794 VPWR.t1137 XThR.TB6 XThR.Tn[13].t2 VPWR.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1795 VPWR.t406 XThR.TB3.t11 a_n1049_7493# VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1802 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1797 VPWR.t1833 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1832 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1798 VGND.t2439 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t2438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1799 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t307 VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1800 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t268 VPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 VPWR.t564 data[4].t3 XThR.TA3 VPWR.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1802 VGND.t1647 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1803 VGND.t2441 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t2440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1804 VGND.t1129 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t1128 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1805 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t1131 VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t663 VGND.t662 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XThC.Tn[6].t9 XThC.TBN.t80 VGND.t820 VGND.t819 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1808 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t551 VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1809 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t548 VPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1810 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t138 VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 VPWR.t1078 VGND.t2699 XA.XIR[0].XIC[6].icell.PUM VPWR.t1077 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1812 VPWR.t1056 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t1055 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 XThR.Tn[5].t1 XThR.TB6 VGND.t1955 VGND.t1620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1814 VPWR.t286 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1815 VPWR.t1267 XThC.TB5 a_5155_9615# VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1816 VPWR.t1555 VPWR.t1553 XA.XIR[3].XIC_15.icell.PUM VPWR.t1554 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1817 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1818 VPWR.t1552 VPWR.t1550 XA.XIR[7].XIC_15.icell.PUM VPWR.t1551 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1819 VGND.t2443 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t2442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1820 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1821 XThR.Tn[4].t2 XThR.TB5 VGND.t1625 VGND.t1624 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1822 a_4861_9615# XThC.TB4.t13 VPWR.t933 VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1823 a_5949_9615# XThC.TBN.t81 XThC.Tn[5].t5 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1824 VGND.t2445 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t2444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1825 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t340 VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1826 VGND.t1133 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t1132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t195 VGND.t1720 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1828 VGND.t821 XThC.TBN.t82 XThC.Tn[2].t9 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1829 VGND.t1135 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t1134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1830 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t102 VGND.t765 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1831 VPWR.t1298 XThC.TB1.t14 XThC.Tn[8].t9 VPWR.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1832 VGND.t433 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1833 a_5155_10571# XThC.TAN XThC.TB5 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1834 a_10915_9569# XThC.TBN.t83 VGND.t823 VGND.t822 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1835 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t521 VPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1836 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1355 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1837 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t631 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 VPWR.t1835 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1834 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1839 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t1165 VPWR.t1164 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1840 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t450 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1841 VGND.t2447 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t2446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1842 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t270 VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1843 XThC.Tn[3].t8 XThC.TB4.t14 VGND.t1580 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1844 VGND.t2449 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t2448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1845 VGND.t1649 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1846 VGND.t2239 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t2238 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t2325 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t550 VPWR.t549 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1849 VGND.t857 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t856 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1850 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t1776 VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1852 XThR.Tn[3].t8 XThR.TBN.t79 VGND.t1559 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1853 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1854 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t309 VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1855 VGND.t2451 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t2450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1856 VGND.t2453 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t2452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t272 VPWR.t271 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1858 VGND.t2455 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t2454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1859 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1548 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1549 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1860 a_10915_9569# XThC.TB7 XThC.Tn[14].t1 VGND.t1018 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1861 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1862 a_4387_10575# XThC.TAN VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1863 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t482 VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1864 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t108 VGND.t847 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1865 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t140 VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1866 VPWR.t1076 VGND.t2700 XA.XIR[0].XIC[1].icell.PUM VPWR.t1075 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1867 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t1058 VPWR.t1057 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1868 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t2250 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1869 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t213 VGND.t2064 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1870 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1871 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 a_10051_9569# XThC.TBN.t84 VGND.t824 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1876 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t2492 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1877 XThC.TB1.t2 XThC.TAN VPWR.t558 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1878 a_n1049_6699# XThR.TBN.t80 XThR.Tn[3].t5 VPWR.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1879 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t158 VGND.t1332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1880 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t193 VGND.t1712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 VGND.t1216 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t1215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1882 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1545 VPWR.t1547 VPWR.t1546 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1883 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t1179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1884 a_n1049_8581# XThR.TBN.t81 XThR.Tn[0].t5 VPWR.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1885 a_7651_9569# XThC.TBN.t85 VGND.t825 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1886 VGND.t1841 VGND.t1839 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1840 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1887 VGND.t1587 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1888 VPWR.t1155 XThC.TA3 a_6243_10571# VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1889 VPWR.t1544 VPWR.t1542 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1543 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1890 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t1960 VGND.t1959 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1891 VPWR.t1837 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1836 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1892 XThC.Tn[10].t4 XThC.TB3.t13 a_8739_9569# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1893 VGND.t1218 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t1217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1894 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t34 VGND.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1895 VGND.t1250 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t1249 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1896 VGND.t1561 XThR.TBN.t82 XThR.Tn[2].t6 VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1897 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t94 VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1898 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t96 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t30 VGND.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1900 XThR.TA1 data[5].t3 VGND.t1283 VGND.t1282 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1901 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t79 VGND.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1902 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1540 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1541 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1903 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t1778 VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t359 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1905 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XThR.Tn[12].t9 XThR.TBN.t83 VPWR.t913 VPWR.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1907 VGND.t1138 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t1137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1908 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t376 VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t1199 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XThR.Tn[12].t1 XThR.TB5 a_n997_1803# VGND.t1623 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1911 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t32 VGND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1912 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t1200 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1913 XThR.Tn[3].t1 XThR.TB4 VGND.t2281 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1914 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t205 VGND.t1972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1915 VGND.t1562 XThR.TBN.t84 a_n997_2667# VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1916 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t1140 VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1917 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1918 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t27 VGND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1919 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1920 VGND.t1220 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t1219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1921 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1537 VPWR.t1539 VPWR.t1538 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1922 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t944 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1923 VGND.t290 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1924 VGND.t2007 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t2006 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1925 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1926 a_5155_9615# XThC.TB5 VPWR.t1266 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1927 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t619 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1928 VPWR.t1265 XThC.TB5 XThC.Tn[12].t8 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1929 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t1779 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1930 VPWR.t523 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1931 XA.XIR[7].XIC_15.icell.PUM VPWR.t1535 XA.XIR[7].XIC_15.icell.Ien VPWR.t1536 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1932 VPWR.t408 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1933 VPWR.t1534 VPWR.t1532 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1533 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VGND.t492 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1935 XThC.Tn[5].t4 XThC.TBN.t86 a_5949_9615# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1936 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t97 VGND.t758 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1937 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t361 VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1938 VGND.t2095 XThC.TB5 XThC.Tn[4].t8 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1939 a_n1049_6405# XThR.TBN.t85 XThR.Tn[4].t5 VPWR.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1940 VPWR.t680 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t679 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1941 VPWR.t1145 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t1144 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1942 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t127 VGND.t1157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1943 XThC.Tn[2].t8 XThC.TBN.t87 VGND.t826 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1944 VPWR.t1387 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1945 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t1444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1947 a_5155_9615# XThC.TBN.t88 XThC.Tn[4].t1 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1948 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1962 VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1949 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t363 VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t381 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1951 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t183 VGND.t1607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1952 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1953 VPWR.t1406 XThR.TAN XThR.TB2 VPWR.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1954 Vbias.t0 bias[2].t0 VPWR.t517 VPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1955 XThC.Tn[8].t4 XThC.TB1.t15 a_7651_9569# VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t98 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1957 VGND.t718 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t85 VGND.t665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t1447 VGND.t1446 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t611 XThC.TA1 XThC.TB5 VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t1838 VGND.t1836 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 VGND.t1308 XThR.TB7 XThR.Tn[6].t0 VGND.t1307 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t2270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t215 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1966 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1171 VGND.t1170 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 VPWR.t525 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1969 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t452 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[4].XIC_15.icell.PUM VPWR.t1530 XA.XIR[4].XIC_15.icell.Ien VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t2272 VGND.t2271 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t28 VGND.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1973 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t1449 VGND.t1448 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[15].XIC[9].icell.Ien VPWR.t1527 VPWR.t1529 VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1975 VGND.t859 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1976 XThR.Tn[9].t0 XThR.TBN.t86 VPWR.t914 VPWR.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 VGND.t2126 XThC.TBN.t89 a_9827_9569# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1978 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1356 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t682 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 VGND.t567 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1981 VGND.t1451 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t1450 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t142 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t1222 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t1221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1984 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t527 VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1985 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1524 VPWR.t1526 VPWR.t1525 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1986 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1987 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1522 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1523 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1988 XThC.Tn[0].t11 XThC.TB1.t16 VGND.t2117 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t1224 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t1223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 VGND.t1226 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t1225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1991 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t2568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1992 VGND.t1651 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t1650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1993 a_10051_9569# XThC.TB6 XThC.Tn[13].t0 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t1701 VGND.t1700 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1995 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t743 VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VGND.t1228 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t1227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1997 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t418 VPWR.t417 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1998 VPWR.t684 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t683 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1999 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t100 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2000 VGND.t40 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2001 VPWR.t1147 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t1146 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t1400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2003 XThR.Tn[14].t9 XThR.TBN.t87 VPWR.t915 VPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1389 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1388 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 VPWR.t1521 VPWR.t1519 XA.XIR[0].XIC_15.icell.PUM VPWR.t1520 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2006 VPWR.t410 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2007 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t1452 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2008 a_n997_3755# XThR.TBN.t88 VGND.t1564 VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 XThR.Tn[8].t7 XThR.TB1.t13 VPWR.t1113 VPWR.t1112 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2010 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t1149 VPWR.t1148 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2012 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1173 VGND.t1172 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2013 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t148 VGND.t1289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 VGND.t1230 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t1229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2015 a_n1049_7787# XThR.TB2 VPWR.t1901 VPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t196 VGND.t1722 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t1589 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t1588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2018 VPWR.t93 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2019 a_n1331_2891# data[5].t4 VGND.t2289 VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND.t1232 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t1231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2021 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2022 VPWR.t1518 VPWR.t1516 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1517 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t779 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t778 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2024 VPWR.t529 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2025 XThR.TAN data[6].t1 VGND.t481 VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 XThR.Tn[2].t7 XThR.TBN.t89 a_n1049_7493# VPWR.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2027 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t737 VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t2260 VGND.t2259 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2029 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t741 VPWR.t740 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2030 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t229 VGND.t2286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2031 VGND.t187 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 VGND.t42 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2033 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t1453 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t1454 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VGND.t1234 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t1233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2036 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 VPWR.t1308 XThC.TBN.t90 XThC.Tn[8].t2 VPWR.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2038 XThR.Tn[10].t6 XThR.TB3.t12 VPWR.t1143 VPWR.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2039 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t979 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XThR.Tn[4].t9 XThR.TBN.t90 VGND.t1566 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2043 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1514 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1515 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t739 VPWR.t738 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t22 VGND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t2294 XThR.TAN XThR.TB5 VGND.t2293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t1236 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t1235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t292 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2049 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t1780 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2050 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t531 VPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2051 VGND.t2009 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t2008 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 VPWR.t412 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t411 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t594 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2054 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2055 VPWR.t97 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 VPWR.t1371 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t1370 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t59 VGND.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2060 VPWR.t1839 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2061 a_n997_3755# XThR.TB2 XThR.Tn[9].t5 VGND.t1429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 XThC.Tn[4].t0 XThC.TBN.t91 a_5155_9615# VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2063 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t414 VPWR.t413 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2064 VGND.t1238 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t1237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2065 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t209 VGND.t2003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2066 VGND.t1240 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t1239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t248 VGND.t2608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2068 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1511 VPWR.t1513 VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 VGND.t2166 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t2165 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 VGND.t2185 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t2184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2071 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t1963 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2072 VPWR.t1060 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t1059 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2073 VGND.t2495 XThR.TBN.t91 a_n997_1579# VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2074 VPWR.t50 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2075 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t1456 VGND.t1455 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2076 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2077 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2078 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t2262 VGND.t2261 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t88 VGND.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t110 VGND.t850 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2082 a_9827_9569# XThC.TB5 XThC.Tn[12].t5 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2083 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t712 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t17 VGND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1509 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1510 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t157 VGND.t1331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2087 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t532 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t2274 VGND.t2273 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[0].XIC[5].icell.PDM VGND.t1833 VGND.t1835 VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 VPWR.t1373 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t1372 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2091 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t1782 VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t222 VGND.t2111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2093 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t2494 VGND.t2493 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2094 VGND.t569 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t335 VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2096 XThR.TBN.t2 XThR.TAN2 VPWR.t995 VPWR.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2097 VGND.t2187 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t2186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2098 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1123 VPWR.t1122 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 VPWR.t987 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t986 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2100 VGND.t294 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2101 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t1964 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2102 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t632 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2103 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2104 VGND.t2011 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t2010 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2105 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1506 VPWR.t1508 VPWR.t1507 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VPWR.t52 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2107 XA.XIR[0].XIC_15.icell.PUM VPWR.t1504 XA.XIR[0].XIC_15.icell.Ien VPWR.t1505 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2109 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t686 VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2110 VGND.t2189 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t2188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 VGND.t2241 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t2240 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2112 VGND.t2327 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t2326 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t1842 XThR.TBN.t92 XThR.Tn[11].t9 VPWR.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1391 VPWR.t1390 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2115 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t2264 VGND.t2263 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t1909 data[1].t4 XThC.TA3 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 VPWR.t1062 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t1061 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2118 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1841 VPWR.t1840 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2119 a_8739_9569# XThC.TBN.t92 VGND.t2127 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 VGND.t1706 XThR.TAN2 XThR.TBN.t0 VGND.t1705 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XThC.Tn[6].t2 XThC.TB7 VGND.t1017 VGND.t1016 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1803 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t1346 VGND.t1345 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t383 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t0 XThR.TB5 a_n997_1803# VGND.t1622 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t1458 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t1457 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t2191 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t2190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2130 VGND.t720 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 VGND.t781 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t780 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t2193 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t2192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 a_n997_3979# XThR.TBN.t93 VGND.t2496 VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 XThC.TB7 XThC.TAN VGND.t750 VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 XA.XIR[0].XIC[0].icell.PDM VGND.t1830 VGND.t1832 VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2136 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1501 VPWR.t1503 VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2137 VGND.t2195 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t2194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2138 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t688 VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2139 VGND.t2197 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t2196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2140 XThC.Tn[8].t1 XThC.TBN.t93 VPWR.t1310 VPWR.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2141 VGND.t2243 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2142 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t2000 VGND.t1999 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2143 VGND.t861 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t860 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 VGND.t2199 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t2198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2145 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t672 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t369 VPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2147 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t1460 VGND.t1459 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2148 VGND.t571 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2150 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1188 VPWR.t1187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2151 a_n1049_6699# XThR.TB4 VPWR.t1396 VPWR.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2152 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t130 VGND.t1193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2153 VPWR.t54 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2154 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t2265 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2155 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t980 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2156 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t492 VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2157 VGND.t2201 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t2200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2158 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1499 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1500 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2159 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t173 VGND.t1399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2160 VGND.t1252 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1497 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1498 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1393 VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2163 VGND.t2203 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t2202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t2205 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t2204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VGND.t44 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2167 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t1461 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 VGND.t1463 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t1462 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2171 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t1709 data[1].t5 XThC.TA2 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 VPWR.t337 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2176 VPWR.t1496 VPWR.t1494 XA.XIR[14].XIC_15.icell.PUM VPWR.t1495 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2177 a_n997_2891# XThR.TBN.t94 VGND.t2498 VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 VGND.t2207 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t2206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2179 VGND.t2209 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t2208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2180 VGND.t1591 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t1590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2181 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 VPWR.t274 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2183 VPWR.t1493 VPWR.t1491 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1492 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2184 VGND.t1256 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t1255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2185 VGND.t1829 VGND.t1827 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2186 VGND.t1151 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t1490 VPWR.t1488 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1489 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VPWR.t99 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2189 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t1464 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2190 XThR.Tn[11].t1 XThR.TB4 a_n997_2667# VGND.t1319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2191 VGND.t1258 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t1257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2192 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t534 VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2193 VPWR.t1264 XThC.TB5 a_5155_9615# VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t713 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2195 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t93 VGND.t745 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t594 VGND.t593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t592 VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 VGND.t1260 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t1259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2199 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2201 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1190 VPWR.t1189 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t2407 VGND.t2406 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2203 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t2267 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2204 VGND.t2329 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t2500 XThR.TBN.t95 XThR.Tn[0].t9 VGND.t2499 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2207 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2208 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 a_n1049_6405# XThR.TB5 VPWR.t958 VPWR.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2210 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t214 VGND.t2065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2211 XThR.Tn[8].t0 XThR.TB1.t14 VPWR.t868 VPWR.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t239 VGND.t2486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2213 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2214 VGND.t1262 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t1261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t402 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t235 VGND.t2482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t1466 VGND.t1465 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t1264 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t1263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t86 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 VGND.t296 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2223 VGND.t1266 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t1265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2224 XThR.Tn[1].t9 XThR.TB2 VGND.t2605 VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2225 VGND.t298 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 VGND.t88 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2227 VPWR.t254 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t253 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2228 VGND.t2128 XThC.TBN.t94 a_8739_9569# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t339 VPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2230 VGND.t1268 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t1267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2231 VPWR.t1487 VPWR.t1485 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 XThC.Tn[1].t2 XThC.TB2 VGND.t513 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 VGND.t1015 XThC.TB7 XThC.Tn[6].t1 VGND.t1014 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t1467 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2235 VPWR.t1375 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t1374 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 VPWR.t1484 VPWR.t1482 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1483 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2237 a_6243_9615# XThC.TBN.t95 XThC.Tn[6].t5 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2238 VGND.t1270 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2239 VGND.t1272 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t1271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2240 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t56 VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[2].t10 XThR.TBN.t96 a_n1049_7493# VPWR.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t1469 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2243 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t255 VGND.t2688 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2244 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t1125 VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t220 VGND.t2104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2246 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t1348 VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XThR.Tn[13].t8 XThR.TBN.t97 VPWR.t1843 VPWR.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2248 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2249 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t538 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2250 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t826 VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t141 VGND.t1206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2252 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t385 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t590 VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XThR.Tn[10].t3 XThR.TB3.t13 VPWR.t783 VPWR.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t1336 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2256 XThR.Tn[4].t8 XThR.TBN.t98 VGND.t2501 VGND.t1576 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 VPWR.t101 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2258 VGND.t1826 VGND.t1824 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2259 VGND.t1954 XThR.TB6 XThR.Tn[5].t0 VGND.t1618 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 VGND.t1026 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t1025 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2261 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 VGND.t1274 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t1273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 a_4861_9615# XThC.TBN.t96 XThC.Tn[3].t1 VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t404 VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t254 VGND.t2677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2266 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t1945 VGND.t1944 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t1471 VGND.t1470 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 a_n997_3755# XThR.TB2 XThR.Tn[9].t4 VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 VGND.t2030 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t2029 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2270 VGND.t1276 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t1275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t1315 VPWR.t1314 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t171 VGND.t1397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t2032 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t1278 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t1277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t989 VPWR.t988 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 VPWR.t828 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t827 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2277 VGND.t1473 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t1472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1479 VPWR.t1481 VPWR.t1480 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2279 VGND.t1280 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t1279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VPWR.t1224 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1223 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t269 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t945 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2283 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t633 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t588 VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2286 VGND.t1475 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t1474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t166 VGND.t1392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 VGND.t494 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VPWR.t1129 XThR.TB3.t14 a_n1049_7493# VPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2290 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t194 VGND.t1719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2291 VPWR.t1377 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2292 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2293 VPWR.t1192 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2294 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t830 VPWR.t829 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2295 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1804 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2296 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2297 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t217 VGND.t2088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2298 VGND.t2457 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t2456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2299 VGND.t1153 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 VPWR.t103 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2301 XThC.TB2 XThC.TA2 a_3523_10575# VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VPWR.t1478 VPWR.t1476 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1477 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2303 VGND.t1155 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t1154 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VGND.t2459 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t2458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2305 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t991 VPWR.t990 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2306 XThR.Tn[4].t1 XThR.TB5 VGND.t1621 VGND.t1620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2307 VPWR.t1844 XThR.TBN.t99 XThR.Tn[14].t8 VPWR.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2308 VPWR.t1317 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2309 XThC.Tn[13].t5 XThC.TB6 VPWR.t391 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2310 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t1946 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2311 VGND.t501 XThC.TB6 XThC.Tn[5].t0 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2312 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t1948 VGND.t1947 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2313 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t112 VGND.t862 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2314 VPWR.t1845 XThR.TBN.t100 XThR.Tn[11].t8 VPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 VGND.t2461 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t2460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2316 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t1319 VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2317 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t153 VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2318 VGND.t1823 VGND.t1821 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1822 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2319 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t2002 VGND.t2001 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2320 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t201 VGND.t1952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2321 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2322 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t981 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XThC.Tn[9].t0 XThC.TB2 a_7875_9569# VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t1477 VGND.t1476 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2325 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 VGND.t1254 XThC.TA2 XThC.TB6 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 VGND.t512 XThC.TB2 XThC.Tn[1].t1 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t155 VGND.t1306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2330 VGND.t2463 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t2462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2331 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1474 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1475 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2332 XThC.Tn[6].t4 XThC.TBN.t97 a_6243_9615# VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2333 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t5 VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t2465 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t2464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 VGND.t2467 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t2466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t189 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2337 VGND.t1653 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2339 VPWR.t807 XThR.TB7 a_n1049_5317# VPWR.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 VPWR.t1379 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t1378 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2341 VGND.t1479 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t1478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 VPWR.t390 XThC.TB6 XThC.Tn[13].t4 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2343 VPWR.t1194 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2344 a_n997_3979# XThR.TBN.t101 VGND.t2502 VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t256 VPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2346 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t1381 VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2348 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t125 VGND.t1149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2349 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1471 VPWR.t1473 VPWR.t1472 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 VGND.t2469 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t2468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t2471 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t2470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t71 VGND.t553 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t2280 XThR.TB4 XThR.Tn[3].t0 VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t135 VGND.t1198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t650 VPWR.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# XThC.TBN.t98 XThC.Tn[2].t5 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 VPWR.t737 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t736 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2358 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t155 VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t86 VGND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1196 VPWR.t1195 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2361 VGND.t2473 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t2472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VGND.t1820 VGND.t1818 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2363 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t993 VPWR.t992 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2364 VPWR.t420 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2365 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t392 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2366 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t244 VGND.t2600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t1480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2368 VPWR.t258 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 a_n1049_6699# XThR.TBN.t102 XThR.Tn[3].t4 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 XA.XIR[0].XIC[11].icell.PDM VGND.t1815 VGND.t1817 VGND.t1816 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2372 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t1482 VGND.t1481 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2373 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t70 VGND.t519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2374 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t247 VGND.t2603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XThC.Tn[3].t0 XThC.TBN.t99 a_4861_9615# VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t119 VGND.t1023 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1469 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1470 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 VPWR.t719 bias[0].t0 Vbias.t3 VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X2379 XThC.TA1 data[0].t3 VGND.t981 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VGND.t2168 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t2167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2381 VPWR.t1395 XThR.TB4 XThR.Tn[11].t5 VPWR.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2382 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t2422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2383 XA.XIR[0].XIC[2].icell.PDM VGND.t1812 VGND.t1814 VGND.t1813 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2384 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t151 VGND.t1293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2385 VGND.t722 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2386 VGND.t2504 XThR.TBN.t103 a_n997_715# VGND.t2503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 a_n997_2891# XThR.TBN.t104 VGND.t2505 VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2388 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t1704 VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2389 VGND.t1811 VGND.t1809 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2390 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t260 VPWR.t259 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2391 VPWR.t1815 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t1814 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2392 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t1383 VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2393 VPWR.t735 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2394 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1466 VPWR.t1468 VPWR.t1467 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2395 VPWR.t422 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2396 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2397 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t946 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2398 XThR.Tn[11].t0 XThR.TB4 a_n997_2667# VGND.t2103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2399 VPWR.t1465 VPWR.t1463 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1464 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2400 VGND.t283 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2401 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2402 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t51 VGND.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2403 VPWR.t398 XThC.TB2 XThC.Tn[9].t4 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2404 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t1817 VPWR.t1816 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2405 a_n997_3979# XThR.TB1.t15 XThR.Tn[8].t1 VGND.t1429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2406 VGND.t1484 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t1483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2407 VGND.t496 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2408 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t208 VGND.t1986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2409 VPWR.t1312 XThC.TBN.t100 XThC.Tn[8].t0 VPWR.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2410 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t68 VGND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2411 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2412 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t2042 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2413 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t1330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2414 a_n1335_8331# XThR.TA1 XThR.TB1.t1 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2415 VPWR.t341 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t340 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2416 XA.XIR[0].XIC[6].icell.PDM VGND.t1806 VGND.t1808 VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2417 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t1995 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2418 a_n1049_6405# XThR.TBN.t105 XThR.Tn[4].t4 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2419 XA.XIR[15].XIC[7].icell.Ien VPWR.t1460 VPWR.t1462 VPWR.t1461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2420 XThR.Tn[7].t4 XThR.TBN.t106 VPWR.t12 VPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2421 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t1486 VGND.t1485 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2422 VPWR.t262 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2423 VGND.t1805 VGND.t1803 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2424 VPWR.t371 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t370 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2425 XThC.Tn[9].t8 XThC.TBN.t101 VPWR.t1313 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2426 XThR.Tn[1].t5 XThR.TBN.t107 VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2427 VPWR.t1459 VPWR.t1457 XA.XIR[13].XIC_15.icell.PUM VPWR.t1458 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2428 VGND.t2475 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t2474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2429 VGND.t1593 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t1592 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t534 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t1997 VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t1582 VGND.t1581 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t1488 VGND.t1487 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2434 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1226 VPWR.t1225 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t1819 VPWR.t1818 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2436 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t2130 VGND.t2129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2437 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t21 VGND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2438 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2439 VPWR.t73 XThC.TBN.t102 XThC.Tn[11].t9 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2440 VPWR.t733 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t732 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2441 VPWR.t1136 XThR.TB6 a_n1049_5611# VPWR.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2442 VGND.t1490 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2443 a_n997_2891# XThR.TB3.t15 XThR.Tn[10].t1 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2444 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2445 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t92 VGND.t744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2446 VPWR.t424 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2447 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2448 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1455 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1456 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2449 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t62 VGND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2450 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t624 VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t626 VGND.t625 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2453 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2454 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t439 VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2456 VGND.t2477 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t2476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2457 XA.XIR[15].XIC[11].icell.Ien VPWR.t1452 VPWR.t1454 VPWR.t1453 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2458 VGND.t1599 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 VGND.t1492 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[11].XIC_15.icell.PUM VPWR.t1450 XA.XIR[11].XIC_15.icell.Ien VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2461 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2462 VGND.t2479 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t2478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2463 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2464 VGND.t2331 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 VGND.t1494 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2466 XThC.Tn[2].t4 XThC.TBN.t103 a_4067_9615# VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2467 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t2043 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2468 VPWR.t494 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 VPWR.t343 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2470 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2471 VGND.t2292 XThR.TAN XThR.TB4 VGND.t2291 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2472 VPWR.t1449 VPWR.t1447 XA.XIR[10].XIC_15.icell.PUM VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2473 VGND.t2481 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t2480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2474 XA.XIR[15].XIC[2].icell.Ien VPWR.t1444 VPWR.t1446 VPWR.t1445 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2475 VGND.t983 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t982 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2476 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t1321 VPWR.t1320 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2477 VGND.t1431 XThR.TB1.t16 XThR.Tn[0].t0 VGND.t1430 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2478 VPWR.t504 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t503 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2479 VPWR.t264 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2480 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t333 VPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2481 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t9 VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2482 VPWR.t496 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2483 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2484 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2485 VGND.t724 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t723 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2486 VGND.t985 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2487 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1441 VPWR.t1443 VPWR.t1442 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2488 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t38 VGND.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2489 a_8739_9569# XThC.TBN.t104 VGND.t121 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2490 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t629 VGND.t628 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2491 XThC.Tn[6].t0 XThC.TB7 VGND.t1013 VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2492 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t1821 VPWR.t1820 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2493 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t2132 VGND.t2131 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t334 VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2495 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2496 VGND.t987 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2497 VGND.t123 XThC.TBN.t105 XThC.Tn[7].t0 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2498 XThC.Tn[12].t0 XThC.TBN.t106 VPWR.t75 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2499 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t107 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2500 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t2044 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2501 VGND.t285 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2502 XThC.Tn[12].t4 XThC.TB5 a_9827_9569# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2503 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t199 VGND.t1949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2504 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t633 VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1337 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2507 a_8963_9569# XThC.TB4.t15 XThC.Tn[11].t5 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2508 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t154 VGND.t1305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2509 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2510 VGND.t989 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2511 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1439 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2512 VGND.t991 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t990 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2513 VGND.t90 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 VGND.t864 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2515 XThR.Tn[13].t1 XThR.TB6 VPWR.t1135 VPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2516 VGND.t993 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t992 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2517 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t109 VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2518 VGND.t1028 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t1027 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2519 VGND.t995 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2520 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t936 VPWR.t935 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2521 VGND.t191 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2522 VPWR.t506 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t505 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2523 VGND.t46 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t1243 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2525 VGND.t125 XThC.TBN.t107 a_7875_9569# VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2526 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1496 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2528 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2529 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t731 VPWR.t730 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2530 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2531 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t115 VGND.t928 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2532 VGND.t997 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2533 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t426 VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t266 VPWR.t265 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2535 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t230 VGND.t2287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2536 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t1385 VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2537 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2538 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2539 VPWR.t1074 VGND.t2701 XA.XIR[0].XIC[12].icell.PUM VPWR.t1073 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2540 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2541 a_8963_9569# XThC.TBN.t108 VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2542 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2543 VGND.t1595 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t1594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2545 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t635 VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2546 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2547 VPWR.t1438 VPWR.t1436 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1437 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2548 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t1350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2552 VPWR.t938 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t937 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2553 VGND.t2170 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t2169 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2554 XThC.Tn[11].t8 XThC.TBN.t109 VPWR.t76 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2555 VPWR.t1323 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2556 VGND.t999 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t998 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2557 XThR.Tn[6].t5 XThR.TBN.t108 a_n1049_5317# VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2558 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1805 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2559 VPWR.t934 XThC.TB4.t16 XThC.Tn[11].t6 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2560 XThR.TB7 XThR.TAN a_n1319_5317# VPWR.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2561 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2562 VGND.t1001 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t1000 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2563 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t411 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t397 VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t2269 VGND.t2268 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t1499 VGND.t1498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 VGND.t2034 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t2033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2568 VGND.t1003 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t1002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2569 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t428 VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t729 VPWR.t728 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2571 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t1501 VGND.t1500 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2572 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t111 VGND.t851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2573 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t167 VGND.t1393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2574 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t189 VGND.t1654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2575 VPWR.t1072 VGND.t2702 XA.XIR[0].XIC[10].icell.PUM VPWR.t1071 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2576 VPWR.t646 XThC.TB3.t14 a_4067_9615# VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2577 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2578 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2579 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2580 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2581 VGND.t26 XThR.TBN.t109 a_n997_1803# VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2582 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t1583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2583 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2584 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1215 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t1244 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2586 XA.XIR[10].XIC_15.icell.PUM VPWR.t1434 XA.XIR[10].XIC_15.icell.Ien VPWR.t1435 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2587 a_3773_9615# XThC.TB2 VPWR.t396 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2588 VPWR.t1433 VPWR.t1431 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2589 VGND.t1005 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t1004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2590 VGND.t63 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 VGND.t2333 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t2332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2592 VPWR.t940 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t939 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2593 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t949 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2594 VPWR.t1394 XThR.TB4 XThR.Tn[11].t4 VPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2595 a_n997_715# XThR.TBN.t110 VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2596 VGND.t1007 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t1006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2597 VPWR.t870 XThR.TB1.t17 a_n1049_8581# VPWR.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2598 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1806 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2599 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t276 VPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2600 XThR.Tn[14].t5 XThR.TB7 VPWR.t805 VPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2601 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t842 VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2602 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t1911 VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2603 VGND.t1657 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t1656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2604 VGND.t129 XThC.TBN.t110 XThC.Tn[3].t5 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2605 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t498 VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2606 VGND.t2062 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t2061 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2607 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t1503 VGND.t1502 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2608 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2609 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t848 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2610 VPWR.t942 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2611 XThC.Tn[1].t0 XThC.TB2 VGND.t511 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2612 VPWR.t727 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t726 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2613 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2614 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1182 VPWR.t1181 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2615 VPWR.t1251 XThC.TAN2 XThC.TBN.t2 VPWR.t1250 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2616 VPWR.t1218 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1217 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2617 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t2664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2618 VPWR.t430 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2619 VGND.t1659 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t1658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2620 VPWR.t1430 VPWR.t1428 XA.XIR[6].XIC_15.icell.PUM VPWR.t1429 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2621 VGND.t1661 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t1660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2622 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2623 XThR.Tn[2].t2 XThR.TB3.t16 VGND.t313 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2624 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t2666 VGND.t2665 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2625 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t536 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2626 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t191 VGND.t1682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2627 VGND.t1663 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t1662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2628 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t432 VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2629 VGND.t1802 VGND.t1800 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 VGND.t1665 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t1664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2631 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t740 VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2632 a_n997_3979# XThR.TB1.t18 XThR.Tn[8].t2 VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2633 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t87 VGND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2634 a_3299_10575# XThC.TAN VGND.t748 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2635 VGND.t1505 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t1504 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2636 VGND.t30 XThR.TBN.t111 XThR.Tn[6].t8 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 VPWR.t1070 VGND.t2703 XA.XIR[0].XIC[5].icell.PUM VPWR.t1069 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2638 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2639 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2640 VPWR.t1184 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2641 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2642 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1425 VPWR.t1427 VPWR.t1426 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2643 VGND.t1667 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t1666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VGND.t1669 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t1668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2645 VGND.t1030 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t1029 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 VGND.t1601 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2647 VGND.t1671 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t1670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2648 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t500 VPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2649 VGND.t271 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2650 VGND.t1673 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t1672 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2651 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2652 VGND.t2335 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t2334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2653 VPWR.t78 XThC.TBN.t111 XThC.Tn[10].t0 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2654 VGND.t48 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2655 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t1506 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2656 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2657 VGND.t130 XThC.TBN.t112 a_8963_9569# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2658 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t278 VPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2659 VGND.t1675 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t1674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2660 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t541 VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2661 VPWR.t462 XThC.TA1 a_5155_10571# VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2662 VPWR.t651 XThC.TB7 XThC.Tn[14].t4 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2663 XThR.Tn[1].t4 XThR.TBN.t112 VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2664 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t508 VPWR.t507 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t1913 VPWR.t1912 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2666 VGND.t1677 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t1676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2667 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t502 VPWR.t501 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2668 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t1823 VPWR.t1822 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2669 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t160 VGND.t1344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2670 VPWR.t1154 XThC.TA3 XThC.TB3.t2 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2671 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1186 VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2672 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2673 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t124 VGND.t1148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2674 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t240 VGND.t2487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2675 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2676 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t2667 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2677 XThR.Tn[8].t8 XThR.TBN.t113 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2678 VPWR.t510 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t509 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2679 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t1507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2680 XThR.Tn[5].t4 XThR.TBN.t114 a_n1049_5611# VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2681 a_n997_2891# XThR.TB3.t17 XThR.Tn[10].t2 VGND.t1183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2682 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2683 XThR.TB6 XThR.TAN a_n1319_5611# VPWR.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2684 VPWR.t1424 VPWR.t1422 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1423 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2685 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t18 VGND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2686 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t83 VGND.t603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2687 a_n1049_7787# XThR.TBN.t115 XThR.Tn[1].t0 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2688 a_3773_9615# XThC.TBN.t113 XThC.Tn[1].t5 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2689 VPWR.t1404 XThR.TAN XThR.TB3.t0 VPWR.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2690 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t1508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2691 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1339 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2692 a_4067_9615# XThC.TB3.t15 VPWR.t647 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2693 VGND.t1679 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t1678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2694 VPWR.t648 XThC.TB3.t16 XThC.Tn[10].t5 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2695 VPWR.t80 XThC.TBN.t114 XThC.Tn[14].t9 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2696 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t484 VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2697 VGND.t1799 VGND.t1797 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2698 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t950 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2699 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t1510 VGND.t1509 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2700 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t161 VGND.t1351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2701 VGND.t1032 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t1031 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2702 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t15 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2703 VGND.t34 XThR.TBN.t116 XThR.Tn[0].t8 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2704 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t187 VGND.t1630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2705 VGND.t927 XThC.TB3.t17 XThC.Tn[2].t0 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2706 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t1245 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2707 XThR.Tn[10].t8 XThR.TBN.t117 VPWR.t18 VPWR.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2708 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t543 VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t1512 VGND.t1511 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2710 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2711 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t242 VGND.t2598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2712 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t48 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2713 VGND.t1681 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t1680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2714 VPWR.t389 XThC.TB6 a_5949_9615# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2715 XThR.Tn[1].t8 XThR.TB2 VGND.t2604 VGND.t1934 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2716 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t131 VGND.t1194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2717 VGND.t36 XThR.TBN.t118 a_n997_3755# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2718 VPWR.t367 data[3].t1 XThC.TAN2 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2719 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t90 VGND.t738 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2720 a_2979_9615# XThC.TB1.t17 VPWR.t438 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2721 XThC.Tn[3].t4 XThC.TBN.t115 VGND.t162 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2722 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t725 VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2723 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t218 VGND.t2089 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2724 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t869 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2725 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t2408 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2726 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t635 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2727 VPWR.t623 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t622 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2728 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t52 VGND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2729 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1220 VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2730 a_5949_10571# XThC.TAN XThC.TB6 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2731 VPWR.t486 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t485 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2732 VPWR.t146 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2733 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2036 VGND.t2035 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2734 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2735 XThR.Tn[13].t0 XThR.TB6 VPWR.t1134 VPWR.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2736 VPWR.t1228 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1227 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2737 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t139 VGND.t1204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2738 a_n1049_7493# XThR.TB3.t18 VPWR.t1133 VPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2739 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1807 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2741 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t538 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t742 VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2743 VGND.t1796 VGND.t1794 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2744 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t2424 VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2745 VGND.t903 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t902 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2746 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t2038 VGND.t2037 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2747 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t14 VGND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2748 VPWR.t440 XThC.TB1.t18 XThC.Tn[8].t8 VPWR.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2749 VGND.t726 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t725 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2750 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t12 VGND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2751 VGND.t1619 XThR.TB5 XThR.Tn[4].t0 VGND.t1618 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2752 XThC.Tn[10].t1 XThC.TBN.t116 VPWR.t110 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2753 VGND.t164 XThC.TBN.t117 XThC.Tn[6].t8 VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2754 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t2409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2755 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2756 VPWR.t345 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2757 VPWR.t625 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2758 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2759 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t636 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[3].XIC_15.icell.PUM VPWR.t1420 XA.XIR[3].XIC_15.icell.Ien VPWR.t1421 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t1568 VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2763 VGND.t905 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t904 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2764 VGND.t273 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t1514 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t1513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t2337 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t2336 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 VGND.t287 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VGND.t498 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2769 VPWR.t148 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2770 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t554 VPWR.t553 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2771 VPWR.t1402 XThC.TB4.t17 a_4861_9615# VPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2772 VPWR.t917 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t916 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2773 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t347 VPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2774 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t1515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2775 VGND.t1517 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t1516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2777 VGND.t907 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2778 XThR.Tn[6].t4 XThR.TBN.t119 a_n1049_5317# VPWR.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2779 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1418 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1419 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2780 a_10915_9569# XThC.TB7 XThC.Tn[14].t0 VGND.t1011 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2781 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t723 VPWR.t722 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2782 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1222 VPWR.t1221 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2783 VGND.t909 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2784 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t1006 VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2785 VGND.t166 XThC.TBN.t118 a_10915_9569# VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2786 VPWR.t488 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t487 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2787 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t280 VPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2788 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t2040 VGND.t2039 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2789 VGND.t103 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2790 VGND.t911 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2791 VPWR.t150 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2792 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t1915 VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2793 VPWR.t919 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t918 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 VPWR.t1068 VGND.t2704 XA.XIR[0].XIC[14].icell.PUM VPWR.t1067 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2795 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t1518 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t2428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2797 XThC.Tn[1].t4 XThC.TBN.t119 a_3773_9615# VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2798 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t116 VGND.t1008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2799 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2800 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t2427 VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2801 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t1570 VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2802 VGND.t913 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2803 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t136 VGND.t1201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2804 XThC.Tn[14].t8 XThC.TBN.t120 VPWR.t111 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2805 VGND.t915 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2806 VGND.t917 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t916 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2807 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t1519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2808 VGND.t1597 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t1596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2809 VGND.t2136 XThR.TBN.t120 a_n997_715# VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2810 VPWR.t1417 VPWR.t1415 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1416 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2811 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t349 VPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2812 VPWR.t627 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2813 VPWR.t803 XThR.TB7 XThR.Tn[14].t4 VPWR.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2814 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2815 VGND.t1793 VGND.t1791 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2816 VGND.t919 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t918 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2817 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t106 VGND.t845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2818 XThR.TA2 data[5].t5 VGND.t2113 VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2819 XThR.Tn[0].t4 XThR.TBN.t121 a_n1049_8581# VPWR.t1325 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2820 VGND.t1034 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t1033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2822 a_5949_9615# XThC.TB6 VPWR.t388 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2823 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t2139 VGND.t2138 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2824 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t198 VGND.t1752 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2825 VGND.t1036 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t1035 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 VGND.t2172 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t2171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2827 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t556 VPWR.t555 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2828 VGND.t168 XThC.TBN.t121 a_10051_9569# VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2829 VGND.t921 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t920 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2830 VGND.t105 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 VGND.t2156 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t2155 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15

*** ANTON
* X2832 Vbias.t260 VGND.t922 sky130_fd_pr__cap_mim_m3_1 l=4.81 w=11.82
*X2832 Vbias.t260 VGND.t922 sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
*CVb Vbias.t260 VGND.t922 120f


X2833 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t1520 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2834 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t1521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2835 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t2140 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2836 XA.XIR[0].XIC[9].icell.PDM VGND.t1788 VGND.t1790 VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2837 VPWR.t112 XThC.TBN.t122 XThC.Tn[11].t7 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2838 VGND.t170 XThC.TBN.t123 a_7651_9569# VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2839 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t721 VPWR.t720 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2840 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t35 VGND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2841 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t490 VPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2842 XThR.Tn[2].t9 XThR.TBN.t122 VGND.t2137 VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2843 VPWR.t801 XThR.TB7 a_n1049_5317# VPWR.t800 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2844 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t1182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2845 VGND.t924 Vbias.t261 XA.XIR[15].XIC_15.icell.SM VGND.t923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2846 a_8739_9569# XThC.TB3.t18 XThC.Tn[10].t2 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2847 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t948 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2848 VGND.t866 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t865 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2849 VGND.t92 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2850 VPWR.t1327 XThR.TBN.t123 XThR.Tn[12].t8 VPWR.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2851 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t2425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2852 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t1721 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2853 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2854 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t40 VGND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2855 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t2668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2856 VPWR.t1414 VPWR.t1412 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1413 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2857 VGND.t65 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2858 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t104 VGND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2859 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t2670 VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2860 VGND.t926 Vbias.t262 XA.XIR[13].XIC[2].icell.SM VGND.t925 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2861 VPWR.t1825 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n2840 VGND.n7 32072.7
R1 VGND.n3018 VGND.n3017 21075.4
R2 VGND.n2876 VGND.n2844 13477
R3 VGND.n2844 VGND.n2843 11635.6
R4 VGND.n3011 VGND.n3010 9309.26
R5 VGND.n2909 VGND.n2876 9223.7
R6 VGND.n2910 VGND.n2909 9223.7
R7 VGND.n2963 VGND.n34 9223.7
R8 VGND.n2996 VGND.n2963 9223.7
R9 VGND.n2997 VGND.n2996 7447.41
R10 VGND.n1509 VGND.n1508 7387.65
R11 VGND.n1508 VGND.n1507 7387.65
R12 VGND.n2834 VGND.n147 7387.65
R13 VGND.n3016 VGND.n3015 7387.65
R14 VGND.n3015 VGND.n3014 7387.65
R15 VGND.n3014 VGND.n3013 7387.65
R16 VGND.n3013 VGND.n3012 7387.65
R17 VGND.n3012 VGND.n3011 7387.65
R18 VGND.n2839 VGND.n2834 7048.53
R19 VGND.n1511 VGND.t1168 6324.96
R20 VGND.n3017 VGND.n3016 5925.05
R21 VGND.n2910 VGND.n34 5231.11
R22 VGND.n1291 VGND.t1124 5131.29
R23 VGND.n3010 VGND.n3009 5074.71
R24 VGND.n2843 VGND.n7 4937.78
R25 VGND.n3017 VGND.n7 4804.6
R26 VGND.n1110 VGND.n578 4542.17
R27 VGND.n2840 VGND.n2839 4343.1
R28 VGND.n3010 VGND 4240.58
R29 VGND.n2415 VGND.n273 4110.84
R30 VGND.n1295 VGND.n1293 3417.39
R31 VGND.n1295 VGND.n1294 3417.39
R32 VGND.n1513 VGND.n1512 3417.39
R33 VGND.n960 VGND.n580 3417.39
R34 VGND.n635 VGND.n177 3417.39
R35 VGND.n2833 VGND.n114 3417.39
R36 VGND.n2842 VGND.n2841 3417.39
R37 VGND.n2416 VGND.n2415 3331.79
R38 VGND.n2417 VGND.n2416 3331.79
R39 VGND.n2418 VGND.n2417 3331.79
R40 VGND.n2419 VGND.n2418 3331.79
R41 VGND.n2420 VGND.n2419 3331.79
R42 VGND.n2421 VGND.n2420 3331.79
R43 VGND.n2422 VGND.n2421 3331.79
R44 VGND.n2423 VGND.n2422 3331.79
R45 VGND.n2424 VGND.n2423 3331.79
R46 VGND.n2425 VGND.n2424 3331.79
R47 VGND.n2426 VGND.n2425 3331.79
R48 VGND.n2427 VGND.n2426 3331.79
R49 VGND.n2428 VGND.n2427 3331.79
R50 VGND.n2428 VGND.n32 3331.79
R51 VGND.n2999 VGND.n32 3331.79
R52 VGND.n2999 VGND.n2998 3331.79
R53 VGND.n1294 VGND.n578 3273.91
R54 VGND.n961 VGND.n579 3265.22
R55 VGND.n2840 VGND.n114 2756.52
R56 VGND.n2876 VGND.t135 2655.17
R57 VGND.n2909 VGND.t2490 2655.17
R58 VGND.n2998 VGND.n2997 2602.7
R59 VGND.n2834 VGND.n2833 2517.39
R60 VGND.n2837 VGND.n5 2229.43
R61 VGND.n3019 VGND.n5 2229.43
R62 VGND.n3019 VGND.n6 2229.43
R63 VGND.n2837 VGND.n6 2229.43
R64 VGND.n1293 VGND.n1292 2130.43
R65 VGND.n2843 VGND.n2842 2082.61
R66 VGND VGND.n34 1997.7
R67 VGND.n2963 VGND 1997.7
R68 VGND.n2996 VGND 1997.7
R69 VGND.n1506 VGND.n147 1831.57
R70 VGND.t29 VGND.n2910 1807.04
R71 VGND.n2994 VGND.t318 1785.51
R72 VGND.n1507 VGND.n580 1691.3
R73 VGND.n2922 VGND.t1784 1618.39
R74 VGND.t1319 VGND.n2962 1618.39
R75 VGND.t1623 VGND.n2995 1618.39
R76 VGND.n2844 VGND.t2499 1517.24
R77 VGND.n1510 VGND.n1509 1513.49
R78 VGND.n1511 VGND.n1510 1370.36
R79 VGND.n1292 VGND.n1291 1286.96
R80 VGND.n1510 VGND.t1789 1270.28
R81 VGND.n1083 VGND.t167 1268.93
R82 VGND.n1083 VGND.t70 1268.93
R83 VGND.n146 VGND.t128 1253.59
R84 VGND.t751 VGND.n146 1253.59
R85 VGND.n614 VGND.t500 1253.59
R86 VGND.t610 VGND.n614 1253.59
R87 VGND.n1021 VGND.t124 1253.59
R88 VGND.n1021 VGND.t169 1253.59
R89 VGND.n1052 VGND.t126 1253.59
R90 VGND.n1052 VGND.t68 1253.59
R91 VGND.n176 VGND.t510 1253.59
R92 VGND.t66 VGND.n176 1253.59
R93 VGND.n1506 VGND.t1834 1237.71
R94 VGND.n2839 VGND.n2838 1217.3
R95 VGND.n2922 VGND.t1328 1213.79
R96 VGND.n1111 VGND.n1110 1198.25
R97 VGND.n3009 VGND.n3008 1198.25
R98 VGND.n2652 VGND.n33 1180.79
R99 VGND.n3001 VGND.n3000 1180.79
R100 VGND.n2491 VGND.n2490 1180.79
R101 VGND.n2430 VGND.n2429 1180.79
R102 VGND.n2313 VGND.n261 1180.79
R103 VGND.n2127 VGND.n262 1180.79
R104 VGND.n2122 VGND.n263 1180.79
R105 VGND.n2338 VGND.n264 1180.79
R106 VGND.n1953 VGND.n265 1180.79
R107 VGND.n1948 VGND.n266 1180.79
R108 VGND.n2363 VGND.n267 1180.79
R109 VGND.n1779 VGND.n268 1180.79
R110 VGND.n1774 VGND.n269 1180.79
R111 VGND.n2388 VGND.n270 1180.79
R112 VGND.n1605 VGND.n271 1180.79
R113 VGND.n2408 VGND.n272 1180.79
R114 VGND.n1233 VGND.n273 1180.79
R115 VGND.n2414 VGND.n2413 1180.79
R116 VGND.n1290 VGND.n1289 1180.46
R117 VGND.n720 VGND.n679 1180.46
R118 VGND.n725 VGND.n724 1180.46
R119 VGND.n730 VGND.n729 1180.46
R120 VGND.n735 VGND.n734 1180.46
R121 VGND.n740 VGND.n739 1180.46
R122 VGND.n745 VGND.n744 1180.46
R123 VGND.n750 VGND.n749 1180.46
R124 VGND.n755 VGND.n754 1180.46
R125 VGND.n760 VGND.n759 1180.46
R126 VGND.n765 VGND.n764 1180.46
R127 VGND.n770 VGND.n769 1180.46
R128 VGND.n775 VGND.n774 1180.46
R129 VGND.n780 VGND.n779 1180.46
R130 VGND.n782 VGND.n781 1180.46
R131 VGND.n1230 VGND.n1229 1180.46
R132 VGND.n1228 VGND.n1227 1180.46
R133 VGND.n1211 VGND.n1210 1180.46
R134 VGND.n1209 VGND.n1208 1180.46
R135 VGND.n1198 VGND.n1197 1180.46
R136 VGND.n1196 VGND.n1195 1180.46
R137 VGND.n1179 VGND.n1178 1180.46
R138 VGND.n1177 VGND.n1176 1180.46
R139 VGND.n1166 VGND.n1165 1180.46
R140 VGND.n1164 VGND.n1163 1180.46
R141 VGND.n1147 VGND.n1146 1180.46
R142 VGND.n1145 VGND.n1144 1180.46
R143 VGND.n1134 VGND.n1133 1180.46
R144 VGND.n1132 VGND.n1131 1180.46
R145 VGND.n1124 VGND.n1123 1180.46
R146 VGND.n2579 VGND.n2578 1180.46
R147 VGND.n2707 VGND.n2706 1180.46
R148 VGND.n2705 VGND.n2704 1180.46
R149 VGND.n2699 VGND.n2698 1180.46
R150 VGND.n2697 VGND.n2696 1180.46
R151 VGND.n2691 VGND.n2690 1180.46
R152 VGND.n2689 VGND.n2688 1180.46
R153 VGND.n2683 VGND.n2682 1180.46
R154 VGND.n2681 VGND.n2680 1180.46
R155 VGND.n2675 VGND.n2674 1180.46
R156 VGND.n2673 VGND.n2672 1180.46
R157 VGND.n2667 VGND.n2666 1180.46
R158 VGND.n2665 VGND.n2664 1180.46
R159 VGND.n2659 VGND.n2658 1180.46
R160 VGND.n2657 VGND.n2656 1180.46
R161 VGND.n234 VGND.n233 1180.46
R162 VGND.n2720 VGND.n2719 1180.46
R163 VGND.n2725 VGND.n2724 1180.46
R164 VGND.n2730 VGND.n2729 1180.46
R165 VGND.n2735 VGND.n2734 1180.46
R166 VGND.n2740 VGND.n2739 1180.46
R167 VGND.n2745 VGND.n2744 1180.46
R168 VGND.n2750 VGND.n2749 1180.46
R169 VGND.n2755 VGND.n2754 1180.46
R170 VGND.n2760 VGND.n2759 1180.46
R171 VGND.n2765 VGND.n2764 1180.46
R172 VGND.n2770 VGND.n2769 1180.46
R173 VGND.n2775 VGND.n2774 1180.46
R174 VGND.n2780 VGND.n2779 1180.46
R175 VGND.n2782 VGND.n2781 1180.46
R176 VGND.n2516 VGND.n2515 1180.46
R177 VGND.n2514 VGND.n2513 1180.46
R178 VGND.n2509 VGND.n2508 1180.46
R179 VGND.n2434 VGND.n244 1180.46
R180 VGND.n2439 VGND.n2438 1180.46
R181 VGND.n2444 VGND.n2443 1180.46
R182 VGND.n2449 VGND.n2448 1180.46
R183 VGND.n2454 VGND.n2453 1180.46
R184 VGND.n2459 VGND.n2458 1180.46
R185 VGND.n2464 VGND.n2463 1180.46
R186 VGND.n2469 VGND.n2468 1180.46
R187 VGND.n2474 VGND.n2473 1180.46
R188 VGND.n2479 VGND.n2478 1180.46
R189 VGND.n2484 VGND.n2483 1180.46
R190 VGND.n2489 VGND.n2488 1180.46
R191 VGND.n2832 VGND.n2831 1180.46
R192 VGND.n371 VGND.n182 1180.46
R193 VGND.n373 VGND.n372 1180.46
R194 VGND.n2172 VGND.n2171 1180.46
R195 VGND.n2174 VGND.n2173 1180.46
R196 VGND.n2198 VGND.n2197 1180.46
R197 VGND.n2200 VGND.n2199 1180.46
R198 VGND.n2224 VGND.n2223 1180.46
R199 VGND.n2226 VGND.n2225 1180.46
R200 VGND.n2250 VGND.n2249 1180.46
R201 VGND.n2252 VGND.n2251 1180.46
R202 VGND.n2281 VGND.n2280 1180.46
R203 VGND.n2286 VGND.n2285 1180.46
R204 VGND.n2291 VGND.n2290 1180.46
R205 VGND.n2293 VGND.n2292 1180.46
R206 VGND.n1429 VGND.n1428 1180.46
R207 VGND.n1431 VGND.n1430 1180.46
R208 VGND.n2159 VGND.n2158 1180.46
R209 VGND.n2161 VGND.n2160 1180.46
R210 VGND.n2185 VGND.n2184 1180.46
R211 VGND.n2187 VGND.n2186 1180.46
R212 VGND.n2211 VGND.n2210 1180.46
R213 VGND.n2213 VGND.n2212 1180.46
R214 VGND.n2237 VGND.n2236 1180.46
R215 VGND.n2239 VGND.n2238 1180.46
R216 VGND.n2263 VGND.n2262 1180.46
R217 VGND.n2270 VGND.n2269 1180.46
R218 VGND.n2268 VGND.n2267 1180.46
R219 VGND.n2308 VGND.n2307 1180.46
R220 VGND.n2310 VGND.n2309 1180.46
R221 VGND.n1443 VGND.n1442 1180.46
R222 VGND.n1495 VGND.n1494 1180.46
R223 VGND.n1493 VGND.n1492 1180.46
R224 VGND.n1488 VGND.n1487 1180.46
R225 VGND.n1483 VGND.n1482 1180.46
R226 VGND.n1478 VGND.n1477 1180.46
R227 VGND.n1473 VGND.n1472 1180.46
R228 VGND.n1468 VGND.n1467 1180.46
R229 VGND.n1463 VGND.n1462 1180.46
R230 VGND.n1458 VGND.n1457 1180.46
R231 VGND.n1453 VGND.n1452 1180.46
R232 VGND.n1448 VGND.n1447 1180.46
R233 VGND.n2138 VGND.n2137 1180.46
R234 VGND.n2136 VGND.n2135 1180.46
R235 VGND.n2131 VGND.n2130 1180.46
R236 VGND.n1505 VGND.n1504 1180.46
R237 VGND.n626 VGND.n619 1180.46
R238 VGND.n628 VGND.n627 1180.46
R239 VGND.n1998 VGND.n1997 1180.46
R240 VGND.n2000 VGND.n1999 1180.46
R241 VGND.n2024 VGND.n2023 1180.46
R242 VGND.n2026 VGND.n2025 1180.46
R243 VGND.n2050 VGND.n2049 1180.46
R244 VGND.n2052 VGND.n2051 1180.46
R245 VGND.n2076 VGND.n2075 1180.46
R246 VGND.n2078 VGND.n2077 1180.46
R247 VGND.n2107 VGND.n2106 1180.46
R248 VGND.n2112 VGND.n2111 1180.46
R249 VGND.n2117 VGND.n2116 1180.46
R250 VGND.n2119 VGND.n2118 1180.46
R251 VGND.n652 VGND.n651 1180.46
R252 VGND.n654 VGND.n653 1180.46
R253 VGND.n1985 VGND.n1984 1180.46
R254 VGND.n1987 VGND.n1986 1180.46
R255 VGND.n2011 VGND.n2010 1180.46
R256 VGND.n2013 VGND.n2012 1180.46
R257 VGND.n2037 VGND.n2036 1180.46
R258 VGND.n2039 VGND.n2038 1180.46
R259 VGND.n2063 VGND.n2062 1180.46
R260 VGND.n2065 VGND.n2064 1180.46
R261 VGND.n2089 VGND.n2088 1180.46
R262 VGND.n2096 VGND.n2095 1180.46
R263 VGND.n2094 VGND.n2093 1180.46
R264 VGND.n2333 VGND.n2332 1180.46
R265 VGND.n2335 VGND.n2334 1180.46
R266 VGND.n959 VGND.n958 1180.46
R267 VGND.n954 VGND.n953 1180.46
R268 VGND.n949 VGND.n948 1180.46
R269 VGND.n944 VGND.n943 1180.46
R270 VGND.n939 VGND.n938 1180.46
R271 VGND.n934 VGND.n933 1180.46
R272 VGND.n929 VGND.n928 1180.46
R273 VGND.n924 VGND.n923 1180.46
R274 VGND.n919 VGND.n918 1180.46
R275 VGND.n914 VGND.n913 1180.46
R276 VGND.n909 VGND.n908 1180.46
R277 VGND.n904 VGND.n903 1180.46
R278 VGND.n1964 VGND.n1963 1180.46
R279 VGND.n1962 VGND.n1961 1180.46
R280 VGND.n1957 VGND.n1956 1180.46
R281 VGND.n1396 VGND.n1395 1180.46
R282 VGND.n1401 VGND.n1400 1180.46
R283 VGND.n1403 VGND.n1402 1180.46
R284 VGND.n1824 VGND.n1823 1180.46
R285 VGND.n1826 VGND.n1825 1180.46
R286 VGND.n1850 VGND.n1849 1180.46
R287 VGND.n1852 VGND.n1851 1180.46
R288 VGND.n1876 VGND.n1875 1180.46
R289 VGND.n1878 VGND.n1877 1180.46
R290 VGND.n1902 VGND.n1901 1180.46
R291 VGND.n1904 VGND.n1903 1180.46
R292 VGND.n1933 VGND.n1932 1180.46
R293 VGND.n1938 VGND.n1937 1180.46
R294 VGND.n1943 VGND.n1942 1180.46
R295 VGND.n1945 VGND.n1944 1180.46
R296 VGND.n1381 VGND.n1380 1180.46
R297 VGND.n1383 VGND.n1382 1180.46
R298 VGND.n1811 VGND.n1810 1180.46
R299 VGND.n1813 VGND.n1812 1180.46
R300 VGND.n1837 VGND.n1836 1180.46
R301 VGND.n1839 VGND.n1838 1180.46
R302 VGND.n1863 VGND.n1862 1180.46
R303 VGND.n1865 VGND.n1864 1180.46
R304 VGND.n1889 VGND.n1888 1180.46
R305 VGND.n1891 VGND.n1890 1180.46
R306 VGND.n1915 VGND.n1914 1180.46
R307 VGND.n1922 VGND.n1921 1180.46
R308 VGND.n1920 VGND.n1919 1180.46
R309 VGND.n2358 VGND.n2357 1180.46
R310 VGND.n2360 VGND.n2359 1180.46
R311 VGND.n1313 VGND.n1312 1180.46
R312 VGND.n1365 VGND.n1364 1180.46
R313 VGND.n1363 VGND.n1362 1180.46
R314 VGND.n1358 VGND.n1357 1180.46
R315 VGND.n1353 VGND.n1352 1180.46
R316 VGND.n1348 VGND.n1347 1180.46
R317 VGND.n1343 VGND.n1342 1180.46
R318 VGND.n1338 VGND.n1337 1180.46
R319 VGND.n1333 VGND.n1332 1180.46
R320 VGND.n1328 VGND.n1327 1180.46
R321 VGND.n1323 VGND.n1322 1180.46
R322 VGND.n1318 VGND.n1317 1180.46
R323 VGND.n1790 VGND.n1789 1180.46
R324 VGND.n1788 VGND.n1787 1180.46
R325 VGND.n1783 VGND.n1782 1180.46
R326 VGND.n1518 VGND.n1517 1180.46
R327 VGND.n1523 VGND.n1522 1180.46
R328 VGND.n1525 VGND.n1524 1180.46
R329 VGND.n1650 VGND.n1649 1180.46
R330 VGND.n1652 VGND.n1651 1180.46
R331 VGND.n1676 VGND.n1675 1180.46
R332 VGND.n1678 VGND.n1677 1180.46
R333 VGND.n1702 VGND.n1701 1180.46
R334 VGND.n1704 VGND.n1703 1180.46
R335 VGND.n1728 VGND.n1727 1180.46
R336 VGND.n1730 VGND.n1729 1180.46
R337 VGND.n1759 VGND.n1758 1180.46
R338 VGND.n1764 VGND.n1763 1180.46
R339 VGND.n1769 VGND.n1768 1180.46
R340 VGND.n1771 VGND.n1770 1180.46
R341 VGND.n1538 VGND.n1537 1180.46
R342 VGND.n1540 VGND.n1539 1180.46
R343 VGND.n1637 VGND.n1636 1180.46
R344 VGND.n1639 VGND.n1638 1180.46
R345 VGND.n1663 VGND.n1662 1180.46
R346 VGND.n1665 VGND.n1664 1180.46
R347 VGND.n1689 VGND.n1688 1180.46
R348 VGND.n1691 VGND.n1690 1180.46
R349 VGND.n1715 VGND.n1714 1180.46
R350 VGND.n1717 VGND.n1716 1180.46
R351 VGND.n1741 VGND.n1740 1180.46
R352 VGND.n1748 VGND.n1747 1180.46
R353 VGND.n1746 VGND.n1745 1180.46
R354 VGND.n2383 VGND.n2382 1180.46
R355 VGND.n2385 VGND.n2384 1180.46
R356 VGND.n1297 VGND.n1296 1180.46
R357 VGND.n1551 VGND.n1550 1180.46
R358 VGND.n1556 VGND.n1555 1180.46
R359 VGND.n1561 VGND.n1560 1180.46
R360 VGND.n1566 VGND.n1565 1180.46
R361 VGND.n1571 VGND.n1570 1180.46
R362 VGND.n1576 VGND.n1575 1180.46
R363 VGND.n1581 VGND.n1580 1180.46
R364 VGND.n1586 VGND.n1585 1180.46
R365 VGND.n1591 VGND.n1590 1180.46
R366 VGND.n1596 VGND.n1595 1180.46
R367 VGND.n1601 VGND.n1600 1180.46
R368 VGND.n1616 VGND.n1615 1180.46
R369 VGND.n1614 VGND.n1613 1180.46
R370 VGND.n1609 VGND.n1608 1180.46
R371 VGND.n835 VGND.n834 1180.46
R372 VGND.n840 VGND.n839 1180.46
R373 VGND.n892 VGND.n891 1180.46
R374 VGND.n890 VGND.n889 1180.46
R375 VGND.n885 VGND.n884 1180.46
R376 VGND.n880 VGND.n879 1180.46
R377 VGND.n875 VGND.n874 1180.46
R378 VGND.n870 VGND.n869 1180.46
R379 VGND.n865 VGND.n864 1180.46
R380 VGND.n860 VGND.n859 1180.46
R381 VGND.n855 VGND.n854 1180.46
R382 VGND.n850 VGND.n849 1180.46
R383 VGND.n845 VGND.n844 1180.46
R384 VGND.n2403 VGND.n2402 1180.46
R385 VGND.n2405 VGND.n2404 1180.46
R386 VGND.n2962 VGND.t1327 1180.08
R387 VGND.n1512 VGND.n1511 1169.57
R388 VGND.n3014 VGND.t59 1146.36
R389 VGND.n3016 VGND.t58 1112.64
R390 VGND.n3015 VGND.t2672 1112.64
R391 VGND.n2997 VGND 1055.35
R392 VGND.n1507 VGND.n1506 1052.29
R393 VGND.t2056 VGND.n961 1032.59
R394 VGND.t2359 VGND.n2579 988.926
R395 VGND.n2706 VGND.t1455 988.926
R396 VGND.n2705 VGND.t1130 988.926
R397 VGND.n2698 VGND.t2357 988.926
R398 VGND.n2697 VGND.t2346 988.926
R399 VGND.n2690 VGND.t1502 988.926
R400 VGND.n2689 VGND.t1060 988.926
R401 VGND.n2682 VGND.t2404 988.926
R402 VGND.n2681 VGND.t1498 988.926
R403 VGND.n2674 VGND.t1114 988.926
R404 VGND.n2673 VGND.t1102 988.926
R405 VGND.n2666 VGND.t2375 988.926
R406 VGND.n2665 VGND.t1485 988.926
R407 VGND.n2658 VGND.t1090 988.926
R408 VGND.n2657 VGND.t2389 988.926
R409 VGND.n233 VGND.t1717 988.926
R410 VGND.t109 VGND.n2720 988.926
R411 VGND.t2426 VGND.n2725 988.926
R412 VGND.t1982 VGND.n2730 988.926
R413 VGND.t523 VGND.n2735 988.926
R414 VGND.t330 VGND.n2740 988.926
R415 VGND.t529 VGND.n2745 988.926
R416 VGND.t772 VGND.n2750 988.926
R417 VGND.t1336 VGND.n2755 988.926
R418 VGND.t2665 VGND.n2760 988.926
R419 VGND.t2131 VGND.n2765 988.926
R420 VGND.t2509 VGND.n2770 988.926
R421 VGND.t2016 VGND.n2775 988.926
R422 VGND.t1947 VGND.n2780 988.926
R423 VGND.n2781 VGND.t653 988.926
R424 VGND.n2515 VGND.t1347 988.926
R425 VGND.n2514 VGND.t303 988.926
R426 VGND.n2509 VGND.t80 988.926
R427 VGND.t2406 VGND.n2434 988.926
R428 VGND.t2273 VGND.n2439 988.926
R429 VGND.t339 VGND.n2444 988.926
R430 VGND.t415 VGND.n2449 988.926
R431 VGND.t741 VGND.n2454 988.926
R432 VGND.t201 VGND.n2459 988.926
R433 VGND.t1545 VGND.n2464 988.926
R434 VGND.t2340 VGND.n2469 988.926
R435 VGND.t1996 VGND.n2474 988.926
R436 VGND.t2565 VGND.n2479 988.926
R437 VGND.t389 VGND.n2484 988.926
R438 VGND.t410 VGND.n2489 988.926
R439 VGND.n2832 VGND.t608 988.926
R440 VGND.t307 VGND.n371 988.926
R441 VGND.n372 VGND.t1693 988.926
R442 VGND.t1727 VGND.n2172 988.926
R443 VGND.n2173 VGND.t2051 988.926
R444 VGND.t1300 VGND.n2198 988.926
R445 VGND.n2199 VGND.t535 988.926
R446 VGND.t362 VGND.n2224 988.926
R447 VGND.n2225 VGND.t1342 988.926
R448 VGND.t2118 VGND.n2250 988.926
R449 VGND.n2251 VGND.t2037 988.926
R450 VGND.t175 VGND.n2281 988.926
R451 VGND.t2022 VGND.n2286 988.926
R452 VGND.t396 VGND.n2291 988.926
R453 VGND.n2292 VGND.t660 988.926
R454 VGND.t218 VGND.n1429 988.926
R455 VGND.n1430 VGND.t632 988.926
R456 VGND.t589 VGND.n2159 988.926
R457 VGND.n2160 VGND.t835 988.926
R458 VGND.t226 VGND.n2185 988.926
R459 VGND.n2186 VGND.t350 988.926
R460 VGND.t369 VGND.n2211 988.926
R461 VGND.n2212 VGND.t10 988.926
R462 VGND.t871 VGND.n2237 988.926
R463 VGND.n2238 VGND.t2261 988.926
R464 VGND.t97 VGND.n2263 988.926
R465 VGND.n2269 VGND.t1422 988.926
R466 VGND.n2268 VGND.t114 988.926
R467 VGND.t548 VGND.n2308 988.926
R468 VGND.n2309 VGND.t248 988.926
R469 VGND.t1961 VGND.n1443 988.926
R470 VGND.n1494 VGND.t2092 988.926
R471 VGND.n1493 VGND.t1698 988.926
R472 VGND.n1488 VGND.t1777 988.926
R473 VGND.n1483 VGND.t617 988.926
R474 VGND.n1478 VGND.t326 988.926
R475 VGND.n1473 VGND.t542 988.926
R476 VGND.n1468 VGND.t1581 988.926
R477 VGND.n1463 VGND.t1176 988.926
R478 VGND.n1458 VGND.t1540 988.926
R479 VGND.n1453 VGND.t561 988.926
R480 VGND.n1448 VGND.t1999 988.926
R481 VGND.n2137 VGND.t2559 988.926
R482 VGND.n2136 VGND.t19 988.926
R483 VGND.n2131 VGND.t403 988.926
R484 VGND.n1505 VGND.t1715 988.926
R485 VGND.t107 VGND.n626 988.926
R486 VGND.n627 VGND.t2423 988.926
R487 VGND.t1980 VGND.n1998 988.926
R488 VGND.n1999 VGND.t521 988.926
R489 VGND.t328 VGND.n2024 988.926
R490 VGND.n2025 VGND.t375 988.926
R491 VGND.t770 VGND.n2050 988.926
R492 VGND.n2051 VGND.t1334 988.926
R493 VGND.t2268 VGND.n2076 988.926
R494 VGND.n2077 VGND.t2129 988.926
R495 VGND.t2506 VGND.n2107 988.926
R496 VGND.t2014 VGND.n2112 988.926
R497 VGND.t1944 VGND.n2117 988.926
R498 VGND.n2118 VGND.t651 988.926
R499 VGND.t1975 VGND.n652 988.926
R500 VGND.n653 VGND.t309 988.926
R501 VGND.t1691 VGND.n1985 988.926
R502 VGND.n1986 VGND.t1729 988.926
R503 VGND.t2053 VGND.n2011 988.926
R504 VGND.n2012 VGND.t1302 988.926
R505 VGND.t537 VGND.n2037 988.926
R506 VGND.n2038 VGND.t1700 988.926
R507 VGND.t2100 VGND.n2063 988.926
R508 VGND.n2064 VGND.t2120 988.926
R509 VGND.t2039 VGND.n2089 988.926
R510 VGND.n2095 VGND.t177 988.926
R511 VGND.n2094 VGND.t2024 988.926
R512 VGND.t841 VGND.n2333 988.926
R513 VGND.n2334 VGND.t662 988.926
R514 VGND.n959 VGND.t220 988.926
R515 VGND.n954 VGND.t634 988.926
R516 VGND.n949 VGND.t587 988.926
R517 VGND.n944 VGND.t837 988.926
R518 VGND.n939 VGND.t228 988.926
R519 VGND.n934 VGND.t352 988.926
R520 VGND.n929 VGND.t371 988.926
R521 VGND.n924 VGND.t766 988.926
R522 VGND.n919 VGND.t873 988.926
R523 VGND.n914 VGND.t2263 988.926
R524 VGND.n909 VGND.t99 988.926
R525 VGND.n904 VGND.t1424 988.926
R526 VGND.n1963 VGND.t116 988.926
R527 VGND.n1962 VGND.t550 988.926
R528 VGND.n1957 VGND.t250 988.926
R529 VGND.t233 VGND.n1396 988.926
R530 VGND.t623 VGND.n1401 988.926
R531 VGND.n1402 VGND.t593 988.926
R532 VGND.t831 VGND.n1824 988.926
R533 VGND.n1825 VGND.t2079 988.926
R534 VGND.t348 VGND.n1850 988.926
R535 VGND.n1851 VGND.t2595 988.926
R536 VGND.t6 VGND.n1876 988.926
R537 VGND.n1877 VGND.t639 988.926
R538 VGND.t2259 VGND.n1902 988.926
R539 VGND.n1903 VGND.t95 988.926
R540 VGND.t1420 VGND.n1933 988.926
R541 VGND.t2138 VGND.n1938 988.926
R542 VGND.t212 VGND.n1943 988.926
R543 VGND.n1944 VGND.t246 988.926
R544 VGND.t1959 VGND.n1381 988.926
R545 VGND.n1382 VGND.t2090 988.926
R546 VGND.t76 VGND.n1811 988.926
R547 VGND.n1812 VGND.t1775 988.926
R548 VGND.t615 VGND.n1837 988.926
R549 VGND.n1838 VGND.t324 988.926
R550 VGND.t540 VGND.n1863 988.926
R551 VGND.n1864 VGND.t1703 988.926
R552 VGND.t1174 VGND.n1889 988.926
R553 VGND.n1890 VGND.t2124 988.926
R554 VGND.t559 VGND.n1915 988.926
R555 VGND.n1921 VGND.t2493 988.926
R556 VGND.n1920 VGND.t2557 988.926
R557 VGND.t12 VGND.n2358 988.926
R558 VGND.n2359 VGND.t401 988.926
R559 VGND.t811 VGND.n1313 988.926
R560 VGND.n1364 VGND.t1172 988.926
R561 VGND.n1363 VGND.t579 988.926
R562 VGND.n1358 VGND.t1734 988.926
R563 VGND.n1353 VGND.t1569 988.926
R564 VGND.n1348 VGND.t335 988.926
R565 VGND.n1343 VGND.t2588 988.926
R566 VGND.n1338 VGND.t1404 988.926
R567 VGND.n1333 VGND.t628 988.926
R568 VGND.n1328 VGND.t732 988.926
R569 VGND.n1323 VGND.t2245 988.926
R570 VGND.n1318 VGND.t1426 988.926
R571 VGND.n1789 VGND.t154 988.926
R572 VGND.n1788 VGND.t1942 988.926
R573 VGND.n1783 VGND.t381 988.926
R574 VGND.t606 VGND.n1518 988.926
R575 VGND.t305 VGND.n1523 988.926
R576 VGND.n1524 VGND.t1695 988.926
R577 VGND.t1725 VGND.n1650 988.926
R578 VGND.n1651 VGND.t527 988.926
R579 VGND.t1298 VGND.n1676 988.926
R580 VGND.n1677 VGND.t533 988.926
R581 VGND.t360 VGND.n1702 988.926
R582 VGND.n1703 VGND.t1340 988.926
R583 VGND.t2669 VGND.n1728 988.926
R584 VGND.n1729 VGND.t2035 988.926
R585 VGND.t173 VGND.n1759 988.926
R586 VGND.t2020 VGND.n1764 988.926
R587 VGND.t394 VGND.n1769 988.926
R588 VGND.n1770 VGND.t658 988.926
R589 VGND.t809 VGND.n1538 988.926
R590 VGND.n1539 VGND.t1170 988.926
R591 VGND.t581 VGND.n1637 988.926
R592 VGND.n1638 VGND.t1732 988.926
R593 VGND.t1567 VGND.n1663 988.926
R594 VGND.n1664 VGND.t333 988.926
R595 VGND.t2586 VGND.n1689 988.926
R596 VGND.n1690 VGND.t1402 988.926
R597 VGND.t438 VGND.n1715 988.926
R598 VGND.n1716 VGND.t730 988.926
R599 VGND.t193 VGND.n1741 988.926
R600 VGND.n1747 VGND.t1613 988.926
R601 VGND.n1746 VGND.t152 988.926
R602 VGND.t1940 VGND.n2383 988.926
R603 VGND.n2384 VGND.t379 988.926
R604 VGND.n1296 VGND.t1345 988.926
R605 VGND.t301 VGND.n1551 988.926
R606 VGND.t83 VGND.n1556 988.926
R607 VGND.t1781 VGND.n1561 988.926
R608 VGND.t2271 VGND.n1566 988.926
R609 VGND.t337 VGND.n1571 988.926
R610 VGND.t413 VGND.n1576 988.926
R611 VGND.t739 VGND.n1581 988.926
R612 VGND.t199 VGND.n1586 988.926
R613 VGND.t1542 VGND.n1591 988.926
R614 VGND.t2338 VGND.n1596 988.926
R615 VGND.t2001 VGND.n1601 988.926
R616 VGND.n1615 VGND.t2563 988.926
R617 VGND.n1614 VGND.t21 988.926
R618 VGND.n1609 VGND.t407 988.926
R619 VGND.t235 VGND.n835 988.926
R620 VGND.t625 VGND.n840 988.926
R621 VGND.n891 VGND.t591 988.926
R622 VGND.n890 VGND.t833 988.926
R623 VGND.n885 VGND.t2081 988.926
R624 VGND.n880 VGND.t346 988.926
R625 VGND.n875 VGND.t2593 988.926
R626 VGND.n870 VGND.t4 988.926
R627 VGND.n865 VGND.t637 988.926
R628 VGND.n860 VGND.t736 988.926
R629 VGND.n855 VGND.t93 988.926
R630 VGND.n850 VGND.t1418 988.926
R631 VGND.n845 VGND.t159 988.926
R632 VGND.t546 VGND.n2403 988.926
R633 VGND.n2404 VGND.t244 988.926
R634 VGND.n1290 VGND.t1481 988.926
R635 VGND.t1096 VGND.n720 988.926
R636 VGND.t1074 VGND.n725 988.926
R637 VGND.t1476 VGND.n730 988.926
R638 VGND.t1465 VGND.n735 988.926
R639 VGND.t1446 VGND.n740 988.926
R640 VGND.t2369 VGND.n745 988.926
R641 VGND.t2348 VGND.n750 988.926
R642 VGND.t1139 VGND.n755 988.926
R643 VGND.t1062 VGND.n760 988.926
R644 VGND.t1049 VGND.n765 988.926
R645 VGND.t1500 VGND.n770 988.926
R646 VGND.t1122 VGND.n775 988.926
R647 VGND.t2398 VGND.n780 988.926
R648 VGND.n781 VGND.t1509 988.926
R649 VGND.n1509 VGND.n579 934.784
R650 VGND.n2908 VGND 927.203
R651 VGND.n2911 VGND 927.203
R652 VGND.n962 VGND 918.774
R653 VGND.n113 VGND 910.346
R654 VGND.n2875 VGND 910.346
R655 VGND.n3009 VGND.t1316 909.365
R656 VGND.n2834 VGND.n177 900
R657 VGND.n2579 VGND.t2094 852.769
R658 VGND.n2706 VGND.t238 852.769
R659 VGND.t1608 VGND.n2705 852.769
R660 VGND.n2698 VGND.t1400 852.769
R661 VGND.t1711 VGND.n2697 852.769
R662 VGND.n2690 VGND.t601 852.769
R663 VGND.t214 VGND.n2689 852.769
R664 VGND.n2682 VGND.t667 852.769
R665 VGND.t484 VGND.n2681 852.769
R666 VGND.n2674 VGND.t848 852.769
R667 VGND.t50 VGND.n2673 852.769
R668 VGND.n2666 VGND.t467 852.769
R669 VGND.t1951 VGND.n2665 852.769
R670 VGND.n2658 VGND.t1632 852.769
R671 VGND.t1443 VGND.n2657 852.769
R672 VGND.t573 VGND.n33 852.769
R673 VGND.n233 VGND.t2671 852.769
R674 VGND.n2720 VGND.t0 852.769
R675 VGND.n2725 VGND.t507 852.769
R676 VGND.n2730 VGND.t1206 852.769
R677 VGND.n2735 VGND.t1605 852.769
R678 VGND.n2740 VGND.t278 852.769
R679 VGND.n2745 VGND.t2065 852.769
R680 VGND.n2750 VGND.t1607 852.769
R681 VGND.n2755 VGND.t1156 852.769
R682 VGND.n2760 VGND.t2483 852.769
R683 VGND.n2765 VGND.t57 852.769
R684 VGND.n2770 VGND.t315 852.769
R685 VGND.n2775 VGND.t274 852.769
R686 VGND.n2780 VGND.t2663 852.769
R687 VGND.n2781 VGND.t2099 852.769
R688 VGND.n3000 VGND.t1291 852.769
R689 VGND.n2515 VGND.t2599 852.769
R690 VGND.t1949 VGND.n2514 852.769
R691 VGND.t1293 VGND.n2509 852.769
R692 VGND.n2434 VGND.t1602 852.769
R693 VGND.n2439 VGND.t583 852.769
R694 VGND.n2444 VGND.t519 852.769
R695 VGND.n2449 VGND.t747 852.769
R696 VGND.n2454 VGND.t516 852.769
R697 VGND.n2459 VGND.t222 852.769
R698 VGND.n2464 VGND.t850 852.769
R699 VGND.n2469 VGND.t665 852.769
R700 VGND.n2474 VGND.t2285 852.769
R701 VGND.n2479 VGND.t1408 852.769
R702 VGND.n2484 VGND.t55 852.769
R703 VGND.n2489 VGND.t602 852.769
R704 VGND.n2490 VGND.t2429 852.769
R705 VGND.t2410 VGND.n2832 852.769
R706 VGND.n371 VGND.t275 852.769
R707 VGND.n372 VGND.t366 852.769
R708 VGND.n2172 VGND.t1304 852.769
R709 VGND.n2173 VGND.t224 852.769
R710 VGND.n2198 VGND.t2598 852.769
R711 VGND.n2199 VGND.t277 852.769
R712 VGND.n2224 VGND.t2602 852.769
R713 VGND.n2225 VGND.t1401 852.769
R714 VGND.n2250 VGND.t317 852.769
R715 VGND.n2251 VGND.t1392 852.769
R716 VGND.n2281 VGND.t1196 852.769
R717 VGND.n2286 VGND.t18 852.769
R718 VGND.n2291 VGND.t1142 852.769
R719 VGND.n2292 VGND.t2105 852.769
R720 VGND.n2429 VGND.t468 852.769
R721 VGND.n1429 VGND.t1295 852.769
R722 VGND.n1430 VGND.t440 852.769
R723 VGND.n2159 VGND.t758 852.769
R724 VGND.n2160 VGND.t2284 852.769
R725 VGND.n2185 VGND.t782 852.769
R726 VGND.n2186 VGND.t1972 852.769
R727 VGND.n2211 VGND.t1143 852.769
R728 VGND.n2212 VGND.t1616 852.769
R729 VGND.n2237 VGND.t738 852.769
R730 VGND.n2238 VGND.t2277 852.769
R731 VGND.n2263 VGND.t279 852.769
R732 VGND.n2269 VGND.t603 852.769
R733 VGND.t1986 VGND.n2268 852.769
R734 VGND.n2308 VGND.t1719 852.769
R735 VGND.n2309 VGND.t574 852.769
R736 VGND.t1281 VGND.n261 852.769
R737 VGND.n1443 VGND.t1149 852.769
R738 VGND.n1494 VGND.t614 852.769
R739 VGND.t2066 VGND.n1493 852.769
R740 VGND.t207 VGND.n1488 852.769
R741 VGND.t2003 VGND.n1483 852.769
R742 VGND.t16 VGND.n1478 852.769
R743 VGND.t849 VGND.n1473 852.769
R744 VGND.t2089 VGND.n1468 852.769
R745 VGND.t209 VGND.n1463 852.769
R746 VGND.t2027 VGND.n1458 852.769
R747 VGND.t1585 VGND.n1453 852.769
R748 VGND.t1712 VGND.n1448 852.769
R749 VGND.n2137 VGND.t206 852.769
R750 VGND.t288 VGND.n2136 852.769
R751 VGND.t2287 VGND.n2131 852.769
R752 VGND.t515 VGND.n262 852.769
R753 VGND.t14 VGND.n1505 852.769
R754 VGND.n626 VGND.t54 852.769
R755 VGND.n627 VGND.t555 852.769
R756 VGND.n1998 VGND.t745 852.769
R757 VGND.n1999 VGND.t387 852.769
R758 VGND.n2024 VGND.t1203 852.769
R759 VGND.n2025 VGND.t1399 852.769
R760 VGND.n2050 VGND.t253 852.769
R761 VGND.n2051 VGND.t1953 852.769
R762 VGND.n2076 VGND.t845 852.769
R763 VGND.n2077 VGND.t1351 852.769
R764 VGND.n2107 VGND.t2060 852.769
R765 VGND.n2112 VGND.t2601 852.769
R766 VGND.n2117 VGND.t1950 852.769
R767 VGND.n2118 VGND.t1409 852.769
R768 VGND.t1333 VGND.n263 852.769
R769 VGND.n652 VGND.t1141 852.769
R770 VGND.n653 VGND.t499 852.769
R771 VGND.n1985 VGND.t1306 852.769
R772 VGND.n1986 VGND.t868 852.769
R773 VGND.n2011 VGND.t1394 852.769
R774 VGND.n2012 VGND.t862 852.769
R775 VGND.n2037 VGND.t469 852.769
R776 VGND.n2038 VGND.t1326 852.769
R777 VGND.n2063 VGND.t597 852.769
R778 VGND.n2064 VGND.t2286 852.769
R779 VGND.n2089 VGND.t223 852.769
R780 VGND.n2095 VGND.t2067 852.769
R781 VGND.t1752 VGND.n2094 852.769
R782 VGND.n2333 VGND.t1630 852.769
R783 VGND.n2334 VGND.t1958 852.769
R784 VGND.t1352 VGND.n264 852.769
R785 VGND.t276 VGND.n959 852.769
R786 VGND.t1008 VGND.n954 852.769
R787 VGND.t120 VGND.n949 852.769
R788 VGND.t1389 VGND.n944 852.769
R789 VGND.t256 VGND.n939 852.769
R790 VGND.t1344 VGND.n934 852.769
R791 VGND.t2609 VGND.n929 852.769
R792 VGND.t764 VGND.n924 852.769
R793 VGND.t2484 VGND.n919 852.769
R794 VGND.t553 VGND.n914 852.769
R795 VGND.t2688 VGND.n909 852.769
R796 VGND.t1615 VGND.n904 852.769
R797 VGND.n1963 VGND.t1973 852.769
R798 VGND.t757 VGND.n1962 852.769
R799 VGND.t1192 VGND.n1957 852.769
R800 VGND.t1391 VGND.n265 852.769
R801 VGND.n1396 VGND.t670 852.769
R802 VGND.n1401 VGND.t1289 852.769
R803 VGND.n1402 VGND.t1332 852.769
R804 VGND.n1824 VGND.t2675 852.769
R805 VGND.n1825 VGND.t1201 852.769
R806 VGND.n1850 VGND.t847 852.769
R807 VGND.n1851 VGND.t208 852.769
R808 VGND.n1876 VGND.t1974 852.769
R809 VGND.n1877 VGND.t1148 852.769
R810 VGND.n1902 VGND.t2244 852.769
R811 VGND.n1903 VGND.t2676 852.769
R812 VGND.n1933 VGND.t1682 852.769
R813 VGND.n1938 VGND.t666 852.769
R814 VGND.n1943 VGND.t2104 852.769
R815 VGND.n1944 VGND.t1390 852.769
R816 VGND.t1655 VGND.n266 852.769
R817 VGND.n1381 VGND.t2088 852.769
R818 VGND.n1382 VGND.t1396 852.769
R819 VGND.n1811 VGND.t508 852.769
R820 VGND.n1812 VGND.t1158 852.769
R821 VGND.n1837 VGND.t1722 852.769
R822 VGND.n1838 VGND.t1195 852.769
R823 VGND.n1863 VGND.t1284 852.769
R824 VGND.n1864 VGND.t2487 852.769
R825 VGND.n1889 VGND.t2064 852.769
R826 VGND.n1890 VGND.t1710 852.769
R827 VGND.n1915 VGND.t1205 852.769
R828 VGND.n1921 VGND.t1720 852.769
R829 VGND.t875 VGND.n1920 852.769
R830 VGND.n2358 VGND.t505 852.769
R831 VGND.n2359 VGND.t52 852.769
R832 VGND.t2600 VGND.n267 852.769
R833 VGND.n1313 VGND.t2290 852.769
R834 VGND.n1364 VGND.t259 852.769
R835 VGND.t2603 VGND.n1363 852.769
R836 VGND.t49 VGND.n1358 852.769
R837 VGND.t53 VGND.n1353 852.769
R838 VGND.t1198 VGND.n1348 852.769
R839 VGND.t839 VGND.n1343 852.769
R840 VGND.t280 VGND.n1338 852.769
R841 VGND.t509 VGND.n1333 852.769
R842 VGND.t2608 VGND.n1328 852.769
R843 VGND.t1157 VGND.n1323 852.769
R844 VGND.t385 VGND.n1318 852.769
R845 VGND.n1789 VGND.t775 852.769
R846 VGND.t1204 VGND.n1788 852.769
R847 VGND.t599 VGND.n1783 852.769
R848 VGND.t258 VGND.n268 852.769
R849 VGND.n1518 VGND.t2677 852.769
R850 VGND.n1523 VGND.t386 852.769
R851 VGND.n1524 VGND.t1197 852.769
R852 VGND.n1650 VGND.t746 852.769
R853 VGND.n1651 VGND.t215 852.769
R854 VGND.n1676 VGND.t1971 852.769
R855 VGND.n1677 VGND.t1407 852.769
R856 VGND.n1702 VGND.t668 852.769
R857 VGND.n1703 VGND.t765 852.769
R858 VGND.n1728 VGND.t2597 852.769
R859 VGND.n1729 VGND.t195 852.769
R860 VGND.n1759 VGND.t1631 852.769
R861 VGND.n1764 VGND.t1147 852.769
R862 VGND.n1769 VGND.t763 852.769
R863 VGND.n1770 VGND.t196 852.769
R864 VGND.t1952 VGND.n269 852.769
R865 VGND.n1538 VGND.t572 852.769
R866 VGND.n1539 VGND.t2486 852.769
R867 VGND.n1637 VGND.t2111 852.769
R868 VGND.n1638 VGND.t1 852.769
R869 VGND.n1663 VGND.t384 852.769
R870 VGND.n1664 VGND.t669 852.769
R871 VGND.n1689 VGND.t2485 852.769
R872 VGND.n1690 VGND.t1606 852.769
R873 VGND.n1715 VGND.t1290 852.769
R874 VGND.n1716 VGND.t596 852.769
R875 VGND.n1741 VGND.t554 852.769
R876 VGND.n1747 VGND.t254 852.769
R877 VGND.t851 VGND.n1746 852.769
R878 VGND.n2383 VGND.t744 852.769
R879 VGND.n2384 VGND.t281 852.769
R880 VGND.t421 VGND.n270 852.769
R881 VGND.n1296 VGND.t1305 852.769
R882 VGND.n1551 VGND.t600 852.769
R883 VGND.n1556 VGND.t1202 852.769
R884 VGND.n1561 VGND.t2278 852.769
R885 VGND.n1566 VGND.t2482 852.769
R886 VGND.n1571 VGND.t846 852.769
R887 VGND.n1576 VGND.t240 852.769
R888 VGND.n1581 VGND.t1288 852.769
R889 VGND.n1586 VGND.t118 852.769
R890 VGND.n1591 VGND.t1395 852.769
R891 VGND.n1596 VGND.t1617 852.769
R892 VGND.n1601 VGND.t197 852.769
R893 VGND.n1615 VGND.t506 852.769
R894 VGND.t1010 VGND.n1614 852.769
R895 VGND.t74 VGND.n1609 852.769
R896 VGND.t1654 VGND.n271 852.769
R897 VGND.n835 VGND.t1398 852.769
R898 VGND.n840 VGND.t1522 852.769
R899 VGND.n891 VGND.t15 852.769
R900 VGND.t1023 VGND.n890 852.769
R901 VGND.t316 VGND.n885 852.769
R902 VGND.t56 VGND.n880 852.769
R903 VGND.t17 VGND.n875 852.769
R904 VGND.t1331 VGND.n870 852.769
R905 VGND.t760 VGND.n865 852.769
R906 VGND.t51 VGND.n860 852.769
R907 VGND.t1723 VGND.n855 852.769
R908 VGND.t1286 VGND.n850 852.769
R909 VGND.t2063 VGND.n845 852.769
R910 VGND.n2403 VGND.t75 852.769
R911 VGND.n2404 VGND.t598 852.769
R912 VGND.t314 VGND.n272 852.769
R913 VGND.t1009 VGND.n1290 852.769
R914 VGND.n720 VGND.t239 852.769
R915 VGND.n725 VGND.t1287 852.769
R916 VGND.n730 VGND.t743 852.769
R917 VGND.n735 VGND.t1194 852.769
R918 VGND.n740 VGND.t2279 852.769
R919 VGND.n745 VGND.t161 852.769
R920 VGND.n750 VGND.t420 852.769
R921 VGND.n755 VGND.t1393 852.769
R922 VGND.n760 VGND.t2411 852.769
R923 VGND.n765 VGND.t203 852.769
R924 VGND.n770 VGND.t928 852.769
R925 VGND.n775 VGND.t1397 852.769
R926 VGND.n780 VGND.t1193 852.769
R927 VGND.n781 VGND.t759 852.769
R928 VGND.n2414 VGND.t1285 852.769
R929 VGND.n1508 VGND 851.341
R930 VGND.n2842 VGND.t1072 809.773
R931 VGND.n2841 VGND.t1831 809.773
R932 VGND.t1906 VGND.n114 809.773
R933 VGND.n2833 VGND.t1813 809.773
R934 VGND.t1855 VGND.n177 809.773
R935 VGND.t1927 VGND.n635 809.773
R936 VGND.t1807 VGND.n580 809.773
R937 VGND.n960 VGND.t1849 809.773
R938 VGND.t1861 VGND.n579 809.773
R939 VGND.n1512 VGND.t1885 809.773
R940 VGND.t1816 VGND.n1513 809.773
R941 VGND.n1294 VGND.t1888 809.773
R942 VGND.t1918 VGND.n1295 809.773
R943 VGND.n1293 VGND.t1858 809.773
R944 VGND.n1291 VGND.t2384 809.773
R945 VGND.t2499 VGND.t31 708.047
R946 VGND.t31 VGND.t33 708.047
R947 VGND.t33 VGND.t23 708.047
R948 VGND.t23 VGND.t1430 708.047
R949 VGND.t1430 VGND.t1785 708.047
R950 VGND.t1785 VGND.t1936 708.047
R951 VGND.t1936 VGND.t1934 708.047
R952 VGND.t2296 VGND.t58 708.047
R953 VGND.t135 VGND.t137 708.047
R954 VGND.t137 VGND.t1560 708.047
R955 VGND.t1560 VGND.t1574 708.047
R956 VGND.t1574 VGND.t1037 708.047
R957 VGND.t1037 VGND.t312 708.047
R958 VGND.t312 VGND.t1633 708.047
R959 VGND.t1633 VGND.t216 708.047
R960 VGND.t2490 VGND.t1576 708.047
R961 VGND.t1576 VGND.t1523 708.047
R962 VGND.t1523 VGND.t1565 708.047
R963 VGND.t1565 VGND.t1628 708.047
R964 VGND.t1628 VGND.t1624 708.047
R965 VGND.t1624 VGND.t1618 708.047
R966 VGND.t1618 VGND.t1620 708.047
R967 VGND.t2293 VGND.t59 708.047
R968 VGND.t1529 VGND.t1563 708.047
R969 VGND.t1578 VGND.t1529 708.047
R970 VGND.t35 VGND.t1578 708.047
R971 VGND.t1432 VGND.t35 708.047
R972 VGND.t1787 VGND.t1432 708.047
R973 VGND.t1429 VGND.t1787 708.047
R974 VGND.t1784 VGND.t1429 708.047
R975 VGND.t1527 VGND.t1533 708.047
R976 VGND.t1533 VGND.t2497 708.047
R977 VGND.t2497 VGND.t140 708.047
R978 VGND.t140 VGND.t1183 708.047
R979 VGND.t1183 VGND.t2103 708.047
R980 VGND.t2103 VGND.t1024 708.047
R981 VGND.t1024 VGND.t1319 708.047
R982 VGND.t148 VGND.t25 708.047
R983 VGND.t25 VGND.t133 708.047
R984 VGND.t133 VGND.t1525 708.047
R985 VGND.t1525 VGND.t1626 708.047
R986 VGND.t1626 VGND.t1622 708.047
R987 VGND.t1622 VGND.t1627 708.047
R988 VGND.t1627 VGND.t1623 708.047
R989 VGND.n2995 VGND.n2994 708.047
R990 VGND.t2084 VGND.t1969 691.188
R991 VGND.t1705 VGND.t2673 691.188
R992 VGND.n2838 VGND.t544 685.545
R993 VGND.n3018 VGND.t544 685.545
R994 VGND.n2841 VGND.n2840 660.87
R995 VGND.t2304 VGND.t1016 657.471
R996 VGND.t2313 VGND.t1014 657.471
R997 VGND.t122 VGND.t1012 657.471
R998 VGND.t1355 VGND.t817 657.471
R999 VGND.t146 VGND.t1531 657.471
R1000 VGND.t1535 VGND.t1317 657.471
R1001 VGND.t131 VGND.t1313 657.471
R1002 VGND.t1557 VGND.t1307 657.471
R1003 VGND.t817 VGND.t819 654.197
R1004 VGND.t1531 VGND.t142 654.197
R1005 VGND.n962 VGND 640.614
R1006 VGND VGND.n113 640.614
R1007 VGND VGND.n2875 640.614
R1008 VGND VGND.n2908 640.614
R1009 VGND.n2911 VGND 632.184
R1010 VGND.t1461 VGND.t2361 630.62
R1011 VGND.t1084 VGND.t1457 630.62
R1012 VGND.t1076 VGND.t1071 630.62
R1013 VGND.t1520 VGND.t1056 630.62
R1014 VGND.t2354 VGND.t1453 630.62
R1015 VGND.t1058 VGND.t1132 630.62
R1016 VGND.t1118 VGND.t2356 630.62
R1017 VGND.t1508 VGND.t2350 630.62
R1018 VGND.t1504 VGND.t1120 630.62
R1019 VGND.t1059 VGND.t1134 630.62
R1020 VGND.t1039 VGND.t1506 630.62
R1021 VGND.t1496 VGND.t2391 630.62
R1022 VGND.t1116 VGND.t1111 630.62
R1023 VGND.t2395 VGND.t1104 630.62
R1024 VGND.t1088 VGND.t2372 630.62
R1025 VGND.t1489 VGND.t1108 630.62
R1026 VGND.t814 VGND.t1243 630.62
R1027 VGND.t1754 VGND.t621 630.62
R1028 VGND.t595 VGND.t1251 630.62
R1029 VGND.t1979 VGND.t1249 630.62
R1030 VGND.t2077 VGND.t1241 630.62
R1031 VGND.t342 VGND.t1033 630.62
R1032 VGND.t2591 VGND.t1031 630.62
R1033 VGND.t2 VGND.t1760 630.62
R1034 VGND.t869 VGND.t1758 630.62
R1035 VGND.t735 VGND.t1035 630.62
R1036 VGND.t2343 VGND.t1247 630.62
R1037 VGND.t1417 VGND.t1245 630.62
R1038 VGND.t157 VGND.t1029 630.62
R1039 VGND.t211 VGND.t1027 630.62
R1040 VGND.t650 VGND.t1025 630.62
R1041 VGND.t1756 VGND.t1497 630.62
R1042 VGND.t605 VGND.t268 630.62
R1043 VGND.t2555 VGND.t112 630.62
R1044 VGND.t1322 VGND.t563 630.62
R1045 VGND.t1780 VGND.t1320 630.62
R1046 VGND.t526 VGND.t2242 630.62
R1047 VGND.t345 VGND.t2551 630.62
R1048 VGND.t532 VGND.t2549 630.62
R1049 VGND.t359 VGND.t2240 630.62
R1050 VGND.t1339 VGND.t2238 630.62
R1051 VGND.t2122 VGND.t2553 630.62
R1052 VGND.t2250 VGND.t272 630.62
R1053 VGND.t179 VGND.t270 630.62
R1054 VGND.t2019 VGND.t2547 630.62
R1055 VGND.t843 VGND.t2545 630.62
R1056 VGND.t406 VGND.t1324 630.62
R1057 VGND.t1043 VGND.t2236 630.62
R1058 VGND.t854 VGND.t232 630.62
R1059 VGND.t627 VGND.t1159 630.62
R1060 VGND.t585 VGND.t282 630.62
R1061 VGND.t860 VGND.t1985 630.62
R1062 VGND.t2083 VGND.t852 630.62
R1063 VGND.t2072 VGND.t344 630.62
R1064 VGND.t367 VGND.t2070 630.62
R1065 VGND.t1165 VGND.t8 630.62
R1066 VGND.t641 VGND.t1163 630.62
R1067 VGND.t2074 VGND.t2266 630.62
R1068 VGND.t2345 VGND.t858 630.62
R1069 VGND.t856 VGND.t1932 630.62
R1070 VGND.t2140 VGND.t2068 630.62
R1071 VGND.t517 VGND.t286 630.62
R1072 VGND.t656 VGND.t284 630.62
R1073 VGND.t1161 VGND.t1518 630.62
R1074 VGND.t204 VGND.t478 630.62
R1075 VGND.t2109 VGND.t2033 630.62
R1076 VGND.t2543 VGND.t575 630.62
R1077 VGND.t829 VGND.t2541 630.62
R1078 VGND.t476 VGND.t2043 630.62
R1079 VGND.t322 VGND.t2029 630.62
R1080 VGND.t570 VGND.t2584 630.62
R1081 VGND.t612 VGND.t474 630.62
R1082 VGND.t472 VGND.t436 630.62
R1083 VGND.t728 VGND.t2031 630.62
R1084 VGND.t2539 VGND.t557 630.62
R1085 VGND.t1611 VGND.t2537 630.62
R1086 VGND.t568 VGND.t150 630.62
R1087 VGND.t566 VGND.t1146 630.62
R1088 VGND.t242 VGND.t564 630.62
R1089 VGND.t470 VGND.t1452 630.62
R1090 VGND.t1714 VGND.t1650 630.62
R1091 VGND.t106 VGND.t2255 630.62
R1092 VGND.t1929 VGND.t2425 630.62
R1093 VGND.t1600 VGND.t1774 630.62
R1094 VGND.t1648 VGND.t520 630.62
R1095 VGND.t2251 VGND.t356 630.62
R1096 VGND.t1642 VGND.t374 630.62
R1097 VGND.t1646 VGND.t769 630.62
R1098 VGND.t1644 VGND.t762 630.62
R1099 VGND.t2253 VGND.t2667 630.62
R1100 VGND.t1598 VGND.t2248 630.62
R1101 VGND.t1652 VGND.t171 630.62
R1102 VGND.t1640 VGND.t2013 630.62
R1103 VGND.t1638 VGND.t392 630.62
R1104 VGND.t1636 VGND.t400 630.62
R1105 VGND.t2257 VGND.t2382 630.62
R1106 VGND.t2182 VGND.t813 630.62
R1107 VGND.t620 VGND.t418 630.62
R1108 VGND.t584 VGND.t2326 630.62
R1109 VGND.t2324 VGND.t1978 630.62
R1110 VGND.t2076 VGND.t2180 630.62
R1111 VGND.t2336 VGND.t341 630.62
R1112 VGND.t2590 VGND.t2334 630.62
R1113 VGND.t2178 VGND.t1406 630.62
R1114 VGND.t630 VGND.t2176 630.62
R1115 VGND.t497 VGND.t734 630.62
R1116 VGND.t2342 VGND.t2322 630.62
R1117 VGND.t2320 VGND.t1428 630.62
R1118 VGND.t156 VGND.t2332 630.62
R1119 VGND.t210 VGND.t2330 630.62
R1120 VGND.t252 VGND.t2328 630.62
R1121 VGND.t2174 VGND.t1495 630.62
R1122 VGND.t237 VGND.t1772 630.62
R1123 VGND.t631 VGND.t1762 630.62
R1124 VGND.t1592 VGND.t2422 630.62
R1125 VGND.t1724 VGND.t1590 630.62
R1126 VGND.t1770 VGND.t225 630.62
R1127 VGND.t332 VGND.t646 630.62
R1128 VGND.t644 VGND.t368 630.62
R1129 VGND.t9 VGND.t1768 630.62
R1130 VGND.t1766 VGND.t870 630.62
R1131 VGND.t2267 VGND.t648 630.62
R1132 VGND.t1588 VGND.t192 630.62
R1133 VGND.t1933 VGND.t1586 630.62
R1134 VGND.t642 VGND.t113 630.62
R1135 VGND.t1596 VGND.t518 630.62
R1136 VGND.t657 VGND.t1594 630.62
R1137 VGND.t1764 VGND.t1521 630.62
R1138 VGND.t260 VGND.t205 630.62
R1139 VGND.t2061 VGND.t2110 630.62
R1140 VGND.t2275 VGND.t578 630.62
R1141 VGND.t266 VGND.t830 630.62
R1142 VGND.t1993 VGND.t2044 630.62
R1143 VGND.t1152 VGND.t323 630.62
R1144 VGND.t1150 VGND.t2585 630.62
R1145 VGND.t1991 VGND.t613 630.62
R1146 VGND.t1989 VGND.t437 630.62
R1147 VGND.t1154 VGND.t729 630.62
R1148 VGND.t264 VGND.t558 630.62
R1149 VGND.t262 VGND.t1612 630.62
R1150 VGND.t780 VGND.t151 630.62
R1151 VGND.t778 VGND.t1939 630.62
R1152 VGND.t776 VGND.t243 630.62
R1153 VGND.t1987 VGND.t1454 630.62
R1154 VGND.t1349 VGND.t1213 630.62
R1155 VGND.t2108 VGND.t89 630.62
R1156 VGND.t577 VGND.t1555 630.62
R1157 VGND.t1553 VGND.t828 630.62
R1158 VGND.t2041 VGND.t1211 630.62
R1159 VGND.t85 VGND.t320 630.62
R1160 VGND.t2583 VGND.t2010 630.62
R1161 VGND.t1209 VGND.t399 630.62
R1162 VGND.t435 VGND.t1207 630.62
R1163 VGND.t87 VGND.t727 630.62
R1164 VGND.t556 VGND.t1551 630.62
R1165 VGND.t1549 VGND.t1610 630.62
R1166 VGND.t2568 VGND.t2008 630.62
R1167 VGND.t1145 VGND.t2006 630.62
R1168 VGND.t383 VGND.t2004 630.62
R1169 VGND.t91 VGND.t1445 630.62
R1170 VGND.t1713 VGND.t491 630.62
R1171 VGND.t2106 VGND.t2579 630.62
R1172 VGND.t64 VGND.t2428 630.62
R1173 VGND.t1731 VGND.t62 630.62
R1174 VGND.t489 VGND.t840 630.62
R1175 VGND.t355 VGND.t2575 630.62
R1176 VGND.t2573 VGND.t373 630.62
R1177 VGND.t768 VGND.t487 630.62
R1178 VGND.t485 VGND.t761 630.62
R1179 VGND.t2664 VGND.t2577 630.62
R1180 VGND.t495 VGND.t2247 630.62
R1181 VGND.t2508 VGND.t493 630.62
R1182 VGND.t2571 VGND.t2012 630.62
R1183 VGND.t2569 VGND.t1946 630.62
R1184 VGND.t664 VGND.t482 630.62
R1185 VGND.t2581 VGND.t2377 630.62
R1186 VGND.t1964 VGND.t1738 630.62
R1187 VGND.t300 VGND.t2165 630.62
R1188 VGND.t1746 VGND.t79 630.62
R1189 VGND.t1744 VGND.t2409 630.62
R1190 VGND.t1736 VGND.t2270 630.62
R1191 VGND.t2161 VGND.t1297 630.62
R1192 VGND.t2159 VGND.t412 630.62
R1193 VGND.t2171 VGND.t1584 630.62
R1194 VGND.t2169 VGND.t198 630.62
R1195 VGND.t2163 VGND.t1547 630.62
R1196 VGND.t1742 VGND.t2134 630.62
R1197 VGND.t1740 VGND.t1998 630.62
R1198 VGND.t2157 VGND.t2562 630.62
R1199 VGND.t1750 VGND.t391 630.62
R1200 VGND.t1748 VGND.t378 630.62
R1201 VGND.t2167 VGND.t1101 630.62
R1202 VGND.t231 VGND.t430 630.62
R1203 VGND.t622 VGND.t2420 630.62
R1204 VGND.t586 VGND.t721 630.62
R1205 VGND.t719 VGND.t1984 630.62
R1206 VGND.t2078 VGND.t428 630.62
R1207 VGND.t2416 VGND.t343 630.62
R1208 VGND.t2592 VGND.t2414 630.62
R1209 VGND.t426 VGND.t3 630.62
R1210 VGND.t636 VGND.t424 630.62
R1211 VGND.t2418 VGND.t2265 630.62
R1212 VGND.t2344 VGND.t717 630.62
R1213 VGND.t432 VGND.t1931 630.62
R1214 VGND.t158 VGND.t2412 630.62
R1215 VGND.t552 VGND.t725 630.62
R1216 VGND.t655 VGND.t723 630.62
R1217 VGND.t422 VGND.t1515 630.62
R1218 VGND.t2045 VGND.t1963 630.62
R1219 VGND.t299 VGND.t186 630.62
R1220 VGND.t1435 VGND.t82 630.62
R1221 VGND.t2408 VGND.t1433 630.62
R1222 VGND.t104 VGND.t619 630.62
R1223 VGND.t1296 VGND.t182 630.62
R1224 VGND.t180 VGND.t1721 630.62
R1225 VGND.t1583 VGND.t102 630.62
R1226 VGND.t190 VGND.t1178 630.62
R1227 VGND.t1544 VGND.t184 630.62
R1228 VGND.t2049 VGND.t2133 630.62
R1229 VGND.t1995 VGND.t2047 630.62
R1230 VGND.t1441 VGND.t2561 630.62
R1231 VGND.t1439 VGND.t388 630.62
R1232 VGND.t377 VGND.t1437 630.62
R1233 VGND.t188 VGND.t1098 630.62
R1234 VGND.t604 VGND.t43 630.62
R1235 VGND.t2151 VGND.t111 630.62
R1236 VGND.t1697 VGND.t1965 630.62
R1237 VGND.t1779 VGND.t2155 630.62
R1238 VGND.t525 VGND.t41 630.62
R1239 VGND.t357 VGND.t2147 630.62
R1240 VGND.t531 VGND.t2145 630.62
R1241 VGND.t358 VGND.t39 630.62
R1242 VGND.t1338 VGND.t37 630.62
R1243 VGND.t2668 VGND.t2149 630.62
R1244 VGND.t2249 VGND.t47 630.62
R1245 VGND.t172 VGND.t45 630.62
R1246 VGND.t2018 VGND.t2143 630.62
R1247 VGND.t2141 VGND.t393 630.62
R1248 VGND.t1967 VGND.t405 630.62
R1249 VGND.t2153 VGND.t2397 630.62
R1250 VGND.t1350 VGND.t1188 630.62
R1251 VGND.t2107 VGND.t863 630.62
R1252 VGND.t576 VGND.t1687 630.62
R1253 VGND.t1685 VGND.t827 630.62
R1254 VGND.t1186 VGND.t2042 630.62
R1255 VGND.t295 VGND.t321 630.62
R1256 VGND.t293 VGND.t417 630.62
R1257 VGND.t1184 VGND.t398 630.62
R1258 VGND.t1180 VGND.t434 630.62
R1259 VGND.t297 VGND.t1548 630.62
R1260 VGND.t1683 VGND.t1938 630.62
R1261 VGND.t1190 VGND.t1609 630.62
R1262 VGND.t291 VGND.t2567 630.62
R1263 VGND.t289 VGND.t1144 630.62
R1264 VGND.t241 VGND.t1689 630.62
R1265 VGND.t865 VGND.t1444 630.62
R1266 VGND.t1483 VGND.t1977 630.62
R1267 VGND.t311 VGND.t1099 630.62
R1268 VGND.t78 VGND.t2387 630.62
R1269 VGND.t1783 VGND.t2365 630.62
R1270 VGND.t2055 VGND.t1472 630.62
R1271 VGND.t354 VGND.t1080 630.62
R1272 VGND.t539 VGND.t1069 630.62
R1273 VGND.t1702 VGND.t1468 630.62
R1274 VGND.t2102 VGND.t1450 630.62
R1275 VGND.t2123 VGND.t1082 630.62
R1276 VGND.t101 VGND.t2352 630.62
R1277 VGND.t2492 VGND.t1516 630.62
R1278 VGND.t2026 VGND.t1064 630.62
R1279 VGND.t844 VGND.t1051 630.62
R1280 VGND.t409 VGND.t2393 630.62
R1281 VGND.t1126 VGND.t1055 630.62
R1282 VGND.n990 VGND.n962 599.125
R1283 VGND.n113 VGND.n112 599.125
R1284 VGND.n2875 VGND.n2874 599.125
R1285 VGND.n2908 VGND.n2907 599.125
R1286 VGND.n2912 VGND.n2911 599.125
R1287 VGND.n2923 VGND.n2922 599.125
R1288 VGND.n2995 VGND.n2993 599.125
R1289 VGND.n2962 VGND.n2961 599.125
R1290 VGND.t2288 VGND 581.61
R1291 VGND.t1934 VGND 573.181
R1292 VGND.t216 VGND 573.181
R1293 VGND.t1620 VGND 573.181
R1294 VGND VGND.t1309 573.181
R1295 VGND.t1707 VGND 564.751
R1296 VGND.n3013 VGND 564.751
R1297 VGND.n3012 VGND 564.751
R1298 VGND.n3011 VGND 556.322
R1299 VGND VGND.t749 539.465
R1300 VGND.t1282 VGND 539.465
R1301 VGND.n1123 VGND.t1047 500.166
R1302 VGND.t1511 VGND.n1132 500.166
R1303 VGND.n1133 VGND.t1487 500.166
R1304 VGND.t1045 VGND.n1145 500.166
R1305 VGND.n1146 VGND.t2400 500.166
R1306 VGND.t2378 VGND.n1164 500.166
R1307 VGND.n1165 VGND.t1112 500.166
R1308 VGND.t1092 VGND.n1177 500.166
R1309 VGND.n1178 VGND.t2373 500.166
R1310 VGND.t1470 VGND.n1196 500.166
R1311 VGND.n1197 VGND.t1459 500.166
R1312 VGND.t1067 VGND.n1209 500.166
R1313 VGND.n1210 VGND.t2363 500.166
R1314 VGND.t1448 VGND.n1228 500.166
R1315 VGND.n1229 VGND.t1078 500.166
R1316 VGND.t167 VGND.n578 494.779
R1317 VGND.t819 VGND.t163 481.877
R1318 VGND.t163 VGND.t2056 481.877
R1319 VGND.t1538 VGND.t29 481.877
R1320 VGND.t142 VGND.t1538 481.877
R1321 VGND.t1168 VGND 452.382
R1322 VGND.n1123 VGND.t1294 431.301
R1323 VGND.n1132 VGND.t257 431.301
R1324 VGND.n1133 VGND.t1753 431.301
R1325 VGND.n1145 VGND.t255 431.301
R1326 VGND.n1146 VGND.t2028 431.301
R1327 VGND.n1164 VGND.t1182 431.301
R1328 VGND.n1165 VGND.t1179 431.301
R1329 VGND.n1177 VGND.t1604 431.301
R1330 VGND.n1178 VGND.t1167 431.301
R1331 VGND.n1196 VGND.t867 431.301
R1332 VGND.n1197 VGND.t1330 431.301
R1333 VGND.n1209 VGND.t774 431.301
R1334 VGND.n1210 VGND.t119 431.301
R1335 VGND.n1228 VGND.t2488 431.301
R1336 VGND.n1229 VGND.t1635 431.301
R1337 VGND.t2636 VGND.n273 431.301
R1338 VGND.t70 VGND 419.68
R1339 VGND.n635 VGND.n147 413.043
R1340 VGND.t1843 VGND.t1072 408.469
R1341 VGND.t1792 VGND.t2359 408.469
R1342 VGND.t1455 VGND.t1798 408.469
R1343 VGND.t1804 VGND.t1130 408.469
R1344 VGND.t2357 VGND.t1891 408.469
R1345 VGND.t1897 VGND.t2346 408.469
R1346 VGND.t1502 VGND.t1810 408.469
R1347 VGND.t1852 VGND.t1060 408.469
R1348 VGND.t2404 VGND.t1867 408.469
R1349 VGND.t1903 VGND.t1498 408.469
R1350 VGND.t1114 VGND.t1825 408.469
R1351 VGND.t1870 VGND.t1102 408.469
R1352 VGND.t2375 VGND.t1909 408.469
R1353 VGND.t1921 VGND.t1485 408.469
R1354 VGND.t1090 VGND.t1837 408.469
R1355 VGND.t2389 VGND.t1879 408.469
R1356 VGND.t1233 VGND.t1831 408.469
R1357 VGND.t1717 VGND.t945 408.469
R1358 VGND.t683 VGND.t109 408.469
R1359 VGND.t1678 VGND.t2426 408.469
R1360 VGND.t2513 VGND.t1982 408.469
R1361 VGND.t455 VGND.t523 408.469
R1362 VGND.t1674 VGND.t330 408.469
R1363 VGND.t2450 VGND.t529 408.469
R1364 VGND.t785 VGND.t772 408.469
R1365 VGND.t886 VGND.t1336 408.469
R1366 VGND.t988 VGND.t2665 408.469
R1367 VGND.t1379 VGND.t2131 408.469
R1368 VGND.t878 VGND.t2509 408.469
R1369 VGND.t715 VGND.t2016 408.469
R1370 VGND.t1261 VGND.t1947 408.469
R1371 VGND.t653 VGND.t2228 408.469
R1372 VGND.t2616 VGND.t1906 408.469
R1373 VGND.t1347 VGND.t1279 408.469
R1374 VGND.t303 VGND.t2200 408.469
R1375 VGND.t1217 VGND.t80 408.469
R1376 VGND.t947 VGND.t2406 408.469
R1377 VGND.t918 VGND.t2273 408.469
R1378 VGND.t2454 VGND.t339 408.469
R1379 VGND.t2515 VGND.t415 408.469
R1380 VGND.t457 VGND.t741 408.469
R1381 VGND.t1676 VGND.t201 408.469
R1382 VGND.t803 VGND.t1545 408.469
R1383 VGND.t443 VGND.t2340 408.469
R1384 VGND.t1666 VGND.t1996 408.469
R1385 VGND.t992 VGND.t2565 408.469
R1386 VGND.t2230 VGND.t389 408.469
R1387 VGND.t880 VGND.t410 408.469
R1388 VGND.t1813 VGND.t783 408.469
R1389 VGND.t1658 VGND.t608 408.469
R1390 VGND.t984 VGND.t307 408.469
R1391 VGND.t1693 VGND.t1269 408.469
R1392 VGND.t975 VGND.t1727 408.469
R1393 VGND.t2051 VGND.t697 408.469
R1394 VGND.t1257 VGND.t1300 408.469
R1395 VGND.t535 VGND.t2220 408.469
R1396 VGND.t2527 VGND.t362 408.469
R1397 VGND.t1342 VGND.t933 408.469
R1398 VGND.t1237 VGND.t2118 408.469
R1399 VGND.t2037 VGND.t2521 408.469
R1400 VGND.t687 VGND.t175 408.469
R1401 VGND.t925 VGND.t2022 408.469
R1402 VGND.t2432 VGND.t396 408.469
R1403 VGND.t660 VGND.t2649 408.469
R1404 VGND.t451 VGND.t1855 408.469
R1405 VGND.t2442 VGND.t218 408.469
R1406 VGND.t632 VGND.t797 408.469
R1407 VGND.t1363 VGND.t589 408.469
R1408 VGND.t835 VGND.t1660 408.469
R1409 VGND.t2468 VGND.t226 408.469
R1410 VGND.t350 VGND.t2222 408.469
R1411 VGND.t977 VGND.t369 408.469
R1412 VGND.t10 VGND.t699 408.469
R1413 VGND.t1259 VGND.t871 408.469
R1414 VGND.t2261 VGND.t2620 408.469
R1415 VGND.t691 VGND.t97 408.469
R1416 VGND.t1422 VGND.t2206 408.469
R1417 VGND.t114 VGND.t2184 408.469
R1418 VGND.t2651 VGND.t548 408.469
R1419 VGND.t248 VGND.t929 408.469
R1420 VGND.t912 VGND.t1927 408.469
R1421 VGND.t2659 VGND.t1961 408.469
R1422 VGND.t2092 VGND.t2637 408.469
R1423 VGND.t1698 VGND.t890 408.469
R1424 VGND.t1777 VGND.t2444 408.469
R1425 VGND.t617 VGND.t1385 408.469
R1426 VGND.t326 VGND.t979 408.469
R1427 VGND.t542 VGND.t1662 408.469
R1428 VGND.t1581 VGND.t2472 408.469
R1429 VGND.t1176 VGND.t2224 408.469
R1430 VGND.t1540 VGND.t713 408.469
R1431 VGND.t561 VGND.t2460 408.469
R1432 VGND.t1999 VGND.t2218 408.469
R1433 VGND.t2559 VGND.t2622 408.469
R1434 VGND.t19 VGND.t931 408.469
R1435 VGND.t403 VGND.t1255 408.469
R1436 VGND.t1834 VGND.t1223 408.469
R1437 VGND.t937 VGND.t1715 408.469
R1438 VGND.t673 VGND.t107 408.469
R1439 VGND.t2423 VGND.t1668 408.469
R1440 VGND.t2655 VGND.t1980 408.469
R1441 VGND.t521 VGND.t896 408.469
R1442 VGND.t1006 VGND.t328 408.469
R1443 VGND.t375 VGND.t2438 408.469
R1444 VGND.t1373 VGND.t770 408.469
R1445 VGND.t1334 VGND.t971 408.469
R1446 VGND.t2476 VGND.t2268 408.469
R1447 VGND.t2129 VGND.t1367 408.469
R1448 VGND.t967 VGND.t2506 408.469
R1449 VGND.t707 VGND.t2014 408.469
R1450 VGND.t2204 VGND.t1944 408.469
R1451 VGND.t651 VGND.t2212 408.469
R1452 VGND.t2533 VGND.t1807 408.469
R1453 VGND.t1267 VGND.t1975 408.469
R1454 VGND.t309 VGND.t2188 408.469
R1455 VGND.t2448 VGND.t1691 408.469
R1456 VGND.t1729 VGND.t939 408.469
R1457 VGND.t904 VGND.t2053 408.469
R1458 VGND.t1302 VGND.t2440 408.469
R1459 VGND.t2657 VGND.t537 408.469
R1460 VGND.t1700 VGND.t441 408.469
R1461 VGND.t1656 VGND.t2100 408.469
R1462 VGND.t2120 VGND.t791 408.469
R1463 VGND.t892 VGND.t2039 408.469
R1464 VGND.t177 VGND.t1004 408.469
R1465 VGND.t2024 VGND.t2478 408.469
R1466 VGND.t2214 VGND.t841 408.469
R1467 VGND.t662 VGND.t969 408.469
R1468 VGND.t1849 VGND.t1371 408.469
R1469 VGND.t220 VGND.t998 408.469
R1470 VGND.t634 VGND.t2474 408.469
R1471 VGND.t587 VGND.t2208 408.469
R1472 VGND.t837 VGND.t959 408.469
R1473 VGND.t228 VGND.t951 408.469
R1474 VGND.t352 VGND.t2194 408.469
R1475 VGND.t371 VGND.t2632 408.469
R1476 VGND.t766 VGND.t2519 408.469
R1477 VGND.t873 VGND.t681 408.469
R1478 VGND.t2263 VGND.t1229 408.469
R1479 VGND.t99 VGND.t2661 408.469
R1480 VGND.t1424 VGND.t675 408.469
R1481 VGND.t116 VGND.t916 408.469
R1482 VGND.t550 VGND.t799 408.469
R1483 VGND.t250 VGND.t2639 408.469
R1484 VGND.t894 VGND.t1861 408.469
R1485 VGND.t2434 VGND.t233 408.469
R1486 VGND.t789 VGND.t623 408.469
R1487 VGND.t593 VGND.t2216 408.469
R1488 VGND.t1000 VGND.t831 408.469
R1489 VGND.t2079 VGND.t2456 408.469
R1490 VGND.t2634 VGND.t348 408.469
R1491 VGND.t2595 VGND.t961 408.469
R1492 VGND.t953 VGND.t6 408.469
R1493 VGND.t639 VGND.t2198 408.469
R1494 VGND.t2610 VGND.t2259 408.469
R1495 VGND.t95 VGND.t943 408.469
R1496 VGND.t2190 VGND.t1420 408.469
R1497 VGND.t1231 VGND.t2138 408.469
R1498 VGND.t2641 VGND.t212 408.469
R1499 VGND.t246 VGND.t677 408.469
R1500 VGND.t902 VGND.t1789 408.469
R1501 VGND.t2653 VGND.t1959 408.469
R1502 VGND.t2090 VGND.t465 408.469
R1503 VGND.t973 VGND.t76 408.469
R1504 VGND.t1775 VGND.t2436 408.469
R1505 VGND.t1369 VGND.t615 408.469
R1506 VGND.t324 VGND.t963 408.469
R1507 VGND.t1002 VGND.t540 408.469
R1508 VGND.t1703 VGND.t2458 408.469
R1509 VGND.t2210 VGND.t1174 408.469
R1510 VGND.t2124 VGND.t705 408.469
R1511 VGND.t1275 VGND.t559 408.469
R1512 VGND.t2493 VGND.t2630 408.469
R1513 VGND.t2557 VGND.t2612 408.469
R1514 VGND.t679 VGND.t12 408.469
R1515 VGND.t401 VGND.t2192 408.469
R1516 VGND.t2614 VGND.t1885 408.469
R1517 VGND.t1273 VGND.t811 408.469
R1518 VGND.t1172 VGND.t2196 408.469
R1519 VGND.t579 VGND.t1215 408.469
R1520 VGND.t1734 VGND.t941 408.469
R1521 VGND.t1569 VGND.t914 408.469
R1522 VGND.t335 VGND.t2446 408.469
R1523 VGND.t2588 VGND.t2511 408.469
R1524 VGND.t1404 VGND.t453 408.469
R1525 VGND.t628 VGND.t1670 408.469
R1526 VGND.t732 VGND.t801 408.469
R1527 VGND.t2245 VGND.t898 408.469
R1528 VGND.t1426 VGND.t1664 408.469
R1529 VGND.t154 VGND.t986 408.469
R1530 VGND.t1942 VGND.t2226 408.469
R1531 VGND.t381 VGND.t876 408.469
R1532 VGND.t1680 VGND.t1816 408.469
R1533 VGND.t2645 VGND.t606 408.469
R1534 VGND.t461 VGND.t305 408.469
R1535 VGND.t1695 VGND.t965 408.469
R1536 VGND.t2430 VGND.t1725 408.469
R1537 VGND.t527 VGND.t1365 408.469
R1538 VGND.t957 VGND.t1298 408.469
R1539 VGND.t533 VGND.t996 408.469
R1540 VGND.t1277 VGND.t360 408.469
R1541 VGND.t1340 VGND.t2628 408.469
R1542 VGND.t701 VGND.t2669 408.469
R1543 VGND.t2035 VGND.t1271 408.469
R1544 VGND.t2626 VGND.t173 408.469
R1545 VGND.t2529 VGND.t2020 408.469
R1546 VGND.t671 VGND.t394 408.469
R1547 VGND.t658 VGND.t2186 408.469
R1548 VGND.t1888 VGND.t2647 408.469
R1549 VGND.t1221 VGND.t809 408.469
R1550 VGND.t1170 VGND.t2452 408.469
R1551 VGND.t787 VGND.t581 408.469
R1552 VGND.t1732 VGND.t906 408.469
R1553 VGND.t990 VGND.t1567 408.469
R1554 VGND.t333 VGND.t1383 408.469
R1555 VGND.t445 VGND.t2586 408.469
R1556 VGND.t1402 VGND.t955 408.469
R1557 VGND.t2470 VGND.t438 408.469
R1558 VGND.t730 VGND.t2232 408.469
R1559 VGND.t709 VGND.t193 408.469
R1560 VGND.t1613 VGND.t2462 408.469
R1561 VGND.t152 VGND.t1265 408.469
R1562 VGND.t2523 VGND.t1940 408.469
R1563 VGND.t379 VGND.t693 408.469
R1564 VGND.t685 VGND.t1918 408.469
R1565 VGND.t1345 VGND.t2531 408.469
R1566 VGND.t2517 VGND.t301 408.469
R1567 VGND.t459 VGND.t83 408.469
R1568 VGND.t1225 VGND.t1781 408.469
R1569 VGND.t805 VGND.t2271 408.469
R1570 VGND.t447 VGND.t337 408.469
R1571 VGND.t908 VGND.t413 408.469
R1572 VGND.t994 VGND.t739 408.469
R1573 VGND.t1387 VGND.t199 408.469
R1574 VGND.t882 VGND.t1542 408.469
R1575 VGND.t982 VGND.t2338 408.469
R1576 VGND.t1375 VGND.t2001 408.469
R1577 VGND.t2563 VGND.t2234 408.469
R1578 VGND.t21 VGND.t695 408.469
R1579 VGND.t407 VGND.t2464 408.469
R1580 VGND.t2202 VGND.t1858 408.469
R1581 VGND.t703 VGND.t235 408.469
R1582 VGND.t949 VGND.t625 408.469
R1583 VGND.t591 VGND.t920 408.469
R1584 VGND.t833 VGND.t2535 408.469
R1585 VGND.t2081 VGND.t2643 408.469
R1586 VGND.t346 VGND.t910 408.469
R1587 VGND.t2593 VGND.t1227 408.469
R1588 VGND.t4 VGND.t807 408.469
R1589 VGND.t637 VGND.t449 408.469
R1590 VGND.t736 VGND.t1672 408.469
R1591 VGND.t93 VGND.t795 408.469
R1592 VGND.t1418 VGND.t900 408.469
R1593 VGND.t159 VGND.t884 408.469
R1594 VGND.t2466 VGND.t546 408.469
R1595 VGND.t244 VGND.t1377 408.469
R1596 VGND.t2384 VGND.t888 408.469
R1597 VGND.t793 VGND.t1481 408.469
R1598 VGND.t1381 VGND.t1096 408.469
R1599 VGND.t2624 VGND.t1074 408.469
R1600 VGND.t2480 VGND.t1476 408.469
R1601 VGND.t1263 VGND.t1465 408.469
R1602 VGND.t2618 VGND.t1446 408.469
R1603 VGND.t711 VGND.t2369 408.469
R1604 VGND.t935 VGND.t2348 408.469
R1605 VGND.t1239 VGND.t1139 408.469
R1606 VGND.t2525 VGND.t1062 408.469
R1607 VGND.t689 VGND.t1049 408.469
R1608 VGND.t1235 VGND.t1500 408.469
R1609 VGND.t1219 VGND.t1122 408.469
R1610 VGND.t463 VGND.t2398 408.469
R1611 VGND.t1509 VGND.t923 408.469
R1612 VGND.t144 VGND.t2135 397.848
R1613 VGND.t2135 VGND.t27 397.848
R1614 VGND.t27 VGND.t2503 397.848
R1615 VGND.t2503 VGND.t1311 397.848
R1616 VGND.t1311 VGND.t1312 397.848
R1617 VGND.t1312 VGND.t1315 397.848
R1618 VGND.t1315 VGND.t1316 397.848
R1619 VGND.t2291 VGND.t2672 396.17
R1620 VGND.t1327 VGND.t480 396.17
R1621 VGND.n2998 VGND.n33 394.137
R1622 VGND.n3000 VGND.n2999 394.137
R1623 VGND.n2490 VGND.n32 394.137
R1624 VGND.n2429 VGND.n2428 394.137
R1625 VGND.n2427 VGND.n261 394.137
R1626 VGND.n2426 VGND.n262 394.137
R1627 VGND.n2425 VGND.n263 394.137
R1628 VGND.n2424 VGND.n264 394.137
R1629 VGND.n2423 VGND.n265 394.137
R1630 VGND.n2422 VGND.n266 394.137
R1631 VGND.n2421 VGND.n267 394.137
R1632 VGND.n2420 VGND.n268 394.137
R1633 VGND.n2419 VGND.n269 394.137
R1634 VGND.n2418 VGND.n270 394.137
R1635 VGND.n2417 VGND.n271 394.137
R1636 VGND.n2416 VGND.n272 394.137
R1637 VGND.n2415 VGND.n2414 394.137
R1638 VGND.n147 VGND.t128 387.421
R1639 VGND.n1507 VGND.t500 387.421
R1640 VGND.n1509 VGND.t124 387.421
R1641 VGND.n1511 VGND.t126 387.421
R1642 VGND.n2834 VGND.t510 387.421
R1643 VGND.t1328 VGND.t2112 362.452
R1644 VGND.t2112 VGND.t1282 345.594
R1645 VGND VGND.t751 328.616
R1646 VGND VGND.t610 328.616
R1647 VGND.t169 VGND 328.616
R1648 VGND.t68 VGND 328.616
R1649 VGND VGND.t66 328.616
R1650 VGND.t1519 VGND.t1053 318.947
R1651 VGND.t1513 VGND.t1136 318.947
R1652 VGND.t1121 VGND.t1128 318.947
R1653 VGND.t1106 VGND.t2396 318.947
R1654 VGND.t1507 VGND.t1041 318.947
R1655 VGND.t1491 VGND.t1109 318.947
R1656 VGND.t1044 VGND.t1478 318.947
R1657 VGND.t2402 VGND.t2386 318.947
R1658 VGND.t1480 VGND.t2380 318.947
R1659 VGND.t1493 VGND.t1110 318.947
R1660 VGND.t2383 VGND.t1094 318.947
R1661 VGND.t1085 VGND.t2371 318.947
R1662 VGND.t1467 VGND.t1474 318.947
R1663 VGND.t1462 VGND.t1087 318.947
R1664 VGND.t1066 VGND.t1137 318.947
R1665 VGND.t2367 VGND.t1464 318.947
R1666 VGND.t2300 VGND.t2291 311.877
R1667 VGND.t480 VGND.t2288 311.877
R1668 VGND VGND.t2296 303.449
R1669 VGND VGND.t2300 295.019
R1670 VGND.n70 VGND.t30 287.832
R1671 VGND VGND.t1019 286.591
R1672 VGND.n964 VGND.t2305 282.327
R1673 VGND.n62 VGND.t1558 282.327
R1674 VGND.n969 VGND.t1356 281.13
R1675 VGND.n73 VGND.t147 281.13
R1676 VGND.n126 VGND.t1357 280.978
R1677 VGND.n126 VGND.t162 280.978
R1678 VGND.n594 VGND.t2310 280.978
R1679 VGND.n594 VGND.t1413 280.978
R1680 VGND.n974 VGND.t2057 280.978
R1681 VGND.n156 VGND.t815 280.978
R1682 VGND.n156 VGND.t1416 280.978
R1683 VGND.n96 VGND.t2500 280.978
R1684 VGND.n96 VGND.t2686 280.978
R1685 VGND.n2856 VGND.t1537 280.978
R1686 VGND.n2856 VGND.t136 280.978
R1687 VGND.n2888 VGND.t2679 280.978
R1688 VGND.n2888 VGND.t2491 280.978
R1689 VGND.t2086 VGND 278.161
R1690 VGND.n2994 VGND 271.014
R1691 VGND.n3020 VGND.n4 259.389
R1692 VGND.n2836 VGND.n4 259.389
R1693 VGND.n3021 VGND.n3 252.988
R1694 VGND VGND.t2293 252.875
R1695 VGND VGND.t2298 252.875
R1696 VGND.t1563 VGND 252.875
R1697 VGND VGND.t1527 252.875
R1698 VGND VGND.t148 252.875
R1699 VGND.n676 VGND.t889 241.393
R1700 VGND.n2575 VGND.t1844 241.393
R1701 VGND.n229 VGND.t1234 241.393
R1702 VGND.n239 VGND.t2617 241.393
R1703 VGND.n179 VGND.t784 241.393
R1704 VGND.n1420 VGND.t452 241.393
R1705 VGND.n637 VGND.t913 241.393
R1706 VGND.n616 VGND.t1224 241.393
R1707 VGND.n643 VGND.t2534 241.393
R1708 VGND.n659 VGND.t1372 241.393
R1709 VGND.n668 VGND.t895 241.393
R1710 VGND.n1372 VGND.t903 241.393
R1711 VGND.n1304 VGND.t2615 241.393
R1712 VGND.n572 VGND.t1681 241.393
R1713 VGND.n568 VGND.t2648 241.393
R1714 VGND.n671 VGND.t686 241.393
R1715 VGND.n825 VGND.t2203 241.393
R1716 VGND.n815 VGND.t1847 241.393
R1717 VGND.n1288 VGND.t794 241.284
R1718 VGND.n683 VGND.t1382 241.284
R1719 VGND.n723 VGND.t2625 241.284
R1720 VGND.n728 VGND.t2481 241.284
R1721 VGND.n733 VGND.t1264 241.284
R1722 VGND.n738 VGND.t2619 241.284
R1723 VGND.n743 VGND.t712 241.284
R1724 VGND.n748 VGND.t936 241.284
R1725 VGND.n753 VGND.t1240 241.284
R1726 VGND.n758 VGND.t2526 241.284
R1727 VGND.n763 VGND.t690 241.284
R1728 VGND.n768 VGND.t1236 241.284
R1729 VGND.n773 VGND.t1220 241.284
R1730 VGND.n778 VGND.t464 241.284
R1731 VGND.n1231 VGND.t1883 241.284
R1732 VGND.n1226 VGND.t1841 241.284
R1733 VGND.n794 VGND.t1925 241.284
R1734 VGND.n1207 VGND.t1916 241.284
R1735 VGND.n1199 VGND.t1877 241.284
R1736 VGND.n1194 VGND.t1829 241.284
R1737 VGND.n802 VGND.t1913 241.284
R1738 VGND.n1175 VGND.t1874 241.284
R1739 VGND.n1167 VGND.t1865 241.284
R1740 VGND.n1162 VGND.t1823 241.284
R1741 VGND.n810 VGND.t1901 241.284
R1742 VGND.n1143 VGND.t1895 241.284
R1743 VGND.n1135 VGND.t1820 241.284
R1744 VGND.n1130 VGND.t1802 241.284
R1745 VGND.n1125 VGND.t1796 241.284
R1746 VGND.n2577 VGND.t1793 241.284
R1747 VGND.n2573 VGND.t1799 241.284
R1748 VGND.n2703 VGND.t1805 241.284
R1749 VGND.n2628 VGND.t1892 241.284
R1750 VGND.n2695 VGND.t1898 241.284
R1751 VGND.n2632 VGND.t1811 241.284
R1752 VGND.n2687 VGND.t1853 241.284
R1753 VGND.n2636 VGND.t1868 241.284
R1754 VGND.n2679 VGND.t1904 241.284
R1755 VGND.n2640 VGND.t1826 241.284
R1756 VGND.n2671 VGND.t1871 241.284
R1757 VGND.n2644 VGND.t1910 241.284
R1758 VGND.n2663 VGND.t1922 241.284
R1759 VGND.n2648 VGND.t1838 241.284
R1760 VGND.n2655 VGND.t1880 241.284
R1761 VGND.n232 VGND.t946 241.284
R1762 VGND.n2718 VGND.t684 241.284
R1763 VGND.n2723 VGND.t1679 241.284
R1764 VGND.n2728 VGND.t2514 241.284
R1765 VGND.n2733 VGND.t456 241.284
R1766 VGND.n2738 VGND.t1675 241.284
R1767 VGND.n2743 VGND.t2451 241.284
R1768 VGND.n2748 VGND.t786 241.284
R1769 VGND.n2753 VGND.t887 241.284
R1770 VGND.n2758 VGND.t989 241.284
R1771 VGND.n2763 VGND.t1380 241.284
R1772 VGND.n2768 VGND.t879 241.284
R1773 VGND.n2773 VGND.t716 241.284
R1774 VGND.n2778 VGND.t1262 241.284
R1775 VGND.n227 VGND.t2229 241.284
R1776 VGND.n242 VGND.t1280 241.284
R1777 VGND.n2512 VGND.t2201 241.284
R1778 VGND.n2507 VGND.t1218 241.284
R1779 VGND.n246 VGND.t948 241.284
R1780 VGND.n2437 VGND.t919 241.284
R1781 VGND.n2442 VGND.t2455 241.284
R1782 VGND.n2447 VGND.t2516 241.284
R1783 VGND.n2452 VGND.t458 241.284
R1784 VGND.n2457 VGND.t1677 241.284
R1785 VGND.n2462 VGND.t804 241.284
R1786 VGND.n2467 VGND.t444 241.284
R1787 VGND.n2472 VGND.t1667 241.284
R1788 VGND.n2477 VGND.t993 241.284
R1789 VGND.n2482 VGND.t2231 241.284
R1790 VGND.n2487 VGND.t881 241.284
R1791 VGND.n2830 VGND.t1659 241.284
R1792 VGND.n366 VGND.t985 241.284
R1793 VGND.n370 VGND.t1270 241.284
R1794 VGND.n2170 VGND.t976 241.284
R1795 VGND.n364 VGND.t698 241.284
R1796 VGND.n2196 VGND.t1258 241.284
R1797 VGND.n356 VGND.t2221 241.284
R1798 VGND.n2222 VGND.t2528 241.284
R1799 VGND.n348 VGND.t934 241.284
R1800 VGND.n2248 VGND.t1238 241.284
R1801 VGND.n340 VGND.t2522 241.284
R1802 VGND.n2279 VGND.t688 241.284
R1803 VGND.n2284 VGND.t926 241.284
R1804 VGND.n2289 VGND.t2433 241.284
R1805 VGND.n332 VGND.t2650 241.284
R1806 VGND.n1427 VGND.t2443 241.284
R1807 VGND.n1424 VGND.t798 241.284
R1808 VGND.n2157 VGND.t1364 241.284
R1809 VGND.n379 VGND.t1661 241.284
R1810 VGND.n2183 VGND.t2469 241.284
R1811 VGND.n360 VGND.t2223 241.284
R1812 VGND.n2209 VGND.t978 241.284
R1813 VGND.n352 VGND.t700 241.284
R1814 VGND.n2235 VGND.t1260 241.284
R1815 VGND.n344 VGND.t2621 241.284
R1816 VGND.n2261 VGND.t692 241.284
R1817 VGND.n336 VGND.t2207 241.284
R1818 VGND.n2266 VGND.t2185 241.284
R1819 VGND.n2306 VGND.t2652 241.284
R1820 VGND.n2311 VGND.t930 241.284
R1821 VGND.n1441 VGND.t2660 241.284
R1822 VGND.n634 VGND.t2638 241.284
R1823 VGND.n1491 VGND.t891 241.284
R1824 VGND.n1486 VGND.t2445 241.284
R1825 VGND.n1481 VGND.t1386 241.284
R1826 VGND.n1476 VGND.t980 241.284
R1827 VGND.n1471 VGND.t1663 241.284
R1828 VGND.n1466 VGND.t2473 241.284
R1829 VGND.n1461 VGND.t2225 241.284
R1830 VGND.n1456 VGND.t714 241.284
R1831 VGND.n1451 VGND.t2461 241.284
R1832 VGND.n1446 VGND.t2219 241.284
R1833 VGND.n393 VGND.t2623 241.284
R1834 VGND.n2134 VGND.t932 241.284
R1835 VGND.n2129 VGND.t1256 241.284
R1836 VGND.n1503 VGND.t938 241.284
R1837 VGND.n621 VGND.t674 241.284
R1838 VGND.n625 VGND.t1669 241.284
R1839 VGND.n1996 VGND.t2656 241.284
R1840 VGND.n431 VGND.t897 241.284
R1841 VGND.n2022 VGND.t1007 241.284
R1842 VGND.n423 VGND.t2439 241.284
R1843 VGND.n2048 VGND.t1374 241.284
R1844 VGND.n415 VGND.t972 241.284
R1845 VGND.n2074 VGND.t2477 241.284
R1846 VGND.n407 VGND.t1368 241.284
R1847 VGND.n2105 VGND.t968 241.284
R1848 VGND.n2110 VGND.t708 241.284
R1849 VGND.n2115 VGND.t2205 241.284
R1850 VGND.n2120 VGND.t2213 241.284
R1851 VGND.n650 VGND.t1268 241.284
R1852 VGND.n647 VGND.t2189 241.284
R1853 VGND.n1983 VGND.t2449 241.284
R1854 VGND.n435 VGND.t940 241.284
R1855 VGND.n2009 VGND.t905 241.284
R1856 VGND.n427 VGND.t2441 241.284
R1857 VGND.n2035 VGND.t2658 241.284
R1858 VGND.n419 VGND.t442 241.284
R1859 VGND.n2061 VGND.t1657 241.284
R1860 VGND.n411 VGND.t792 241.284
R1861 VGND.n2087 VGND.t893 241.284
R1862 VGND.n403 VGND.t1005 241.284
R1863 VGND.n2092 VGND.t2479 241.284
R1864 VGND.n2331 VGND.t2215 241.284
R1865 VGND.n2336 VGND.t970 241.284
R1866 VGND.n957 VGND.t999 241.284
R1867 VGND.n952 VGND.t2475 241.284
R1868 VGND.n947 VGND.t2209 241.284
R1869 VGND.n942 VGND.t960 241.284
R1870 VGND.n937 VGND.t952 241.284
R1871 VGND.n932 VGND.t2195 241.284
R1872 VGND.n927 VGND.t2633 241.284
R1873 VGND.n922 VGND.t2520 241.284
R1874 VGND.n917 VGND.t682 241.284
R1875 VGND.n912 VGND.t1230 241.284
R1876 VGND.n907 VGND.t2662 241.284
R1877 VGND.n902 VGND.t676 241.284
R1878 VGND.n449 VGND.t917 241.284
R1879 VGND.n1960 VGND.t800 241.284
R1880 VGND.n1955 VGND.t2640 241.284
R1881 VGND.n1394 VGND.t2435 241.284
R1882 VGND.n1399 VGND.t790 241.284
R1883 VGND.n666 VGND.t2217 241.284
R1884 VGND.n1822 VGND.t1001 241.284
R1885 VGND.n487 VGND.t2457 241.284
R1886 VGND.n1848 VGND.t2635 241.284
R1887 VGND.n479 VGND.t962 241.284
R1888 VGND.n1874 VGND.t954 241.284
R1889 VGND.n471 VGND.t2199 241.284
R1890 VGND.n1900 VGND.t2611 241.284
R1891 VGND.n463 VGND.t944 241.284
R1892 VGND.n1931 VGND.t2191 241.284
R1893 VGND.n1936 VGND.t1232 241.284
R1894 VGND.n1941 VGND.t2642 241.284
R1895 VGND.n1946 VGND.t678 241.284
R1896 VGND.n1379 VGND.t2654 241.284
R1897 VGND.n1376 VGND.t466 241.284
R1898 VGND.n1809 VGND.t974 241.284
R1899 VGND.n491 VGND.t2437 241.284
R1900 VGND.n1835 VGND.t1370 241.284
R1901 VGND.n483 VGND.t964 241.284
R1902 VGND.n1861 VGND.t1003 241.284
R1903 VGND.n475 VGND.t2459 241.284
R1904 VGND.n1887 VGND.t2211 241.284
R1905 VGND.n467 VGND.t706 241.284
R1906 VGND.n1913 VGND.t1276 241.284
R1907 VGND.n459 VGND.t2631 241.284
R1908 VGND.n1918 VGND.t2613 241.284
R1909 VGND.n2356 VGND.t680 241.284
R1910 VGND.n2361 VGND.t2193 241.284
R1911 VGND.n1311 VGND.t1274 241.284
R1912 VGND.n1308 VGND.t2197 241.284
R1913 VGND.n1361 VGND.t1216 241.284
R1914 VGND.n1356 VGND.t942 241.284
R1915 VGND.n1351 VGND.t915 241.284
R1916 VGND.n1346 VGND.t2447 241.284
R1917 VGND.n1341 VGND.t2512 241.284
R1918 VGND.n1336 VGND.t454 241.284
R1919 VGND.n1331 VGND.t1671 241.284
R1920 VGND.n1326 VGND.t802 241.284
R1921 VGND.n1321 VGND.t899 241.284
R1922 VGND.n1316 VGND.t1665 241.284
R1923 VGND.n505 VGND.t987 241.284
R1924 VGND.n1786 VGND.t2227 241.284
R1925 VGND.n1781 VGND.t877 241.284
R1926 VGND.n1516 VGND.t2646 241.284
R1927 VGND.n1521 VGND.t462 241.284
R1928 VGND.n577 VGND.t966 241.284
R1929 VGND.n1648 VGND.t2431 241.284
R1930 VGND.n543 VGND.t1366 241.284
R1931 VGND.n1674 VGND.t958 241.284
R1932 VGND.n535 VGND.t997 241.284
R1933 VGND.n1700 VGND.t1278 241.284
R1934 VGND.n527 VGND.t2629 241.284
R1935 VGND.n1726 VGND.t702 241.284
R1936 VGND.n519 VGND.t1272 241.284
R1937 VGND.n1757 VGND.t2627 241.284
R1938 VGND.n1762 VGND.t2530 241.284
R1939 VGND.n1767 VGND.t672 241.284
R1940 VGND.n1772 VGND.t2187 241.284
R1941 VGND.n1536 VGND.t1222 241.284
R1942 VGND.n566 VGND.t2453 241.284
R1943 VGND.n1635 VGND.t788 241.284
R1944 VGND.n547 VGND.t907 241.284
R1945 VGND.n1661 VGND.t991 241.284
R1946 VGND.n539 VGND.t1384 241.284
R1947 VGND.n1687 VGND.t446 241.284
R1948 VGND.n531 VGND.t956 241.284
R1949 VGND.n1713 VGND.t2471 241.284
R1950 VGND.n523 VGND.t2233 241.284
R1951 VGND.n1739 VGND.t710 241.284
R1952 VGND.n515 VGND.t2463 241.284
R1953 VGND.n1744 VGND.t1266 241.284
R1954 VGND.n2381 VGND.t2524 241.284
R1955 VGND.n2386 VGND.t694 241.284
R1956 VGND.n674 VGND.t2532 241.284
R1957 VGND.n1549 VGND.t2518 241.284
R1958 VGND.n1554 VGND.t460 241.284
R1959 VGND.n1559 VGND.t1226 241.284
R1960 VGND.n1564 VGND.t806 241.284
R1961 VGND.n1569 VGND.t448 241.284
R1962 VGND.n1574 VGND.t909 241.284
R1963 VGND.n1579 VGND.t995 241.284
R1964 VGND.n1584 VGND.t1388 241.284
R1965 VGND.n1589 VGND.t883 241.284
R1966 VGND.n1594 VGND.t983 241.284
R1967 VGND.n1599 VGND.t1376 241.284
R1968 VGND.n561 VGND.t2235 241.284
R1969 VGND.n1612 VGND.t696 241.284
R1970 VGND.n1607 VGND.t2465 241.284
R1971 VGND.n833 VGND.t704 241.284
R1972 VGND.n838 VGND.t950 241.284
R1973 VGND.n830 VGND.t921 241.284
R1974 VGND.n888 VGND.t2536 241.284
R1975 VGND.n883 VGND.t2644 241.284
R1976 VGND.n878 VGND.t911 241.284
R1977 VGND.n873 VGND.t1228 241.284
R1978 VGND.n868 VGND.t808 241.284
R1979 VGND.n863 VGND.t450 241.284
R1980 VGND.n858 VGND.t1673 241.284
R1981 VGND.n853 VGND.t796 241.284
R1982 VGND.n848 VGND.t901 241.284
R1983 VGND.n843 VGND.t885 241.284
R1984 VGND.n2401 VGND.t2467 241.284
R1985 VGND.n2406 VGND.t1378 241.284
R1986 VGND.n719 VGND.t924 241.284
R1987 VGND.t2361 VGND.t1843 222.15
R1988 VGND.t2094 VGND.t1461 222.15
R1989 VGND.t1457 VGND.t1792 222.15
R1990 VGND.t238 VGND.t1084 222.15
R1991 VGND.t1798 VGND.t1076 222.15
R1992 VGND.t1071 VGND.t1608 222.15
R1993 VGND.t1056 VGND.t1804 222.15
R1994 VGND.t1400 VGND.t1520 222.15
R1995 VGND.t1891 VGND.t2354 222.15
R1996 VGND.t1453 VGND.t1711 222.15
R1997 VGND.t1132 VGND.t1897 222.15
R1998 VGND.t601 VGND.t1058 222.15
R1999 VGND.t1810 VGND.t1118 222.15
R2000 VGND.t2356 VGND.t214 222.15
R2001 VGND.t2350 VGND.t1852 222.15
R2002 VGND.t667 VGND.t1508 222.15
R2003 VGND.t1867 VGND.t1504 222.15
R2004 VGND.t1120 VGND.t484 222.15
R2005 VGND.t1134 VGND.t1903 222.15
R2006 VGND.t848 VGND.t1059 222.15
R2007 VGND.t1825 VGND.t1039 222.15
R2008 VGND.t1506 VGND.t50 222.15
R2009 VGND.t2391 VGND.t1870 222.15
R2010 VGND.t467 VGND.t1496 222.15
R2011 VGND.t1909 VGND.t1116 222.15
R2012 VGND.t1111 VGND.t1951 222.15
R2013 VGND.t1104 VGND.t1921 222.15
R2014 VGND.t1632 VGND.t2395 222.15
R2015 VGND.t1837 VGND.t1088 222.15
R2016 VGND.t2372 VGND.t1443 222.15
R2017 VGND.t1879 VGND.t1489 222.15
R2018 VGND.t1108 VGND.t573 222.15
R2019 VGND.t1243 VGND.t1233 222.15
R2020 VGND.t2671 VGND.t814 222.15
R2021 VGND.t945 VGND.t1754 222.15
R2022 VGND.t621 VGND.t0 222.15
R2023 VGND.t1251 VGND.t683 222.15
R2024 VGND.t507 VGND.t595 222.15
R2025 VGND.t1249 VGND.t1678 222.15
R2026 VGND.t1206 VGND.t1979 222.15
R2027 VGND.t1241 VGND.t2513 222.15
R2028 VGND.t1605 VGND.t2077 222.15
R2029 VGND.t1033 VGND.t455 222.15
R2030 VGND.t278 VGND.t342 222.15
R2031 VGND.t1031 VGND.t1674 222.15
R2032 VGND.t2065 VGND.t2591 222.15
R2033 VGND.t1760 VGND.t2450 222.15
R2034 VGND.t1607 VGND.t2 222.15
R2035 VGND.t1758 VGND.t785 222.15
R2036 VGND.t1156 VGND.t869 222.15
R2037 VGND.t1035 VGND.t886 222.15
R2038 VGND.t2483 VGND.t735 222.15
R2039 VGND.t1247 VGND.t988 222.15
R2040 VGND.t57 VGND.t2343 222.15
R2041 VGND.t1245 VGND.t1379 222.15
R2042 VGND.t315 VGND.t1417 222.15
R2043 VGND.t1029 VGND.t878 222.15
R2044 VGND.t274 VGND.t157 222.15
R2045 VGND.t1027 VGND.t715 222.15
R2046 VGND.t2663 VGND.t211 222.15
R2047 VGND.t1025 VGND.t1261 222.15
R2048 VGND.t2099 VGND.t650 222.15
R2049 VGND.t2228 VGND.t1756 222.15
R2050 VGND.t1497 VGND.t1291 222.15
R2051 VGND.t268 VGND.t2616 222.15
R2052 VGND.t2599 VGND.t605 222.15
R2053 VGND.t1279 VGND.t2555 222.15
R2054 VGND.t112 VGND.t1949 222.15
R2055 VGND.t2200 VGND.t1322 222.15
R2056 VGND.t563 VGND.t1293 222.15
R2057 VGND.t1320 VGND.t1217 222.15
R2058 VGND.t1602 VGND.t1780 222.15
R2059 VGND.t2242 VGND.t947 222.15
R2060 VGND.t583 VGND.t526 222.15
R2061 VGND.t2551 VGND.t918 222.15
R2062 VGND.t519 VGND.t345 222.15
R2063 VGND.t2549 VGND.t2454 222.15
R2064 VGND.t747 VGND.t532 222.15
R2065 VGND.t2240 VGND.t2515 222.15
R2066 VGND.t516 VGND.t359 222.15
R2067 VGND.t2238 VGND.t457 222.15
R2068 VGND.t222 VGND.t1339 222.15
R2069 VGND.t2553 VGND.t1676 222.15
R2070 VGND.t850 VGND.t2122 222.15
R2071 VGND.t272 VGND.t803 222.15
R2072 VGND.t665 VGND.t2250 222.15
R2073 VGND.t270 VGND.t443 222.15
R2074 VGND.t2285 VGND.t179 222.15
R2075 VGND.t2547 VGND.t1666 222.15
R2076 VGND.t1408 VGND.t2019 222.15
R2077 VGND.t2545 VGND.t992 222.15
R2078 VGND.t55 VGND.t843 222.15
R2079 VGND.t1324 VGND.t2230 222.15
R2080 VGND.t602 VGND.t406 222.15
R2081 VGND.t2236 VGND.t880 222.15
R2082 VGND.t2429 VGND.t1043 222.15
R2083 VGND.t783 VGND.t854 222.15
R2084 VGND.t232 VGND.t2410 222.15
R2085 VGND.t1159 VGND.t1658 222.15
R2086 VGND.t275 VGND.t627 222.15
R2087 VGND.t282 VGND.t984 222.15
R2088 VGND.t366 VGND.t585 222.15
R2089 VGND.t1269 VGND.t860 222.15
R2090 VGND.t1985 VGND.t1304 222.15
R2091 VGND.t852 VGND.t975 222.15
R2092 VGND.t224 VGND.t2083 222.15
R2093 VGND.t697 VGND.t2072 222.15
R2094 VGND.t344 VGND.t2598 222.15
R2095 VGND.t2070 VGND.t1257 222.15
R2096 VGND.t277 VGND.t367 222.15
R2097 VGND.t2220 VGND.t1165 222.15
R2098 VGND.t8 VGND.t2602 222.15
R2099 VGND.t1163 VGND.t2527 222.15
R2100 VGND.t1401 VGND.t641 222.15
R2101 VGND.t933 VGND.t2074 222.15
R2102 VGND.t2266 VGND.t317 222.15
R2103 VGND.t858 VGND.t1237 222.15
R2104 VGND.t1392 VGND.t2345 222.15
R2105 VGND.t2521 VGND.t856 222.15
R2106 VGND.t1932 VGND.t1196 222.15
R2107 VGND.t2068 VGND.t687 222.15
R2108 VGND.t18 VGND.t2140 222.15
R2109 VGND.t286 VGND.t925 222.15
R2110 VGND.t1142 VGND.t517 222.15
R2111 VGND.t284 VGND.t2432 222.15
R2112 VGND.t2105 VGND.t656 222.15
R2113 VGND.t2649 VGND.t1161 222.15
R2114 VGND.t1518 VGND.t468 222.15
R2115 VGND.t478 VGND.t451 222.15
R2116 VGND.t1295 VGND.t204 222.15
R2117 VGND.t2033 VGND.t2442 222.15
R2118 VGND.t440 VGND.t2109 222.15
R2119 VGND.t797 VGND.t2543 222.15
R2120 VGND.t575 VGND.t758 222.15
R2121 VGND.t2541 VGND.t1363 222.15
R2122 VGND.t2284 VGND.t829 222.15
R2123 VGND.t1660 VGND.t476 222.15
R2124 VGND.t2043 VGND.t782 222.15
R2125 VGND.t2029 VGND.t2468 222.15
R2126 VGND.t1972 VGND.t322 222.15
R2127 VGND.t2222 VGND.t570 222.15
R2128 VGND.t2584 VGND.t1143 222.15
R2129 VGND.t474 VGND.t977 222.15
R2130 VGND.t1616 VGND.t612 222.15
R2131 VGND.t699 VGND.t472 222.15
R2132 VGND.t436 VGND.t738 222.15
R2133 VGND.t2031 VGND.t1259 222.15
R2134 VGND.t2277 VGND.t728 222.15
R2135 VGND.t2620 VGND.t2539 222.15
R2136 VGND.t557 VGND.t279 222.15
R2137 VGND.t2537 VGND.t691 222.15
R2138 VGND.t603 VGND.t1611 222.15
R2139 VGND.t2206 VGND.t568 222.15
R2140 VGND.t150 VGND.t1986 222.15
R2141 VGND.t2184 VGND.t566 222.15
R2142 VGND.t1146 VGND.t1719 222.15
R2143 VGND.t564 VGND.t2651 222.15
R2144 VGND.t574 VGND.t242 222.15
R2145 VGND.t929 VGND.t470 222.15
R2146 VGND.t1452 VGND.t1281 222.15
R2147 VGND.t1650 VGND.t912 222.15
R2148 VGND.t1149 VGND.t1714 222.15
R2149 VGND.t2255 VGND.t2659 222.15
R2150 VGND.t614 VGND.t106 222.15
R2151 VGND.t2637 VGND.t1929 222.15
R2152 VGND.t2425 VGND.t2066 222.15
R2153 VGND.t890 VGND.t1600 222.15
R2154 VGND.t1774 VGND.t207 222.15
R2155 VGND.t2444 VGND.t1648 222.15
R2156 VGND.t520 VGND.t2003 222.15
R2157 VGND.t1385 VGND.t2251 222.15
R2158 VGND.t356 VGND.t16 222.15
R2159 VGND.t979 VGND.t1642 222.15
R2160 VGND.t374 VGND.t849 222.15
R2161 VGND.t1662 VGND.t1646 222.15
R2162 VGND.t769 VGND.t2089 222.15
R2163 VGND.t2472 VGND.t1644 222.15
R2164 VGND.t762 VGND.t209 222.15
R2165 VGND.t2224 VGND.t2253 222.15
R2166 VGND.t2667 VGND.t2027 222.15
R2167 VGND.t713 VGND.t1598 222.15
R2168 VGND.t2248 VGND.t1585 222.15
R2169 VGND.t2460 VGND.t1652 222.15
R2170 VGND.t171 VGND.t1712 222.15
R2171 VGND.t2218 VGND.t1640 222.15
R2172 VGND.t2013 VGND.t206 222.15
R2173 VGND.t2622 VGND.t1638 222.15
R2174 VGND.t392 VGND.t288 222.15
R2175 VGND.t931 VGND.t1636 222.15
R2176 VGND.t400 VGND.t2287 222.15
R2177 VGND.t1255 VGND.t2257 222.15
R2178 VGND.t2382 VGND.t515 222.15
R2179 VGND.t1223 VGND.t2182 222.15
R2180 VGND.t813 VGND.t14 222.15
R2181 VGND.t418 VGND.t937 222.15
R2182 VGND.t54 VGND.t620 222.15
R2183 VGND.t2326 VGND.t673 222.15
R2184 VGND.t555 VGND.t584 222.15
R2185 VGND.t1668 VGND.t2324 222.15
R2186 VGND.t1978 VGND.t745 222.15
R2187 VGND.t2180 VGND.t2655 222.15
R2188 VGND.t387 VGND.t2076 222.15
R2189 VGND.t896 VGND.t2336 222.15
R2190 VGND.t341 VGND.t1203 222.15
R2191 VGND.t2334 VGND.t1006 222.15
R2192 VGND.t1399 VGND.t2590 222.15
R2193 VGND.t2438 VGND.t2178 222.15
R2194 VGND.t1406 VGND.t253 222.15
R2195 VGND.t2176 VGND.t1373 222.15
R2196 VGND.t1953 VGND.t630 222.15
R2197 VGND.t971 VGND.t497 222.15
R2198 VGND.t734 VGND.t845 222.15
R2199 VGND.t2322 VGND.t2476 222.15
R2200 VGND.t1351 VGND.t2342 222.15
R2201 VGND.t1367 VGND.t2320 222.15
R2202 VGND.t1428 VGND.t2060 222.15
R2203 VGND.t2332 VGND.t967 222.15
R2204 VGND.t2601 VGND.t156 222.15
R2205 VGND.t2330 VGND.t707 222.15
R2206 VGND.t1950 VGND.t210 222.15
R2207 VGND.t2328 VGND.t2204 222.15
R2208 VGND.t1409 VGND.t252 222.15
R2209 VGND.t2212 VGND.t2174 222.15
R2210 VGND.t1495 VGND.t1333 222.15
R2211 VGND.t1772 VGND.t2533 222.15
R2212 VGND.t1141 VGND.t237 222.15
R2213 VGND.t1762 VGND.t1267 222.15
R2214 VGND.t499 VGND.t631 222.15
R2215 VGND.t2188 VGND.t1592 222.15
R2216 VGND.t2422 VGND.t1306 222.15
R2217 VGND.t1590 VGND.t2448 222.15
R2218 VGND.t868 VGND.t1724 222.15
R2219 VGND.t939 VGND.t1770 222.15
R2220 VGND.t225 VGND.t1394 222.15
R2221 VGND.t646 VGND.t904 222.15
R2222 VGND.t862 VGND.t332 222.15
R2223 VGND.t2440 VGND.t644 222.15
R2224 VGND.t368 VGND.t469 222.15
R2225 VGND.t1768 VGND.t2657 222.15
R2226 VGND.t1326 VGND.t9 222.15
R2227 VGND.t441 VGND.t1766 222.15
R2228 VGND.t870 VGND.t597 222.15
R2229 VGND.t648 VGND.t1656 222.15
R2230 VGND.t2286 VGND.t2267 222.15
R2231 VGND.t791 VGND.t1588 222.15
R2232 VGND.t192 VGND.t223 222.15
R2233 VGND.t1586 VGND.t892 222.15
R2234 VGND.t2067 VGND.t1933 222.15
R2235 VGND.t1004 VGND.t642 222.15
R2236 VGND.t113 VGND.t1752 222.15
R2237 VGND.t2478 VGND.t1596 222.15
R2238 VGND.t518 VGND.t1630 222.15
R2239 VGND.t1594 VGND.t2214 222.15
R2240 VGND.t1958 VGND.t657 222.15
R2241 VGND.t969 VGND.t1764 222.15
R2242 VGND.t1521 VGND.t1352 222.15
R2243 VGND.t1371 VGND.t260 222.15
R2244 VGND.t205 VGND.t276 222.15
R2245 VGND.t998 VGND.t2061 222.15
R2246 VGND.t2110 VGND.t1008 222.15
R2247 VGND.t2474 VGND.t2275 222.15
R2248 VGND.t578 VGND.t120 222.15
R2249 VGND.t2208 VGND.t266 222.15
R2250 VGND.t830 VGND.t1389 222.15
R2251 VGND.t959 VGND.t1993 222.15
R2252 VGND.t2044 VGND.t256 222.15
R2253 VGND.t951 VGND.t1152 222.15
R2254 VGND.t323 VGND.t1344 222.15
R2255 VGND.t2194 VGND.t1150 222.15
R2256 VGND.t2585 VGND.t2609 222.15
R2257 VGND.t2632 VGND.t1991 222.15
R2258 VGND.t613 VGND.t764 222.15
R2259 VGND.t2519 VGND.t1989 222.15
R2260 VGND.t437 VGND.t2484 222.15
R2261 VGND.t681 VGND.t1154 222.15
R2262 VGND.t729 VGND.t553 222.15
R2263 VGND.t1229 VGND.t264 222.15
R2264 VGND.t558 VGND.t2688 222.15
R2265 VGND.t2661 VGND.t262 222.15
R2266 VGND.t1612 VGND.t1615 222.15
R2267 VGND.t675 VGND.t780 222.15
R2268 VGND.t151 VGND.t1973 222.15
R2269 VGND.t916 VGND.t778 222.15
R2270 VGND.t1939 VGND.t757 222.15
R2271 VGND.t799 VGND.t776 222.15
R2272 VGND.t243 VGND.t1192 222.15
R2273 VGND.t2639 VGND.t1987 222.15
R2274 VGND.t1454 VGND.t1391 222.15
R2275 VGND.t1213 VGND.t894 222.15
R2276 VGND.t670 VGND.t1349 222.15
R2277 VGND.t89 VGND.t2434 222.15
R2278 VGND.t1289 VGND.t2108 222.15
R2279 VGND.t1555 VGND.t789 222.15
R2280 VGND.t1332 VGND.t577 222.15
R2281 VGND.t2216 VGND.t1553 222.15
R2282 VGND.t828 VGND.t2675 222.15
R2283 VGND.t1211 VGND.t1000 222.15
R2284 VGND.t1201 VGND.t2041 222.15
R2285 VGND.t2456 VGND.t85 222.15
R2286 VGND.t320 VGND.t847 222.15
R2287 VGND.t2010 VGND.t2634 222.15
R2288 VGND.t208 VGND.t2583 222.15
R2289 VGND.t961 VGND.t1209 222.15
R2290 VGND.t399 VGND.t1974 222.15
R2291 VGND.t1207 VGND.t953 222.15
R2292 VGND.t1148 VGND.t435 222.15
R2293 VGND.t2198 VGND.t87 222.15
R2294 VGND.t727 VGND.t2244 222.15
R2295 VGND.t1551 VGND.t2610 222.15
R2296 VGND.t2676 VGND.t556 222.15
R2297 VGND.t943 VGND.t1549 222.15
R2298 VGND.t1610 VGND.t1682 222.15
R2299 VGND.t2008 VGND.t2190 222.15
R2300 VGND.t666 VGND.t2568 222.15
R2301 VGND.t2006 VGND.t1231 222.15
R2302 VGND.t2104 VGND.t1145 222.15
R2303 VGND.t2004 VGND.t2641 222.15
R2304 VGND.t1390 VGND.t383 222.15
R2305 VGND.t677 VGND.t91 222.15
R2306 VGND.t1445 VGND.t1655 222.15
R2307 VGND.t491 VGND.t902 222.15
R2308 VGND.t2088 VGND.t1713 222.15
R2309 VGND.t2579 VGND.t2653 222.15
R2310 VGND.t1396 VGND.t2106 222.15
R2311 VGND.t465 VGND.t64 222.15
R2312 VGND.t2428 VGND.t508 222.15
R2313 VGND.t62 VGND.t973 222.15
R2314 VGND.t1158 VGND.t1731 222.15
R2315 VGND.t2436 VGND.t489 222.15
R2316 VGND.t840 VGND.t1722 222.15
R2317 VGND.t2575 VGND.t1369 222.15
R2318 VGND.t1195 VGND.t355 222.15
R2319 VGND.t963 VGND.t2573 222.15
R2320 VGND.t373 VGND.t1284 222.15
R2321 VGND.t487 VGND.t1002 222.15
R2322 VGND.t2487 VGND.t768 222.15
R2323 VGND.t2458 VGND.t485 222.15
R2324 VGND.t761 VGND.t2064 222.15
R2325 VGND.t2577 VGND.t2210 222.15
R2326 VGND.t1710 VGND.t2664 222.15
R2327 VGND.t705 VGND.t495 222.15
R2328 VGND.t2247 VGND.t1205 222.15
R2329 VGND.t493 VGND.t1275 222.15
R2330 VGND.t1720 VGND.t2508 222.15
R2331 VGND.t2630 VGND.t2571 222.15
R2332 VGND.t2012 VGND.t875 222.15
R2333 VGND.t2612 VGND.t2569 222.15
R2334 VGND.t1946 VGND.t505 222.15
R2335 VGND.t482 VGND.t679 222.15
R2336 VGND.t52 VGND.t664 222.15
R2337 VGND.t2192 VGND.t2581 222.15
R2338 VGND.t2377 VGND.t2600 222.15
R2339 VGND.t1738 VGND.t2614 222.15
R2340 VGND.t2290 VGND.t1964 222.15
R2341 VGND.t2165 VGND.t1273 222.15
R2342 VGND.t259 VGND.t300 222.15
R2343 VGND.t2196 VGND.t1746 222.15
R2344 VGND.t79 VGND.t2603 222.15
R2345 VGND.t1215 VGND.t1744 222.15
R2346 VGND.t2409 VGND.t49 222.15
R2347 VGND.t941 VGND.t1736 222.15
R2348 VGND.t2270 VGND.t53 222.15
R2349 VGND.t914 VGND.t2161 222.15
R2350 VGND.t1297 VGND.t1198 222.15
R2351 VGND.t2446 VGND.t2159 222.15
R2352 VGND.t412 VGND.t839 222.15
R2353 VGND.t2511 VGND.t2171 222.15
R2354 VGND.t1584 VGND.t280 222.15
R2355 VGND.t453 VGND.t2169 222.15
R2356 VGND.t198 VGND.t509 222.15
R2357 VGND.t1670 VGND.t2163 222.15
R2358 VGND.t1547 VGND.t2608 222.15
R2359 VGND.t801 VGND.t1742 222.15
R2360 VGND.t2134 VGND.t1157 222.15
R2361 VGND.t898 VGND.t1740 222.15
R2362 VGND.t1998 VGND.t385 222.15
R2363 VGND.t1664 VGND.t2157 222.15
R2364 VGND.t2562 VGND.t775 222.15
R2365 VGND.t986 VGND.t1750 222.15
R2366 VGND.t391 VGND.t1204 222.15
R2367 VGND.t2226 VGND.t1748 222.15
R2368 VGND.t378 VGND.t599 222.15
R2369 VGND.t876 VGND.t2167 222.15
R2370 VGND.t1101 VGND.t258 222.15
R2371 VGND.t430 VGND.t1680 222.15
R2372 VGND.t2677 VGND.t231 222.15
R2373 VGND.t2420 VGND.t2645 222.15
R2374 VGND.t386 VGND.t622 222.15
R2375 VGND.t721 VGND.t461 222.15
R2376 VGND.t1197 VGND.t586 222.15
R2377 VGND.t965 VGND.t719 222.15
R2378 VGND.t1984 VGND.t746 222.15
R2379 VGND.t428 VGND.t2430 222.15
R2380 VGND.t215 VGND.t2078 222.15
R2381 VGND.t1365 VGND.t2416 222.15
R2382 VGND.t343 VGND.t1971 222.15
R2383 VGND.t2414 VGND.t957 222.15
R2384 VGND.t1407 VGND.t2592 222.15
R2385 VGND.t996 VGND.t426 222.15
R2386 VGND.t3 VGND.t668 222.15
R2387 VGND.t424 VGND.t1277 222.15
R2388 VGND.t765 VGND.t636 222.15
R2389 VGND.t2628 VGND.t2418 222.15
R2390 VGND.t2265 VGND.t2597 222.15
R2391 VGND.t717 VGND.t701 222.15
R2392 VGND.t195 VGND.t2344 222.15
R2393 VGND.t1271 VGND.t432 222.15
R2394 VGND.t1931 VGND.t1631 222.15
R2395 VGND.t2412 VGND.t2626 222.15
R2396 VGND.t1147 VGND.t158 222.15
R2397 VGND.t725 VGND.t2529 222.15
R2398 VGND.t763 VGND.t552 222.15
R2399 VGND.t723 VGND.t671 222.15
R2400 VGND.t196 VGND.t655 222.15
R2401 VGND.t2186 VGND.t422 222.15
R2402 VGND.t1515 VGND.t1952 222.15
R2403 VGND.t2647 VGND.t2045 222.15
R2404 VGND.t1963 VGND.t572 222.15
R2405 VGND.t186 VGND.t1221 222.15
R2406 VGND.t2486 VGND.t299 222.15
R2407 VGND.t2452 VGND.t1435 222.15
R2408 VGND.t82 VGND.t2111 222.15
R2409 VGND.t1433 VGND.t787 222.15
R2410 VGND.t1 VGND.t2408 222.15
R2411 VGND.t906 VGND.t104 222.15
R2412 VGND.t619 VGND.t384 222.15
R2413 VGND.t182 VGND.t990 222.15
R2414 VGND.t669 VGND.t1296 222.15
R2415 VGND.t1383 VGND.t180 222.15
R2416 VGND.t1721 VGND.t2485 222.15
R2417 VGND.t102 VGND.t445 222.15
R2418 VGND.t1606 VGND.t1583 222.15
R2419 VGND.t955 VGND.t190 222.15
R2420 VGND.t1178 VGND.t1290 222.15
R2421 VGND.t184 VGND.t2470 222.15
R2422 VGND.t596 VGND.t1544 222.15
R2423 VGND.t2232 VGND.t2049 222.15
R2424 VGND.t2133 VGND.t554 222.15
R2425 VGND.t2047 VGND.t709 222.15
R2426 VGND.t254 VGND.t1995 222.15
R2427 VGND.t2462 VGND.t1441 222.15
R2428 VGND.t2561 VGND.t851 222.15
R2429 VGND.t1265 VGND.t1439 222.15
R2430 VGND.t388 VGND.t744 222.15
R2431 VGND.t1437 VGND.t2523 222.15
R2432 VGND.t281 VGND.t377 222.15
R2433 VGND.t693 VGND.t188 222.15
R2434 VGND.t1098 VGND.t421 222.15
R2435 VGND.t43 VGND.t685 222.15
R2436 VGND.t1305 VGND.t604 222.15
R2437 VGND.t2531 VGND.t2151 222.15
R2438 VGND.t111 VGND.t600 222.15
R2439 VGND.t1965 VGND.t2517 222.15
R2440 VGND.t1202 VGND.t1697 222.15
R2441 VGND.t2155 VGND.t459 222.15
R2442 VGND.t2278 VGND.t1779 222.15
R2443 VGND.t41 VGND.t1225 222.15
R2444 VGND.t2482 VGND.t525 222.15
R2445 VGND.t2147 VGND.t805 222.15
R2446 VGND.t846 VGND.t357 222.15
R2447 VGND.t2145 VGND.t447 222.15
R2448 VGND.t240 VGND.t531 222.15
R2449 VGND.t39 VGND.t908 222.15
R2450 VGND.t1288 VGND.t358 222.15
R2451 VGND.t37 VGND.t994 222.15
R2452 VGND.t118 VGND.t1338 222.15
R2453 VGND.t2149 VGND.t1387 222.15
R2454 VGND.t1395 VGND.t2668 222.15
R2455 VGND.t47 VGND.t882 222.15
R2456 VGND.t1617 VGND.t2249 222.15
R2457 VGND.t45 VGND.t982 222.15
R2458 VGND.t197 VGND.t172 222.15
R2459 VGND.t2143 VGND.t1375 222.15
R2460 VGND.t506 VGND.t2018 222.15
R2461 VGND.t2234 VGND.t2141 222.15
R2462 VGND.t393 VGND.t1010 222.15
R2463 VGND.t695 VGND.t1967 222.15
R2464 VGND.t405 VGND.t74 222.15
R2465 VGND.t2464 VGND.t2153 222.15
R2466 VGND.t2397 VGND.t1654 222.15
R2467 VGND.t1188 VGND.t2202 222.15
R2468 VGND.t1398 VGND.t1350 222.15
R2469 VGND.t863 VGND.t703 222.15
R2470 VGND.t1522 VGND.t2107 222.15
R2471 VGND.t1687 VGND.t949 222.15
R2472 VGND.t15 VGND.t576 222.15
R2473 VGND.t920 VGND.t1685 222.15
R2474 VGND.t827 VGND.t1023 222.15
R2475 VGND.t2535 VGND.t1186 222.15
R2476 VGND.t2042 VGND.t316 222.15
R2477 VGND.t2643 VGND.t295 222.15
R2478 VGND.t321 VGND.t56 222.15
R2479 VGND.t910 VGND.t293 222.15
R2480 VGND.t417 VGND.t17 222.15
R2481 VGND.t1227 VGND.t1184 222.15
R2482 VGND.t398 VGND.t1331 222.15
R2483 VGND.t807 VGND.t1180 222.15
R2484 VGND.t434 VGND.t760 222.15
R2485 VGND.t449 VGND.t297 222.15
R2486 VGND.t1548 VGND.t51 222.15
R2487 VGND.t1672 VGND.t1683 222.15
R2488 VGND.t1938 VGND.t1723 222.15
R2489 VGND.t795 VGND.t1190 222.15
R2490 VGND.t1609 VGND.t1286 222.15
R2491 VGND.t900 VGND.t291 222.15
R2492 VGND.t2567 VGND.t2063 222.15
R2493 VGND.t884 VGND.t289 222.15
R2494 VGND.t1144 VGND.t75 222.15
R2495 VGND.t1689 VGND.t2466 222.15
R2496 VGND.t598 VGND.t241 222.15
R2497 VGND.t1377 VGND.t865 222.15
R2498 VGND.t1444 VGND.t314 222.15
R2499 VGND.t888 VGND.t1483 222.15
R2500 VGND.t1977 VGND.t1009 222.15
R2501 VGND.t1099 VGND.t793 222.15
R2502 VGND.t239 VGND.t311 222.15
R2503 VGND.t2387 VGND.t1381 222.15
R2504 VGND.t1287 VGND.t78 222.15
R2505 VGND.t2365 VGND.t2624 222.15
R2506 VGND.t743 VGND.t1783 222.15
R2507 VGND.t1472 VGND.t2480 222.15
R2508 VGND.t1194 VGND.t2055 222.15
R2509 VGND.t1080 VGND.t1263 222.15
R2510 VGND.t2279 VGND.t354 222.15
R2511 VGND.t1069 VGND.t2618 222.15
R2512 VGND.t161 VGND.t539 222.15
R2513 VGND.t1468 VGND.t711 222.15
R2514 VGND.t420 VGND.t1702 222.15
R2515 VGND.t1450 VGND.t935 222.15
R2516 VGND.t1393 VGND.t2102 222.15
R2517 VGND.t1082 VGND.t1239 222.15
R2518 VGND.t2411 VGND.t2123 222.15
R2519 VGND.t2352 VGND.t2525 222.15
R2520 VGND.t203 VGND.t101 222.15
R2521 VGND.t1516 VGND.t689 222.15
R2522 VGND.t928 VGND.t2492 222.15
R2523 VGND.t1064 VGND.t1235 222.15
R2524 VGND.t1397 VGND.t2026 222.15
R2525 VGND.t1051 VGND.t1219 222.15
R2526 VGND.t1193 VGND.t844 222.15
R2527 VGND.t2393 VGND.t463 222.15
R2528 VGND.t759 VGND.t409 222.15
R2529 VGND.t923 VGND.t1126 222.15
R2530 VGND.t1055 VGND.t1285 222.15
R2531 VGND.n2835 VGND.n3 218.73
R2532 VGND.n133 VGND.n131 214.365
R2533 VGND.n133 VGND.n132 214.365
R2534 VGND.n123 VGND.n121 214.365
R2535 VGND.n123 VGND.n122 214.365
R2536 VGND.n141 VGND.n139 214.365
R2537 VGND.n141 VGND.n140 214.365
R2538 VGND.n601 VGND.n599 214.365
R2539 VGND.n601 VGND.n600 214.365
R2540 VGND.n591 VGND.n589 214.365
R2541 VGND.n591 VGND.n590 214.365
R2542 VGND.n609 VGND.n607 214.365
R2543 VGND.n609 VGND.n608 214.365
R2544 VGND.n971 VGND.n970 214.365
R2545 VGND.n163 VGND.n161 214.365
R2546 VGND.n163 VGND.n162 214.365
R2547 VGND.n153 VGND.n151 214.365
R2548 VGND.n153 VGND.n152 214.365
R2549 VGND.n171 VGND.n169 214.365
R2550 VGND.n171 VGND.n170 214.365
R2551 VGND.n1096 VGND.n1095 213.613
R2552 VGND.n1098 VGND.n1097 213.613
R2553 VGND.n1068 VGND.n1066 213.613
R2554 VGND.n1068 VGND.n1067 213.613
R2555 VGND.n1071 VGND.n1069 213.613
R2556 VGND.n1071 VGND.n1070 213.613
R2557 VGND.n1006 VGND.n1004 213.613
R2558 VGND.n1006 VGND.n1005 213.613
R2559 VGND.n1009 VGND.n1007 213.613
R2560 VGND.n1009 VGND.n1008 213.613
R2561 VGND.n1037 VGND.n1035 213.613
R2562 VGND.n1037 VGND.n1036 213.613
R2563 VGND.n1040 VGND.n1038 213.613
R2564 VGND.n1040 VGND.n1039 213.613
R2565 VGND.n1110 VGND.t1011 212.422
R2566 VGND.n968 VGND.n967 207.965
R2567 VGND.n985 VGND.n965 207.965
R2568 VGND.n98 VGND.n94 207.965
R2569 VGND.n98 VGND.n95 207.965
R2570 VGND.n92 VGND.n90 207.965
R2571 VGND.n92 VGND.n91 207.965
R2572 VGND.n105 VGND.n88 207.965
R2573 VGND.n105 VGND.n89 207.965
R2574 VGND.n2858 VGND.n2854 207.965
R2575 VGND.n2858 VGND.n2855 207.965
R2576 VGND.n2852 VGND.n2850 207.965
R2577 VGND.n2852 VGND.n2851 207.965
R2578 VGND.n2865 VGND.n2848 207.965
R2579 VGND.n2865 VGND.n2849 207.965
R2580 VGND.n2890 VGND.n2886 207.965
R2581 VGND.n2890 VGND.n2887 207.965
R2582 VGND.n2884 VGND.n2882 207.965
R2583 VGND.n2884 VGND.n2883 207.965
R2584 VGND.n2897 VGND.n2880 207.965
R2585 VGND.n2897 VGND.n2881 207.965
R2586 VGND.n67 VGND.n66 207.965
R2587 VGND.n79 VGND.n64 207.965
R2588 VGND.n71 VGND.n69 207.965
R2589 VGND.n984 VGND.n966 207.213
R2590 VGND.n14 VGND.n13 207.213
R2591 VGND.n18 VGND.n12 207.213
R2592 VGND.n43 VGND.n41 207.213
R2593 VGND.n43 VGND.n42 207.213
R2594 VGND.n47 VGND.n39 207.213
R2595 VGND.n47 VGND.n40 207.213
R2596 VGND.n78 VGND.n65 207.213
R2597 VGND.n2932 VGND.n2930 207.213
R2598 VGND.n2932 VGND.n2931 207.213
R2599 VGND.n2936 VGND.n2927 207.213
R2600 VGND.n2936 VGND.n2928 207.213
R2601 VGND.n2972 VGND.n2970 207.213
R2602 VGND.n2972 VGND.n2971 207.213
R2603 VGND.n2976 VGND.n2968 207.213
R2604 VGND.n2976 VGND.n2969 207.213
R2605 VGND.t1846 VGND.t1124 206.59
R2606 VGND.t1047 VGND.t1795 206.59
R2607 VGND.t1801 VGND.t1511 206.59
R2608 VGND.t1487 VGND.t1819 206.59
R2609 VGND.t1894 VGND.t1045 206.59
R2610 VGND.t2400 VGND.t1900 206.59
R2611 VGND.t1822 VGND.t2378 206.59
R2612 VGND.t1112 VGND.t1864 206.59
R2613 VGND.t1873 VGND.t1092 206.59
R2614 VGND.t2373 VGND.t1912 206.59
R2615 VGND.t1828 VGND.t1470 206.59
R2616 VGND.t1459 VGND.t1876 206.59
R2617 VGND.t1915 VGND.t1067 206.59
R2618 VGND.t2363 VGND.t1924 206.59
R2619 VGND.t1840 VGND.t1448 206.59
R2620 VGND.t1078 VGND.t1882 206.59
R2621 VGND VGND.n2653 194.419
R2622 VGND VGND.n2649 194.419
R2623 VGND VGND.n2661 194.419
R2624 VGND VGND.n2645 194.419
R2625 VGND VGND.n2669 194.419
R2626 VGND VGND.n2641 194.419
R2627 VGND VGND.n2677 194.419
R2628 VGND VGND.n2637 194.419
R2629 VGND VGND.n2685 194.419
R2630 VGND VGND.n2633 194.419
R2631 VGND VGND.n2693 194.419
R2632 VGND VGND.n2629 194.419
R2633 VGND VGND.n2701 194.419
R2634 VGND VGND.n2580 194.419
R2635 VGND VGND.n2571 194.419
R2636 VGND.n676 VGND.n675 194.391
R2637 VGND.n1287 VGND.n678 194.391
R2638 VGND.n684 VGND.n682 194.391
R2639 VGND.n722 VGND.n721 194.391
R2640 VGND.n727 VGND.n726 194.391
R2641 VGND.n732 VGND.n731 194.391
R2642 VGND.n737 VGND.n736 194.391
R2643 VGND.n742 VGND.n741 194.391
R2644 VGND.n747 VGND.n746 194.391
R2645 VGND.n752 VGND.n751 194.391
R2646 VGND.n757 VGND.n756 194.391
R2647 VGND.n762 VGND.n761 194.391
R2648 VGND.n767 VGND.n766 194.391
R2649 VGND.n772 VGND.n771 194.391
R2650 VGND.n777 VGND.n776 194.391
R2651 VGND.n1232 VGND.n787 194.391
R2652 VGND.n1225 VGND.n1224 194.391
R2653 VGND.n793 VGND.n792 194.391
R2654 VGND.n1206 VGND.n1205 194.391
R2655 VGND.n1200 VGND.n795 194.391
R2656 VGND.n1193 VGND.n1192 194.391
R2657 VGND.n801 VGND.n800 194.391
R2658 VGND.n1174 VGND.n1173 194.391
R2659 VGND.n1168 VGND.n803 194.391
R2660 VGND.n1161 VGND.n1160 194.391
R2661 VGND.n809 VGND.n808 194.391
R2662 VGND.n1142 VGND.n1141 194.391
R2663 VGND.n1136 VGND.n811 194.391
R2664 VGND.n1129 VGND.n1128 194.391
R2665 VGND.n1126 VGND.n813 194.391
R2666 VGND.n2575 VGND.n2574 194.391
R2667 VGND.n229 VGND.n228 194.391
R2668 VGND.n231 VGND.n230 194.391
R2669 VGND.n2717 VGND.n2716 194.391
R2670 VGND.n2722 VGND.n2721 194.391
R2671 VGND.n2727 VGND.n2726 194.391
R2672 VGND.n2732 VGND.n2731 194.391
R2673 VGND.n2737 VGND.n2736 194.391
R2674 VGND.n2742 VGND.n2741 194.391
R2675 VGND.n2747 VGND.n2746 194.391
R2676 VGND.n2752 VGND.n2751 194.391
R2677 VGND.n2757 VGND.n2756 194.391
R2678 VGND.n2762 VGND.n2761 194.391
R2679 VGND.n2767 VGND.n2766 194.391
R2680 VGND.n2772 VGND.n2771 194.391
R2681 VGND.n2777 VGND.n2776 194.391
R2682 VGND.n226 VGND.n225 194.391
R2683 VGND.n239 VGND.n238 194.391
R2684 VGND.n241 VGND.n240 194.391
R2685 VGND.n2511 VGND.n2510 194.391
R2686 VGND.n2506 VGND.n243 194.391
R2687 VGND.n247 VGND.n245 194.391
R2688 VGND.n2436 VGND.n2435 194.391
R2689 VGND.n2441 VGND.n2440 194.391
R2690 VGND.n2446 VGND.n2445 194.391
R2691 VGND.n2451 VGND.n2450 194.391
R2692 VGND.n2456 VGND.n2455 194.391
R2693 VGND.n2461 VGND.n2460 194.391
R2694 VGND.n2466 VGND.n2465 194.391
R2695 VGND.n2471 VGND.n2470 194.391
R2696 VGND.n2476 VGND.n2475 194.391
R2697 VGND.n2481 VGND.n2480 194.391
R2698 VGND.n2486 VGND.n2485 194.391
R2699 VGND.n179 VGND.n178 194.391
R2700 VGND.n2829 VGND.n181 194.391
R2701 VGND.n367 VGND.n365 194.391
R2702 VGND.n369 VGND.n368 194.391
R2703 VGND.n2169 VGND.n2168 194.391
R2704 VGND.n363 VGND.n362 194.391
R2705 VGND.n2195 VGND.n2194 194.391
R2706 VGND.n355 VGND.n354 194.391
R2707 VGND.n2221 VGND.n2220 194.391
R2708 VGND.n347 VGND.n346 194.391
R2709 VGND.n2247 VGND.n2246 194.391
R2710 VGND.n339 VGND.n338 194.391
R2711 VGND.n2278 VGND.n2277 194.391
R2712 VGND.n2283 VGND.n2282 194.391
R2713 VGND.n2288 VGND.n2287 194.391
R2714 VGND.n331 VGND.n330 194.391
R2715 VGND.n1420 VGND.n1419 194.391
R2716 VGND.n1426 VGND.n1425 194.391
R2717 VGND.n1423 VGND.n1422 194.391
R2718 VGND.n2156 VGND.n2155 194.391
R2719 VGND.n378 VGND.n377 194.391
R2720 VGND.n2182 VGND.n2181 194.391
R2721 VGND.n359 VGND.n358 194.391
R2722 VGND.n2208 VGND.n2207 194.391
R2723 VGND.n351 VGND.n350 194.391
R2724 VGND.n2234 VGND.n2233 194.391
R2725 VGND.n343 VGND.n342 194.391
R2726 VGND.n2260 VGND.n2259 194.391
R2727 VGND.n335 VGND.n334 194.391
R2728 VGND.n2265 VGND.n2264 194.391
R2729 VGND.n2305 VGND.n2304 194.391
R2730 VGND.n2312 VGND.n326 194.391
R2731 VGND.n637 VGND.n636 194.391
R2732 VGND.n1440 VGND.n1439 194.391
R2733 VGND.n633 VGND.n632 194.391
R2734 VGND.n1490 VGND.n1489 194.391
R2735 VGND.n1485 VGND.n1484 194.391
R2736 VGND.n1480 VGND.n1479 194.391
R2737 VGND.n1475 VGND.n1474 194.391
R2738 VGND.n1470 VGND.n1469 194.391
R2739 VGND.n1465 VGND.n1464 194.391
R2740 VGND.n1460 VGND.n1459 194.391
R2741 VGND.n1455 VGND.n1454 194.391
R2742 VGND.n1450 VGND.n1449 194.391
R2743 VGND.n1445 VGND.n1444 194.391
R2744 VGND.n392 VGND.n391 194.391
R2745 VGND.n2133 VGND.n2132 194.391
R2746 VGND.n2128 VGND.n394 194.391
R2747 VGND.n616 VGND.n615 194.391
R2748 VGND.n1502 VGND.n618 194.391
R2749 VGND.n622 VGND.n620 194.391
R2750 VGND.n624 VGND.n623 194.391
R2751 VGND.n1995 VGND.n1994 194.391
R2752 VGND.n430 VGND.n429 194.391
R2753 VGND.n2021 VGND.n2020 194.391
R2754 VGND.n422 VGND.n421 194.391
R2755 VGND.n2047 VGND.n2046 194.391
R2756 VGND.n414 VGND.n413 194.391
R2757 VGND.n2073 VGND.n2072 194.391
R2758 VGND.n406 VGND.n405 194.391
R2759 VGND.n2104 VGND.n2103 194.391
R2760 VGND.n2109 VGND.n2108 194.391
R2761 VGND.n2114 VGND.n2113 194.391
R2762 VGND.n2121 VGND.n397 194.391
R2763 VGND.n643 VGND.n642 194.391
R2764 VGND.n649 VGND.n648 194.391
R2765 VGND.n646 VGND.n645 194.391
R2766 VGND.n1982 VGND.n1981 194.391
R2767 VGND.n434 VGND.n433 194.391
R2768 VGND.n2008 VGND.n2007 194.391
R2769 VGND.n426 VGND.n425 194.391
R2770 VGND.n2034 VGND.n2033 194.391
R2771 VGND.n418 VGND.n417 194.391
R2772 VGND.n2060 VGND.n2059 194.391
R2773 VGND.n410 VGND.n409 194.391
R2774 VGND.n2086 VGND.n2085 194.391
R2775 VGND.n402 VGND.n401 194.391
R2776 VGND.n2091 VGND.n2090 194.391
R2777 VGND.n2330 VGND.n2329 194.391
R2778 VGND.n2337 VGND.n315 194.391
R2779 VGND.n659 VGND.n658 194.391
R2780 VGND.n956 VGND.n955 194.391
R2781 VGND.n951 VGND.n950 194.391
R2782 VGND.n946 VGND.n945 194.391
R2783 VGND.n941 VGND.n940 194.391
R2784 VGND.n936 VGND.n935 194.391
R2785 VGND.n931 VGND.n930 194.391
R2786 VGND.n926 VGND.n925 194.391
R2787 VGND.n921 VGND.n920 194.391
R2788 VGND.n916 VGND.n915 194.391
R2789 VGND.n911 VGND.n910 194.391
R2790 VGND.n906 VGND.n905 194.391
R2791 VGND.n901 VGND.n900 194.391
R2792 VGND.n448 VGND.n447 194.391
R2793 VGND.n1959 VGND.n1958 194.391
R2794 VGND.n1954 VGND.n450 194.391
R2795 VGND.n668 VGND.n667 194.391
R2796 VGND.n1393 VGND.n1392 194.391
R2797 VGND.n1398 VGND.n1397 194.391
R2798 VGND.n665 VGND.n664 194.391
R2799 VGND.n1821 VGND.n1820 194.391
R2800 VGND.n486 VGND.n485 194.391
R2801 VGND.n1847 VGND.n1846 194.391
R2802 VGND.n478 VGND.n477 194.391
R2803 VGND.n1873 VGND.n1872 194.391
R2804 VGND.n470 VGND.n469 194.391
R2805 VGND.n1899 VGND.n1898 194.391
R2806 VGND.n462 VGND.n461 194.391
R2807 VGND.n1930 VGND.n1929 194.391
R2808 VGND.n1935 VGND.n1934 194.391
R2809 VGND.n1940 VGND.n1939 194.391
R2810 VGND.n1947 VGND.n453 194.391
R2811 VGND.n1372 VGND.n1371 194.391
R2812 VGND.n1378 VGND.n1377 194.391
R2813 VGND.n1375 VGND.n1374 194.391
R2814 VGND.n1808 VGND.n1807 194.391
R2815 VGND.n490 VGND.n489 194.391
R2816 VGND.n1834 VGND.n1833 194.391
R2817 VGND.n482 VGND.n481 194.391
R2818 VGND.n1860 VGND.n1859 194.391
R2819 VGND.n474 VGND.n473 194.391
R2820 VGND.n1886 VGND.n1885 194.391
R2821 VGND.n466 VGND.n465 194.391
R2822 VGND.n1912 VGND.n1911 194.391
R2823 VGND.n458 VGND.n457 194.391
R2824 VGND.n1917 VGND.n1916 194.391
R2825 VGND.n2355 VGND.n2354 194.391
R2826 VGND.n2362 VGND.n303 194.391
R2827 VGND.n1304 VGND.n1303 194.391
R2828 VGND.n1310 VGND.n1309 194.391
R2829 VGND.n1307 VGND.n1306 194.391
R2830 VGND.n1360 VGND.n1359 194.391
R2831 VGND.n1355 VGND.n1354 194.391
R2832 VGND.n1350 VGND.n1349 194.391
R2833 VGND.n1345 VGND.n1344 194.391
R2834 VGND.n1340 VGND.n1339 194.391
R2835 VGND.n1335 VGND.n1334 194.391
R2836 VGND.n1330 VGND.n1329 194.391
R2837 VGND.n1325 VGND.n1324 194.391
R2838 VGND.n1320 VGND.n1319 194.391
R2839 VGND.n1315 VGND.n1314 194.391
R2840 VGND.n504 VGND.n503 194.391
R2841 VGND.n1785 VGND.n1784 194.391
R2842 VGND.n1780 VGND.n506 194.391
R2843 VGND.n572 VGND.n571 194.391
R2844 VGND.n1515 VGND.n1514 194.391
R2845 VGND.n1520 VGND.n1519 194.391
R2846 VGND.n576 VGND.n575 194.391
R2847 VGND.n1647 VGND.n1646 194.391
R2848 VGND.n542 VGND.n541 194.391
R2849 VGND.n1673 VGND.n1672 194.391
R2850 VGND.n534 VGND.n533 194.391
R2851 VGND.n1699 VGND.n1698 194.391
R2852 VGND.n526 VGND.n525 194.391
R2853 VGND.n1725 VGND.n1724 194.391
R2854 VGND.n518 VGND.n517 194.391
R2855 VGND.n1756 VGND.n1755 194.391
R2856 VGND.n1761 VGND.n1760 194.391
R2857 VGND.n1766 VGND.n1765 194.391
R2858 VGND.n1773 VGND.n509 194.391
R2859 VGND.n568 VGND.n567 194.391
R2860 VGND.n1535 VGND.n1534 194.391
R2861 VGND.n565 VGND.n564 194.391
R2862 VGND.n1634 VGND.n1633 194.391
R2863 VGND.n546 VGND.n545 194.391
R2864 VGND.n1660 VGND.n1659 194.391
R2865 VGND.n538 VGND.n537 194.391
R2866 VGND.n1686 VGND.n1685 194.391
R2867 VGND.n530 VGND.n529 194.391
R2868 VGND.n1712 VGND.n1711 194.391
R2869 VGND.n522 VGND.n521 194.391
R2870 VGND.n1738 VGND.n1737 194.391
R2871 VGND.n514 VGND.n513 194.391
R2872 VGND.n1743 VGND.n1742 194.391
R2873 VGND.n2380 VGND.n2379 194.391
R2874 VGND.n2387 VGND.n290 194.391
R2875 VGND.n671 VGND.n670 194.391
R2876 VGND.n673 VGND.n672 194.391
R2877 VGND.n1548 VGND.n1547 194.391
R2878 VGND.n1553 VGND.n1552 194.391
R2879 VGND.n1558 VGND.n1557 194.391
R2880 VGND.n1563 VGND.n1562 194.391
R2881 VGND.n1568 VGND.n1567 194.391
R2882 VGND.n1573 VGND.n1572 194.391
R2883 VGND.n1578 VGND.n1577 194.391
R2884 VGND.n1583 VGND.n1582 194.391
R2885 VGND.n1588 VGND.n1587 194.391
R2886 VGND.n1593 VGND.n1592 194.391
R2887 VGND.n1598 VGND.n1597 194.391
R2888 VGND.n560 VGND.n559 194.391
R2889 VGND.n1611 VGND.n1610 194.391
R2890 VGND.n1606 VGND.n1602 194.391
R2891 VGND.n825 VGND.n824 194.391
R2892 VGND.n832 VGND.n831 194.391
R2893 VGND.n837 VGND.n836 194.391
R2894 VGND.n829 VGND.n828 194.391
R2895 VGND.n887 VGND.n886 194.391
R2896 VGND.n882 VGND.n881 194.391
R2897 VGND.n877 VGND.n876 194.391
R2898 VGND.n872 VGND.n871 194.391
R2899 VGND.n867 VGND.n866 194.391
R2900 VGND.n862 VGND.n861 194.391
R2901 VGND.n857 VGND.n856 194.391
R2902 VGND.n852 VGND.n851 194.391
R2903 VGND.n847 VGND.n846 194.391
R2904 VGND.n842 VGND.n841 194.391
R2905 VGND.n2400 VGND.n2399 194.391
R2906 VGND.n2407 VGND.n278 194.391
R2907 VGND.n815 VGND.n814 194.391
R2908 VGND.n718 VGND.n717 194.391
R2909 VGND.n2565 VGND.n2564 161.308
R2910 VGND.n2562 VGND.n2561 161.308
R2911 VGND.n2559 VGND.n2558 161.308
R2912 VGND.n2556 VGND.n2555 161.308
R2913 VGND.n2553 VGND.n2552 161.308
R2914 VGND.n2550 VGND.n2549 161.308
R2915 VGND.n2547 VGND.n2546 161.308
R2916 VGND.n2544 VGND.n2543 161.308
R2917 VGND.n2541 VGND.n2540 161.308
R2918 VGND.n2538 VGND.n2537 161.308
R2919 VGND.n2535 VGND.n2534 161.308
R2920 VGND.n2532 VGND.n2531 161.308
R2921 VGND.n2529 VGND.n2528 161.308
R2922 VGND.n2526 VGND.n2525 161.308
R2923 VGND.n2523 VGND.n2522 161.308
R2924 VGND.n2564 VGND.t2696 159.978
R2925 VGND.n2561 VGND.t2700 159.978
R2926 VGND.n2558 VGND.t2694 159.978
R2927 VGND.n2555 VGND.t2690 159.978
R2928 VGND.n2552 VGND.t2695 159.978
R2929 VGND.n2549 VGND.t2703 159.978
R2930 VGND.n2546 VGND.t2699 159.978
R2931 VGND.n2543 VGND.t2692 159.978
R2932 VGND.n2540 VGND.t2689 159.978
R2933 VGND.n2537 VGND.t2691 159.978
R2934 VGND.n2534 VGND.t2702 159.978
R2935 VGND.n2531 VGND.t2693 159.978
R2936 VGND.n2528 VGND.t2701 159.978
R2937 VGND.n2525 VGND.t2698 159.978
R2938 VGND.n2522 VGND.t2704 159.978
R2939 VGND.n996 VGND.t2087 159.315
R2940 VGND.n2918 VGND.t1708 159.315
R2941 VGND.n1088 VGND.t1169 158.361
R2942 VGND.n2988 VGND.t319 158.361
R2943 VGND.n898 VGND.t2085 157.291
R2944 VGND.n2916 VGND.t1706 157.291
R2945 VGND.n582 VGND.t756 156.915
R2946 VGND.n2878 VGND.t2294 156.915
R2947 VGND.n582 VGND.t754 156.915
R2948 VGND.n2878 VGND.t2295 156.915
R2949 VGND.n584 VGND.t611 154.131
R2950 VGND.n584 VGND.t1254 154.131
R2951 VGND.n996 VGND.t1970 154.131
R2952 VGND.n999 VGND.t981 154.131
R2953 VGND.n2902 VGND.t61 154.131
R2954 VGND.n2902 VGND.t60 154.131
R2955 VGND.n2918 VGND.t2674 154.131
R2956 VGND.n2948 VGND.t1329 154.131
R2957 VGND.n118 VGND.t753 153.631
R2958 VGND.n1026 VGND.t1709 153.631
R2959 VGND.n1057 VGND.t2114 153.631
R2960 VGND.n2870 VGND.t2292 153.631
R2961 VGND.n2950 VGND.t2113 153.631
R2962 VGND.n2955 VGND.t481 153.631
R2963 VGND.n1027 VGND.t1253 152.757
R2964 VGND.n2951 VGND.t1283 152.757
R2965 VGND.n991 VGND.t750 152.381
R2966 VGND.n61 VGND.t2299 152.381
R2967 VGND.n961 VGND.n960 152.174
R2968 VGND.n149 VGND.t755 150.922
R2969 VGND.n149 VGND.t748 150.922
R2970 VGND.n86 VGND.t2302 150.922
R2971 VGND.n86 VGND.t2297 150.922
R2972 VGND.n116 VGND.t2173 150.922
R2973 VGND.n581 VGND.t501 150.922
R2974 VGND.n148 VGND.t514 150.922
R2975 VGND.n85 VGND.t2604 150.922
R2976 VGND.n2845 VGND.t2281 150.922
R2977 VGND.n2877 VGND.t1955 150.922
R2978 VGND.n116 VGND.t927 150.922
R2979 VGND.n581 VGND.t2095 150.922
R2980 VGND.n148 VGND.t1292 150.922
R2981 VGND.n85 VGND.t1935 150.922
R2982 VGND.n2845 VGND.t217 150.922
R2983 VGND.n2877 VGND.t1621 150.922
R2984 VGND.n117 VGND.t752 147.411
R2985 VGND.n1058 VGND.t230 147.411
R2986 VGND.n2869 VGND.t2301 147.411
R2987 VGND.n2956 VGND.t2289 147.411
R2988 VGND.n899 VGND.t1020 146.964
R2989 VGND.n84 VGND.t1310 146.964
R2990 VGND.n2564 VGND.t1830 143.911
R2991 VGND.n2561 VGND.t1905 143.911
R2992 VGND.n2558 VGND.t1812 143.911
R2993 VGND.n2555 VGND.t1854 143.911
R2994 VGND.n2552 VGND.t1926 143.911
R2995 VGND.n2549 VGND.t1833 143.911
R2996 VGND.n2546 VGND.t1806 143.911
R2997 VGND.n2543 VGND.t1848 143.911
R2998 VGND.n2540 VGND.t1860 143.911
R2999 VGND.n2537 VGND.t1788 143.911
R3000 VGND.n2534 VGND.t1884 143.911
R3001 VGND.n2531 VGND.t1815 143.911
R3002 VGND.n2528 VGND.t1887 143.911
R3003 VGND.n2525 VGND.t1917 143.911
R3004 VGND.n2522 VGND.t1857 143.911
R3005 VGND.n1513 VGND.n578 143.478
R3006 VGND VGND.t144 142.089
R3007 VGND.n822 VGND.t1845 119.309
R3008 VGND.n785 VGND.t1881 119.309
R3009 VGND.n2586 VGND.t1878 119.309
R3010 VGND.n2583 VGND.t1842 119.309
R3011 VGND.n2569 VGND.t1791 119.309
R3012 VGND.n2582 VGND.t1797 119.309
R3013 VGND.n2621 VGND.t1803 119.309
R3014 VGND.n2618 VGND.t1890 119.309
R3015 VGND.n2615 VGND.t1896 119.309
R3016 VGND.n2612 VGND.t1809 119.309
R3017 VGND.n2609 VGND.t1851 119.309
R3018 VGND.n2606 VGND.t1866 119.309
R3019 VGND.n2603 VGND.t1902 119.309
R3020 VGND.n2600 VGND.t1824 119.309
R3021 VGND.n2597 VGND.t1869 119.309
R3022 VGND.n2594 VGND.t1908 119.309
R3023 VGND.n2591 VGND.t1920 119.309
R3024 VGND.n2588 VGND.t1836 119.309
R3025 VGND.n819 VGND.t1794 119.309
R3026 VGND.n816 VGND.t1800 119.309
R3027 VGND.n1137 VGND.t1818 119.309
R3028 VGND.n807 VGND.t1893 119.309
R3029 VGND.n805 VGND.t1899 119.309
R3030 VGND.n1152 VGND.t1821 119.309
R3031 VGND.n1169 VGND.t1863 119.309
R3032 VGND.n799 VGND.t1872 119.309
R3033 VGND.n797 VGND.t1911 119.309
R3034 VGND.n1184 VGND.t1827 119.309
R3035 VGND.n1201 VGND.t1875 119.309
R3036 VGND.n791 VGND.t1914 119.309
R3037 VGND.n789 VGND.t1923 119.309
R3038 VGND.n1216 VGND.t1839 119.309
R3039 VGND.n6 VGND.n4 117.001
R3040 VGND.t544 VGND.n6 117.001
R3041 VGND.n5 VGND.n3 117.001
R3042 VGND.t544 VGND.n5 117.001
R3043 VGND.t1053 VGND.t1846 112.356
R3044 VGND.t1294 VGND.t1519 112.356
R3045 VGND.t1795 VGND.t1513 112.356
R3046 VGND.t1136 VGND.t257 112.356
R3047 VGND.t1128 VGND.t1801 112.356
R3048 VGND.t1753 VGND.t1121 112.356
R3049 VGND.t1819 VGND.t1106 112.356
R3050 VGND.t2396 VGND.t255 112.356
R3051 VGND.t1041 VGND.t1894 112.356
R3052 VGND.t2028 VGND.t1507 112.356
R3053 VGND.t1900 VGND.t1491 112.356
R3054 VGND.t1109 VGND.t1182 112.356
R3055 VGND.t1478 VGND.t1822 112.356
R3056 VGND.t1179 VGND.t1044 112.356
R3057 VGND.t1864 VGND.t2402 112.356
R3058 VGND.t2386 VGND.t1604 112.356
R3059 VGND.t2380 VGND.t1873 112.356
R3060 VGND.t1167 VGND.t1480 112.356
R3061 VGND.t1912 VGND.t1493 112.356
R3062 VGND.t1110 VGND.t867 112.356
R3063 VGND.t1094 VGND.t1828 112.356
R3064 VGND.t1330 VGND.t2383 112.356
R3065 VGND.t1876 VGND.t1085 112.356
R3066 VGND.t2371 VGND.t774 112.356
R3067 VGND.t1474 VGND.t1915 112.356
R3068 VGND.t119 VGND.t1467 112.356
R3069 VGND.t1924 VGND.t1462 112.356
R3070 VGND.t1087 VGND.t2488 112.356
R3071 VGND.t1137 VGND.t1840 112.356
R3072 VGND.t1635 VGND.t1066 112.356
R3073 VGND.t1882 VGND.t2367 112.356
R3074 VGND.t1464 VGND.t2636 112.356
R3075 VGND.t1011 VGND.t1021 92.9349
R3076 VGND.t1021 VGND.t1018 92.9349
R3077 VGND.t1018 VGND.t1022 92.9349
R3078 VGND.t1022 VGND.t2306 92.9349
R3079 VGND.t2306 VGND.t2315 92.9349
R3080 VGND.t2315 VGND.t822 92.9349
R3081 VGND.t822 VGND.t165 92.9349
R3082 VGND VGND.n578 80.9529
R3083 VGND.n1292 VGND 75.2331
R3084 VGND VGND.n578 75.1009
R3085 VGND.t165 VGND 70.8076
R3086 VGND.n147 VGND 58.8055
R3087 VGND.n1507 VGND 58.8055
R3088 VGND.n1509 VGND 58.8055
R3089 VGND.n1511 VGND 58.8055
R3090 VGND.n2834 VGND 58.8055
R3091 VGND.n2837 VGND.n2836 53.1823
R3092 VGND.n2838 VGND.n2837 53.1823
R3093 VGND.n3020 VGND.n3019 53.1823
R3094 VGND.n3019 VGND.n3018 53.1823
R3095 VGND.t1019 VGND.t2304 50.5752
R3096 VGND.t1016 VGND.t2313 50.5752
R3097 VGND.t1014 VGND.t122 50.5752
R3098 VGND.t1012 VGND.t1355 50.5752
R3099 VGND.t1317 VGND.t146 50.5752
R3100 VGND.t1313 VGND.t1535 50.5752
R3101 VGND.t1307 VGND.t131 50.5752
R3102 VGND.t1309 VGND.t1557 50.5752
R3103 VGND VGND.n14 43.2063
R3104 VGND VGND.n43 43.2063
R3105 VGND VGND.n2932 43.2063
R3106 VGND VGND.n2972 43.2063
R3107 VGND.n2836 VGND.n2835 40.6593
R3108 VGND.n675 VGND.t2385 34.8005
R3109 VGND.n675 VGND.t1484 34.8005
R3110 VGND.n678 VGND.t1482 34.8005
R3111 VGND.n678 VGND.t1100 34.8005
R3112 VGND.n682 VGND.t1097 34.8005
R3113 VGND.n682 VGND.t2388 34.8005
R3114 VGND.n721 VGND.t1075 34.8005
R3115 VGND.n721 VGND.t2366 34.8005
R3116 VGND.n726 VGND.t1477 34.8005
R3117 VGND.n726 VGND.t1473 34.8005
R3118 VGND.n731 VGND.t1466 34.8005
R3119 VGND.n731 VGND.t1081 34.8005
R3120 VGND.n736 VGND.t1447 34.8005
R3121 VGND.n736 VGND.t1070 34.8005
R3122 VGND.n741 VGND.t2370 34.8005
R3123 VGND.n741 VGND.t1469 34.8005
R3124 VGND.n746 VGND.t2349 34.8005
R3125 VGND.n746 VGND.t1451 34.8005
R3126 VGND.n751 VGND.t1140 34.8005
R3127 VGND.n751 VGND.t1083 34.8005
R3128 VGND.n756 VGND.t1063 34.8005
R3129 VGND.n756 VGND.t2353 34.8005
R3130 VGND.n761 VGND.t1050 34.8005
R3131 VGND.n761 VGND.t1517 34.8005
R3132 VGND.n766 VGND.t1501 34.8005
R3133 VGND.n766 VGND.t1065 34.8005
R3134 VGND.n771 VGND.t1123 34.8005
R3135 VGND.n771 VGND.t1052 34.8005
R3136 VGND.n776 VGND.t2399 34.8005
R3137 VGND.n776 VGND.t2394 34.8005
R3138 VGND.n787 VGND.t1079 34.8005
R3139 VGND.n787 VGND.t2368 34.8005
R3140 VGND.n1224 VGND.t1449 34.8005
R3141 VGND.n1224 VGND.t1138 34.8005
R3142 VGND.n792 VGND.t2364 34.8005
R3143 VGND.n792 VGND.t1463 34.8005
R3144 VGND.n1205 VGND.t1068 34.8005
R3145 VGND.n1205 VGND.t1475 34.8005
R3146 VGND.n795 VGND.t1460 34.8005
R3147 VGND.n795 VGND.t1086 34.8005
R3148 VGND.n1192 VGND.t1471 34.8005
R3149 VGND.n1192 VGND.t1095 34.8005
R3150 VGND.n800 VGND.t2374 34.8005
R3151 VGND.n800 VGND.t1494 34.8005
R3152 VGND.n1173 VGND.t1093 34.8005
R3153 VGND.n1173 VGND.t2381 34.8005
R3154 VGND.n803 VGND.t1113 34.8005
R3155 VGND.n803 VGND.t2403 34.8005
R3156 VGND.n1160 VGND.t2379 34.8005
R3157 VGND.n1160 VGND.t1479 34.8005
R3158 VGND.n808 VGND.t2401 34.8005
R3159 VGND.n808 VGND.t1492 34.8005
R3160 VGND.n1141 VGND.t1046 34.8005
R3161 VGND.n1141 VGND.t1042 34.8005
R3162 VGND.n811 VGND.t1488 34.8005
R3163 VGND.n811 VGND.t1107 34.8005
R3164 VGND.n1128 VGND.t1512 34.8005
R3165 VGND.n1128 VGND.t1129 34.8005
R3166 VGND.n813 VGND.t1048 34.8005
R3167 VGND.n813 VGND.t1514 34.8005
R3168 VGND.n2574 VGND.t1073 34.8005
R3169 VGND.n2574 VGND.t2362 34.8005
R3170 VGND.n2653 VGND.t2390 34.8005
R3171 VGND.n2653 VGND.t1490 34.8005
R3172 VGND.n2649 VGND.t1091 34.8005
R3173 VGND.n2649 VGND.t1089 34.8005
R3174 VGND.n2661 VGND.t1486 34.8005
R3175 VGND.n2661 VGND.t1105 34.8005
R3176 VGND.n2645 VGND.t2376 34.8005
R3177 VGND.n2645 VGND.t1117 34.8005
R3178 VGND.n2669 VGND.t1103 34.8005
R3179 VGND.n2669 VGND.t2392 34.8005
R3180 VGND.n2641 VGND.t1115 34.8005
R3181 VGND.n2641 VGND.t1040 34.8005
R3182 VGND.n2677 VGND.t1499 34.8005
R3183 VGND.n2677 VGND.t1135 34.8005
R3184 VGND.n2637 VGND.t2405 34.8005
R3185 VGND.n2637 VGND.t1505 34.8005
R3186 VGND.n2685 VGND.t1061 34.8005
R3187 VGND.n2685 VGND.t2351 34.8005
R3188 VGND.n2633 VGND.t1503 34.8005
R3189 VGND.n2633 VGND.t1119 34.8005
R3190 VGND.n2693 VGND.t2347 34.8005
R3191 VGND.n2693 VGND.t1133 34.8005
R3192 VGND.n2629 VGND.t2358 34.8005
R3193 VGND.n2629 VGND.t2355 34.8005
R3194 VGND.n2701 VGND.t1131 34.8005
R3195 VGND.n2701 VGND.t1057 34.8005
R3196 VGND.n2580 VGND.t1456 34.8005
R3197 VGND.n2580 VGND.t1077 34.8005
R3198 VGND.n2571 VGND.t2360 34.8005
R3199 VGND.n2571 VGND.t1458 34.8005
R3200 VGND.n228 VGND.t1832 34.8005
R3201 VGND.n228 VGND.t1244 34.8005
R3202 VGND.n230 VGND.t1718 34.8005
R3203 VGND.n230 VGND.t1755 34.8005
R3204 VGND.n2716 VGND.t110 34.8005
R3205 VGND.n2716 VGND.t1252 34.8005
R3206 VGND.n2721 VGND.t2427 34.8005
R3207 VGND.n2721 VGND.t1250 34.8005
R3208 VGND.n2726 VGND.t1983 34.8005
R3209 VGND.n2726 VGND.t1242 34.8005
R3210 VGND.n2731 VGND.t524 34.8005
R3211 VGND.n2731 VGND.t1034 34.8005
R3212 VGND.n2736 VGND.t331 34.8005
R3213 VGND.n2736 VGND.t1032 34.8005
R3214 VGND.n2741 VGND.t530 34.8005
R3215 VGND.n2741 VGND.t1761 34.8005
R3216 VGND.n2746 VGND.t773 34.8005
R3217 VGND.n2746 VGND.t1759 34.8005
R3218 VGND.n2751 VGND.t1337 34.8005
R3219 VGND.n2751 VGND.t1036 34.8005
R3220 VGND.n2756 VGND.t2666 34.8005
R3221 VGND.n2756 VGND.t1248 34.8005
R3222 VGND.n2761 VGND.t2132 34.8005
R3223 VGND.n2761 VGND.t1246 34.8005
R3224 VGND.n2766 VGND.t2510 34.8005
R3225 VGND.n2766 VGND.t1030 34.8005
R3226 VGND.n2771 VGND.t2017 34.8005
R3227 VGND.n2771 VGND.t1028 34.8005
R3228 VGND.n2776 VGND.t1948 34.8005
R3229 VGND.n2776 VGND.t1026 34.8005
R3230 VGND.n225 VGND.t654 34.8005
R3231 VGND.n225 VGND.t1757 34.8005
R3232 VGND.n238 VGND.t1907 34.8005
R3233 VGND.n238 VGND.t269 34.8005
R3234 VGND.n240 VGND.t1348 34.8005
R3235 VGND.n240 VGND.t2556 34.8005
R3236 VGND.n2510 VGND.t304 34.8005
R3237 VGND.n2510 VGND.t1323 34.8005
R3238 VGND.n243 VGND.t81 34.8005
R3239 VGND.n243 VGND.t1321 34.8005
R3240 VGND.n245 VGND.t2407 34.8005
R3241 VGND.n245 VGND.t2243 34.8005
R3242 VGND.n2435 VGND.t2274 34.8005
R3243 VGND.n2435 VGND.t2552 34.8005
R3244 VGND.n2440 VGND.t340 34.8005
R3245 VGND.n2440 VGND.t2550 34.8005
R3246 VGND.n2445 VGND.t416 34.8005
R3247 VGND.n2445 VGND.t2241 34.8005
R3248 VGND.n2450 VGND.t742 34.8005
R3249 VGND.n2450 VGND.t2239 34.8005
R3250 VGND.n2455 VGND.t202 34.8005
R3251 VGND.n2455 VGND.t2554 34.8005
R3252 VGND.n2460 VGND.t1546 34.8005
R3253 VGND.n2460 VGND.t273 34.8005
R3254 VGND.n2465 VGND.t2341 34.8005
R3255 VGND.n2465 VGND.t271 34.8005
R3256 VGND.n2470 VGND.t1997 34.8005
R3257 VGND.n2470 VGND.t2548 34.8005
R3258 VGND.n2475 VGND.t2566 34.8005
R3259 VGND.n2475 VGND.t2546 34.8005
R3260 VGND.n2480 VGND.t390 34.8005
R3261 VGND.n2480 VGND.t1325 34.8005
R3262 VGND.n2485 VGND.t411 34.8005
R3263 VGND.n2485 VGND.t2237 34.8005
R3264 VGND.n178 VGND.t1814 34.8005
R3265 VGND.n178 VGND.t855 34.8005
R3266 VGND.n181 VGND.t609 34.8005
R3267 VGND.n181 VGND.t1160 34.8005
R3268 VGND.n365 VGND.t308 34.8005
R3269 VGND.n365 VGND.t283 34.8005
R3270 VGND.n368 VGND.t1694 34.8005
R3271 VGND.n368 VGND.t861 34.8005
R3272 VGND.n2168 VGND.t1728 34.8005
R3273 VGND.n2168 VGND.t853 34.8005
R3274 VGND.n362 VGND.t2052 34.8005
R3275 VGND.n362 VGND.t2073 34.8005
R3276 VGND.n2194 VGND.t1301 34.8005
R3277 VGND.n2194 VGND.t2071 34.8005
R3278 VGND.n354 VGND.t536 34.8005
R3279 VGND.n354 VGND.t1166 34.8005
R3280 VGND.n2220 VGND.t363 34.8005
R3281 VGND.n2220 VGND.t1164 34.8005
R3282 VGND.n346 VGND.t1343 34.8005
R3283 VGND.n346 VGND.t2075 34.8005
R3284 VGND.n2246 VGND.t2119 34.8005
R3285 VGND.n2246 VGND.t859 34.8005
R3286 VGND.n338 VGND.t2038 34.8005
R3287 VGND.n338 VGND.t857 34.8005
R3288 VGND.n2277 VGND.t176 34.8005
R3289 VGND.n2277 VGND.t2069 34.8005
R3290 VGND.n2282 VGND.t2023 34.8005
R3291 VGND.n2282 VGND.t287 34.8005
R3292 VGND.n2287 VGND.t397 34.8005
R3293 VGND.n2287 VGND.t285 34.8005
R3294 VGND.n330 VGND.t661 34.8005
R3295 VGND.n330 VGND.t1162 34.8005
R3296 VGND.n1419 VGND.t1856 34.8005
R3297 VGND.n1419 VGND.t479 34.8005
R3298 VGND.n1425 VGND.t219 34.8005
R3299 VGND.n1425 VGND.t2034 34.8005
R3300 VGND.n1422 VGND.t633 34.8005
R3301 VGND.n1422 VGND.t2544 34.8005
R3302 VGND.n2155 VGND.t590 34.8005
R3303 VGND.n2155 VGND.t2542 34.8005
R3304 VGND.n377 VGND.t836 34.8005
R3305 VGND.n377 VGND.t477 34.8005
R3306 VGND.n2181 VGND.t227 34.8005
R3307 VGND.n2181 VGND.t2030 34.8005
R3308 VGND.n358 VGND.t351 34.8005
R3309 VGND.n358 VGND.t571 34.8005
R3310 VGND.n2207 VGND.t370 34.8005
R3311 VGND.n2207 VGND.t475 34.8005
R3312 VGND.n350 VGND.t11 34.8005
R3313 VGND.n350 VGND.t473 34.8005
R3314 VGND.n2233 VGND.t872 34.8005
R3315 VGND.n2233 VGND.t2032 34.8005
R3316 VGND.n342 VGND.t2262 34.8005
R3317 VGND.n342 VGND.t2540 34.8005
R3318 VGND.n2259 VGND.t98 34.8005
R3319 VGND.n2259 VGND.t2538 34.8005
R3320 VGND.n334 VGND.t1423 34.8005
R3321 VGND.n334 VGND.t569 34.8005
R3322 VGND.n2264 VGND.t115 34.8005
R3323 VGND.n2264 VGND.t567 34.8005
R3324 VGND.n2304 VGND.t549 34.8005
R3325 VGND.n2304 VGND.t565 34.8005
R3326 VGND.n326 VGND.t249 34.8005
R3327 VGND.n326 VGND.t471 34.8005
R3328 VGND.n636 VGND.t1928 34.8005
R3329 VGND.n636 VGND.t1651 34.8005
R3330 VGND.n1439 VGND.t1962 34.8005
R3331 VGND.n1439 VGND.t2256 34.8005
R3332 VGND.n632 VGND.t2093 34.8005
R3333 VGND.n632 VGND.t1930 34.8005
R3334 VGND.n1489 VGND.t1699 34.8005
R3335 VGND.n1489 VGND.t1601 34.8005
R3336 VGND.n1484 VGND.t1778 34.8005
R3337 VGND.n1484 VGND.t1649 34.8005
R3338 VGND.n1479 VGND.t618 34.8005
R3339 VGND.n1479 VGND.t2252 34.8005
R3340 VGND.n1474 VGND.t327 34.8005
R3341 VGND.n1474 VGND.t1643 34.8005
R3342 VGND.n1469 VGND.t543 34.8005
R3343 VGND.n1469 VGND.t1647 34.8005
R3344 VGND.n1464 VGND.t1582 34.8005
R3345 VGND.n1464 VGND.t1645 34.8005
R3346 VGND.n1459 VGND.t1177 34.8005
R3347 VGND.n1459 VGND.t2254 34.8005
R3348 VGND.n1454 VGND.t1541 34.8005
R3349 VGND.n1454 VGND.t1599 34.8005
R3350 VGND.n1449 VGND.t562 34.8005
R3351 VGND.n1449 VGND.t1653 34.8005
R3352 VGND.n1444 VGND.t2000 34.8005
R3353 VGND.n1444 VGND.t1641 34.8005
R3354 VGND.n391 VGND.t2560 34.8005
R3355 VGND.n391 VGND.t1639 34.8005
R3356 VGND.n2132 VGND.t20 34.8005
R3357 VGND.n2132 VGND.t1637 34.8005
R3358 VGND.n394 VGND.t404 34.8005
R3359 VGND.n394 VGND.t2258 34.8005
R3360 VGND.n615 VGND.t1835 34.8005
R3361 VGND.n615 VGND.t2183 34.8005
R3362 VGND.n618 VGND.t1716 34.8005
R3363 VGND.n618 VGND.t419 34.8005
R3364 VGND.n620 VGND.t108 34.8005
R3365 VGND.n620 VGND.t2327 34.8005
R3366 VGND.n623 VGND.t2424 34.8005
R3367 VGND.n623 VGND.t2325 34.8005
R3368 VGND.n1994 VGND.t1981 34.8005
R3369 VGND.n1994 VGND.t2181 34.8005
R3370 VGND.n429 VGND.t522 34.8005
R3371 VGND.n429 VGND.t2337 34.8005
R3372 VGND.n2020 VGND.t329 34.8005
R3373 VGND.n2020 VGND.t2335 34.8005
R3374 VGND.n421 VGND.t376 34.8005
R3375 VGND.n421 VGND.t2179 34.8005
R3376 VGND.n2046 VGND.t771 34.8005
R3377 VGND.n2046 VGND.t2177 34.8005
R3378 VGND.n413 VGND.t1335 34.8005
R3379 VGND.n413 VGND.t498 34.8005
R3380 VGND.n2072 VGND.t2269 34.8005
R3381 VGND.n2072 VGND.t2323 34.8005
R3382 VGND.n405 VGND.t2130 34.8005
R3383 VGND.n405 VGND.t2321 34.8005
R3384 VGND.n2103 VGND.t2507 34.8005
R3385 VGND.n2103 VGND.t2333 34.8005
R3386 VGND.n2108 VGND.t2015 34.8005
R3387 VGND.n2108 VGND.t2331 34.8005
R3388 VGND.n2113 VGND.t1945 34.8005
R3389 VGND.n2113 VGND.t2329 34.8005
R3390 VGND.n397 VGND.t652 34.8005
R3391 VGND.n397 VGND.t2175 34.8005
R3392 VGND.n642 VGND.t1808 34.8005
R3393 VGND.n642 VGND.t1773 34.8005
R3394 VGND.n648 VGND.t1976 34.8005
R3395 VGND.n648 VGND.t1763 34.8005
R3396 VGND.n645 VGND.t310 34.8005
R3397 VGND.n645 VGND.t1593 34.8005
R3398 VGND.n1981 VGND.t1692 34.8005
R3399 VGND.n1981 VGND.t1591 34.8005
R3400 VGND.n433 VGND.t1730 34.8005
R3401 VGND.n433 VGND.t1771 34.8005
R3402 VGND.n2007 VGND.t2054 34.8005
R3403 VGND.n2007 VGND.t647 34.8005
R3404 VGND.n425 VGND.t1303 34.8005
R3405 VGND.n425 VGND.t645 34.8005
R3406 VGND.n2033 VGND.t538 34.8005
R3407 VGND.n2033 VGND.t1769 34.8005
R3408 VGND.n417 VGND.t1701 34.8005
R3409 VGND.n417 VGND.t1767 34.8005
R3410 VGND.n2059 VGND.t2101 34.8005
R3411 VGND.n2059 VGND.t649 34.8005
R3412 VGND.n409 VGND.t2121 34.8005
R3413 VGND.n409 VGND.t1589 34.8005
R3414 VGND.n2085 VGND.t2040 34.8005
R3415 VGND.n2085 VGND.t1587 34.8005
R3416 VGND.n401 VGND.t178 34.8005
R3417 VGND.n401 VGND.t643 34.8005
R3418 VGND.n2090 VGND.t2025 34.8005
R3419 VGND.n2090 VGND.t1597 34.8005
R3420 VGND.n2329 VGND.t842 34.8005
R3421 VGND.n2329 VGND.t1595 34.8005
R3422 VGND.n315 VGND.t663 34.8005
R3423 VGND.n315 VGND.t1765 34.8005
R3424 VGND.n658 VGND.t1850 34.8005
R3425 VGND.n658 VGND.t261 34.8005
R3426 VGND.n955 VGND.t221 34.8005
R3427 VGND.n955 VGND.t2062 34.8005
R3428 VGND.n950 VGND.t635 34.8005
R3429 VGND.n950 VGND.t2276 34.8005
R3430 VGND.n945 VGND.t588 34.8005
R3431 VGND.n945 VGND.t267 34.8005
R3432 VGND.n940 VGND.t838 34.8005
R3433 VGND.n940 VGND.t1994 34.8005
R3434 VGND.n935 VGND.t229 34.8005
R3435 VGND.n935 VGND.t1153 34.8005
R3436 VGND.n930 VGND.t353 34.8005
R3437 VGND.n930 VGND.t1151 34.8005
R3438 VGND.n925 VGND.t372 34.8005
R3439 VGND.n925 VGND.t1992 34.8005
R3440 VGND.n920 VGND.t767 34.8005
R3441 VGND.n920 VGND.t1990 34.8005
R3442 VGND.n915 VGND.t874 34.8005
R3443 VGND.n915 VGND.t1155 34.8005
R3444 VGND.n910 VGND.t2264 34.8005
R3445 VGND.n910 VGND.t265 34.8005
R3446 VGND.n905 VGND.t100 34.8005
R3447 VGND.n905 VGND.t263 34.8005
R3448 VGND.n900 VGND.t1425 34.8005
R3449 VGND.n900 VGND.t781 34.8005
R3450 VGND.n447 VGND.t117 34.8005
R3451 VGND.n447 VGND.t779 34.8005
R3452 VGND.n1958 VGND.t551 34.8005
R3453 VGND.n1958 VGND.t777 34.8005
R3454 VGND.n450 VGND.t251 34.8005
R3455 VGND.n450 VGND.t1988 34.8005
R3456 VGND.n667 VGND.t1862 34.8005
R3457 VGND.n667 VGND.t1214 34.8005
R3458 VGND.n1392 VGND.t234 34.8005
R3459 VGND.n1392 VGND.t90 34.8005
R3460 VGND.n1397 VGND.t624 34.8005
R3461 VGND.n1397 VGND.t1556 34.8005
R3462 VGND.n664 VGND.t594 34.8005
R3463 VGND.n664 VGND.t1554 34.8005
R3464 VGND.n1820 VGND.t832 34.8005
R3465 VGND.n1820 VGND.t1212 34.8005
R3466 VGND.n485 VGND.t2080 34.8005
R3467 VGND.n485 VGND.t86 34.8005
R3468 VGND.n1846 VGND.t349 34.8005
R3469 VGND.n1846 VGND.t2011 34.8005
R3470 VGND.n477 VGND.t2596 34.8005
R3471 VGND.n477 VGND.t1210 34.8005
R3472 VGND.n1872 VGND.t7 34.8005
R3473 VGND.n1872 VGND.t1208 34.8005
R3474 VGND.n469 VGND.t640 34.8005
R3475 VGND.n469 VGND.t88 34.8005
R3476 VGND.n1898 VGND.t2260 34.8005
R3477 VGND.n1898 VGND.t1552 34.8005
R3478 VGND.n461 VGND.t96 34.8005
R3479 VGND.n461 VGND.t1550 34.8005
R3480 VGND.n1929 VGND.t1421 34.8005
R3481 VGND.n1929 VGND.t2009 34.8005
R3482 VGND.n1934 VGND.t2139 34.8005
R3483 VGND.n1934 VGND.t2007 34.8005
R3484 VGND.n1939 VGND.t213 34.8005
R3485 VGND.n1939 VGND.t2005 34.8005
R3486 VGND.n453 VGND.t247 34.8005
R3487 VGND.n453 VGND.t92 34.8005
R3488 VGND.n1371 VGND.t1790 34.8005
R3489 VGND.n1371 VGND.t492 34.8005
R3490 VGND.n1377 VGND.t1960 34.8005
R3491 VGND.n1377 VGND.t2580 34.8005
R3492 VGND.n1374 VGND.t2091 34.8005
R3493 VGND.n1374 VGND.t65 34.8005
R3494 VGND.n1807 VGND.t77 34.8005
R3495 VGND.n1807 VGND.t63 34.8005
R3496 VGND.n489 VGND.t1776 34.8005
R3497 VGND.n489 VGND.t490 34.8005
R3498 VGND.n1833 VGND.t616 34.8005
R3499 VGND.n1833 VGND.t2576 34.8005
R3500 VGND.n481 VGND.t325 34.8005
R3501 VGND.n481 VGND.t2574 34.8005
R3502 VGND.n1859 VGND.t541 34.8005
R3503 VGND.n1859 VGND.t488 34.8005
R3504 VGND.n473 VGND.t1704 34.8005
R3505 VGND.n473 VGND.t486 34.8005
R3506 VGND.n1885 VGND.t1175 34.8005
R3507 VGND.n1885 VGND.t2578 34.8005
R3508 VGND.n465 VGND.t2125 34.8005
R3509 VGND.n465 VGND.t496 34.8005
R3510 VGND.n1911 VGND.t560 34.8005
R3511 VGND.n1911 VGND.t494 34.8005
R3512 VGND.n457 VGND.t2494 34.8005
R3513 VGND.n457 VGND.t2572 34.8005
R3514 VGND.n1916 VGND.t2558 34.8005
R3515 VGND.n1916 VGND.t2570 34.8005
R3516 VGND.n2354 VGND.t13 34.8005
R3517 VGND.n2354 VGND.t483 34.8005
R3518 VGND.n303 VGND.t402 34.8005
R3519 VGND.n303 VGND.t2582 34.8005
R3520 VGND.n1303 VGND.t1886 34.8005
R3521 VGND.n1303 VGND.t1739 34.8005
R3522 VGND.n1309 VGND.t812 34.8005
R3523 VGND.n1309 VGND.t2166 34.8005
R3524 VGND.n1306 VGND.t1173 34.8005
R3525 VGND.n1306 VGND.t1747 34.8005
R3526 VGND.n1359 VGND.t580 34.8005
R3527 VGND.n1359 VGND.t1745 34.8005
R3528 VGND.n1354 VGND.t1735 34.8005
R3529 VGND.n1354 VGND.t1737 34.8005
R3530 VGND.n1349 VGND.t1570 34.8005
R3531 VGND.n1349 VGND.t2162 34.8005
R3532 VGND.n1344 VGND.t336 34.8005
R3533 VGND.n1344 VGND.t2160 34.8005
R3534 VGND.n1339 VGND.t2589 34.8005
R3535 VGND.n1339 VGND.t2172 34.8005
R3536 VGND.n1334 VGND.t1405 34.8005
R3537 VGND.n1334 VGND.t2170 34.8005
R3538 VGND.n1329 VGND.t629 34.8005
R3539 VGND.n1329 VGND.t2164 34.8005
R3540 VGND.n1324 VGND.t733 34.8005
R3541 VGND.n1324 VGND.t1743 34.8005
R3542 VGND.n1319 VGND.t2246 34.8005
R3543 VGND.n1319 VGND.t1741 34.8005
R3544 VGND.n1314 VGND.t1427 34.8005
R3545 VGND.n1314 VGND.t2158 34.8005
R3546 VGND.n503 VGND.t155 34.8005
R3547 VGND.n503 VGND.t1751 34.8005
R3548 VGND.n1784 VGND.t1943 34.8005
R3549 VGND.n1784 VGND.t1749 34.8005
R3550 VGND.n506 VGND.t382 34.8005
R3551 VGND.n506 VGND.t2168 34.8005
R3552 VGND.n571 VGND.t1817 34.8005
R3553 VGND.n571 VGND.t431 34.8005
R3554 VGND.n1514 VGND.t607 34.8005
R3555 VGND.n1514 VGND.t2421 34.8005
R3556 VGND.n1519 VGND.t306 34.8005
R3557 VGND.n1519 VGND.t722 34.8005
R3558 VGND.n575 VGND.t1696 34.8005
R3559 VGND.n575 VGND.t720 34.8005
R3560 VGND.n1646 VGND.t1726 34.8005
R3561 VGND.n1646 VGND.t429 34.8005
R3562 VGND.n541 VGND.t528 34.8005
R3563 VGND.n541 VGND.t2417 34.8005
R3564 VGND.n1672 VGND.t1299 34.8005
R3565 VGND.n1672 VGND.t2415 34.8005
R3566 VGND.n533 VGND.t534 34.8005
R3567 VGND.n533 VGND.t427 34.8005
R3568 VGND.n1698 VGND.t361 34.8005
R3569 VGND.n1698 VGND.t425 34.8005
R3570 VGND.n525 VGND.t1341 34.8005
R3571 VGND.n525 VGND.t2419 34.8005
R3572 VGND.n1724 VGND.t2670 34.8005
R3573 VGND.n1724 VGND.t718 34.8005
R3574 VGND.n517 VGND.t2036 34.8005
R3575 VGND.n517 VGND.t433 34.8005
R3576 VGND.n1755 VGND.t174 34.8005
R3577 VGND.n1755 VGND.t2413 34.8005
R3578 VGND.n1760 VGND.t2021 34.8005
R3579 VGND.n1760 VGND.t726 34.8005
R3580 VGND.n1765 VGND.t395 34.8005
R3581 VGND.n1765 VGND.t724 34.8005
R3582 VGND.n509 VGND.t659 34.8005
R3583 VGND.n509 VGND.t423 34.8005
R3584 VGND.n567 VGND.t1889 34.8005
R3585 VGND.n567 VGND.t2046 34.8005
R3586 VGND.n1534 VGND.t810 34.8005
R3587 VGND.n1534 VGND.t187 34.8005
R3588 VGND.n564 VGND.t1171 34.8005
R3589 VGND.n564 VGND.t1436 34.8005
R3590 VGND.n1633 VGND.t582 34.8005
R3591 VGND.n1633 VGND.t1434 34.8005
R3592 VGND.n545 VGND.t1733 34.8005
R3593 VGND.n545 VGND.t105 34.8005
R3594 VGND.n1659 VGND.t1568 34.8005
R3595 VGND.n1659 VGND.t183 34.8005
R3596 VGND.n537 VGND.t334 34.8005
R3597 VGND.n537 VGND.t181 34.8005
R3598 VGND.n1685 VGND.t2587 34.8005
R3599 VGND.n1685 VGND.t103 34.8005
R3600 VGND.n529 VGND.t1403 34.8005
R3601 VGND.n529 VGND.t191 34.8005
R3602 VGND.n1711 VGND.t439 34.8005
R3603 VGND.n1711 VGND.t185 34.8005
R3604 VGND.n521 VGND.t731 34.8005
R3605 VGND.n521 VGND.t2050 34.8005
R3606 VGND.n1737 VGND.t194 34.8005
R3607 VGND.n1737 VGND.t2048 34.8005
R3608 VGND.n513 VGND.t1614 34.8005
R3609 VGND.n513 VGND.t1442 34.8005
R3610 VGND.n1742 VGND.t153 34.8005
R3611 VGND.n1742 VGND.t1440 34.8005
R3612 VGND.n2379 VGND.t1941 34.8005
R3613 VGND.n2379 VGND.t1438 34.8005
R3614 VGND.n290 VGND.t380 34.8005
R3615 VGND.n290 VGND.t189 34.8005
R3616 VGND.n670 VGND.t1919 34.8005
R3617 VGND.n670 VGND.t44 34.8005
R3618 VGND.n672 VGND.t1346 34.8005
R3619 VGND.n672 VGND.t2152 34.8005
R3620 VGND.n1547 VGND.t302 34.8005
R3621 VGND.n1547 VGND.t1966 34.8005
R3622 VGND.n1552 VGND.t84 34.8005
R3623 VGND.n1552 VGND.t2156 34.8005
R3624 VGND.n1557 VGND.t1782 34.8005
R3625 VGND.n1557 VGND.t42 34.8005
R3626 VGND.n1562 VGND.t2272 34.8005
R3627 VGND.n1562 VGND.t2148 34.8005
R3628 VGND.n1567 VGND.t338 34.8005
R3629 VGND.n1567 VGND.t2146 34.8005
R3630 VGND.n1572 VGND.t414 34.8005
R3631 VGND.n1572 VGND.t40 34.8005
R3632 VGND.n1577 VGND.t740 34.8005
R3633 VGND.n1577 VGND.t38 34.8005
R3634 VGND.n1582 VGND.t200 34.8005
R3635 VGND.n1582 VGND.t2150 34.8005
R3636 VGND.n1587 VGND.t1543 34.8005
R3637 VGND.n1587 VGND.t48 34.8005
R3638 VGND.n1592 VGND.t2339 34.8005
R3639 VGND.n1592 VGND.t46 34.8005
R3640 VGND.n1597 VGND.t2002 34.8005
R3641 VGND.n1597 VGND.t2144 34.8005
R3642 VGND.n559 VGND.t2564 34.8005
R3643 VGND.n559 VGND.t2142 34.8005
R3644 VGND.n1610 VGND.t22 34.8005
R3645 VGND.n1610 VGND.t1968 34.8005
R3646 VGND.n1602 VGND.t408 34.8005
R3647 VGND.n1602 VGND.t2154 34.8005
R3648 VGND.n824 VGND.t1859 34.8005
R3649 VGND.n824 VGND.t1189 34.8005
R3650 VGND.n831 VGND.t236 34.8005
R3651 VGND.n831 VGND.t864 34.8005
R3652 VGND.n836 VGND.t626 34.8005
R3653 VGND.n836 VGND.t1688 34.8005
R3654 VGND.n828 VGND.t592 34.8005
R3655 VGND.n828 VGND.t1686 34.8005
R3656 VGND.n886 VGND.t834 34.8005
R3657 VGND.n886 VGND.t1187 34.8005
R3658 VGND.n881 VGND.t2082 34.8005
R3659 VGND.n881 VGND.t296 34.8005
R3660 VGND.n876 VGND.t347 34.8005
R3661 VGND.n876 VGND.t294 34.8005
R3662 VGND.n871 VGND.t2594 34.8005
R3663 VGND.n871 VGND.t1185 34.8005
R3664 VGND.n866 VGND.t5 34.8005
R3665 VGND.n866 VGND.t1181 34.8005
R3666 VGND.n861 VGND.t638 34.8005
R3667 VGND.n861 VGND.t298 34.8005
R3668 VGND.n856 VGND.t737 34.8005
R3669 VGND.n856 VGND.t1684 34.8005
R3670 VGND.n851 VGND.t94 34.8005
R3671 VGND.n851 VGND.t1191 34.8005
R3672 VGND.n846 VGND.t1419 34.8005
R3673 VGND.n846 VGND.t292 34.8005
R3674 VGND.n841 VGND.t160 34.8005
R3675 VGND.n841 VGND.t290 34.8005
R3676 VGND.n2399 VGND.t547 34.8005
R3677 VGND.n2399 VGND.t1690 34.8005
R3678 VGND.n278 VGND.t245 34.8005
R3679 VGND.n278 VGND.t866 34.8005
R3680 VGND.n814 VGND.t1125 34.8005
R3681 VGND.n814 VGND.t1054 34.8005
R3682 VGND.n717 VGND.t1510 34.8005
R3683 VGND.n717 VGND.t1127 34.8005
R3684 VGND.n74 VGND.n72 34.6358
R3685 VGND.n1109 VGND.n1091 34.6358
R3686 VGND.n1105 VGND.n1091 34.6358
R3687 VGND.n1105 VGND.n1104 34.6358
R3688 VGND.n1104 VGND.n1103 34.6358
R3689 VGND.n1103 VGND.n1093 34.6358
R3690 VGND.n1087 VGND.n1061 34.6358
R3691 VGND.n1082 VGND.n1062 34.6358
R3692 VGND.n1078 VGND.n1062 34.6358
R3693 VGND.n1078 VGND.n1077 34.6358
R3694 VGND.n1077 VGND.n1076 34.6358
R3695 VGND.n1076 VGND.n1064 34.6358
R3696 VGND.n130 VGND.n125 34.6358
R3697 VGND.n135 VGND.n134 34.6358
R3698 VGND.n598 VGND.n593 34.6358
R3699 VGND.n603 VGND.n602 34.6358
R3700 VGND.n976 VGND.n975 34.6358
R3701 VGND.n984 VGND.n983 34.6358
R3702 VGND.n980 VGND.n979 34.6358
R3703 VGND.n1020 VGND.n1000 34.6358
R3704 VGND.n1016 VGND.n1000 34.6358
R3705 VGND.n1016 VGND.n1015 34.6358
R3706 VGND.n1015 VGND.n1014 34.6358
R3707 VGND.n1014 VGND.n1002 34.6358
R3708 VGND.n1056 VGND.n1030 34.6358
R3709 VGND.n1051 VGND.n1031 34.6358
R3710 VGND.n1047 VGND.n1031 34.6358
R3711 VGND.n1047 VGND.n1046 34.6358
R3712 VGND.n1046 VGND.n1045 34.6358
R3713 VGND.n1045 VGND.n1033 34.6358
R3714 VGND.n160 VGND.n155 34.6358
R3715 VGND.n165 VGND.n164 34.6358
R3716 VGND.n17 VGND.n16 34.6358
R3717 VGND.n19 VGND.n10 34.6358
R3718 VGND.n23 VGND.n10 34.6358
R3719 VGND.n24 VGND.n23 34.6358
R3720 VGND.n25 VGND.n24 34.6358
R3721 VGND.n25 VGND.n8 34.6358
R3722 VGND.n46 VGND.n45 34.6358
R3723 VGND.n48 VGND.n37 34.6358
R3724 VGND.n52 VGND.n37 34.6358
R3725 VGND.n53 VGND.n52 34.6358
R3726 VGND.n54 VGND.n53 34.6358
R3727 VGND.n54 VGND.n35 34.6358
R3728 VGND.n100 VGND.n99 34.6358
R3729 VGND.n104 VGND.n103 34.6358
R3730 VGND.n2860 VGND.n2859 34.6358
R3731 VGND.n2864 VGND.n2863 34.6358
R3732 VGND.n2892 VGND.n2891 34.6358
R3733 VGND.n2896 VGND.n2895 34.6358
R3734 VGND.n78 VGND.n77 34.6358
R3735 VGND.n2935 VGND.n2929 34.6358
R3736 VGND.n2938 VGND.n2937 34.6358
R3737 VGND.n2938 VGND.n2925 34.6358
R3738 VGND.n2942 VGND.n2925 34.6358
R3739 VGND.n2943 VGND.n2942 34.6358
R3740 VGND.n2944 VGND.n2943 34.6358
R3741 VGND.n2960 VGND.n58 34.6358
R3742 VGND.n2975 VGND.n2974 34.6358
R3743 VGND.n2977 VGND.n2966 34.6358
R3744 VGND.n2981 VGND.n2966 34.6358
R3745 VGND.n2982 VGND.n2981 34.6358
R3746 VGND.n2983 VGND.n2982 34.6358
R3747 VGND.n2983 VGND.n2964 34.6358
R3748 VGND.n2992 VGND.n2987 34.6358
R3749 VGND.n2 VGND.t545 34.4422
R3750 VGND.n995 VGND.n898 33.1299
R3751 VGND.n2917 VGND.n2916 33.1299
R3752 VGND.n80 VGND.n62 32.377
R3753 VGND.n986 VGND.n985 32.377
R3754 VGND.n106 VGND.n105 32.377
R3755 VGND.n2866 VGND.n2865 32.377
R3756 VGND.n2898 VGND.n2897 32.377
R3757 VGND.n80 VGND.n79 32.377
R3758 VGND.n986 VGND.n964 32.0005
R3759 VGND.n141 VGND.n138 30.4946
R3760 VGND.n609 VGND.n606 30.4946
R3761 VGND.n171 VGND.n168 30.4946
R3762 VGND.n109 VGND.n86 29.8709
R3763 VGND.n1099 VGND.n1098 28.9887
R3764 VGND.n1072 VGND.n1071 28.9887
R3765 VGND.n1010 VGND.n1009 28.9887
R3766 VGND.n1041 VGND.n1040 28.9887
R3767 VGND.n18 VGND.n17 27.8593
R3768 VGND.n47 VGND.n46 27.8593
R3769 VGND.n2936 VGND.n2935 27.8593
R3770 VGND.n2976 VGND.n2975 27.8593
R3771 VGND.n119 VGND.n118 27.0003
R3772 VGND.n2871 VGND.n2870 26.8591
R3773 VGND.n983 VGND.n968 26.3534
R3774 VGND.n103 VGND.n92 26.3534
R3775 VGND.n2863 VGND.n2852 26.3534
R3776 VGND.n2895 VGND.n2884 26.3534
R3777 VGND.n77 VGND.n67 26.3534
R3778 VGND.n142 VGND.n141 25.977
R3779 VGND.n610 VGND.n609 25.977
R3780 VGND.n585 VGND.n582 25.977
R3781 VGND.n172 VGND.n171 25.977
R3782 VGND.n2903 VGND.n2878 25.977
R3783 VGND.n1095 VGND.t2307 24.9236
R3784 VGND.n1095 VGND.t2316 24.9236
R3785 VGND.n1097 VGND.t823 24.9236
R3786 VGND.n1097 VGND.t166 24.9236
R3787 VGND.n1067 VGND.t71 24.9236
R3788 VGND.n1067 VGND.t72 24.9236
R3789 VGND.n1066 VGND.t2308 24.9236
R3790 VGND.n1066 VGND.t2318 24.9236
R3791 VGND.n1070 VGND.t73 24.9236
R3792 VGND.n1070 VGND.t2126 24.9236
R3793 VGND.n1069 VGND.t824 24.9236
R3794 VGND.n1069 VGND.t168 24.9236
R3795 VGND.n132 VGND.t826 24.9236
R3796 VGND.n132 VGND.t2059 24.9236
R3797 VGND.n131 VGND.t816 24.9236
R3798 VGND.n131 VGND.t129 24.9236
R3799 VGND.n122 VGND.t1200 24.9236
R3800 VGND.n122 VGND.t821 24.9236
R3801 VGND.n121 VGND.t1580 24.9236
R3802 VGND.n121 VGND.t2312 24.9236
R3803 VGND.n140 VGND.t1603 24.9236
R3804 VGND.n140 VGND.t1199 24.9236
R3805 VGND.n139 VGND.t364 24.9236
R3806 VGND.n139 VGND.t365 24.9236
R3807 VGND.n600 VGND.t1361 24.9236
R3808 VGND.n600 VGND.t2303 24.9236
R3809 VGND.n599 VGND.t1354 24.9236
R3810 VGND.n599 VGND.t1411 24.9236
R3811 VGND.n590 VGND.t2096 24.9236
R3812 VGND.n590 VGND.t1360 24.9236
R3813 VGND.n589 VGND.t502 24.9236
R3814 VGND.n589 VGND.t2058 24.9236
R3815 VGND.n608 VGND.t2098 24.9236
R3816 VGND.n608 VGND.t2097 24.9236
R3817 VGND.n607 VGND.t504 24.9236
R3818 VGND.n607 VGND.t503 24.9236
R3819 VGND.n966 VGND.t2314 24.9236
R3820 VGND.n966 VGND.t123 24.9236
R3821 VGND.n967 VGND.t1013 24.9236
R3822 VGND.n967 VGND.t818 24.9236
R3823 VGND.n965 VGND.t1017 24.9236
R3824 VGND.n965 VGND.t1015 24.9236
R3825 VGND.n970 VGND.t820 24.9236
R3826 VGND.n970 VGND.t164 24.9236
R3827 VGND.n1005 VGND.t2309 24.9236
R3828 VGND.n1005 VGND.t2319 24.9236
R3829 VGND.n1004 VGND.t1412 24.9236
R3830 VGND.n1004 VGND.t1415 24.9236
R3831 VGND.n1008 VGND.t825 24.9236
R3832 VGND.n1008 VGND.t170 24.9236
R3833 VGND.n1007 VGND.t2317 24.9236
R3834 VGND.n1007 VGND.t125 24.9236
R3835 VGND.n1036 VGND.t2127 24.9236
R3836 VGND.n1036 VGND.t2128 24.9236
R3837 VGND.n1035 VGND.t127 24.9236
R3838 VGND.n1035 VGND.t130 24.9236
R3839 VGND.n1039 VGND.t121 24.9236
R3840 VGND.n1039 VGND.t69 24.9236
R3841 VGND.n1038 VGND.t1353 24.9236
R3842 VGND.n1038 VGND.t1410 24.9236
R3843 VGND.n162 VGND.t67 24.9236
R3844 VGND.n162 VGND.t2311 24.9236
R3845 VGND.n161 VGND.t1359 24.9236
R3846 VGND.n161 VGND.t1414 24.9236
R3847 VGND.n152 VGND.t2117 24.9236
R3848 VGND.n152 VGND.t1362 24.9236
R3849 VGND.n151 VGND.t511 24.9236
R3850 VGND.n151 VGND.t1358 24.9236
R3851 VGND.n170 VGND.t2115 24.9236
R3852 VGND.n170 VGND.t2116 24.9236
R3853 VGND.n169 VGND.t513 24.9236
R3854 VGND.n169 VGND.t512 24.9236
R3855 VGND.n13 VGND.t145 24.9236
R3856 VGND.n13 VGND.t2136 24.9236
R3857 VGND.n12 VGND.t28 24.9236
R3858 VGND.n12 VGND.t2504 24.9236
R3859 VGND.n42 VGND.t1528 24.9236
R3860 VGND.n42 VGND.t2489 24.9236
R3861 VGND.n41 VGND.t2505 24.9236
R3862 VGND.n41 VGND.t1534 24.9236
R3863 VGND.n40 VGND.t2685 24.9236
R3864 VGND.n40 VGND.t1562 24.9236
R3865 VGND.n39 VGND.t2498 24.9236
R3866 VGND.n39 VGND.t141 24.9236
R3867 VGND.n95 VGND.t32 24.9236
R3868 VGND.n95 VGND.t1571 24.9236
R3869 VGND.n94 VGND.t2687 24.9236
R3870 VGND.n94 VGND.t34 24.9236
R3871 VGND.n91 VGND.t24 24.9236
R3872 VGND.n91 VGND.t2606 24.9236
R3873 VGND.n90 VGND.t2682 24.9236
R3874 VGND.n90 VGND.t1431 24.9236
R3875 VGND.n89 VGND.t2605 24.9236
R3876 VGND.n89 VGND.t2607 24.9236
R3877 VGND.n88 VGND.t1786 24.9236
R3878 VGND.n88 VGND.t1937 24.9236
R3879 VGND.n2855 VGND.t1559 24.9236
R3880 VGND.n2855 VGND.t2681 24.9236
R3881 VGND.n2854 VGND.t138 24.9236
R3882 VGND.n2854 VGND.t1561 24.9236
R3883 VGND.n2851 VGND.t1575 24.9236
R3884 VGND.n2851 VGND.t2283 24.9236
R3885 VGND.n2850 VGND.t2137 24.9236
R3886 VGND.n2850 VGND.t1038 24.9236
R3887 VGND.n2849 VGND.t2282 24.9236
R3888 VGND.n2849 VGND.t2280 24.9236
R3889 VGND.n2848 VGND.t313 24.9236
R3890 VGND.n2848 VGND.t1634 24.9236
R3891 VGND.n2887 VGND.t1577 24.9236
R3892 VGND.n2887 VGND.t2678 24.9236
R3893 VGND.n2886 VGND.t2501 24.9236
R3894 VGND.n2886 VGND.t1524 24.9236
R3895 VGND.n2883 VGND.t1572 24.9236
R3896 VGND.n2883 VGND.t1957 24.9236
R3897 VGND.n2882 VGND.t1566 24.9236
R3898 VGND.n2882 VGND.t1629 24.9236
R3899 VGND.n2881 VGND.t1956 24.9236
R3900 VGND.n2881 VGND.t1954 24.9236
R3901 VGND.n2880 VGND.t1625 24.9236
R3902 VGND.n2880 VGND.t1619 24.9236
R3903 VGND.n65 VGND.t1536 24.9236
R3904 VGND.n65 VGND.t132 24.9236
R3905 VGND.n66 VGND.t1532 24.9236
R3906 VGND.n66 VGND.t1318 24.9236
R3907 VGND.n64 VGND.t1314 24.9236
R3908 VGND.n64 VGND.t1308 24.9236
R3909 VGND.n69 VGND.t1539 24.9236
R3910 VGND.n69 VGND.t143 24.9236
R3911 VGND.n2931 VGND.t1564 24.9236
R3912 VGND.n2931 VGND.t2683 24.9236
R3913 VGND.n2930 VGND.t2502 24.9236
R3914 VGND.n2930 VGND.t1530 24.9236
R3915 VGND.n2928 VGND.t1579 24.9236
R3916 VGND.n2928 VGND.t36 24.9236
R3917 VGND.n2927 VGND.t2496 24.9236
R3918 VGND.n2927 VGND.t139 24.9236
R3919 VGND.n2971 VGND.t149 24.9236
R3920 VGND.n2971 VGND.t2495 24.9236
R3921 VGND.n2970 VGND.t2684 24.9236
R3922 VGND.n2970 VGND.t26 24.9236
R3923 VGND.n2969 VGND.t134 24.9236
R3924 VGND.n2969 VGND.t1526 24.9236
R3925 VGND.n2968 VGND.t2680 24.9236
R3926 VGND.n2968 VGND.t1573 24.9236
R3927 VGND.n142 VGND.n116 24.4711
R3928 VGND.n610 VGND.n581 24.4711
R3929 VGND.n585 VGND.n584 24.4711
R3930 VGND.n996 VGND.n995 24.4711
R3931 VGND.n1025 VGND.n999 24.4711
R3932 VGND.n172 VGND.n148 24.4711
R3933 VGND.n106 VGND.n85 24.4711
R3934 VGND.n2866 VGND.n2845 24.4711
R3935 VGND.n2898 VGND.n2877 24.4711
R3936 VGND.n2903 VGND.n2902 24.4711
R3937 VGND.n2918 VGND.n2917 24.4711
R3938 VGND.n2949 VGND.n2948 24.4711
R3939 VGND.n2874 VGND.n2846 23.7181
R3940 VGND.n1111 VGND.n1109 23.7181
R3941 VGND.n1083 VGND.n1061 23.7181
R3942 VGND.n1083 VGND.n1082 23.7181
R3943 VGND.n146 VGND.n115 23.7181
R3944 VGND.n990 VGND.n899 23.7181
R3945 VGND.n1021 VGND.n1020 23.7181
R3946 VGND.n1052 VGND.n1030 23.7181
R3947 VGND.n1052 VGND.n1051 23.7181
R3948 VGND.n3008 VGND.n8 23.7181
R3949 VGND.n2961 VGND.n35 23.7181
R3950 VGND.n2944 VGND.n2923 23.7181
R3951 VGND.n2961 VGND.n2960 23.7181
R3952 VGND.n2993 VGND.n2964 23.7181
R3953 VGND.n2993 VGND.n2992 23.7181
R3954 VGND.n991 VGND.n990 23.3417
R3955 VGND.n2912 VGND.n84 23.3417
R3956 VGND.n2912 VGND.n61 23.3417
R3957 VGND.n1099 VGND.n1096 21.4593
R3958 VGND.n1072 VGND.n1068 21.4593
R3959 VGND.n1010 VGND.n1006 21.4593
R3960 VGND.n1041 VGND.n1037 21.4593
R3961 VGND.n98 VGND.n97 21.0905
R3962 VGND.n2858 VGND.n2857 21.0905
R3963 VGND.n2890 VGND.n2889 21.0905
R3964 VGND.n71 VGND.n70 21.0905
R3965 VGND.n99 VGND.n98 20.3299
R3966 VGND.n2859 VGND.n2858 20.3299
R3967 VGND.n2891 VGND.n2890 20.3299
R3968 VGND.n72 VGND.n71 20.3299
R3969 VGND.n138 VGND.n123 19.9534
R3970 VGND.n606 VGND.n591 19.9534
R3971 VGND.n168 VGND.n153 19.9534
R3972 VGND.n1026 VGND.n1025 19.2005
R3973 VGND.n1057 VGND.n1056 19.2005
R3974 VGND.n2950 VGND.n2949 19.2005
R3975 VGND.n2955 VGND.n58 19.2005
R3976 VGND.t1969 VGND.t2086 16.8587
R3977 VGND.t749 VGND.t2084 16.8587
R3978 VGND.t2298 VGND.t1705 16.8587
R3979 VGND.t2673 VGND.t1707 16.8587
R3980 VGND.n1089 VGND.n1088 16.077
R3981 VGND.n2989 VGND.n2988 16.077
R3982 VGND.n1027 VGND.n1026 15.4358
R3983 VGND.n2951 VGND.n2950 15.4358
R3984 VGND.n118 VGND.n117 14.6829
R3985 VGND.n1058 VGND.n1057 14.6829
R3986 VGND.n2870 VGND.n2869 14.6829
R3987 VGND.n2956 VGND.n2955 14.6829
R3988 VGND.n127 VGND.n126 14.5711
R3989 VGND.n595 VGND.n594 14.5711
R3990 VGND.n974 VGND.n973 14.5711
R3991 VGND.n157 VGND.n156 14.5711
R3992 VGND.n614 VGND.n582 14.3064
R3993 VGND.n2907 VGND.n2878 14.3064
R3994 VGND.n134 VGND.n133 13.9299
R3995 VGND.n602 VGND.n601 13.9299
R3996 VGND.n979 VGND.n971 13.9299
R3997 VGND.n164 VGND.n163 13.9299
R3998 VGND.n1021 VGND.n999 13.5534
R3999 VGND.n2948 VGND.n2923 13.5534
R4000 VGND.n146 VGND.n116 13.177
R4001 VGND.n614 VGND.n581 13.177
R4002 VGND.n176 VGND.n148 13.177
R4003 VGND.n112 VGND.n85 13.177
R4004 VGND.n2874 VGND.n2845 13.177
R4005 VGND.n2907 VGND.n2877 13.177
R4006 VGND.n176 VGND.n149 12.8005
R4007 VGND.n112 VGND.n86 12.8005
R4008 VGND.n3022 VGND.t2697 12.5645
R4009 VGND.n1088 VGND.n1087 10.5417
R4010 VGND.n2988 VGND.n2987 10.5417
R4011 VGND.n1059 VGND.n1058 10.0534
R4012 VGND.n2957 VGND.n2956 10.0534
R4013 VGND.n1100 VGND.n1099 9.3005
R4014 VGND.n1101 VGND.n1093 9.3005
R4015 VGND.n1103 VGND.n1102 9.3005
R4016 VGND.n1104 VGND.n1092 9.3005
R4017 VGND.n1106 VGND.n1105 9.3005
R4018 VGND.n1107 VGND.n1091 9.3005
R4019 VGND.n1109 VGND.n1108 9.3005
R4020 VGND.n1112 VGND.n1111 9.3005
R4021 VGND.n1073 VGND.n1072 9.3005
R4022 VGND.n1074 VGND.n1064 9.3005
R4023 VGND.n1076 VGND.n1075 9.3005
R4024 VGND.n1077 VGND.n1063 9.3005
R4025 VGND.n1079 VGND.n1078 9.3005
R4026 VGND.n1080 VGND.n1062 9.3005
R4027 VGND.n1082 VGND.n1081 9.3005
R4028 VGND.n1085 VGND.n1061 9.3005
R4029 VGND.n1087 VGND.n1086 9.3005
R4030 VGND.n1084 VGND.n1083 9.3005
R4031 VGND.n144 VGND.n116 9.3005
R4032 VGND.n128 VGND.n125 9.3005
R4033 VGND.n130 VGND.n129 9.3005
R4034 VGND.n134 VGND.n124 9.3005
R4035 VGND.n136 VGND.n135 9.3005
R4036 VGND.n138 VGND.n137 9.3005
R4037 VGND.n141 VGND.n120 9.3005
R4038 VGND.n143 VGND.n142 9.3005
R4039 VGND.n119 VGND.n115 9.3005
R4040 VGND.n146 VGND.n145 9.3005
R4041 VGND.n584 VGND.n583 9.3005
R4042 VGND.n587 VGND.n582 9.3005
R4043 VGND.n612 VGND.n581 9.3005
R4044 VGND.n596 VGND.n593 9.3005
R4045 VGND.n598 VGND.n597 9.3005
R4046 VGND.n602 VGND.n592 9.3005
R4047 VGND.n604 VGND.n603 9.3005
R4048 VGND.n606 VGND.n605 9.3005
R4049 VGND.n609 VGND.n588 9.3005
R4050 VGND.n611 VGND.n610 9.3005
R4051 VGND.n586 VGND.n585 9.3005
R4052 VGND.n614 VGND.n613 9.3005
R4053 VGND.n997 VGND.n996 9.3005
R4054 VGND.n988 VGND.n899 9.3005
R4055 VGND.n975 VGND.n972 9.3005
R4056 VGND.n977 VGND.n976 9.3005
R4057 VGND.n979 VGND.n978 9.3005
R4058 VGND.n981 VGND.n980 9.3005
R4059 VGND.n983 VGND.n982 9.3005
R4060 VGND.n984 VGND.n963 9.3005
R4061 VGND.n987 VGND.n986 9.3005
R4062 VGND.n993 VGND.n992 9.3005
R4063 VGND.n995 VGND.n994 9.3005
R4064 VGND.n990 VGND.n989 9.3005
R4065 VGND.n1011 VGND.n1010 9.3005
R4066 VGND.n1012 VGND.n1002 9.3005
R4067 VGND.n1014 VGND.n1013 9.3005
R4068 VGND.n1015 VGND.n1001 9.3005
R4069 VGND.n1017 VGND.n1016 9.3005
R4070 VGND.n1018 VGND.n1000 9.3005
R4071 VGND.n1020 VGND.n1019 9.3005
R4072 VGND.n1023 VGND.n999 9.3005
R4073 VGND.n1025 VGND.n1024 9.3005
R4074 VGND.n1028 VGND.n1027 9.3005
R4075 VGND.n1022 VGND.n1021 9.3005
R4076 VGND.n1042 VGND.n1041 9.3005
R4077 VGND.n1043 VGND.n1033 9.3005
R4078 VGND.n1045 VGND.n1044 9.3005
R4079 VGND.n1046 VGND.n1032 9.3005
R4080 VGND.n1048 VGND.n1047 9.3005
R4081 VGND.n1049 VGND.n1031 9.3005
R4082 VGND.n1051 VGND.n1050 9.3005
R4083 VGND.n1054 VGND.n1030 9.3005
R4084 VGND.n1056 VGND.n1055 9.3005
R4085 VGND.n1053 VGND.n1052 9.3005
R4086 VGND.n174 VGND.n148 9.3005
R4087 VGND.n158 VGND.n155 9.3005
R4088 VGND.n160 VGND.n159 9.3005
R4089 VGND.n164 VGND.n154 9.3005
R4090 VGND.n166 VGND.n165 9.3005
R4091 VGND.n168 VGND.n167 9.3005
R4092 VGND.n171 VGND.n150 9.3005
R4093 VGND.n173 VGND.n172 9.3005
R4094 VGND.n176 VGND.n175 9.3005
R4095 VGND.n3008 VGND.n3007 9.3005
R4096 VGND.n16 VGND.n15 9.3005
R4097 VGND.n17 VGND.n11 9.3005
R4098 VGND.n20 VGND.n19 9.3005
R4099 VGND.n21 VGND.n10 9.3005
R4100 VGND.n23 VGND.n22 9.3005
R4101 VGND.n24 VGND.n9 9.3005
R4102 VGND.n26 VGND.n25 9.3005
R4103 VGND.n27 VGND.n8 9.3005
R4104 VGND.n110 VGND.n86 9.3005
R4105 VGND.n99 VGND.n93 9.3005
R4106 VGND.n101 VGND.n100 9.3005
R4107 VGND.n103 VGND.n102 9.3005
R4108 VGND.n104 VGND.n87 9.3005
R4109 VGND.n107 VGND.n106 9.3005
R4110 VGND.n108 VGND.n85 9.3005
R4111 VGND.n112 VGND.n111 9.3005
R4112 VGND.n2872 VGND.n2846 9.3005
R4113 VGND.n2859 VGND.n2853 9.3005
R4114 VGND.n2861 VGND.n2860 9.3005
R4115 VGND.n2863 VGND.n2862 9.3005
R4116 VGND.n2864 VGND.n2847 9.3005
R4117 VGND.n2867 VGND.n2866 9.3005
R4118 VGND.n2868 VGND.n2845 9.3005
R4119 VGND.n2874 VGND.n2873 9.3005
R4120 VGND.n2902 VGND.n2901 9.3005
R4121 VGND.n2891 VGND.n2885 9.3005
R4122 VGND.n2893 VGND.n2892 9.3005
R4123 VGND.n2895 VGND.n2894 9.3005
R4124 VGND.n2896 VGND.n2879 9.3005
R4125 VGND.n2899 VGND.n2898 9.3005
R4126 VGND.n2900 VGND.n2877 9.3005
R4127 VGND.n2905 VGND.n2878 9.3005
R4128 VGND.n2904 VGND.n2903 9.3005
R4129 VGND.n2907 VGND.n2906 9.3005
R4130 VGND.n2919 VGND.n2918 9.3005
R4131 VGND.n72 VGND.n68 9.3005
R4132 VGND.n75 VGND.n74 9.3005
R4133 VGND.n77 VGND.n76 9.3005
R4134 VGND.n78 VGND.n63 9.3005
R4135 VGND.n81 VGND.n80 9.3005
R4136 VGND.n83 VGND.n82 9.3005
R4137 VGND.n2915 VGND.n2914 9.3005
R4138 VGND.n2917 VGND.n60 9.3005
R4139 VGND.n2913 VGND.n2912 9.3005
R4140 VGND.n2952 VGND.n2951 9.3005
R4141 VGND.n2933 VGND.n2929 9.3005
R4142 VGND.n2935 VGND.n2934 9.3005
R4143 VGND.n2937 VGND.n2926 9.3005
R4144 VGND.n2939 VGND.n2938 9.3005
R4145 VGND.n2940 VGND.n2925 9.3005
R4146 VGND.n2942 VGND.n2941 9.3005
R4147 VGND.n2943 VGND.n2924 9.3005
R4148 VGND.n2945 VGND.n2944 9.3005
R4149 VGND.n2948 VGND.n2947 9.3005
R4150 VGND.n2949 VGND.n2921 9.3005
R4151 VGND.n2946 VGND.n2923 9.3005
R4152 VGND.n45 VGND.n44 9.3005
R4153 VGND.n46 VGND.n38 9.3005
R4154 VGND.n49 VGND.n48 9.3005
R4155 VGND.n50 VGND.n37 9.3005
R4156 VGND.n52 VGND.n51 9.3005
R4157 VGND.n53 VGND.n36 9.3005
R4158 VGND.n55 VGND.n54 9.3005
R4159 VGND.n56 VGND.n35 9.3005
R4160 VGND.n2961 VGND.n57 9.3005
R4161 VGND.n2960 VGND.n2959 9.3005
R4162 VGND.n2958 VGND.n58 9.3005
R4163 VGND.n2974 VGND.n2973 9.3005
R4164 VGND.n2975 VGND.n2967 9.3005
R4165 VGND.n2978 VGND.n2977 9.3005
R4166 VGND.n2979 VGND.n2966 9.3005
R4167 VGND.n2981 VGND.n2980 9.3005
R4168 VGND.n2982 VGND.n2965 9.3005
R4169 VGND.n2984 VGND.n2983 9.3005
R4170 VGND.n2985 VGND.n2964 9.3005
R4171 VGND.n2993 VGND.n2986 9.3005
R4172 VGND.n2992 VGND.n2991 9.3005
R4173 VGND.n2990 VGND.n2987 9.3005
R4174 VGND.n100 VGND.n92 8.28285
R4175 VGND.n2860 VGND.n2852 8.28285
R4176 VGND.n2892 VGND.n2884 8.28285
R4177 VGND.n2713 VGND.n235 7.9105
R4178 VGND.n2715 VGND.n2714 7.9105
R4179 VGND.n2820 VGND.n189 7.9105
R4180 VGND.n2819 VGND.n190 7.9105
R4181 VGND.n2814 VGND.n195 7.9105
R4182 VGND.n2813 VGND.n196 7.9105
R4183 VGND.n2808 VGND.n201 7.9105
R4184 VGND.n2807 VGND.n202 7.9105
R4185 VGND.n2802 VGND.n207 7.9105
R4186 VGND.n2801 VGND.n208 7.9105
R4187 VGND.n2796 VGND.n213 7.9105
R4188 VGND.n2795 VGND.n214 7.9105
R4189 VGND.n2790 VGND.n219 7.9105
R4190 VGND.n2789 VGND.n220 7.9105
R4191 VGND.n2784 VGND.n2783 7.9105
R4192 VGND.n3002 VGND.n3001 7.9105
R4193 VGND.n2518 VGND.n2517 7.9105
R4194 VGND.n2824 VGND.n185 7.9105
R4195 VGND.n2823 VGND.n186 7.9105
R4196 VGND.n2505 VGND.n2504 7.9105
R4197 VGND.n2503 VGND.n248 7.9105
R4198 VGND.n2502 VGND.n249 7.9105
R4199 VGND.n2501 VGND.n250 7.9105
R4200 VGND.n2500 VGND.n251 7.9105
R4201 VGND.n2499 VGND.n252 7.9105
R4202 VGND.n2498 VGND.n253 7.9105
R4203 VGND.n2497 VGND.n254 7.9105
R4204 VGND.n2496 VGND.n255 7.9105
R4205 VGND.n2495 VGND.n256 7.9105
R4206 VGND.n2494 VGND.n257 7.9105
R4207 VGND.n2493 VGND.n258 7.9105
R4208 VGND.n2492 VGND.n2491 7.9105
R4209 VGND.n639 VGND.n180 7.9105
R4210 VGND.n2828 VGND.n2827 7.9105
R4211 VGND.n375 VGND.n374 7.9105
R4212 VGND.n2167 VGND.n2166 7.9105
R4213 VGND.n2176 VGND.n2175 7.9105
R4214 VGND.n2193 VGND.n2192 7.9105
R4215 VGND.n2202 VGND.n2201 7.9105
R4216 VGND.n2219 VGND.n2218 7.9105
R4217 VGND.n2228 VGND.n2227 7.9105
R4218 VGND.n2245 VGND.n2244 7.9105
R4219 VGND.n2254 VGND.n2253 7.9105
R4220 VGND.n2276 VGND.n2275 7.9105
R4221 VGND.n2298 VGND.n328 7.9105
R4222 VGND.n2297 VGND.n329 7.9105
R4223 VGND.n2295 VGND.n2294 7.9105
R4224 VGND.n2431 VGND.n2430 7.9105
R4225 VGND.n1434 VGND.n1421 7.9105
R4226 VGND.n1433 VGND.n1432 7.9105
R4227 VGND.n2154 VGND.n2153 7.9105
R4228 VGND.n2163 VGND.n2162 7.9105
R4229 VGND.n2180 VGND.n2179 7.9105
R4230 VGND.n2189 VGND.n2188 7.9105
R4231 VGND.n2206 VGND.n2205 7.9105
R4232 VGND.n2215 VGND.n2214 7.9105
R4233 VGND.n2232 VGND.n2231 7.9105
R4234 VGND.n2241 VGND.n2240 7.9105
R4235 VGND.n2258 VGND.n2257 7.9105
R4236 VGND.n2272 VGND.n2271 7.9105
R4237 VGND.n2301 VGND.n327 7.9105
R4238 VGND.n2303 VGND.n2302 7.9105
R4239 VGND.n2315 VGND.n324 7.9105
R4240 VGND.n2314 VGND.n2313 7.9105
R4241 VGND.n1438 VGND.n1437 7.9105
R4242 VGND.n1497 VGND.n1496 7.9105
R4243 VGND.n2150 VGND.n381 7.9105
R4244 VGND.n2149 VGND.n382 7.9105
R4245 VGND.n2148 VGND.n383 7.9105
R4246 VGND.n2147 VGND.n384 7.9105
R4247 VGND.n2146 VGND.n385 7.9105
R4248 VGND.n2145 VGND.n386 7.9105
R4249 VGND.n2144 VGND.n387 7.9105
R4250 VGND.n2143 VGND.n388 7.9105
R4251 VGND.n2142 VGND.n389 7.9105
R4252 VGND.n2141 VGND.n390 7.9105
R4253 VGND.n2140 VGND.n2139 7.9105
R4254 VGND.n2319 VGND.n321 7.9105
R4255 VGND.n2318 VGND.n322 7.9105
R4256 VGND.n2127 VGND.n2126 7.9105
R4257 VGND.n1415 VGND.n617 7.9105
R4258 VGND.n1501 VGND.n1500 7.9105
R4259 VGND.n630 VGND.n629 7.9105
R4260 VGND.n1993 VGND.n1992 7.9105
R4261 VGND.n2002 VGND.n2001 7.9105
R4262 VGND.n2019 VGND.n2018 7.9105
R4263 VGND.n2028 VGND.n2027 7.9105
R4264 VGND.n2045 VGND.n2044 7.9105
R4265 VGND.n2054 VGND.n2053 7.9105
R4266 VGND.n2071 VGND.n2070 7.9105
R4267 VGND.n2080 VGND.n2079 7.9105
R4268 VGND.n2102 VGND.n2101 7.9105
R4269 VGND.n2323 VGND.n318 7.9105
R4270 VGND.n2322 VGND.n319 7.9105
R4271 VGND.n399 VGND.n398 7.9105
R4272 VGND.n2123 VGND.n2122 7.9105
R4273 VGND.n1413 VGND.n644 7.9105
R4274 VGND.n656 VGND.n655 7.9105
R4275 VGND.n1980 VGND.n1979 7.9105
R4276 VGND.n1989 VGND.n1988 7.9105
R4277 VGND.n2006 VGND.n2005 7.9105
R4278 VGND.n2015 VGND.n2014 7.9105
R4279 VGND.n2032 VGND.n2031 7.9105
R4280 VGND.n2041 VGND.n2040 7.9105
R4281 VGND.n2058 VGND.n2057 7.9105
R4282 VGND.n2067 VGND.n2066 7.9105
R4283 VGND.n2084 VGND.n2083 7.9105
R4284 VGND.n2098 VGND.n2097 7.9105
R4285 VGND.n2326 VGND.n316 7.9105
R4286 VGND.n2328 VGND.n2327 7.9105
R4287 VGND.n2340 VGND.n312 7.9105
R4288 VGND.n2339 VGND.n2338 7.9105
R4289 VGND.n1410 VGND.n660 7.9105
R4290 VGND.n1409 VGND.n661 7.9105
R4291 VGND.n1976 VGND.n437 7.9105
R4292 VGND.n1975 VGND.n438 7.9105
R4293 VGND.n1974 VGND.n439 7.9105
R4294 VGND.n1973 VGND.n440 7.9105
R4295 VGND.n1972 VGND.n441 7.9105
R4296 VGND.n1971 VGND.n442 7.9105
R4297 VGND.n1970 VGND.n443 7.9105
R4298 VGND.n1969 VGND.n444 7.9105
R4299 VGND.n1968 VGND.n445 7.9105
R4300 VGND.n1967 VGND.n446 7.9105
R4301 VGND.n1966 VGND.n1965 7.9105
R4302 VGND.n2344 VGND.n309 7.9105
R4303 VGND.n2343 VGND.n310 7.9105
R4304 VGND.n1953 VGND.n1952 7.9105
R4305 VGND.n1391 VGND.n1390 7.9105
R4306 VGND.n1406 VGND.n663 7.9105
R4307 VGND.n1405 VGND.n1404 7.9105
R4308 VGND.n1819 VGND.n1818 7.9105
R4309 VGND.n1828 VGND.n1827 7.9105
R4310 VGND.n1845 VGND.n1844 7.9105
R4311 VGND.n1854 VGND.n1853 7.9105
R4312 VGND.n1871 VGND.n1870 7.9105
R4313 VGND.n1880 VGND.n1879 7.9105
R4314 VGND.n1897 VGND.n1896 7.9105
R4315 VGND.n1906 VGND.n1905 7.9105
R4316 VGND.n1928 VGND.n1927 7.9105
R4317 VGND.n2348 VGND.n306 7.9105
R4318 VGND.n2347 VGND.n307 7.9105
R4319 VGND.n455 VGND.n454 7.9105
R4320 VGND.n1949 VGND.n1948 7.9105
R4321 VGND.n1387 VGND.n1373 7.9105
R4322 VGND.n1385 VGND.n1384 7.9105
R4323 VGND.n1806 VGND.n1805 7.9105
R4324 VGND.n1815 VGND.n1814 7.9105
R4325 VGND.n1832 VGND.n1831 7.9105
R4326 VGND.n1841 VGND.n1840 7.9105
R4327 VGND.n1858 VGND.n1857 7.9105
R4328 VGND.n1867 VGND.n1866 7.9105
R4329 VGND.n1884 VGND.n1883 7.9105
R4330 VGND.n1893 VGND.n1892 7.9105
R4331 VGND.n1910 VGND.n1909 7.9105
R4332 VGND.n1924 VGND.n1923 7.9105
R4333 VGND.n2351 VGND.n304 7.9105
R4334 VGND.n2353 VGND.n2352 7.9105
R4335 VGND.n2365 VGND.n300 7.9105
R4336 VGND.n2364 VGND.n2363 7.9105
R4337 VGND.n1369 VGND.n1305 7.9105
R4338 VGND.n1368 VGND.n1366 7.9105
R4339 VGND.n1802 VGND.n493 7.9105
R4340 VGND.n1801 VGND.n494 7.9105
R4341 VGND.n1800 VGND.n495 7.9105
R4342 VGND.n1799 VGND.n496 7.9105
R4343 VGND.n1798 VGND.n497 7.9105
R4344 VGND.n1797 VGND.n498 7.9105
R4345 VGND.n1796 VGND.n499 7.9105
R4346 VGND.n1795 VGND.n500 7.9105
R4347 VGND.n1794 VGND.n501 7.9105
R4348 VGND.n1793 VGND.n502 7.9105
R4349 VGND.n1792 VGND.n1791 7.9105
R4350 VGND.n2369 VGND.n297 7.9105
R4351 VGND.n2368 VGND.n298 7.9105
R4352 VGND.n1779 VGND.n1778 7.9105
R4353 VGND.n1529 VGND.n573 7.9105
R4354 VGND.n1528 VGND.n574 7.9105
R4355 VGND.n1527 VGND.n1526 7.9105
R4356 VGND.n1645 VGND.n1644 7.9105
R4357 VGND.n1654 VGND.n1653 7.9105
R4358 VGND.n1671 VGND.n1670 7.9105
R4359 VGND.n1680 VGND.n1679 7.9105
R4360 VGND.n1697 VGND.n1696 7.9105
R4361 VGND.n1706 VGND.n1705 7.9105
R4362 VGND.n1723 VGND.n1722 7.9105
R4363 VGND.n1732 VGND.n1731 7.9105
R4364 VGND.n1754 VGND.n1753 7.9105
R4365 VGND.n2373 VGND.n294 7.9105
R4366 VGND.n2372 VGND.n295 7.9105
R4367 VGND.n511 VGND.n510 7.9105
R4368 VGND.n1775 VGND.n1774 7.9105
R4369 VGND.n1533 VGND.n1532 7.9105
R4370 VGND.n1542 VGND.n1541 7.9105
R4371 VGND.n1632 VGND.n1631 7.9105
R4372 VGND.n1641 VGND.n1640 7.9105
R4373 VGND.n1658 VGND.n1657 7.9105
R4374 VGND.n1667 VGND.n1666 7.9105
R4375 VGND.n1684 VGND.n1683 7.9105
R4376 VGND.n1693 VGND.n1692 7.9105
R4377 VGND.n1710 VGND.n1709 7.9105
R4378 VGND.n1719 VGND.n1718 7.9105
R4379 VGND.n1736 VGND.n1735 7.9105
R4380 VGND.n1750 VGND.n1749 7.9105
R4381 VGND.n2376 VGND.n291 7.9105
R4382 VGND.n2378 VGND.n2377 7.9105
R4383 VGND.n2390 VGND.n287 7.9105
R4384 VGND.n2389 VGND.n2388 7.9105
R4385 VGND.n1299 VGND.n1298 7.9105
R4386 VGND.n1546 VGND.n1545 7.9105
R4387 VGND.n1628 VGND.n549 7.9105
R4388 VGND.n1627 VGND.n550 7.9105
R4389 VGND.n1626 VGND.n551 7.9105
R4390 VGND.n1625 VGND.n552 7.9105
R4391 VGND.n1624 VGND.n553 7.9105
R4392 VGND.n1623 VGND.n554 7.9105
R4393 VGND.n1622 VGND.n555 7.9105
R4394 VGND.n1621 VGND.n556 7.9105
R4395 VGND.n1620 VGND.n557 7.9105
R4396 VGND.n1619 VGND.n558 7.9105
R4397 VGND.n1618 VGND.n1617 7.9105
R4398 VGND.n2394 VGND.n282 7.9105
R4399 VGND.n2393 VGND.n283 7.9105
R4400 VGND.n1605 VGND.n1604 7.9105
R4401 VGND.n896 VGND.n826 7.9105
R4402 VGND.n895 VGND.n827 7.9105
R4403 VGND.n894 VGND.n893 7.9105
R4404 VGND.n1276 VGND.n688 7.9105
R4405 VGND.n1275 VGND.n689 7.9105
R4406 VGND.n1268 VGND.n694 7.9105
R4407 VGND.n1267 VGND.n695 7.9105
R4408 VGND.n1260 VGND.n700 7.9105
R4409 VGND.n1259 VGND.n701 7.9105
R4410 VGND.n1252 VGND.n706 7.9105
R4411 VGND.n1251 VGND.n707 7.9105
R4412 VGND.n1244 VGND.n712 7.9105
R4413 VGND.n1243 VGND.n713 7.9105
R4414 VGND.n2398 VGND.n2397 7.9105
R4415 VGND.n284 VGND.n279 7.9105
R4416 VGND.n2409 VGND.n2408 7.9105
R4417 VGND.n1118 VGND.n677 7.9105
R4418 VGND.n1286 VGND.n1285 7.9105
R4419 VGND.n1280 VGND.n685 7.9105
R4420 VGND.n1279 VGND.n686 7.9105
R4421 VGND.n1272 VGND.n691 7.9105
R4422 VGND.n1271 VGND.n692 7.9105
R4423 VGND.n1264 VGND.n697 7.9105
R4424 VGND.n1263 VGND.n698 7.9105
R4425 VGND.n1256 VGND.n703 7.9105
R4426 VGND.n1255 VGND.n704 7.9105
R4427 VGND.n1248 VGND.n709 7.9105
R4428 VGND.n1247 VGND.n710 7.9105
R4429 VGND.n1240 VGND.n715 7.9105
R4430 VGND.n1239 VGND.n716 7.9105
R4431 VGND.n1238 VGND.n783 7.9105
R4432 VGND.n2413 VGND.n2412 7.9105
R4433 VGND.n133 VGND.n130 7.90638
R4434 VGND.n126 VGND.n125 7.90638
R4435 VGND.n601 VGND.n598 7.90638
R4436 VGND.n594 VGND.n593 7.90638
R4437 VGND.n976 VGND.n971 7.90638
R4438 VGND.n975 VGND.n974 7.90638
R4439 VGND.n163 VGND.n160 7.90638
R4440 VGND.n156 VGND.n155 7.90638
R4441 VGND.n1098 VGND.n1094 7.4049
R4442 VGND.n1071 VGND.n1065 7.4049
R4443 VGND.n1009 VGND.n1003 7.4049
R4444 VGND.n1040 VGND.n1034 7.4049
R4445 VGND VGND.n149 7.12482
R4446 VGND.n97 VGND.n96 6.85473
R4447 VGND.n2857 VGND.n2856 6.85473
R4448 VGND.n2889 VGND.n2888 6.85473
R4449 VGND.n19 VGND.n18 6.77697
R4450 VGND.n48 VGND.n47 6.77697
R4451 VGND.n2937 VGND.n2936 6.77697
R4452 VGND.n2977 VGND.n2976 6.77697
R4453 VGND.n3021 VGND.n3020 6.4005
R4454 VGND.n969 VGND.n968 5.27109
R4455 VGND.n73 VGND.n67 5.27109
R4456 VGND.n2570 VGND.n2569 4.5005
R4457 VGND.n2625 VGND.n2582 4.5005
R4458 VGND.n2622 VGND.n2621 4.5005
R4459 VGND.n2619 VGND.n2618 4.5005
R4460 VGND.n2616 VGND.n2615 4.5005
R4461 VGND.n2613 VGND.n2612 4.5005
R4462 VGND.n2610 VGND.n2609 4.5005
R4463 VGND.n2607 VGND.n2606 4.5005
R4464 VGND.n2604 VGND.n2603 4.5005
R4465 VGND.n2601 VGND.n2600 4.5005
R4466 VGND.n2598 VGND.n2597 4.5005
R4467 VGND.n2595 VGND.n2594 4.5005
R4468 VGND.n2592 VGND.n2591 4.5005
R4469 VGND.n2589 VGND.n2588 4.5005
R4470 VGND.n2651 VGND.n223 4.5005
R4471 VGND.n2660 VGND.n222 4.5005
R4472 VGND.n2647 VGND.n217 4.5005
R4473 VGND.n2668 VGND.n216 4.5005
R4474 VGND.n2643 VGND.n211 4.5005
R4475 VGND.n2676 VGND.n210 4.5005
R4476 VGND.n2639 VGND.n205 4.5005
R4477 VGND.n2684 VGND.n204 4.5005
R4478 VGND.n2635 VGND.n199 4.5005
R4479 VGND.n2692 VGND.n198 4.5005
R4480 VGND.n2631 VGND.n193 4.5005
R4481 VGND.n2700 VGND.n192 4.5005
R4482 VGND.n2627 VGND.n2626 4.5005
R4483 VGND.n2709 VGND.n2708 4.5005
R4484 VGND.n2524 VGND.n2523 4.5005
R4485 VGND.n2527 VGND.n2526 4.5005
R4486 VGND.n2530 VGND.n2529 4.5005
R4487 VGND.n2533 VGND.n2532 4.5005
R4488 VGND.n2536 VGND.n2535 4.5005
R4489 VGND.n2539 VGND.n2538 4.5005
R4490 VGND.n2542 VGND.n2541 4.5005
R4491 VGND.n2545 VGND.n2544 4.5005
R4492 VGND.n2548 VGND.n2547 4.5005
R4493 VGND.n2551 VGND.n2550 4.5005
R4494 VGND.n2554 VGND.n2553 4.5005
R4495 VGND.n2557 VGND.n2556 4.5005
R4496 VGND.n2560 VGND.n2559 4.5005
R4497 VGND.n2563 VGND.n2562 4.5005
R4498 VGND.n2566 VGND.n2565 4.5005
R4499 VGND.n2576 VGND.n2568 4.5005
R4500 VGND.n2584 VGND.n2583 4.5005
R4501 VGND.n2587 VGND.n2586 4.5005
R4502 VGND.n2652 VGND.n30 4.5005
R4503 VGND.n820 VGND.n819 4.5005
R4504 VGND.n817 VGND.n816 4.5005
R4505 VGND.n1138 VGND.n1137 4.5005
R4506 VGND.n1150 VGND.n807 4.5005
R4507 VGND.n1157 VGND.n805 4.5005
R4508 VGND.n1154 VGND.n1152 4.5005
R4509 VGND.n1170 VGND.n1169 4.5005
R4510 VGND.n1182 VGND.n799 4.5005
R4511 VGND.n1189 VGND.n797 4.5005
R4512 VGND.n1186 VGND.n1184 4.5005
R4513 VGND.n1202 VGND.n1201 4.5005
R4514 VGND.n1214 VGND.n791 4.5005
R4515 VGND.n1220 VGND.n789 4.5005
R4516 VGND.n1217 VGND.n1216 4.5005
R4517 VGND.n786 VGND.n785 4.5005
R4518 VGND.n823 VGND.n822 4.5005
R4519 VGND.n1122 VGND.n1121 4.5005
R4520 VGND.n1127 VGND.n680 4.5005
R4521 VGND.n812 VGND.n681 4.5005
R4522 VGND.n1140 VGND.n1139 4.5005
R4523 VGND.n1149 VGND.n1148 4.5005
R4524 VGND.n1159 VGND.n1158 4.5005
R4525 VGND.n1153 VGND.n804 4.5005
R4526 VGND.n1172 VGND.n1171 4.5005
R4527 VGND.n1181 VGND.n1180 4.5005
R4528 VGND.n1191 VGND.n1190 4.5005
R4529 VGND.n1185 VGND.n796 4.5005
R4530 VGND.n1204 VGND.n1203 4.5005
R4531 VGND.n1213 VGND.n1212 4.5005
R4532 VGND.n1223 VGND.n1222 4.5005
R4533 VGND.n788 VGND.n784 4.5005
R4534 VGND.n1234 VGND.n1233 4.5005
R4535 VGND.n1113 VGND.n1112 4.41365
R4536 VGND VGND.n3006 4.35375
R4537 VGND.n1090 VGND.n1089 4.05427
R4538 VGND.n583 VGND.n0 4.05427
R4539 VGND.n998 VGND.n997 4.05427
R4540 VGND.n1029 VGND.n1028 4.05427
R4541 VGND.n1060 VGND.n1059 4.05427
R4542 VGND VGND.n59 3.99438
R4543 VGND.n2920 VGND 3.99438
R4544 VGND.n2953 VGND 3.99438
R4545 VGND VGND.n2954 3.99437
R4546 VGND VGND.n28 3.99437
R4547 VGND.n1235 VGND.n274 3.77268
R4548 VGND.n3004 VGND.n3003 3.77268
R4549 VGND.n1120 VGND.n1119 3.77268
R4550 VGND.n2712 VGND.n2711 3.77268
R4551 VGND.n1282 VGND.n1281 3.77268
R4552 VGND.n2821 VGND.n188 3.77268
R4553 VGND.n1278 VGND.n687 3.77268
R4554 VGND.n2818 VGND.n2817 3.77268
R4555 VGND.n1273 VGND.n690 3.77268
R4556 VGND.n2816 VGND.n2815 3.77268
R4557 VGND.n1270 VGND.n693 3.77268
R4558 VGND.n2812 VGND.n2811 3.77268
R4559 VGND.n1265 VGND.n696 3.77268
R4560 VGND.n2810 VGND.n2809 3.77268
R4561 VGND.n1262 VGND.n699 3.77268
R4562 VGND.n2806 VGND.n2805 3.77268
R4563 VGND.n1257 VGND.n702 3.77268
R4564 VGND.n2804 VGND.n2803 3.77268
R4565 VGND.n1254 VGND.n705 3.77268
R4566 VGND.n2800 VGND.n2799 3.77268
R4567 VGND.n1249 VGND.n708 3.77268
R4568 VGND.n2798 VGND.n2797 3.77268
R4569 VGND.n1246 VGND.n711 3.77268
R4570 VGND.n2794 VGND.n2793 3.77268
R4571 VGND.n1241 VGND.n714 3.77268
R4572 VGND.n2792 VGND.n2791 3.77268
R4573 VGND.n1221 VGND.n280 3.77268
R4574 VGND.n2788 VGND.n2787 3.77268
R4575 VGND.n1237 VGND.n1236 3.77268
R4576 VGND.n2786 VGND.n2785 3.77268
R4577 VGND.n1284 VGND.n1283 3.77268
R4578 VGND.n2710 VGND.n184 3.77268
R4579 VGND.n2585 VGND.n2584 3.75914
R4580 VGND.n2590 VGND.n2587 3.75914
R4581 VGND.n1218 VGND.n786 3.75914
R4582 VGND.n823 VGND.n821 3.75914
R4583 VGND.n2585 VGND.n2570 3.4105
R4584 VGND.n2625 VGND.n2624 3.4105
R4585 VGND.n2623 VGND.n2622 3.4105
R4586 VGND.n2620 VGND.n2619 3.4105
R4587 VGND.n2617 VGND.n2616 3.4105
R4588 VGND.n2614 VGND.n2613 3.4105
R4589 VGND.n2611 VGND.n2610 3.4105
R4590 VGND.n2608 VGND.n2607 3.4105
R4591 VGND.n2605 VGND.n2604 3.4105
R4592 VGND.n2602 VGND.n2601 3.4105
R4593 VGND.n2599 VGND.n2598 3.4105
R4594 VGND.n2596 VGND.n2595 3.4105
R4595 VGND.n2593 VGND.n2592 3.4105
R4596 VGND.n2590 VGND.n2589 3.4105
R4597 VGND.n3004 VGND.n30 3.4105
R4598 VGND.n2786 VGND.n223 3.4105
R4599 VGND.n2787 VGND.n222 3.4105
R4600 VGND.n2792 VGND.n217 3.4105
R4601 VGND.n2793 VGND.n216 3.4105
R4602 VGND.n2798 VGND.n211 3.4105
R4603 VGND.n2799 VGND.n210 3.4105
R4604 VGND.n2804 VGND.n205 3.4105
R4605 VGND.n2805 VGND.n204 3.4105
R4606 VGND.n2810 VGND.n199 3.4105
R4607 VGND.n2811 VGND.n198 3.4105
R4608 VGND.n2816 VGND.n193 3.4105
R4609 VGND.n2817 VGND.n192 3.4105
R4610 VGND.n2626 VGND.n188 3.4105
R4611 VGND.n2710 VGND.n2709 3.4105
R4612 VGND.n2711 VGND.n2568 3.4105
R4613 VGND.n3003 VGND.n3002 3.4105
R4614 VGND.n2713 VGND.n2712 3.4105
R4615 VGND.n2518 VGND.n236 3.4105
R4616 VGND.n2492 VGND.n31 3.4105
R4617 VGND.n2823 VGND.n2822 3.4105
R4618 VGND.n2821 VGND.n2820 3.4105
R4619 VGND.n375 VGND.n187 3.4105
R4620 VGND.n640 VGND.n639 3.4105
R4621 VGND.n2431 VGND.n260 3.4105
R4622 VGND.n2166 VGND.n2165 3.4105
R4623 VGND.n2504 VGND.n191 3.4105
R4624 VGND.n2819 VGND.n2818 3.4105
R4625 VGND.n2164 VGND.n2163 3.4105
R4626 VGND.n2153 VGND.n2152 3.4105
R4627 VGND.n1435 VGND.n1434 3.4105
R4628 VGND.n2314 VGND.n325 3.4105
R4629 VGND.n2179 VGND.n2178 3.4105
R4630 VGND.n2177 VGND.n2176 3.4105
R4631 VGND.n2503 VGND.n194 3.4105
R4632 VGND.n2815 VGND.n2814 3.4105
R4633 VGND.n2148 VGND.n361 3.4105
R4634 VGND.n2149 VGND.n376 3.4105
R4635 VGND.n2151 VGND.n2150 3.4105
R4636 VGND.n1437 VGND.n1436 3.4105
R4637 VGND.n2126 VGND.n395 3.4105
R4638 VGND.n2147 VGND.n357 3.4105
R4639 VGND.n2190 VGND.n2189 3.4105
R4640 VGND.n2192 VGND.n2191 3.4105
R4641 VGND.n2502 VGND.n197 3.4105
R4642 VGND.n2813 VGND.n2812 3.4105
R4643 VGND.n2018 VGND.n2017 3.4105
R4644 VGND.n2003 VGND.n2002 3.4105
R4645 VGND.n1992 VGND.n1991 3.4105
R4646 VGND.n630 VGND.n380 3.4105
R4647 VGND.n1415 VGND.n638 3.4105
R4648 VGND.n2123 VGND.n396 3.4105
R4649 VGND.n2029 VGND.n2028 3.4105
R4650 VGND.n2146 VGND.n353 3.4105
R4651 VGND.n2205 VGND.n2204 3.4105
R4652 VGND.n2203 VGND.n2202 3.4105
R4653 VGND.n2501 VGND.n200 3.4105
R4654 VGND.n2809 VGND.n2808 3.4105
R4655 VGND.n2031 VGND.n2030 3.4105
R4656 VGND.n2016 VGND.n2015 3.4105
R4657 VGND.n2005 VGND.n2004 3.4105
R4658 VGND.n1990 VGND.n1989 3.4105
R4659 VGND.n1979 VGND.n1978 3.4105
R4660 VGND.n1413 VGND.n1412 3.4105
R4661 VGND.n2339 VGND.n313 3.4105
R4662 VGND.n2042 VGND.n2041 3.4105
R4663 VGND.n2044 VGND.n2043 3.4105
R4664 VGND.n2145 VGND.n349 3.4105
R4665 VGND.n2216 VGND.n2215 3.4105
R4666 VGND.n2218 VGND.n2217 3.4105
R4667 VGND.n2500 VGND.n203 3.4105
R4668 VGND.n2807 VGND.n2806 3.4105
R4669 VGND.n1971 VGND.n416 3.4105
R4670 VGND.n1972 VGND.n420 3.4105
R4671 VGND.n1973 VGND.n424 3.4105
R4672 VGND.n1974 VGND.n428 3.4105
R4673 VGND.n1975 VGND.n432 3.4105
R4674 VGND.n1977 VGND.n1976 3.4105
R4675 VGND.n1411 VGND.n1410 3.4105
R4676 VGND.n1952 VGND.n451 3.4105
R4677 VGND.n1970 VGND.n412 3.4105
R4678 VGND.n2057 VGND.n2056 3.4105
R4679 VGND.n2055 VGND.n2054 3.4105
R4680 VGND.n2144 VGND.n345 3.4105
R4681 VGND.n2231 VGND.n2230 3.4105
R4682 VGND.n2229 VGND.n2228 3.4105
R4683 VGND.n2499 VGND.n206 3.4105
R4684 VGND.n2803 VGND.n2802 3.4105
R4685 VGND.n1881 VGND.n1880 3.4105
R4686 VGND.n1870 VGND.n1869 3.4105
R4687 VGND.n1855 VGND.n1854 3.4105
R4688 VGND.n1844 VGND.n1843 3.4105
R4689 VGND.n1829 VGND.n1828 3.4105
R4690 VGND.n1818 VGND.n1817 3.4105
R4691 VGND.n1405 VGND.n436 3.4105
R4692 VGND.n1390 VGND.n657 3.4105
R4693 VGND.n1949 VGND.n452 3.4105
R4694 VGND.n1896 VGND.n1895 3.4105
R4695 VGND.n1969 VGND.n408 3.4105
R4696 VGND.n2068 VGND.n2067 3.4105
R4697 VGND.n2070 VGND.n2069 3.4105
R4698 VGND.n2143 VGND.n341 3.4105
R4699 VGND.n2242 VGND.n2241 3.4105
R4700 VGND.n2244 VGND.n2243 3.4105
R4701 VGND.n2498 VGND.n209 3.4105
R4702 VGND.n2801 VGND.n2800 3.4105
R4703 VGND.n1894 VGND.n1893 3.4105
R4704 VGND.n1883 VGND.n1882 3.4105
R4705 VGND.n1868 VGND.n1867 3.4105
R4706 VGND.n1857 VGND.n1856 3.4105
R4707 VGND.n1842 VGND.n1841 3.4105
R4708 VGND.n1831 VGND.n1830 3.4105
R4709 VGND.n1816 VGND.n1815 3.4105
R4710 VGND.n1805 VGND.n1804 3.4105
R4711 VGND.n1387 VGND.n1386 3.4105
R4712 VGND.n2364 VGND.n301 3.4105
R4713 VGND.n1909 VGND.n1908 3.4105
R4714 VGND.n1907 VGND.n1906 3.4105
R4715 VGND.n1968 VGND.n404 3.4105
R4716 VGND.n2083 VGND.n2082 3.4105
R4717 VGND.n2081 VGND.n2080 3.4105
R4718 VGND.n2142 VGND.n337 3.4105
R4719 VGND.n2257 VGND.n2256 3.4105
R4720 VGND.n2255 VGND.n2254 3.4105
R4721 VGND.n2497 VGND.n212 3.4105
R4722 VGND.n2797 VGND.n2796 3.4105
R4723 VGND.n1794 VGND.n460 3.4105
R4724 VGND.n1795 VGND.n464 3.4105
R4725 VGND.n1796 VGND.n468 3.4105
R4726 VGND.n1797 VGND.n472 3.4105
R4727 VGND.n1798 VGND.n476 3.4105
R4728 VGND.n1799 VGND.n480 3.4105
R4729 VGND.n1800 VGND.n484 3.4105
R4730 VGND.n1801 VGND.n488 3.4105
R4731 VGND.n1803 VGND.n1802 3.4105
R4732 VGND.n1369 VGND.n570 3.4105
R4733 VGND.n1778 VGND.n507 3.4105
R4734 VGND.n1793 VGND.n456 3.4105
R4735 VGND.n1925 VGND.n1924 3.4105
R4736 VGND.n1927 VGND.n1926 3.4105
R4737 VGND.n1967 VGND.n400 3.4105
R4738 VGND.n2099 VGND.n2098 3.4105
R4739 VGND.n2101 VGND.n2100 3.4105
R4740 VGND.n2141 VGND.n333 3.4105
R4741 VGND.n2273 VGND.n2272 3.4105
R4742 VGND.n2275 VGND.n2274 3.4105
R4743 VGND.n2496 VGND.n215 3.4105
R4744 VGND.n2795 VGND.n2794 3.4105
R4745 VGND.n1753 VGND.n1752 3.4105
R4746 VGND.n1733 VGND.n1732 3.4105
R4747 VGND.n1722 VGND.n1721 3.4105
R4748 VGND.n1707 VGND.n1706 3.4105
R4749 VGND.n1696 VGND.n1695 3.4105
R4750 VGND.n1681 VGND.n1680 3.4105
R4751 VGND.n1670 VGND.n1669 3.4105
R4752 VGND.n1655 VGND.n1654 3.4105
R4753 VGND.n1644 VGND.n1643 3.4105
R4754 VGND.n1527 VGND.n492 3.4105
R4755 VGND.n1530 VGND.n1529 3.4105
R4756 VGND.n1775 VGND.n508 3.4105
R4757 VGND.n2374 VGND.n2373 3.4105
R4758 VGND.n1792 VGND.n293 3.4105
R4759 VGND.n2351 VGND.n2350 3.4105
R4760 VGND.n2349 VGND.n2348 3.4105
R4761 VGND.n1966 VGND.n305 3.4105
R4762 VGND.n2326 VGND.n2325 3.4105
R4763 VGND.n2324 VGND.n2323 3.4105
R4764 VGND.n2140 VGND.n317 3.4105
R4765 VGND.n2301 VGND.n2300 3.4105
R4766 VGND.n2299 VGND.n2298 3.4105
R4767 VGND.n2495 VGND.n218 3.4105
R4768 VGND.n2791 VGND.n2790 3.4105
R4769 VGND.n2376 VGND.n2375 3.4105
R4770 VGND.n1751 VGND.n1750 3.4105
R4771 VGND.n1735 VGND.n1734 3.4105
R4772 VGND.n1720 VGND.n1719 3.4105
R4773 VGND.n1709 VGND.n1708 3.4105
R4774 VGND.n1694 VGND.n1693 3.4105
R4775 VGND.n1683 VGND.n1682 3.4105
R4776 VGND.n1668 VGND.n1667 3.4105
R4777 VGND.n1657 VGND.n1656 3.4105
R4778 VGND.n1642 VGND.n1641 3.4105
R4779 VGND.n1631 VGND.n1630 3.4105
R4780 VGND.n1532 VGND.n1531 3.4105
R4781 VGND.n2389 VGND.n288 3.4105
R4782 VGND.n2377 VGND.n281 3.4105
R4783 VGND.n2372 VGND.n2371 3.4105
R4784 VGND.n2370 VGND.n2369 3.4105
R4785 VGND.n2352 VGND.n296 3.4105
R4786 VGND.n2347 VGND.n2346 3.4105
R4787 VGND.n2345 VGND.n2344 3.4105
R4788 VGND.n2327 VGND.n308 3.4105
R4789 VGND.n2322 VGND.n2321 3.4105
R4790 VGND.n2320 VGND.n2319 3.4105
R4791 VGND.n2302 VGND.n320 3.4105
R4792 VGND.n2297 VGND.n2296 3.4105
R4793 VGND.n2494 VGND.n221 3.4105
R4794 VGND.n2789 VGND.n2788 3.4105
R4795 VGND.n2395 VGND.n2394 3.4105
R4796 VGND.n1618 VGND.n292 3.4105
R4797 VGND.n1619 VGND.n512 3.4105
R4798 VGND.n1620 VGND.n516 3.4105
R4799 VGND.n1621 VGND.n520 3.4105
R4800 VGND.n1622 VGND.n524 3.4105
R4801 VGND.n1623 VGND.n528 3.4105
R4802 VGND.n1624 VGND.n532 3.4105
R4803 VGND.n1625 VGND.n536 3.4105
R4804 VGND.n1626 VGND.n540 3.4105
R4805 VGND.n1627 VGND.n544 3.4105
R4806 VGND.n1629 VGND.n1628 3.4105
R4807 VGND.n1299 VGND.n569 3.4105
R4808 VGND.n1604 VGND.n1603 3.4105
R4809 VGND.n2393 VGND.n2392 3.4105
R4810 VGND.n2391 VGND.n2390 3.4105
R4811 VGND.n510 VGND.n286 3.4105
R4812 VGND.n2368 VGND.n2367 3.4105
R4813 VGND.n2366 VGND.n2365 3.4105
R4814 VGND.n454 VGND.n299 3.4105
R4815 VGND.n2343 VGND.n2342 3.4105
R4816 VGND.n2341 VGND.n2340 3.4105
R4817 VGND.n398 VGND.n311 3.4105
R4818 VGND.n2318 VGND.n2317 3.4105
R4819 VGND.n2316 VGND.n2315 3.4105
R4820 VGND.n2295 VGND.n323 3.4105
R4821 VGND.n2493 VGND.n224 3.4105
R4822 VGND.n2785 VGND.n2784 3.4105
R4823 VGND.n285 VGND.n284 3.4105
R4824 VGND.n2397 VGND.n2396 3.4105
R4825 VGND.n1243 VGND.n1242 3.4105
R4826 VGND.n1245 VGND.n1244 3.4105
R4827 VGND.n1251 VGND.n1250 3.4105
R4828 VGND.n1253 VGND.n1252 3.4105
R4829 VGND.n1259 VGND.n1258 3.4105
R4830 VGND.n1261 VGND.n1260 3.4105
R4831 VGND.n1267 VGND.n1266 3.4105
R4832 VGND.n1269 VGND.n1268 3.4105
R4833 VGND.n1275 VGND.n1274 3.4105
R4834 VGND.n1277 VGND.n1276 3.4105
R4835 VGND.n894 VGND.n548 3.4105
R4836 VGND.n897 VGND.n896 3.4105
R4837 VGND.n2409 VGND.n277 3.4105
R4838 VGND.n895 VGND.n562 3.4105
R4839 VGND.n1545 VGND.n1544 3.4105
R4840 VGND.n1543 VGND.n1542 3.4105
R4841 VGND.n1528 VGND.n563 3.4105
R4842 VGND.n1368 VGND.n1367 3.4105
R4843 VGND.n1385 VGND.n662 3.4105
R4844 VGND.n1407 VGND.n1406 3.4105
R4845 VGND.n1409 VGND.n1408 3.4105
R4846 VGND.n656 VGND.n631 3.4105
R4847 VGND.n1500 VGND.n1499 3.4105
R4848 VGND.n1498 VGND.n1497 3.4105
R4849 VGND.n1433 VGND.n183 3.4105
R4850 VGND.n2827 VGND.n2826 3.4105
R4851 VGND.n2825 VGND.n2824 3.4105
R4852 VGND.n2714 VGND.n184 3.4105
R4853 VGND.n1236 VGND.n784 3.4105
R4854 VGND.n1222 VGND.n1221 3.4105
R4855 VGND.n1213 VGND.n714 3.4105
R4856 VGND.n1203 VGND.n711 3.4105
R4857 VGND.n1185 VGND.n708 3.4105
R4858 VGND.n1190 VGND.n705 3.4105
R4859 VGND.n1181 VGND.n702 3.4105
R4860 VGND.n1171 VGND.n699 3.4105
R4861 VGND.n1153 VGND.n696 3.4105
R4862 VGND.n1158 VGND.n693 3.4105
R4863 VGND.n1149 VGND.n690 3.4105
R4864 VGND.n1139 VGND.n687 3.4105
R4865 VGND.n1282 VGND.n681 3.4105
R4866 VGND.n1283 VGND.n680 3.4105
R4867 VGND.n1235 VGND.n1234 3.4105
R4868 VGND.n1218 VGND.n1217 3.4105
R4869 VGND.n1220 VGND.n1219 3.4105
R4870 VGND.n1215 VGND.n1214 3.4105
R4871 VGND.n1202 VGND.n790 3.4105
R4872 VGND.n1187 VGND.n1186 3.4105
R4873 VGND.n1189 VGND.n1188 3.4105
R4874 VGND.n1183 VGND.n1182 3.4105
R4875 VGND.n1170 VGND.n798 3.4105
R4876 VGND.n1155 VGND.n1154 3.4105
R4877 VGND.n1157 VGND.n1156 3.4105
R4878 VGND.n1151 VGND.n1150 3.4105
R4879 VGND.n1138 VGND.n806 3.4105
R4880 VGND.n818 VGND.n817 3.4105
R4881 VGND.n821 VGND.n820 3.4105
R4882 VGND.n1121 VGND.n1120 3.4105
R4883 VGND.n1238 VGND.n1237 3.4105
R4884 VGND.n1239 VGND.n280 3.4105
R4885 VGND.n1241 VGND.n1240 3.4105
R4886 VGND.n1247 VGND.n1246 3.4105
R4887 VGND.n1249 VGND.n1248 3.4105
R4888 VGND.n1255 VGND.n1254 3.4105
R4889 VGND.n1257 VGND.n1256 3.4105
R4890 VGND.n1263 VGND.n1262 3.4105
R4891 VGND.n1265 VGND.n1264 3.4105
R4892 VGND.n1271 VGND.n1270 3.4105
R4893 VGND.n1273 VGND.n1272 3.4105
R4894 VGND.n1279 VGND.n1278 3.4105
R4895 VGND.n1281 VGND.n1280 3.4105
R4896 VGND.n1285 VGND.n1284 3.4105
R4897 VGND.n1119 VGND.n1118 3.4105
R4898 VGND.n2412 VGND.n274 3.4105
R4899 VGND.n980 VGND.n969 3.01226
R4900 VGND.n74 VGND.n73 3.01226
R4901 VGND.n964 VGND.n899 2.63579
R4902 VGND.n2524 VGND 2.52282
R4903 VGND.n2527 VGND 2.52282
R4904 VGND.n2530 VGND 2.52282
R4905 VGND.n2533 VGND 2.52282
R4906 VGND.n2536 VGND 2.52282
R4907 VGND.n2539 VGND 2.52282
R4908 VGND.n2542 VGND 2.52282
R4909 VGND.n2545 VGND 2.52282
R4910 VGND.n2548 VGND 2.52282
R4911 VGND.n2551 VGND 2.52282
R4912 VGND.n2554 VGND 2.52282
R4913 VGND.n2557 VGND 2.52282
R4914 VGND.n2560 VGND 2.52282
R4915 VGND.n2563 VGND 2.52282
R4916 VGND.n2566 VGND 2.52282
R4917 VGND.n985 VGND.n984 2.25932
R4918 VGND.n105 VGND.n104 2.25932
R4919 VGND.n2865 VGND.n2864 2.25932
R4920 VGND.n2897 VGND.n2896 2.25932
R4921 VGND.n83 VGND.n62 2.25932
R4922 VGND.n79 VGND.n78 2.25932
R4923 VGND.n135 VGND.n123 1.88285
R4924 VGND.n603 VGND.n591 1.88285
R4925 VGND.n165 VGND.n153 1.88285
R4926 VGND.n2567 VGND 1.79514
R4927 VGND.n1115 VGND.n275 1.75987
R4928 VGND.n2567 VGND 1.57193
R4929 VGND.n3005 VGND.n3004 1.54254
R4930 VGND.n3002 VGND.n29 1.54254
R4931 VGND.n2492 VGND.n2433 1.54254
R4932 VGND.n2432 VGND.n2431 1.54254
R4933 VGND.n2314 VGND.n259 1.54254
R4934 VGND.n2126 VGND.n2125 1.54254
R4935 VGND.n2124 VGND.n2123 1.54254
R4936 VGND.n2339 VGND.n314 1.54254
R4937 VGND.n1952 VGND.n1951 1.54254
R4938 VGND.n1950 VGND.n1949 1.54254
R4939 VGND.n2364 VGND.n302 1.54254
R4940 VGND.n1778 VGND.n1777 1.54254
R4941 VGND.n1776 VGND.n1775 1.54254
R4942 VGND.n2389 VGND.n289 1.54254
R4943 VGND.n1604 VGND.n276 1.54254
R4944 VGND.n2410 VGND.n2409 1.54254
R4945 VGND.n1235 VGND.n275 1.54254
R4946 VGND.n2412 VGND.n2411 1.54254
R4947 VGND.n992 VGND.n898 1.50638
R4948 VGND.n2916 VGND.n2915 1.50638
R4949 VGND VGND.n2521 1.3946
R4950 VGND.n2520 VGND 1.3946
R4951 VGND.n2519 VGND 1.3946
R4952 VGND VGND.n237 1.3946
R4953 VGND VGND.n1418 1.3946
R4954 VGND.n1417 VGND 1.3946
R4955 VGND.n1416 VGND 1.3946
R4956 VGND.n1414 VGND 1.3946
R4957 VGND VGND.n641 1.3946
R4958 VGND VGND.n1389 1.3946
R4959 VGND.n1388 VGND 1.3946
R4960 VGND.n1370 VGND 1.3946
R4961 VGND.n1302 VGND 1.3946
R4962 VGND.n1301 VGND 1.3946
R4963 VGND.n1300 VGND 1.3946
R4964 VGND VGND.n669 1.3946
R4965 VGND.n1116 VGND 1.3946
R4966 VGND VGND.n1117 1.3946
R4967 VGND.n2709 VGND.n2570 1.00149
R4968 VGND.n2626 VGND.n2625 1.00149
R4969 VGND.n2622 VGND.n192 1.00149
R4970 VGND.n2619 VGND.n193 1.00149
R4971 VGND.n2616 VGND.n198 1.00149
R4972 VGND.n2613 VGND.n199 1.00149
R4973 VGND.n2610 VGND.n204 1.00149
R4974 VGND.n2607 VGND.n205 1.00149
R4975 VGND.n2604 VGND.n210 1.00149
R4976 VGND.n2601 VGND.n211 1.00149
R4977 VGND.n2598 VGND.n216 1.00149
R4978 VGND.n2595 VGND.n217 1.00149
R4979 VGND.n2592 VGND.n222 1.00149
R4980 VGND.n2589 VGND.n223 1.00149
R4981 VGND.n2587 VGND.n30 1.00149
R4982 VGND.n820 VGND.n680 1.00149
R4983 VGND.n817 VGND.n681 1.00149
R4984 VGND.n1139 VGND.n1138 1.00149
R4985 VGND.n1150 VGND.n1149 1.00149
R4986 VGND.n1158 VGND.n1157 1.00149
R4987 VGND.n1154 VGND.n1153 1.00149
R4988 VGND.n1171 VGND.n1170 1.00149
R4989 VGND.n1182 VGND.n1181 1.00149
R4990 VGND.n1190 VGND.n1189 1.00149
R4991 VGND.n1186 VGND.n1185 1.00149
R4992 VGND.n1203 VGND.n1202 1.00149
R4993 VGND.n1214 VGND.n1213 1.00149
R4994 VGND.n1222 VGND.n1220 1.00149
R4995 VGND.n1217 VGND.n784 1.00149
R4996 VGND.n1234 VGND.n786 1.00149
R4997 VGND.n1121 VGND.n823 1.00149
R4998 VGND.n2584 VGND.n2568 0.973133
R4999 VGND.n2835 VGND.n2 0.9305
R5000 VGND.n97 VGND.n93 0.929432
R5001 VGND.n2857 VGND.n2853 0.929432
R5002 VGND.n2889 VGND.n2885 0.929432
R5003 VGND.n70 VGND.n68 0.929432
R5004 VGND.n59 VGND.n1 0.916608
R5005 VGND VGND.n2524 0.839786
R5006 VGND VGND.n2527 0.839786
R5007 VGND VGND.n2530 0.839786
R5008 VGND VGND.n2533 0.839786
R5009 VGND VGND.n2536 0.839786
R5010 VGND VGND.n2539 0.839786
R5011 VGND VGND.n2542 0.839786
R5012 VGND VGND.n2545 0.839786
R5013 VGND VGND.n2548 0.839786
R5014 VGND VGND.n2551 0.839786
R5015 VGND VGND.n2554 0.839786
R5016 VGND VGND.n2557 0.839786
R5017 VGND VGND.n2560 0.839786
R5018 VGND VGND.n2563 0.839786
R5019 VGND VGND.n2566 0.839786
R5020 VGND.n3022 VGND.n3021 0.7755
R5021 VGND.n3023 VGND.n3022 0.774207
R5022 VGND.n117 VGND.n115 0.753441
R5023 VGND.n16 VGND.n14 0.753441
R5024 VGND.n45 VGND.n43 0.753441
R5025 VGND.n2869 VGND.n2846 0.753441
R5026 VGND.n2932 VGND.n2929 0.753441
R5027 VGND.n2974 VGND.n2972 0.753441
R5028 VGND.n1114 VGND.t922 0.632121
R5029 VGND.n1114 VGND.n1113 0.579775
R5030 VGND.n3025 VGND.n3024 0.573119
R5031 VGND VGND.n0 0.542567
R5032 VGND.n3025 VGND.n1 0.507317
R5033 VGND.n1115 VGND.n1114 0.4658
R5034 VGND.n3006 VGND.n3005 0.404308
R5035 VGND.n1096 VGND.n1093 0.376971
R5036 VGND.n1068 VGND.n1064 0.376971
R5037 VGND.n992 VGND.n991 0.376971
R5038 VGND.n1006 VGND.n1002 0.376971
R5039 VGND.n1037 VGND.n1033 0.376971
R5040 VGND.n84 VGND.n83 0.376971
R5041 VGND.n2915 VGND.n61 0.376971
R5042 VGND VGND.n3025 0.37415
R5043 VGND.n277 VGND.n274 0.362676
R5044 VGND.n1603 VGND.n277 0.362676
R5045 VGND.n1603 VGND.n288 0.362676
R5046 VGND.n508 VGND.n288 0.362676
R5047 VGND.n508 VGND.n507 0.362676
R5048 VGND.n507 VGND.n301 0.362676
R5049 VGND.n452 VGND.n301 0.362676
R5050 VGND.n452 VGND.n451 0.362676
R5051 VGND.n451 VGND.n313 0.362676
R5052 VGND.n396 VGND.n313 0.362676
R5053 VGND.n396 VGND.n395 0.362676
R5054 VGND.n395 VGND.n325 0.362676
R5055 VGND.n325 VGND.n260 0.362676
R5056 VGND.n260 VGND.n31 0.362676
R5057 VGND.n3003 VGND.n31 0.362676
R5058 VGND.n1119 VGND.n897 0.362676
R5059 VGND.n897 VGND.n569 0.362676
R5060 VGND.n1531 VGND.n569 0.362676
R5061 VGND.n1531 VGND.n1530 0.362676
R5062 VGND.n1530 VGND.n570 0.362676
R5063 VGND.n1386 VGND.n570 0.362676
R5064 VGND.n1386 VGND.n657 0.362676
R5065 VGND.n1411 VGND.n657 0.362676
R5066 VGND.n1412 VGND.n1411 0.362676
R5067 VGND.n1412 VGND.n638 0.362676
R5068 VGND.n1436 VGND.n638 0.362676
R5069 VGND.n1436 VGND.n1435 0.362676
R5070 VGND.n1435 VGND.n640 0.362676
R5071 VGND.n640 VGND.n236 0.362676
R5072 VGND.n2712 VGND.n236 0.362676
R5073 VGND.n1281 VGND.n548 0.362676
R5074 VGND.n1629 VGND.n548 0.362676
R5075 VGND.n1630 VGND.n1629 0.362676
R5076 VGND.n1630 VGND.n492 0.362676
R5077 VGND.n1803 VGND.n492 0.362676
R5078 VGND.n1804 VGND.n1803 0.362676
R5079 VGND.n1804 VGND.n436 0.362676
R5080 VGND.n1977 VGND.n436 0.362676
R5081 VGND.n1978 VGND.n1977 0.362676
R5082 VGND.n1978 VGND.n380 0.362676
R5083 VGND.n2151 VGND.n380 0.362676
R5084 VGND.n2152 VGND.n2151 0.362676
R5085 VGND.n2152 VGND.n187 0.362676
R5086 VGND.n2822 VGND.n187 0.362676
R5087 VGND.n2822 VGND.n2821 0.362676
R5088 VGND.n1278 VGND.n1277 0.362676
R5089 VGND.n1277 VGND.n544 0.362676
R5090 VGND.n1642 VGND.n544 0.362676
R5091 VGND.n1643 VGND.n1642 0.362676
R5092 VGND.n1643 VGND.n488 0.362676
R5093 VGND.n1816 VGND.n488 0.362676
R5094 VGND.n1817 VGND.n1816 0.362676
R5095 VGND.n1817 VGND.n432 0.362676
R5096 VGND.n1990 VGND.n432 0.362676
R5097 VGND.n1991 VGND.n1990 0.362676
R5098 VGND.n1991 VGND.n376 0.362676
R5099 VGND.n2164 VGND.n376 0.362676
R5100 VGND.n2165 VGND.n2164 0.362676
R5101 VGND.n2165 VGND.n191 0.362676
R5102 VGND.n2818 VGND.n191 0.362676
R5103 VGND.n1274 VGND.n1273 0.362676
R5104 VGND.n1274 VGND.n540 0.362676
R5105 VGND.n1656 VGND.n540 0.362676
R5106 VGND.n1656 VGND.n1655 0.362676
R5107 VGND.n1655 VGND.n484 0.362676
R5108 VGND.n1830 VGND.n484 0.362676
R5109 VGND.n1830 VGND.n1829 0.362676
R5110 VGND.n1829 VGND.n428 0.362676
R5111 VGND.n2004 VGND.n428 0.362676
R5112 VGND.n2004 VGND.n2003 0.362676
R5113 VGND.n2003 VGND.n361 0.362676
R5114 VGND.n2178 VGND.n361 0.362676
R5115 VGND.n2178 VGND.n2177 0.362676
R5116 VGND.n2177 VGND.n194 0.362676
R5117 VGND.n2815 VGND.n194 0.362676
R5118 VGND.n1270 VGND.n1269 0.362676
R5119 VGND.n1269 VGND.n536 0.362676
R5120 VGND.n1668 VGND.n536 0.362676
R5121 VGND.n1669 VGND.n1668 0.362676
R5122 VGND.n1669 VGND.n480 0.362676
R5123 VGND.n1842 VGND.n480 0.362676
R5124 VGND.n1843 VGND.n1842 0.362676
R5125 VGND.n1843 VGND.n424 0.362676
R5126 VGND.n2016 VGND.n424 0.362676
R5127 VGND.n2017 VGND.n2016 0.362676
R5128 VGND.n2017 VGND.n357 0.362676
R5129 VGND.n2190 VGND.n357 0.362676
R5130 VGND.n2191 VGND.n2190 0.362676
R5131 VGND.n2191 VGND.n197 0.362676
R5132 VGND.n2812 VGND.n197 0.362676
R5133 VGND.n1266 VGND.n1265 0.362676
R5134 VGND.n1266 VGND.n532 0.362676
R5135 VGND.n1682 VGND.n532 0.362676
R5136 VGND.n1682 VGND.n1681 0.362676
R5137 VGND.n1681 VGND.n476 0.362676
R5138 VGND.n1856 VGND.n476 0.362676
R5139 VGND.n1856 VGND.n1855 0.362676
R5140 VGND.n1855 VGND.n420 0.362676
R5141 VGND.n2030 VGND.n420 0.362676
R5142 VGND.n2030 VGND.n2029 0.362676
R5143 VGND.n2029 VGND.n353 0.362676
R5144 VGND.n2204 VGND.n353 0.362676
R5145 VGND.n2204 VGND.n2203 0.362676
R5146 VGND.n2203 VGND.n200 0.362676
R5147 VGND.n2809 VGND.n200 0.362676
R5148 VGND.n1262 VGND.n1261 0.362676
R5149 VGND.n1261 VGND.n528 0.362676
R5150 VGND.n1694 VGND.n528 0.362676
R5151 VGND.n1695 VGND.n1694 0.362676
R5152 VGND.n1695 VGND.n472 0.362676
R5153 VGND.n1868 VGND.n472 0.362676
R5154 VGND.n1869 VGND.n1868 0.362676
R5155 VGND.n1869 VGND.n416 0.362676
R5156 VGND.n2042 VGND.n416 0.362676
R5157 VGND.n2043 VGND.n2042 0.362676
R5158 VGND.n2043 VGND.n349 0.362676
R5159 VGND.n2216 VGND.n349 0.362676
R5160 VGND.n2217 VGND.n2216 0.362676
R5161 VGND.n2217 VGND.n203 0.362676
R5162 VGND.n2806 VGND.n203 0.362676
R5163 VGND.n1258 VGND.n1257 0.362676
R5164 VGND.n1258 VGND.n524 0.362676
R5165 VGND.n1708 VGND.n524 0.362676
R5166 VGND.n1708 VGND.n1707 0.362676
R5167 VGND.n1707 VGND.n468 0.362676
R5168 VGND.n1882 VGND.n468 0.362676
R5169 VGND.n1882 VGND.n1881 0.362676
R5170 VGND.n1881 VGND.n412 0.362676
R5171 VGND.n2056 VGND.n412 0.362676
R5172 VGND.n2056 VGND.n2055 0.362676
R5173 VGND.n2055 VGND.n345 0.362676
R5174 VGND.n2230 VGND.n345 0.362676
R5175 VGND.n2230 VGND.n2229 0.362676
R5176 VGND.n2229 VGND.n206 0.362676
R5177 VGND.n2803 VGND.n206 0.362676
R5178 VGND.n1254 VGND.n1253 0.362676
R5179 VGND.n1253 VGND.n520 0.362676
R5180 VGND.n1720 VGND.n520 0.362676
R5181 VGND.n1721 VGND.n1720 0.362676
R5182 VGND.n1721 VGND.n464 0.362676
R5183 VGND.n1894 VGND.n464 0.362676
R5184 VGND.n1895 VGND.n1894 0.362676
R5185 VGND.n1895 VGND.n408 0.362676
R5186 VGND.n2068 VGND.n408 0.362676
R5187 VGND.n2069 VGND.n2068 0.362676
R5188 VGND.n2069 VGND.n341 0.362676
R5189 VGND.n2242 VGND.n341 0.362676
R5190 VGND.n2243 VGND.n2242 0.362676
R5191 VGND.n2243 VGND.n209 0.362676
R5192 VGND.n2800 VGND.n209 0.362676
R5193 VGND.n1250 VGND.n1249 0.362676
R5194 VGND.n1250 VGND.n516 0.362676
R5195 VGND.n1734 VGND.n516 0.362676
R5196 VGND.n1734 VGND.n1733 0.362676
R5197 VGND.n1733 VGND.n460 0.362676
R5198 VGND.n1908 VGND.n460 0.362676
R5199 VGND.n1908 VGND.n1907 0.362676
R5200 VGND.n1907 VGND.n404 0.362676
R5201 VGND.n2082 VGND.n404 0.362676
R5202 VGND.n2082 VGND.n2081 0.362676
R5203 VGND.n2081 VGND.n337 0.362676
R5204 VGND.n2256 VGND.n337 0.362676
R5205 VGND.n2256 VGND.n2255 0.362676
R5206 VGND.n2255 VGND.n212 0.362676
R5207 VGND.n2797 VGND.n212 0.362676
R5208 VGND.n1246 VGND.n1245 0.362676
R5209 VGND.n1245 VGND.n512 0.362676
R5210 VGND.n1751 VGND.n512 0.362676
R5211 VGND.n1752 VGND.n1751 0.362676
R5212 VGND.n1752 VGND.n456 0.362676
R5213 VGND.n1925 VGND.n456 0.362676
R5214 VGND.n1926 VGND.n1925 0.362676
R5215 VGND.n1926 VGND.n400 0.362676
R5216 VGND.n2099 VGND.n400 0.362676
R5217 VGND.n2100 VGND.n2099 0.362676
R5218 VGND.n2100 VGND.n333 0.362676
R5219 VGND.n2273 VGND.n333 0.362676
R5220 VGND.n2274 VGND.n2273 0.362676
R5221 VGND.n2274 VGND.n215 0.362676
R5222 VGND.n2794 VGND.n215 0.362676
R5223 VGND.n1242 VGND.n1241 0.362676
R5224 VGND.n1242 VGND.n292 0.362676
R5225 VGND.n2375 VGND.n292 0.362676
R5226 VGND.n2375 VGND.n2374 0.362676
R5227 VGND.n2374 VGND.n293 0.362676
R5228 VGND.n2350 VGND.n293 0.362676
R5229 VGND.n2350 VGND.n2349 0.362676
R5230 VGND.n2349 VGND.n305 0.362676
R5231 VGND.n2325 VGND.n305 0.362676
R5232 VGND.n2325 VGND.n2324 0.362676
R5233 VGND.n2324 VGND.n317 0.362676
R5234 VGND.n2300 VGND.n317 0.362676
R5235 VGND.n2300 VGND.n2299 0.362676
R5236 VGND.n2299 VGND.n218 0.362676
R5237 VGND.n2791 VGND.n218 0.362676
R5238 VGND.n2396 VGND.n280 0.362676
R5239 VGND.n2396 VGND.n2395 0.362676
R5240 VGND.n2395 VGND.n281 0.362676
R5241 VGND.n2371 VGND.n281 0.362676
R5242 VGND.n2371 VGND.n2370 0.362676
R5243 VGND.n2370 VGND.n296 0.362676
R5244 VGND.n2346 VGND.n296 0.362676
R5245 VGND.n2346 VGND.n2345 0.362676
R5246 VGND.n2345 VGND.n308 0.362676
R5247 VGND.n2321 VGND.n308 0.362676
R5248 VGND.n2321 VGND.n2320 0.362676
R5249 VGND.n2320 VGND.n320 0.362676
R5250 VGND.n2296 VGND.n320 0.362676
R5251 VGND.n2296 VGND.n221 0.362676
R5252 VGND.n2788 VGND.n221 0.362676
R5253 VGND.n1237 VGND.n285 0.362676
R5254 VGND.n2392 VGND.n285 0.362676
R5255 VGND.n2392 VGND.n2391 0.362676
R5256 VGND.n2391 VGND.n286 0.362676
R5257 VGND.n2367 VGND.n286 0.362676
R5258 VGND.n2367 VGND.n2366 0.362676
R5259 VGND.n2366 VGND.n299 0.362676
R5260 VGND.n2342 VGND.n299 0.362676
R5261 VGND.n2342 VGND.n2341 0.362676
R5262 VGND.n2341 VGND.n311 0.362676
R5263 VGND.n2317 VGND.n311 0.362676
R5264 VGND.n2317 VGND.n2316 0.362676
R5265 VGND.n2316 VGND.n323 0.362676
R5266 VGND.n323 VGND.n224 0.362676
R5267 VGND.n2785 VGND.n224 0.362676
R5268 VGND.n1284 VGND.n562 0.362676
R5269 VGND.n1544 VGND.n562 0.362676
R5270 VGND.n1544 VGND.n1543 0.362676
R5271 VGND.n1543 VGND.n563 0.362676
R5272 VGND.n1367 VGND.n563 0.362676
R5273 VGND.n1367 VGND.n662 0.362676
R5274 VGND.n1407 VGND.n662 0.362676
R5275 VGND.n1408 VGND.n1407 0.362676
R5276 VGND.n1408 VGND.n631 0.362676
R5277 VGND.n1499 VGND.n631 0.362676
R5278 VGND.n1499 VGND.n1498 0.362676
R5279 VGND.n1498 VGND.n183 0.362676
R5280 VGND.n2826 VGND.n183 0.362676
R5281 VGND.n2826 VGND.n2825 0.362676
R5282 VGND.n2825 VGND.n184 0.362676
R5283 VGND.n2624 VGND.n2585 0.349144
R5284 VGND.n2624 VGND.n2623 0.349144
R5285 VGND.n2623 VGND.n2620 0.349144
R5286 VGND.n2620 VGND.n2617 0.349144
R5287 VGND.n2617 VGND.n2614 0.349144
R5288 VGND.n2614 VGND.n2611 0.349144
R5289 VGND.n2611 VGND.n2608 0.349144
R5290 VGND.n2608 VGND.n2605 0.349144
R5291 VGND.n2605 VGND.n2602 0.349144
R5292 VGND.n2602 VGND.n2599 0.349144
R5293 VGND.n2599 VGND.n2596 0.349144
R5294 VGND.n2596 VGND.n2593 0.349144
R5295 VGND.n2593 VGND.n2590 0.349144
R5296 VGND.n1219 VGND.n1218 0.349144
R5297 VGND.n1219 VGND.n1215 0.349144
R5298 VGND.n1215 VGND.n790 0.349144
R5299 VGND.n1187 VGND.n790 0.349144
R5300 VGND.n1188 VGND.n1187 0.349144
R5301 VGND.n1188 VGND.n1183 0.349144
R5302 VGND.n1183 VGND.n798 0.349144
R5303 VGND.n1155 VGND.n798 0.349144
R5304 VGND.n1156 VGND.n1155 0.349144
R5305 VGND.n1156 VGND.n1151 0.349144
R5306 VGND.n1151 VGND.n806 0.349144
R5307 VGND.n818 VGND.n806 0.349144
R5308 VGND.n821 VGND.n818 0.349144
R5309 VGND.n2656 VGND.n2651 0.327628
R5310 VGND.n2660 VGND.n2659 0.327628
R5311 VGND.n2664 VGND.n2647 0.327628
R5312 VGND.n2668 VGND.n2667 0.327628
R5313 VGND.n2672 VGND.n2643 0.327628
R5314 VGND.n2676 VGND.n2675 0.327628
R5315 VGND.n2680 VGND.n2639 0.327628
R5316 VGND.n2684 VGND.n2683 0.327628
R5317 VGND.n2688 VGND.n2635 0.327628
R5318 VGND.n2692 VGND.n2691 0.327628
R5319 VGND.n2696 VGND.n2631 0.327628
R5320 VGND.n2700 VGND.n2699 0.327628
R5321 VGND.n2704 VGND.n2627 0.327628
R5322 VGND.n2708 VGND.n2707 0.327628
R5323 VGND.n2578 VGND.n2576 0.327628
R5324 VGND.n2783 VGND.n2782 0.327628
R5325 VGND.n2779 VGND.n220 0.327628
R5326 VGND.n2774 VGND.n219 0.327628
R5327 VGND.n2769 VGND.n214 0.327628
R5328 VGND.n2764 VGND.n213 0.327628
R5329 VGND.n2759 VGND.n208 0.327628
R5330 VGND.n2754 VGND.n207 0.327628
R5331 VGND.n2749 VGND.n202 0.327628
R5332 VGND.n2744 VGND.n201 0.327628
R5333 VGND.n2739 VGND.n196 0.327628
R5334 VGND.n2734 VGND.n195 0.327628
R5335 VGND.n2729 VGND.n190 0.327628
R5336 VGND.n2724 VGND.n189 0.327628
R5337 VGND.n2719 VGND.n2715 0.327628
R5338 VGND.n235 VGND.n234 0.327628
R5339 VGND.n2488 VGND.n258 0.327628
R5340 VGND.n2483 VGND.n257 0.327628
R5341 VGND.n2478 VGND.n256 0.327628
R5342 VGND.n2473 VGND.n255 0.327628
R5343 VGND.n2468 VGND.n254 0.327628
R5344 VGND.n2463 VGND.n253 0.327628
R5345 VGND.n2458 VGND.n252 0.327628
R5346 VGND.n2453 VGND.n251 0.327628
R5347 VGND.n2448 VGND.n250 0.327628
R5348 VGND.n2443 VGND.n249 0.327628
R5349 VGND.n2438 VGND.n248 0.327628
R5350 VGND.n2505 VGND.n244 0.327628
R5351 VGND.n2508 VGND.n186 0.327628
R5352 VGND.n2513 VGND.n185 0.327628
R5353 VGND.n2517 VGND.n2516 0.327628
R5354 VGND.n2294 VGND.n2293 0.327628
R5355 VGND.n2290 VGND.n329 0.327628
R5356 VGND.n2285 VGND.n328 0.327628
R5357 VGND.n2280 VGND.n2276 0.327628
R5358 VGND.n2253 VGND.n2252 0.327628
R5359 VGND.n2249 VGND.n2245 0.327628
R5360 VGND.n2227 VGND.n2226 0.327628
R5361 VGND.n2223 VGND.n2219 0.327628
R5362 VGND.n2201 VGND.n2200 0.327628
R5363 VGND.n2197 VGND.n2193 0.327628
R5364 VGND.n2175 VGND.n2174 0.327628
R5365 VGND.n2171 VGND.n2167 0.327628
R5366 VGND.n374 VGND.n373 0.327628
R5367 VGND.n2828 VGND.n182 0.327628
R5368 VGND.n2831 VGND.n180 0.327628
R5369 VGND.n2310 VGND.n324 0.327628
R5370 VGND.n2307 VGND.n2303 0.327628
R5371 VGND.n2267 VGND.n327 0.327628
R5372 VGND.n2271 VGND.n2270 0.327628
R5373 VGND.n2262 VGND.n2258 0.327628
R5374 VGND.n2240 VGND.n2239 0.327628
R5375 VGND.n2236 VGND.n2232 0.327628
R5376 VGND.n2214 VGND.n2213 0.327628
R5377 VGND.n2210 VGND.n2206 0.327628
R5378 VGND.n2188 VGND.n2187 0.327628
R5379 VGND.n2184 VGND.n2180 0.327628
R5380 VGND.n2162 VGND.n2161 0.327628
R5381 VGND.n2158 VGND.n2154 0.327628
R5382 VGND.n1432 VGND.n1431 0.327628
R5383 VGND.n1428 VGND.n1421 0.327628
R5384 VGND.n2130 VGND.n322 0.327628
R5385 VGND.n2135 VGND.n321 0.327628
R5386 VGND.n2139 VGND.n2138 0.327628
R5387 VGND.n1447 VGND.n390 0.327628
R5388 VGND.n1452 VGND.n389 0.327628
R5389 VGND.n1457 VGND.n388 0.327628
R5390 VGND.n1462 VGND.n387 0.327628
R5391 VGND.n1467 VGND.n386 0.327628
R5392 VGND.n1472 VGND.n385 0.327628
R5393 VGND.n1477 VGND.n384 0.327628
R5394 VGND.n1482 VGND.n383 0.327628
R5395 VGND.n1487 VGND.n382 0.327628
R5396 VGND.n1492 VGND.n381 0.327628
R5397 VGND.n1496 VGND.n1495 0.327628
R5398 VGND.n1442 VGND.n1438 0.327628
R5399 VGND.n2119 VGND.n399 0.327628
R5400 VGND.n2116 VGND.n319 0.327628
R5401 VGND.n2111 VGND.n318 0.327628
R5402 VGND.n2106 VGND.n2102 0.327628
R5403 VGND.n2079 VGND.n2078 0.327628
R5404 VGND.n2075 VGND.n2071 0.327628
R5405 VGND.n2053 VGND.n2052 0.327628
R5406 VGND.n2049 VGND.n2045 0.327628
R5407 VGND.n2027 VGND.n2026 0.327628
R5408 VGND.n2023 VGND.n2019 0.327628
R5409 VGND.n2001 VGND.n2000 0.327628
R5410 VGND.n1997 VGND.n1993 0.327628
R5411 VGND.n629 VGND.n628 0.327628
R5412 VGND.n1501 VGND.n619 0.327628
R5413 VGND.n1504 VGND.n617 0.327628
R5414 VGND.n2335 VGND.n312 0.327628
R5415 VGND.n2332 VGND.n2328 0.327628
R5416 VGND.n2093 VGND.n316 0.327628
R5417 VGND.n2097 VGND.n2096 0.327628
R5418 VGND.n2088 VGND.n2084 0.327628
R5419 VGND.n2066 VGND.n2065 0.327628
R5420 VGND.n2062 VGND.n2058 0.327628
R5421 VGND.n2040 VGND.n2039 0.327628
R5422 VGND.n2036 VGND.n2032 0.327628
R5423 VGND.n2014 VGND.n2013 0.327628
R5424 VGND.n2010 VGND.n2006 0.327628
R5425 VGND.n1988 VGND.n1987 0.327628
R5426 VGND.n1984 VGND.n1980 0.327628
R5427 VGND.n655 VGND.n654 0.327628
R5428 VGND.n651 VGND.n644 0.327628
R5429 VGND.n1956 VGND.n310 0.327628
R5430 VGND.n1961 VGND.n309 0.327628
R5431 VGND.n1965 VGND.n1964 0.327628
R5432 VGND.n903 VGND.n446 0.327628
R5433 VGND.n908 VGND.n445 0.327628
R5434 VGND.n913 VGND.n444 0.327628
R5435 VGND.n918 VGND.n443 0.327628
R5436 VGND.n923 VGND.n442 0.327628
R5437 VGND.n928 VGND.n441 0.327628
R5438 VGND.n933 VGND.n440 0.327628
R5439 VGND.n938 VGND.n439 0.327628
R5440 VGND.n943 VGND.n438 0.327628
R5441 VGND.n948 VGND.n437 0.327628
R5442 VGND.n953 VGND.n661 0.327628
R5443 VGND.n958 VGND.n660 0.327628
R5444 VGND.n1945 VGND.n455 0.327628
R5445 VGND.n1942 VGND.n307 0.327628
R5446 VGND.n1937 VGND.n306 0.327628
R5447 VGND.n1932 VGND.n1928 0.327628
R5448 VGND.n1905 VGND.n1904 0.327628
R5449 VGND.n1901 VGND.n1897 0.327628
R5450 VGND.n1879 VGND.n1878 0.327628
R5451 VGND.n1875 VGND.n1871 0.327628
R5452 VGND.n1853 VGND.n1852 0.327628
R5453 VGND.n1849 VGND.n1845 0.327628
R5454 VGND.n1827 VGND.n1826 0.327628
R5455 VGND.n1823 VGND.n1819 0.327628
R5456 VGND.n1404 VGND.n1403 0.327628
R5457 VGND.n1400 VGND.n663 0.327628
R5458 VGND.n1395 VGND.n1391 0.327628
R5459 VGND.n2360 VGND.n300 0.327628
R5460 VGND.n2357 VGND.n2353 0.327628
R5461 VGND.n1919 VGND.n304 0.327628
R5462 VGND.n1923 VGND.n1922 0.327628
R5463 VGND.n1914 VGND.n1910 0.327628
R5464 VGND.n1892 VGND.n1891 0.327628
R5465 VGND.n1888 VGND.n1884 0.327628
R5466 VGND.n1866 VGND.n1865 0.327628
R5467 VGND.n1862 VGND.n1858 0.327628
R5468 VGND.n1840 VGND.n1839 0.327628
R5469 VGND.n1836 VGND.n1832 0.327628
R5470 VGND.n1814 VGND.n1813 0.327628
R5471 VGND.n1810 VGND.n1806 0.327628
R5472 VGND.n1384 VGND.n1383 0.327628
R5473 VGND.n1380 VGND.n1373 0.327628
R5474 VGND.n1782 VGND.n298 0.327628
R5475 VGND.n1787 VGND.n297 0.327628
R5476 VGND.n1791 VGND.n1790 0.327628
R5477 VGND.n1317 VGND.n502 0.327628
R5478 VGND.n1322 VGND.n501 0.327628
R5479 VGND.n1327 VGND.n500 0.327628
R5480 VGND.n1332 VGND.n499 0.327628
R5481 VGND.n1337 VGND.n498 0.327628
R5482 VGND.n1342 VGND.n497 0.327628
R5483 VGND.n1347 VGND.n496 0.327628
R5484 VGND.n1352 VGND.n495 0.327628
R5485 VGND.n1357 VGND.n494 0.327628
R5486 VGND.n1362 VGND.n493 0.327628
R5487 VGND.n1366 VGND.n1365 0.327628
R5488 VGND.n1312 VGND.n1305 0.327628
R5489 VGND.n1771 VGND.n511 0.327628
R5490 VGND.n1768 VGND.n295 0.327628
R5491 VGND.n1763 VGND.n294 0.327628
R5492 VGND.n1758 VGND.n1754 0.327628
R5493 VGND.n1731 VGND.n1730 0.327628
R5494 VGND.n1727 VGND.n1723 0.327628
R5495 VGND.n1705 VGND.n1704 0.327628
R5496 VGND.n1701 VGND.n1697 0.327628
R5497 VGND.n1679 VGND.n1678 0.327628
R5498 VGND.n1675 VGND.n1671 0.327628
R5499 VGND.n1653 VGND.n1652 0.327628
R5500 VGND.n1649 VGND.n1645 0.327628
R5501 VGND.n1526 VGND.n1525 0.327628
R5502 VGND.n1522 VGND.n574 0.327628
R5503 VGND.n1517 VGND.n573 0.327628
R5504 VGND.n2385 VGND.n287 0.327628
R5505 VGND.n2382 VGND.n2378 0.327628
R5506 VGND.n1745 VGND.n291 0.327628
R5507 VGND.n1749 VGND.n1748 0.327628
R5508 VGND.n1740 VGND.n1736 0.327628
R5509 VGND.n1718 VGND.n1717 0.327628
R5510 VGND.n1714 VGND.n1710 0.327628
R5511 VGND.n1692 VGND.n1691 0.327628
R5512 VGND.n1688 VGND.n1684 0.327628
R5513 VGND.n1666 VGND.n1665 0.327628
R5514 VGND.n1662 VGND.n1658 0.327628
R5515 VGND.n1640 VGND.n1639 0.327628
R5516 VGND.n1636 VGND.n1632 0.327628
R5517 VGND.n1541 VGND.n1540 0.327628
R5518 VGND.n1537 VGND.n1533 0.327628
R5519 VGND.n1608 VGND.n283 0.327628
R5520 VGND.n1613 VGND.n282 0.327628
R5521 VGND.n1617 VGND.n1616 0.327628
R5522 VGND.n1600 VGND.n558 0.327628
R5523 VGND.n1595 VGND.n557 0.327628
R5524 VGND.n1590 VGND.n556 0.327628
R5525 VGND.n1585 VGND.n555 0.327628
R5526 VGND.n1580 VGND.n554 0.327628
R5527 VGND.n1575 VGND.n553 0.327628
R5528 VGND.n1570 VGND.n552 0.327628
R5529 VGND.n1565 VGND.n551 0.327628
R5530 VGND.n1560 VGND.n550 0.327628
R5531 VGND.n1555 VGND.n549 0.327628
R5532 VGND.n1550 VGND.n1546 0.327628
R5533 VGND.n1298 VGND.n1297 0.327628
R5534 VGND.n2405 VGND.n279 0.327628
R5535 VGND.n2402 VGND.n2398 0.327628
R5536 VGND.n844 VGND.n713 0.327628
R5537 VGND.n849 VGND.n712 0.327628
R5538 VGND.n854 VGND.n707 0.327628
R5539 VGND.n859 VGND.n706 0.327628
R5540 VGND.n864 VGND.n701 0.327628
R5541 VGND.n869 VGND.n700 0.327628
R5542 VGND.n874 VGND.n695 0.327628
R5543 VGND.n879 VGND.n694 0.327628
R5544 VGND.n884 VGND.n689 0.327628
R5545 VGND.n889 VGND.n688 0.327628
R5546 VGND.n893 VGND.n892 0.327628
R5547 VGND.n839 VGND.n827 0.327628
R5548 VGND.n834 VGND.n826 0.327628
R5549 VGND.n1124 VGND.n1122 0.327628
R5550 VGND.n1131 VGND.n1127 0.327628
R5551 VGND.n1134 VGND.n812 0.327628
R5552 VGND.n1144 VGND.n1140 0.327628
R5553 VGND.n1148 VGND.n1147 0.327628
R5554 VGND.n1163 VGND.n1159 0.327628
R5555 VGND.n1166 VGND.n804 0.327628
R5556 VGND.n1176 VGND.n1172 0.327628
R5557 VGND.n1180 VGND.n1179 0.327628
R5558 VGND.n1195 VGND.n1191 0.327628
R5559 VGND.n1198 VGND.n796 0.327628
R5560 VGND.n1208 VGND.n1204 0.327628
R5561 VGND.n1212 VGND.n1211 0.327628
R5562 VGND.n1227 VGND.n1223 0.327628
R5563 VGND.n1230 VGND.n788 0.327628
R5564 VGND.n783 VGND.n782 0.327628
R5565 VGND.n779 VGND.n716 0.327628
R5566 VGND.n774 VGND.n715 0.327628
R5567 VGND.n769 VGND.n710 0.327628
R5568 VGND.n764 VGND.n709 0.327628
R5569 VGND.n759 VGND.n704 0.327628
R5570 VGND.n754 VGND.n703 0.327628
R5571 VGND.n749 VGND.n698 0.327628
R5572 VGND.n744 VGND.n697 0.327628
R5573 VGND.n739 VGND.n692 0.327628
R5574 VGND.n734 VGND.n691 0.327628
R5575 VGND.n729 VGND.n686 0.327628
R5576 VGND.n724 VGND.n685 0.327628
R5577 VGND.n1286 VGND.n679 0.327628
R5578 VGND.n1289 VGND.n677 0.327628
R5579 VGND.n3024 VGND.n2 0.247202
R5580 VGND.n2920 VGND.n59 0.213567
R5581 VGND.n2953 VGND.n2920 0.213567
R5582 VGND.n2954 VGND.n2953 0.213567
R5583 VGND.n2954 VGND.n28 0.213567
R5584 VGND.n1113 VGND.n1090 0.213567
R5585 VGND.n1090 VGND.n1060 0.213567
R5586 VGND.n1060 VGND.n1029 0.213567
R5587 VGND.n1029 VGND.n998 0.213567
R5588 VGND.n998 VGND.n0 0.213567
R5589 VGND.n3006 VGND.n28 0.2073
R5590 VGND.n1116 VGND.n1115 0.17205
R5591 VGND.n2711 VGND 0.169807
R5592 VGND.n2710 VGND 0.169807
R5593 VGND VGND.n188 0.169807
R5594 VGND.n2817 VGND 0.169807
R5595 VGND.n2816 VGND 0.169807
R5596 VGND.n2811 VGND 0.169807
R5597 VGND.n2810 VGND 0.169807
R5598 VGND.n2805 VGND 0.169807
R5599 VGND.n2804 VGND 0.169807
R5600 VGND.n2799 VGND 0.169807
R5601 VGND.n2798 VGND 0.169807
R5602 VGND.n2793 VGND 0.169807
R5603 VGND.n2792 VGND 0.169807
R5604 VGND.n2787 VGND 0.169807
R5605 VGND.n2786 VGND 0.169807
R5606 VGND VGND.n2713 0.169807
R5607 VGND.n2714 VGND 0.169807
R5608 VGND.n2820 VGND 0.169807
R5609 VGND.n2819 VGND 0.169807
R5610 VGND.n2814 VGND 0.169807
R5611 VGND.n2813 VGND 0.169807
R5612 VGND.n2808 VGND 0.169807
R5613 VGND.n2807 VGND 0.169807
R5614 VGND.n2802 VGND 0.169807
R5615 VGND.n2801 VGND 0.169807
R5616 VGND.n2796 VGND 0.169807
R5617 VGND.n2795 VGND 0.169807
R5618 VGND.n2790 VGND 0.169807
R5619 VGND.n2789 VGND 0.169807
R5620 VGND.n2784 VGND 0.169807
R5621 VGND.n2518 VGND 0.169807
R5622 VGND.n2824 VGND 0.169807
R5623 VGND.n2823 VGND 0.169807
R5624 VGND.n2504 VGND 0.169807
R5625 VGND.n2503 VGND 0.169807
R5626 VGND.n2502 VGND 0.169807
R5627 VGND.n2501 VGND 0.169807
R5628 VGND.n2500 VGND 0.169807
R5629 VGND.n2499 VGND 0.169807
R5630 VGND.n2498 VGND 0.169807
R5631 VGND.n2497 VGND 0.169807
R5632 VGND.n2496 VGND 0.169807
R5633 VGND.n2495 VGND 0.169807
R5634 VGND.n2494 VGND 0.169807
R5635 VGND.n2493 VGND 0.169807
R5636 VGND.n639 VGND 0.169807
R5637 VGND.n2827 VGND 0.169807
R5638 VGND VGND.n375 0.169807
R5639 VGND.n2166 VGND 0.169807
R5640 VGND.n2176 VGND 0.169807
R5641 VGND.n2192 VGND 0.169807
R5642 VGND.n2202 VGND 0.169807
R5643 VGND.n2218 VGND 0.169807
R5644 VGND.n2228 VGND 0.169807
R5645 VGND.n2244 VGND 0.169807
R5646 VGND.n2254 VGND 0.169807
R5647 VGND.n2275 VGND 0.169807
R5648 VGND.n2298 VGND 0.169807
R5649 VGND.n2297 VGND 0.169807
R5650 VGND.n2295 VGND 0.169807
R5651 VGND.n1434 VGND 0.169807
R5652 VGND.n1433 VGND 0.169807
R5653 VGND.n2153 VGND 0.169807
R5654 VGND.n2163 VGND 0.169807
R5655 VGND.n2179 VGND 0.169807
R5656 VGND.n2189 VGND 0.169807
R5657 VGND.n2205 VGND 0.169807
R5658 VGND.n2215 VGND 0.169807
R5659 VGND.n2231 VGND 0.169807
R5660 VGND.n2241 VGND 0.169807
R5661 VGND.n2257 VGND 0.169807
R5662 VGND.n2272 VGND 0.169807
R5663 VGND VGND.n2301 0.169807
R5664 VGND.n2302 VGND 0.169807
R5665 VGND.n2315 VGND 0.169807
R5666 VGND.n1437 VGND 0.169807
R5667 VGND.n1497 VGND 0.169807
R5668 VGND.n2150 VGND 0.169807
R5669 VGND.n2149 VGND 0.169807
R5670 VGND.n2148 VGND 0.169807
R5671 VGND.n2147 VGND 0.169807
R5672 VGND.n2146 VGND 0.169807
R5673 VGND.n2145 VGND 0.169807
R5674 VGND.n2144 VGND 0.169807
R5675 VGND.n2143 VGND 0.169807
R5676 VGND.n2142 VGND 0.169807
R5677 VGND.n2141 VGND 0.169807
R5678 VGND.n2140 VGND 0.169807
R5679 VGND.n2319 VGND 0.169807
R5680 VGND.n2318 VGND 0.169807
R5681 VGND.n1415 VGND 0.169807
R5682 VGND.n1500 VGND 0.169807
R5683 VGND.n630 VGND 0.169807
R5684 VGND.n1992 VGND 0.169807
R5685 VGND.n2002 VGND 0.169807
R5686 VGND.n2018 VGND 0.169807
R5687 VGND.n2028 VGND 0.169807
R5688 VGND.n2044 VGND 0.169807
R5689 VGND.n2054 VGND 0.169807
R5690 VGND.n2070 VGND 0.169807
R5691 VGND.n2080 VGND 0.169807
R5692 VGND.n2101 VGND 0.169807
R5693 VGND.n2323 VGND 0.169807
R5694 VGND.n2322 VGND 0.169807
R5695 VGND.n398 VGND 0.169807
R5696 VGND.n1413 VGND 0.169807
R5697 VGND.n656 VGND 0.169807
R5698 VGND.n1979 VGND 0.169807
R5699 VGND.n1989 VGND 0.169807
R5700 VGND.n2005 VGND 0.169807
R5701 VGND.n2015 VGND 0.169807
R5702 VGND.n2031 VGND 0.169807
R5703 VGND.n2041 VGND 0.169807
R5704 VGND.n2057 VGND 0.169807
R5705 VGND.n2067 VGND 0.169807
R5706 VGND.n2083 VGND 0.169807
R5707 VGND.n2098 VGND 0.169807
R5708 VGND VGND.n2326 0.169807
R5709 VGND.n2327 VGND 0.169807
R5710 VGND.n2340 VGND 0.169807
R5711 VGND.n1410 VGND 0.169807
R5712 VGND.n1409 VGND 0.169807
R5713 VGND.n1976 VGND 0.169807
R5714 VGND.n1975 VGND 0.169807
R5715 VGND.n1974 VGND 0.169807
R5716 VGND.n1973 VGND 0.169807
R5717 VGND.n1972 VGND 0.169807
R5718 VGND.n1971 VGND 0.169807
R5719 VGND.n1970 VGND 0.169807
R5720 VGND.n1969 VGND 0.169807
R5721 VGND.n1968 VGND 0.169807
R5722 VGND.n1967 VGND 0.169807
R5723 VGND.n1966 VGND 0.169807
R5724 VGND.n2344 VGND 0.169807
R5725 VGND.n2343 VGND 0.169807
R5726 VGND.n1390 VGND 0.169807
R5727 VGND.n1406 VGND 0.169807
R5728 VGND.n1405 VGND 0.169807
R5729 VGND.n1818 VGND 0.169807
R5730 VGND.n1828 VGND 0.169807
R5731 VGND.n1844 VGND 0.169807
R5732 VGND.n1854 VGND 0.169807
R5733 VGND.n1870 VGND 0.169807
R5734 VGND.n1880 VGND 0.169807
R5735 VGND.n1896 VGND 0.169807
R5736 VGND.n1906 VGND 0.169807
R5737 VGND.n1927 VGND 0.169807
R5738 VGND.n2348 VGND 0.169807
R5739 VGND.n2347 VGND 0.169807
R5740 VGND.n454 VGND 0.169807
R5741 VGND.n1387 VGND 0.169807
R5742 VGND.n1385 VGND 0.169807
R5743 VGND.n1805 VGND 0.169807
R5744 VGND.n1815 VGND 0.169807
R5745 VGND.n1831 VGND 0.169807
R5746 VGND.n1841 VGND 0.169807
R5747 VGND.n1857 VGND 0.169807
R5748 VGND.n1867 VGND 0.169807
R5749 VGND.n1883 VGND 0.169807
R5750 VGND.n1893 VGND 0.169807
R5751 VGND.n1909 VGND 0.169807
R5752 VGND.n1924 VGND 0.169807
R5753 VGND VGND.n2351 0.169807
R5754 VGND.n2352 VGND 0.169807
R5755 VGND.n2365 VGND 0.169807
R5756 VGND.n1369 VGND 0.169807
R5757 VGND.n1368 VGND 0.169807
R5758 VGND.n1802 VGND 0.169807
R5759 VGND.n1801 VGND 0.169807
R5760 VGND.n1800 VGND 0.169807
R5761 VGND.n1799 VGND 0.169807
R5762 VGND.n1798 VGND 0.169807
R5763 VGND.n1797 VGND 0.169807
R5764 VGND.n1796 VGND 0.169807
R5765 VGND.n1795 VGND 0.169807
R5766 VGND.n1794 VGND 0.169807
R5767 VGND.n1793 VGND 0.169807
R5768 VGND.n1792 VGND 0.169807
R5769 VGND.n2369 VGND 0.169807
R5770 VGND.n2368 VGND 0.169807
R5771 VGND.n1529 VGND 0.169807
R5772 VGND.n1528 VGND 0.169807
R5773 VGND.n1527 VGND 0.169807
R5774 VGND.n1644 VGND 0.169807
R5775 VGND.n1654 VGND 0.169807
R5776 VGND.n1670 VGND 0.169807
R5777 VGND.n1680 VGND 0.169807
R5778 VGND.n1696 VGND 0.169807
R5779 VGND.n1706 VGND 0.169807
R5780 VGND.n1722 VGND 0.169807
R5781 VGND.n1732 VGND 0.169807
R5782 VGND.n1753 VGND 0.169807
R5783 VGND.n2373 VGND 0.169807
R5784 VGND.n2372 VGND 0.169807
R5785 VGND.n510 VGND 0.169807
R5786 VGND.n1532 VGND 0.169807
R5787 VGND.n1542 VGND 0.169807
R5788 VGND.n1631 VGND 0.169807
R5789 VGND.n1641 VGND 0.169807
R5790 VGND.n1657 VGND 0.169807
R5791 VGND.n1667 VGND 0.169807
R5792 VGND.n1683 VGND 0.169807
R5793 VGND.n1693 VGND 0.169807
R5794 VGND.n1709 VGND 0.169807
R5795 VGND.n1719 VGND 0.169807
R5796 VGND.n1735 VGND 0.169807
R5797 VGND.n1750 VGND 0.169807
R5798 VGND VGND.n2376 0.169807
R5799 VGND.n2377 VGND 0.169807
R5800 VGND.n2390 VGND 0.169807
R5801 VGND.n1299 VGND 0.169807
R5802 VGND.n1545 VGND 0.169807
R5803 VGND.n1628 VGND 0.169807
R5804 VGND.n1627 VGND 0.169807
R5805 VGND.n1626 VGND 0.169807
R5806 VGND.n1625 VGND 0.169807
R5807 VGND.n1624 VGND 0.169807
R5808 VGND.n1623 VGND 0.169807
R5809 VGND.n1622 VGND 0.169807
R5810 VGND.n1621 VGND 0.169807
R5811 VGND.n1620 VGND 0.169807
R5812 VGND.n1619 VGND 0.169807
R5813 VGND.n1618 VGND 0.169807
R5814 VGND.n2394 VGND 0.169807
R5815 VGND.n2393 VGND 0.169807
R5816 VGND.n896 VGND 0.169807
R5817 VGND.n895 VGND 0.169807
R5818 VGND.n894 VGND 0.169807
R5819 VGND.n1276 VGND 0.169807
R5820 VGND.n1275 VGND 0.169807
R5821 VGND.n1268 VGND 0.169807
R5822 VGND.n1267 VGND 0.169807
R5823 VGND.n1260 VGND 0.169807
R5824 VGND.n1259 VGND 0.169807
R5825 VGND.n1252 VGND 0.169807
R5826 VGND.n1251 VGND 0.169807
R5827 VGND.n1244 VGND 0.169807
R5828 VGND.n1243 VGND 0.169807
R5829 VGND.n2397 VGND 0.169807
R5830 VGND.n284 VGND 0.169807
R5831 VGND.n1120 VGND 0.169807
R5832 VGND.n1283 VGND 0.169807
R5833 VGND.n1282 VGND 0.169807
R5834 VGND VGND.n687 0.169807
R5835 VGND VGND.n690 0.169807
R5836 VGND VGND.n693 0.169807
R5837 VGND VGND.n696 0.169807
R5838 VGND VGND.n699 0.169807
R5839 VGND VGND.n702 0.169807
R5840 VGND VGND.n705 0.169807
R5841 VGND VGND.n708 0.169807
R5842 VGND VGND.n711 0.169807
R5843 VGND VGND.n714 0.169807
R5844 VGND.n1221 VGND 0.169807
R5845 VGND.n1236 VGND 0.169807
R5846 VGND.n1118 VGND 0.169807
R5847 VGND.n1285 VGND 0.169807
R5848 VGND.n1280 VGND 0.169807
R5849 VGND.n1279 VGND 0.169807
R5850 VGND.n1272 VGND 0.169807
R5851 VGND.n1271 VGND 0.169807
R5852 VGND.n1264 VGND 0.169807
R5853 VGND.n1263 VGND 0.169807
R5854 VGND.n1256 VGND 0.169807
R5855 VGND.n1255 VGND 0.169807
R5856 VGND.n1248 VGND 0.169807
R5857 VGND.n1247 VGND 0.169807
R5858 VGND.n1240 VGND 0.169807
R5859 VGND.n1239 VGND 0.169807
R5860 VGND.n1238 VGND 0.169807
R5861 VGND.n109 VGND 0.159538
R5862 VGND.n2871 VGND 0.159538
R5863 VGND.n2411 VGND.n275 0.154425
R5864 VGND.n2411 VGND.n2410 0.154425
R5865 VGND.n2410 VGND.n276 0.154425
R5866 VGND.n289 VGND.n276 0.154425
R5867 VGND.n1776 VGND.n289 0.154425
R5868 VGND.n1777 VGND.n1776 0.154425
R5869 VGND.n1777 VGND.n302 0.154425
R5870 VGND.n1950 VGND.n302 0.154425
R5871 VGND.n1951 VGND.n1950 0.154425
R5872 VGND.n1951 VGND.n314 0.154425
R5873 VGND.n2124 VGND.n314 0.154425
R5874 VGND.n2125 VGND.n2124 0.154425
R5875 VGND.n2125 VGND.n259 0.154425
R5876 VGND.n2432 VGND.n259 0.154425
R5877 VGND.n2433 VGND.n2432 0.154425
R5878 VGND.n2433 VGND.n29 0.154425
R5879 VGND.n3005 VGND.n29 0.154425
R5880 VGND.n1117 VGND.n1116 0.154425
R5881 VGND.n1117 VGND.n669 0.154425
R5882 VGND.n1300 VGND.n669 0.154425
R5883 VGND.n1301 VGND.n1300 0.154425
R5884 VGND.n1302 VGND.n1301 0.154425
R5885 VGND.n1370 VGND.n1302 0.154425
R5886 VGND.n1388 VGND.n1370 0.154425
R5887 VGND.n1389 VGND.n1388 0.154425
R5888 VGND.n1389 VGND.n641 0.154425
R5889 VGND.n1414 VGND.n641 0.154425
R5890 VGND.n1416 VGND.n1414 0.154425
R5891 VGND.n1417 VGND.n1416 0.154425
R5892 VGND.n1418 VGND.n1417 0.154425
R5893 VGND.n1418 VGND.n237 0.154425
R5894 VGND.n2519 VGND.n237 0.154425
R5895 VGND.n2520 VGND.n2519 0.154425
R5896 VGND.n2521 VGND.n2520 0.154425
R5897 VGND.n1100 VGND.n1094 0.144904
R5898 VGND.n1073 VGND.n1065 0.144904
R5899 VGND.n1011 VGND.n1003 0.144904
R5900 VGND.n1042 VGND.n1034 0.144904
R5901 VGND.n2568 VGND.n2567 0.138284
R5902 VGND.n2656 VGND.n2655 0.13638
R5903 VGND.n2659 VGND.n2648 0.13638
R5904 VGND.n2664 VGND.n2663 0.13638
R5905 VGND.n2667 VGND.n2644 0.13638
R5906 VGND.n2672 VGND.n2671 0.13638
R5907 VGND.n2675 VGND.n2640 0.13638
R5908 VGND.n2680 VGND.n2679 0.13638
R5909 VGND.n2683 VGND.n2636 0.13638
R5910 VGND.n2688 VGND.n2687 0.13638
R5911 VGND.n2691 VGND.n2632 0.13638
R5912 VGND.n2696 VGND.n2695 0.13638
R5913 VGND.n2699 VGND.n2628 0.13638
R5914 VGND.n2704 VGND.n2703 0.13638
R5915 VGND.n2707 VGND.n2573 0.13638
R5916 VGND.n2578 VGND.n2577 0.13638
R5917 VGND.n2782 VGND.n227 0.13638
R5918 VGND.n2779 VGND.n2778 0.13638
R5919 VGND.n2774 VGND.n2773 0.13638
R5920 VGND.n2769 VGND.n2768 0.13638
R5921 VGND.n2764 VGND.n2763 0.13638
R5922 VGND.n2759 VGND.n2758 0.13638
R5923 VGND.n2754 VGND.n2753 0.13638
R5924 VGND.n2749 VGND.n2748 0.13638
R5925 VGND.n2744 VGND.n2743 0.13638
R5926 VGND.n2739 VGND.n2738 0.13638
R5927 VGND.n2734 VGND.n2733 0.13638
R5928 VGND.n2729 VGND.n2728 0.13638
R5929 VGND.n2724 VGND.n2723 0.13638
R5930 VGND.n2719 VGND.n2718 0.13638
R5931 VGND.n234 VGND.n232 0.13638
R5932 VGND.n2488 VGND.n2487 0.13638
R5933 VGND.n2483 VGND.n2482 0.13638
R5934 VGND.n2478 VGND.n2477 0.13638
R5935 VGND.n2473 VGND.n2472 0.13638
R5936 VGND.n2468 VGND.n2467 0.13638
R5937 VGND.n2463 VGND.n2462 0.13638
R5938 VGND.n2458 VGND.n2457 0.13638
R5939 VGND.n2453 VGND.n2452 0.13638
R5940 VGND.n2448 VGND.n2447 0.13638
R5941 VGND.n2443 VGND.n2442 0.13638
R5942 VGND.n2438 VGND.n2437 0.13638
R5943 VGND.n246 VGND.n244 0.13638
R5944 VGND.n2508 VGND.n2507 0.13638
R5945 VGND.n2513 VGND.n2512 0.13638
R5946 VGND.n2516 VGND.n242 0.13638
R5947 VGND.n2293 VGND.n332 0.13638
R5948 VGND.n2290 VGND.n2289 0.13638
R5949 VGND.n2285 VGND.n2284 0.13638
R5950 VGND.n2280 VGND.n2279 0.13638
R5951 VGND.n2252 VGND.n340 0.13638
R5952 VGND.n2249 VGND.n2248 0.13638
R5953 VGND.n2226 VGND.n348 0.13638
R5954 VGND.n2223 VGND.n2222 0.13638
R5955 VGND.n2200 VGND.n356 0.13638
R5956 VGND.n2197 VGND.n2196 0.13638
R5957 VGND.n2174 VGND.n364 0.13638
R5958 VGND.n2171 VGND.n2170 0.13638
R5959 VGND.n373 VGND.n370 0.13638
R5960 VGND.n366 VGND.n182 0.13638
R5961 VGND.n2831 VGND.n2830 0.13638
R5962 VGND.n2311 VGND.n2310 0.13638
R5963 VGND.n2307 VGND.n2306 0.13638
R5964 VGND.n2267 VGND.n2266 0.13638
R5965 VGND.n2270 VGND.n336 0.13638
R5966 VGND.n2262 VGND.n2261 0.13638
R5967 VGND.n2239 VGND.n344 0.13638
R5968 VGND.n2236 VGND.n2235 0.13638
R5969 VGND.n2213 VGND.n352 0.13638
R5970 VGND.n2210 VGND.n2209 0.13638
R5971 VGND.n2187 VGND.n360 0.13638
R5972 VGND.n2184 VGND.n2183 0.13638
R5973 VGND.n2161 VGND.n379 0.13638
R5974 VGND.n2158 VGND.n2157 0.13638
R5975 VGND.n1431 VGND.n1424 0.13638
R5976 VGND.n1428 VGND.n1427 0.13638
R5977 VGND.n2130 VGND.n2129 0.13638
R5978 VGND.n2135 VGND.n2134 0.13638
R5979 VGND.n2138 VGND.n393 0.13638
R5980 VGND.n1447 VGND.n1446 0.13638
R5981 VGND.n1452 VGND.n1451 0.13638
R5982 VGND.n1457 VGND.n1456 0.13638
R5983 VGND.n1462 VGND.n1461 0.13638
R5984 VGND.n1467 VGND.n1466 0.13638
R5985 VGND.n1472 VGND.n1471 0.13638
R5986 VGND.n1477 VGND.n1476 0.13638
R5987 VGND.n1482 VGND.n1481 0.13638
R5988 VGND.n1487 VGND.n1486 0.13638
R5989 VGND.n1492 VGND.n1491 0.13638
R5990 VGND.n1495 VGND.n634 0.13638
R5991 VGND.n1442 VGND.n1441 0.13638
R5992 VGND.n2120 VGND.n2119 0.13638
R5993 VGND.n2116 VGND.n2115 0.13638
R5994 VGND.n2111 VGND.n2110 0.13638
R5995 VGND.n2106 VGND.n2105 0.13638
R5996 VGND.n2078 VGND.n407 0.13638
R5997 VGND.n2075 VGND.n2074 0.13638
R5998 VGND.n2052 VGND.n415 0.13638
R5999 VGND.n2049 VGND.n2048 0.13638
R6000 VGND.n2026 VGND.n423 0.13638
R6001 VGND.n2023 VGND.n2022 0.13638
R6002 VGND.n2000 VGND.n431 0.13638
R6003 VGND.n1997 VGND.n1996 0.13638
R6004 VGND.n628 VGND.n625 0.13638
R6005 VGND.n621 VGND.n619 0.13638
R6006 VGND.n1504 VGND.n1503 0.13638
R6007 VGND.n2336 VGND.n2335 0.13638
R6008 VGND.n2332 VGND.n2331 0.13638
R6009 VGND.n2093 VGND.n2092 0.13638
R6010 VGND.n2096 VGND.n403 0.13638
R6011 VGND.n2088 VGND.n2087 0.13638
R6012 VGND.n2065 VGND.n411 0.13638
R6013 VGND.n2062 VGND.n2061 0.13638
R6014 VGND.n2039 VGND.n419 0.13638
R6015 VGND.n2036 VGND.n2035 0.13638
R6016 VGND.n2013 VGND.n427 0.13638
R6017 VGND.n2010 VGND.n2009 0.13638
R6018 VGND.n1987 VGND.n435 0.13638
R6019 VGND.n1984 VGND.n1983 0.13638
R6020 VGND.n654 VGND.n647 0.13638
R6021 VGND.n651 VGND.n650 0.13638
R6022 VGND.n1956 VGND.n1955 0.13638
R6023 VGND.n1961 VGND.n1960 0.13638
R6024 VGND.n1964 VGND.n449 0.13638
R6025 VGND.n903 VGND.n902 0.13638
R6026 VGND.n908 VGND.n907 0.13638
R6027 VGND.n913 VGND.n912 0.13638
R6028 VGND.n918 VGND.n917 0.13638
R6029 VGND.n923 VGND.n922 0.13638
R6030 VGND.n928 VGND.n927 0.13638
R6031 VGND.n933 VGND.n932 0.13638
R6032 VGND.n938 VGND.n937 0.13638
R6033 VGND.n943 VGND.n942 0.13638
R6034 VGND.n948 VGND.n947 0.13638
R6035 VGND.n953 VGND.n952 0.13638
R6036 VGND.n958 VGND.n957 0.13638
R6037 VGND.n1946 VGND.n1945 0.13638
R6038 VGND.n1942 VGND.n1941 0.13638
R6039 VGND.n1937 VGND.n1936 0.13638
R6040 VGND.n1932 VGND.n1931 0.13638
R6041 VGND.n1904 VGND.n463 0.13638
R6042 VGND.n1901 VGND.n1900 0.13638
R6043 VGND.n1878 VGND.n471 0.13638
R6044 VGND.n1875 VGND.n1874 0.13638
R6045 VGND.n1852 VGND.n479 0.13638
R6046 VGND.n1849 VGND.n1848 0.13638
R6047 VGND.n1826 VGND.n487 0.13638
R6048 VGND.n1823 VGND.n1822 0.13638
R6049 VGND.n1403 VGND.n666 0.13638
R6050 VGND.n1400 VGND.n1399 0.13638
R6051 VGND.n1395 VGND.n1394 0.13638
R6052 VGND.n2361 VGND.n2360 0.13638
R6053 VGND.n2357 VGND.n2356 0.13638
R6054 VGND.n1919 VGND.n1918 0.13638
R6055 VGND.n1922 VGND.n459 0.13638
R6056 VGND.n1914 VGND.n1913 0.13638
R6057 VGND.n1891 VGND.n467 0.13638
R6058 VGND.n1888 VGND.n1887 0.13638
R6059 VGND.n1865 VGND.n475 0.13638
R6060 VGND.n1862 VGND.n1861 0.13638
R6061 VGND.n1839 VGND.n483 0.13638
R6062 VGND.n1836 VGND.n1835 0.13638
R6063 VGND.n1813 VGND.n491 0.13638
R6064 VGND.n1810 VGND.n1809 0.13638
R6065 VGND.n1383 VGND.n1376 0.13638
R6066 VGND.n1380 VGND.n1379 0.13638
R6067 VGND.n1782 VGND.n1781 0.13638
R6068 VGND.n1787 VGND.n1786 0.13638
R6069 VGND.n1790 VGND.n505 0.13638
R6070 VGND.n1317 VGND.n1316 0.13638
R6071 VGND.n1322 VGND.n1321 0.13638
R6072 VGND.n1327 VGND.n1326 0.13638
R6073 VGND.n1332 VGND.n1331 0.13638
R6074 VGND.n1337 VGND.n1336 0.13638
R6075 VGND.n1342 VGND.n1341 0.13638
R6076 VGND.n1347 VGND.n1346 0.13638
R6077 VGND.n1352 VGND.n1351 0.13638
R6078 VGND.n1357 VGND.n1356 0.13638
R6079 VGND.n1362 VGND.n1361 0.13638
R6080 VGND.n1365 VGND.n1308 0.13638
R6081 VGND.n1312 VGND.n1311 0.13638
R6082 VGND.n1772 VGND.n1771 0.13638
R6083 VGND.n1768 VGND.n1767 0.13638
R6084 VGND.n1763 VGND.n1762 0.13638
R6085 VGND.n1758 VGND.n1757 0.13638
R6086 VGND.n1730 VGND.n519 0.13638
R6087 VGND.n1727 VGND.n1726 0.13638
R6088 VGND.n1704 VGND.n527 0.13638
R6089 VGND.n1701 VGND.n1700 0.13638
R6090 VGND.n1678 VGND.n535 0.13638
R6091 VGND.n1675 VGND.n1674 0.13638
R6092 VGND.n1652 VGND.n543 0.13638
R6093 VGND.n1649 VGND.n1648 0.13638
R6094 VGND.n1525 VGND.n577 0.13638
R6095 VGND.n1522 VGND.n1521 0.13638
R6096 VGND.n1517 VGND.n1516 0.13638
R6097 VGND.n2386 VGND.n2385 0.13638
R6098 VGND.n2382 VGND.n2381 0.13638
R6099 VGND.n1745 VGND.n1744 0.13638
R6100 VGND.n1748 VGND.n515 0.13638
R6101 VGND.n1740 VGND.n1739 0.13638
R6102 VGND.n1717 VGND.n523 0.13638
R6103 VGND.n1714 VGND.n1713 0.13638
R6104 VGND.n1691 VGND.n531 0.13638
R6105 VGND.n1688 VGND.n1687 0.13638
R6106 VGND.n1665 VGND.n539 0.13638
R6107 VGND.n1662 VGND.n1661 0.13638
R6108 VGND.n1639 VGND.n547 0.13638
R6109 VGND.n1636 VGND.n1635 0.13638
R6110 VGND.n1540 VGND.n566 0.13638
R6111 VGND.n1537 VGND.n1536 0.13638
R6112 VGND.n1608 VGND.n1607 0.13638
R6113 VGND.n1613 VGND.n1612 0.13638
R6114 VGND.n1616 VGND.n561 0.13638
R6115 VGND.n1600 VGND.n1599 0.13638
R6116 VGND.n1595 VGND.n1594 0.13638
R6117 VGND.n1590 VGND.n1589 0.13638
R6118 VGND.n1585 VGND.n1584 0.13638
R6119 VGND.n1580 VGND.n1579 0.13638
R6120 VGND.n1575 VGND.n1574 0.13638
R6121 VGND.n1570 VGND.n1569 0.13638
R6122 VGND.n1565 VGND.n1564 0.13638
R6123 VGND.n1560 VGND.n1559 0.13638
R6124 VGND.n1555 VGND.n1554 0.13638
R6125 VGND.n1550 VGND.n1549 0.13638
R6126 VGND.n1297 VGND.n674 0.13638
R6127 VGND.n2406 VGND.n2405 0.13638
R6128 VGND.n2402 VGND.n2401 0.13638
R6129 VGND.n844 VGND.n843 0.13638
R6130 VGND.n849 VGND.n848 0.13638
R6131 VGND.n854 VGND.n853 0.13638
R6132 VGND.n859 VGND.n858 0.13638
R6133 VGND.n864 VGND.n863 0.13638
R6134 VGND.n869 VGND.n868 0.13638
R6135 VGND.n874 VGND.n873 0.13638
R6136 VGND.n879 VGND.n878 0.13638
R6137 VGND.n884 VGND.n883 0.13638
R6138 VGND.n889 VGND.n888 0.13638
R6139 VGND.n892 VGND.n830 0.13638
R6140 VGND.n839 VGND.n838 0.13638
R6141 VGND.n834 VGND.n833 0.13638
R6142 VGND.n1125 VGND.n1124 0.13638
R6143 VGND.n1131 VGND.n1130 0.13638
R6144 VGND.n1135 VGND.n1134 0.13638
R6145 VGND.n1144 VGND.n1143 0.13638
R6146 VGND.n1147 VGND.n810 0.13638
R6147 VGND.n1163 VGND.n1162 0.13638
R6148 VGND.n1167 VGND.n1166 0.13638
R6149 VGND.n1176 VGND.n1175 0.13638
R6150 VGND.n1179 VGND.n802 0.13638
R6151 VGND.n1195 VGND.n1194 0.13638
R6152 VGND.n1199 VGND.n1198 0.13638
R6153 VGND.n1208 VGND.n1207 0.13638
R6154 VGND.n1211 VGND.n794 0.13638
R6155 VGND.n1227 VGND.n1226 0.13638
R6156 VGND.n1231 VGND.n1230 0.13638
R6157 VGND.n782 VGND.n719 0.13638
R6158 VGND.n779 VGND.n778 0.13638
R6159 VGND.n774 VGND.n773 0.13638
R6160 VGND.n769 VGND.n768 0.13638
R6161 VGND.n764 VGND.n763 0.13638
R6162 VGND.n759 VGND.n758 0.13638
R6163 VGND.n754 VGND.n753 0.13638
R6164 VGND.n749 VGND.n748 0.13638
R6165 VGND.n744 VGND.n743 0.13638
R6166 VGND.n739 VGND.n738 0.13638
R6167 VGND.n734 VGND.n733 0.13638
R6168 VGND.n729 VGND.n728 0.13638
R6169 VGND.n724 VGND.n723 0.13638
R6170 VGND.n683 VGND.n679 0.13638
R6171 VGND.n1289 VGND.n1288 0.13638
R6172 VGND VGND.n109 0.120838
R6173 VGND.n1108 VGND.n1107 0.120292
R6174 VGND.n1107 VGND.n1106 0.120292
R6175 VGND.n1106 VGND.n1092 0.120292
R6176 VGND.n1102 VGND.n1092 0.120292
R6177 VGND.n1102 VGND.n1101 0.120292
R6178 VGND.n1101 VGND.n1100 0.120292
R6179 VGND.n1086 VGND.n1085 0.120292
R6180 VGND.n1081 VGND.n1080 0.120292
R6181 VGND.n1080 VGND.n1079 0.120292
R6182 VGND.n1079 VGND.n1063 0.120292
R6183 VGND.n1075 VGND.n1063 0.120292
R6184 VGND.n1075 VGND.n1074 0.120292
R6185 VGND.n1074 VGND.n1073 0.120292
R6186 VGND.n143 VGND.n120 0.120292
R6187 VGND.n137 VGND.n120 0.120292
R6188 VGND.n137 VGND.n136 0.120292
R6189 VGND.n136 VGND.n124 0.120292
R6190 VGND.n129 VGND.n124 0.120292
R6191 VGND.n129 VGND.n128 0.120292
R6192 VGND.n128 VGND.n127 0.120292
R6193 VGND.n586 VGND.n583 0.120292
R6194 VGND.n587 VGND.n586 0.120292
R6195 VGND.n611 VGND.n588 0.120292
R6196 VGND.n605 VGND.n588 0.120292
R6197 VGND.n605 VGND.n604 0.120292
R6198 VGND.n604 VGND.n592 0.120292
R6199 VGND.n597 VGND.n592 0.120292
R6200 VGND.n597 VGND.n596 0.120292
R6201 VGND.n596 VGND.n595 0.120292
R6202 VGND.n994 VGND.n993 0.120292
R6203 VGND.n987 VGND.n963 0.120292
R6204 VGND.n982 VGND.n963 0.120292
R6205 VGND.n982 VGND.n981 0.120292
R6206 VGND.n978 VGND.n977 0.120292
R6207 VGND.n977 VGND.n972 0.120292
R6208 VGND.n973 VGND.n972 0.120292
R6209 VGND.n1024 VGND.n1023 0.120292
R6210 VGND.n1019 VGND.n1018 0.120292
R6211 VGND.n1018 VGND.n1017 0.120292
R6212 VGND.n1017 VGND.n1001 0.120292
R6213 VGND.n1013 VGND.n1001 0.120292
R6214 VGND.n1013 VGND.n1012 0.120292
R6215 VGND.n1012 VGND.n1011 0.120292
R6216 VGND.n1055 VGND.n1054 0.120292
R6217 VGND.n1050 VGND.n1049 0.120292
R6218 VGND.n1049 VGND.n1048 0.120292
R6219 VGND.n1048 VGND.n1032 0.120292
R6220 VGND.n1044 VGND.n1032 0.120292
R6221 VGND.n1044 VGND.n1043 0.120292
R6222 VGND.n1043 VGND.n1042 0.120292
R6223 VGND.n173 VGND.n150 0.120292
R6224 VGND.n167 VGND.n150 0.120292
R6225 VGND.n167 VGND.n166 0.120292
R6226 VGND.n166 VGND.n154 0.120292
R6227 VGND.n159 VGND.n154 0.120292
R6228 VGND.n159 VGND.n158 0.120292
R6229 VGND.n158 VGND.n157 0.120292
R6230 VGND.n15 VGND.n11 0.120292
R6231 VGND.n20 VGND.n11 0.120292
R6232 VGND.n21 VGND.n20 0.120292
R6233 VGND.n22 VGND.n21 0.120292
R6234 VGND.n22 VGND.n9 0.120292
R6235 VGND.n26 VGND.n9 0.120292
R6236 VGND.n27 VGND.n26 0.120292
R6237 VGND.n101 VGND.n93 0.120292
R6238 VGND.n102 VGND.n101 0.120292
R6239 VGND.n102 VGND.n87 0.120292
R6240 VGND.n107 VGND.n87 0.120292
R6241 VGND.n108 VGND.n107 0.120292
R6242 VGND.n2861 VGND.n2853 0.120292
R6243 VGND.n2862 VGND.n2861 0.120292
R6244 VGND.n2862 VGND.n2847 0.120292
R6245 VGND.n2867 VGND.n2847 0.120292
R6246 VGND.n2868 VGND.n2867 0.120292
R6247 VGND.n2893 VGND.n2885 0.120292
R6248 VGND.n2894 VGND.n2893 0.120292
R6249 VGND.n2894 VGND.n2879 0.120292
R6250 VGND.n2899 VGND.n2879 0.120292
R6251 VGND.n2900 VGND.n2899 0.120292
R6252 VGND.n2904 VGND.n2901 0.120292
R6253 VGND.n75 VGND.n68 0.120292
R6254 VGND.n76 VGND.n75 0.120292
R6255 VGND.n76 VGND.n63 0.120292
R6256 VGND.n81 VGND.n63 0.120292
R6257 VGND.n82 VGND.n81 0.120292
R6258 VGND.n2919 VGND.n60 0.120292
R6259 VGND.n2934 VGND.n2933 0.120292
R6260 VGND.n2934 VGND.n2926 0.120292
R6261 VGND.n2939 VGND.n2926 0.120292
R6262 VGND.n2940 VGND.n2939 0.120292
R6263 VGND.n2941 VGND.n2940 0.120292
R6264 VGND.n2941 VGND.n2924 0.120292
R6265 VGND.n2945 VGND.n2924 0.120292
R6266 VGND.n2947 VGND.n2921 0.120292
R6267 VGND.n2952 VGND.n2921 0.120292
R6268 VGND.n44 VGND.n38 0.120292
R6269 VGND.n49 VGND.n38 0.120292
R6270 VGND.n50 VGND.n49 0.120292
R6271 VGND.n51 VGND.n50 0.120292
R6272 VGND.n51 VGND.n36 0.120292
R6273 VGND.n55 VGND.n36 0.120292
R6274 VGND.n56 VGND.n55 0.120292
R6275 VGND.n2959 VGND.n2958 0.120292
R6276 VGND.n2958 VGND.n2957 0.120292
R6277 VGND.n2973 VGND.n2967 0.120292
R6278 VGND.n2978 VGND.n2967 0.120292
R6279 VGND.n2979 VGND.n2978 0.120292
R6280 VGND.n2980 VGND.n2979 0.120292
R6281 VGND.n2980 VGND.n2965 0.120292
R6282 VGND.n2984 VGND.n2965 0.120292
R6283 VGND.n2985 VGND.n2984 0.120292
R6284 VGND.n2991 VGND.n2990 0.120292
R6285 VGND.n2990 VGND.n2989 0.120292
R6286 VGND VGND.n2871 0.119536
R6287 VGND.n1094 VGND 0.117202
R6288 VGND.n1065 VGND 0.117202
R6289 VGND.n1003 VGND 0.117202
R6290 VGND.n1034 VGND 0.117202
R6291 VGND.n227 VGND.n226 0.110872
R6292 VGND.n2778 VGND.n2777 0.110872
R6293 VGND.n2773 VGND.n2772 0.110872
R6294 VGND.n2768 VGND.n2767 0.110872
R6295 VGND.n2763 VGND.n2762 0.110872
R6296 VGND.n2758 VGND.n2757 0.110872
R6297 VGND.n2753 VGND.n2752 0.110872
R6298 VGND.n2748 VGND.n2747 0.110872
R6299 VGND.n2743 VGND.n2742 0.110872
R6300 VGND.n2738 VGND.n2737 0.110872
R6301 VGND.n2733 VGND.n2732 0.110872
R6302 VGND.n2728 VGND.n2727 0.110872
R6303 VGND.n2723 VGND.n2722 0.110872
R6304 VGND.n2718 VGND.n2717 0.110872
R6305 VGND.n232 VGND.n231 0.110872
R6306 VGND.n2487 VGND.n2486 0.110872
R6307 VGND.n2482 VGND.n2481 0.110872
R6308 VGND.n2477 VGND.n2476 0.110872
R6309 VGND.n2472 VGND.n2471 0.110872
R6310 VGND.n2467 VGND.n2466 0.110872
R6311 VGND.n2462 VGND.n2461 0.110872
R6312 VGND.n2457 VGND.n2456 0.110872
R6313 VGND.n2452 VGND.n2451 0.110872
R6314 VGND.n2447 VGND.n2446 0.110872
R6315 VGND.n2442 VGND.n2441 0.110872
R6316 VGND.n2437 VGND.n2436 0.110872
R6317 VGND.n247 VGND.n246 0.110872
R6318 VGND.n2507 VGND.n2506 0.110872
R6319 VGND.n2512 VGND.n2511 0.110872
R6320 VGND.n242 VGND.n241 0.110872
R6321 VGND.n332 VGND.n331 0.110872
R6322 VGND.n2289 VGND.n2288 0.110872
R6323 VGND.n2284 VGND.n2283 0.110872
R6324 VGND.n2279 VGND.n2278 0.110872
R6325 VGND.n340 VGND.n339 0.110872
R6326 VGND.n2248 VGND.n2247 0.110872
R6327 VGND.n348 VGND.n347 0.110872
R6328 VGND.n2222 VGND.n2221 0.110872
R6329 VGND.n356 VGND.n355 0.110872
R6330 VGND.n2196 VGND.n2195 0.110872
R6331 VGND.n364 VGND.n363 0.110872
R6332 VGND.n2170 VGND.n2169 0.110872
R6333 VGND.n370 VGND.n369 0.110872
R6334 VGND.n367 VGND.n366 0.110872
R6335 VGND.n2830 VGND.n2829 0.110872
R6336 VGND.n2312 VGND.n2311 0.110872
R6337 VGND.n2306 VGND.n2305 0.110872
R6338 VGND.n2266 VGND.n2265 0.110872
R6339 VGND.n336 VGND.n335 0.110872
R6340 VGND.n2261 VGND.n2260 0.110872
R6341 VGND.n344 VGND.n343 0.110872
R6342 VGND.n2235 VGND.n2234 0.110872
R6343 VGND.n352 VGND.n351 0.110872
R6344 VGND.n2209 VGND.n2208 0.110872
R6345 VGND.n360 VGND.n359 0.110872
R6346 VGND.n2183 VGND.n2182 0.110872
R6347 VGND.n379 VGND.n378 0.110872
R6348 VGND.n2157 VGND.n2156 0.110872
R6349 VGND.n1424 VGND.n1423 0.110872
R6350 VGND.n1427 VGND.n1426 0.110872
R6351 VGND.n2129 VGND.n2128 0.110872
R6352 VGND.n2134 VGND.n2133 0.110872
R6353 VGND.n393 VGND.n392 0.110872
R6354 VGND.n1446 VGND.n1445 0.110872
R6355 VGND.n1451 VGND.n1450 0.110872
R6356 VGND.n1456 VGND.n1455 0.110872
R6357 VGND.n1461 VGND.n1460 0.110872
R6358 VGND.n1466 VGND.n1465 0.110872
R6359 VGND.n1471 VGND.n1470 0.110872
R6360 VGND.n1476 VGND.n1475 0.110872
R6361 VGND.n1481 VGND.n1480 0.110872
R6362 VGND.n1486 VGND.n1485 0.110872
R6363 VGND.n1491 VGND.n1490 0.110872
R6364 VGND.n634 VGND.n633 0.110872
R6365 VGND.n1441 VGND.n1440 0.110872
R6366 VGND.n2121 VGND.n2120 0.110872
R6367 VGND.n2115 VGND.n2114 0.110872
R6368 VGND.n2110 VGND.n2109 0.110872
R6369 VGND.n2105 VGND.n2104 0.110872
R6370 VGND.n407 VGND.n406 0.110872
R6371 VGND.n2074 VGND.n2073 0.110872
R6372 VGND.n415 VGND.n414 0.110872
R6373 VGND.n2048 VGND.n2047 0.110872
R6374 VGND.n423 VGND.n422 0.110872
R6375 VGND.n2022 VGND.n2021 0.110872
R6376 VGND.n431 VGND.n430 0.110872
R6377 VGND.n1996 VGND.n1995 0.110872
R6378 VGND.n625 VGND.n624 0.110872
R6379 VGND.n622 VGND.n621 0.110872
R6380 VGND.n1503 VGND.n1502 0.110872
R6381 VGND.n2337 VGND.n2336 0.110872
R6382 VGND.n2331 VGND.n2330 0.110872
R6383 VGND.n2092 VGND.n2091 0.110872
R6384 VGND.n403 VGND.n402 0.110872
R6385 VGND.n2087 VGND.n2086 0.110872
R6386 VGND.n411 VGND.n410 0.110872
R6387 VGND.n2061 VGND.n2060 0.110872
R6388 VGND.n419 VGND.n418 0.110872
R6389 VGND.n2035 VGND.n2034 0.110872
R6390 VGND.n427 VGND.n426 0.110872
R6391 VGND.n2009 VGND.n2008 0.110872
R6392 VGND.n435 VGND.n434 0.110872
R6393 VGND.n1983 VGND.n1982 0.110872
R6394 VGND.n647 VGND.n646 0.110872
R6395 VGND.n650 VGND.n649 0.110872
R6396 VGND.n1955 VGND.n1954 0.110872
R6397 VGND.n1960 VGND.n1959 0.110872
R6398 VGND.n449 VGND.n448 0.110872
R6399 VGND.n902 VGND.n901 0.110872
R6400 VGND.n907 VGND.n906 0.110872
R6401 VGND.n912 VGND.n911 0.110872
R6402 VGND.n917 VGND.n916 0.110872
R6403 VGND.n922 VGND.n921 0.110872
R6404 VGND.n927 VGND.n926 0.110872
R6405 VGND.n932 VGND.n931 0.110872
R6406 VGND.n937 VGND.n936 0.110872
R6407 VGND.n942 VGND.n941 0.110872
R6408 VGND.n947 VGND.n946 0.110872
R6409 VGND.n952 VGND.n951 0.110872
R6410 VGND.n957 VGND.n956 0.110872
R6411 VGND.n1947 VGND.n1946 0.110872
R6412 VGND.n1941 VGND.n1940 0.110872
R6413 VGND.n1936 VGND.n1935 0.110872
R6414 VGND.n1931 VGND.n1930 0.110872
R6415 VGND.n463 VGND.n462 0.110872
R6416 VGND.n1900 VGND.n1899 0.110872
R6417 VGND.n471 VGND.n470 0.110872
R6418 VGND.n1874 VGND.n1873 0.110872
R6419 VGND.n479 VGND.n478 0.110872
R6420 VGND.n1848 VGND.n1847 0.110872
R6421 VGND.n487 VGND.n486 0.110872
R6422 VGND.n1822 VGND.n1821 0.110872
R6423 VGND.n666 VGND.n665 0.110872
R6424 VGND.n1399 VGND.n1398 0.110872
R6425 VGND.n1394 VGND.n1393 0.110872
R6426 VGND.n2362 VGND.n2361 0.110872
R6427 VGND.n2356 VGND.n2355 0.110872
R6428 VGND.n1918 VGND.n1917 0.110872
R6429 VGND.n459 VGND.n458 0.110872
R6430 VGND.n1913 VGND.n1912 0.110872
R6431 VGND.n467 VGND.n466 0.110872
R6432 VGND.n1887 VGND.n1886 0.110872
R6433 VGND.n475 VGND.n474 0.110872
R6434 VGND.n1861 VGND.n1860 0.110872
R6435 VGND.n483 VGND.n482 0.110872
R6436 VGND.n1835 VGND.n1834 0.110872
R6437 VGND.n491 VGND.n490 0.110872
R6438 VGND.n1809 VGND.n1808 0.110872
R6439 VGND.n1376 VGND.n1375 0.110872
R6440 VGND.n1379 VGND.n1378 0.110872
R6441 VGND.n1781 VGND.n1780 0.110872
R6442 VGND.n1786 VGND.n1785 0.110872
R6443 VGND.n505 VGND.n504 0.110872
R6444 VGND.n1316 VGND.n1315 0.110872
R6445 VGND.n1321 VGND.n1320 0.110872
R6446 VGND.n1326 VGND.n1325 0.110872
R6447 VGND.n1331 VGND.n1330 0.110872
R6448 VGND.n1336 VGND.n1335 0.110872
R6449 VGND.n1341 VGND.n1340 0.110872
R6450 VGND.n1346 VGND.n1345 0.110872
R6451 VGND.n1351 VGND.n1350 0.110872
R6452 VGND.n1356 VGND.n1355 0.110872
R6453 VGND.n1361 VGND.n1360 0.110872
R6454 VGND.n1308 VGND.n1307 0.110872
R6455 VGND.n1311 VGND.n1310 0.110872
R6456 VGND.n1773 VGND.n1772 0.110872
R6457 VGND.n1767 VGND.n1766 0.110872
R6458 VGND.n1762 VGND.n1761 0.110872
R6459 VGND.n1757 VGND.n1756 0.110872
R6460 VGND.n519 VGND.n518 0.110872
R6461 VGND.n1726 VGND.n1725 0.110872
R6462 VGND.n527 VGND.n526 0.110872
R6463 VGND.n1700 VGND.n1699 0.110872
R6464 VGND.n535 VGND.n534 0.110872
R6465 VGND.n1674 VGND.n1673 0.110872
R6466 VGND.n543 VGND.n542 0.110872
R6467 VGND.n1648 VGND.n1647 0.110872
R6468 VGND.n577 VGND.n576 0.110872
R6469 VGND.n1521 VGND.n1520 0.110872
R6470 VGND.n1516 VGND.n1515 0.110872
R6471 VGND.n2387 VGND.n2386 0.110872
R6472 VGND.n2381 VGND.n2380 0.110872
R6473 VGND.n1744 VGND.n1743 0.110872
R6474 VGND.n515 VGND.n514 0.110872
R6475 VGND.n1739 VGND.n1738 0.110872
R6476 VGND.n523 VGND.n522 0.110872
R6477 VGND.n1713 VGND.n1712 0.110872
R6478 VGND.n531 VGND.n530 0.110872
R6479 VGND.n1687 VGND.n1686 0.110872
R6480 VGND.n539 VGND.n538 0.110872
R6481 VGND.n1661 VGND.n1660 0.110872
R6482 VGND.n547 VGND.n546 0.110872
R6483 VGND.n1635 VGND.n1634 0.110872
R6484 VGND.n566 VGND.n565 0.110872
R6485 VGND.n1536 VGND.n1535 0.110872
R6486 VGND.n1607 VGND.n1606 0.110872
R6487 VGND.n1612 VGND.n1611 0.110872
R6488 VGND.n561 VGND.n560 0.110872
R6489 VGND.n1599 VGND.n1598 0.110872
R6490 VGND.n1594 VGND.n1593 0.110872
R6491 VGND.n1589 VGND.n1588 0.110872
R6492 VGND.n1584 VGND.n1583 0.110872
R6493 VGND.n1579 VGND.n1578 0.110872
R6494 VGND.n1574 VGND.n1573 0.110872
R6495 VGND.n1569 VGND.n1568 0.110872
R6496 VGND.n1564 VGND.n1563 0.110872
R6497 VGND.n1559 VGND.n1558 0.110872
R6498 VGND.n1554 VGND.n1553 0.110872
R6499 VGND.n1549 VGND.n1548 0.110872
R6500 VGND.n674 VGND.n673 0.110872
R6501 VGND.n2407 VGND.n2406 0.110872
R6502 VGND.n2401 VGND.n2400 0.110872
R6503 VGND.n843 VGND.n842 0.110872
R6504 VGND.n848 VGND.n847 0.110872
R6505 VGND.n853 VGND.n852 0.110872
R6506 VGND.n858 VGND.n857 0.110872
R6507 VGND.n863 VGND.n862 0.110872
R6508 VGND.n868 VGND.n867 0.110872
R6509 VGND.n873 VGND.n872 0.110872
R6510 VGND.n878 VGND.n877 0.110872
R6511 VGND.n883 VGND.n882 0.110872
R6512 VGND.n888 VGND.n887 0.110872
R6513 VGND.n830 VGND.n829 0.110872
R6514 VGND.n838 VGND.n837 0.110872
R6515 VGND.n833 VGND.n832 0.110872
R6516 VGND.n1126 VGND.n1125 0.110872
R6517 VGND.n1130 VGND.n1129 0.110872
R6518 VGND.n1136 VGND.n1135 0.110872
R6519 VGND.n1143 VGND.n1142 0.110872
R6520 VGND.n810 VGND.n809 0.110872
R6521 VGND.n1162 VGND.n1161 0.110872
R6522 VGND.n1168 VGND.n1167 0.110872
R6523 VGND.n1175 VGND.n1174 0.110872
R6524 VGND.n802 VGND.n801 0.110872
R6525 VGND.n1194 VGND.n1193 0.110872
R6526 VGND.n1200 VGND.n1199 0.110872
R6527 VGND.n1207 VGND.n1206 0.110872
R6528 VGND.n794 VGND.n793 0.110872
R6529 VGND.n1226 VGND.n1225 0.110872
R6530 VGND.n1232 VGND.n1231 0.110872
R6531 VGND.n719 VGND.n718 0.110872
R6532 VGND.n778 VGND.n777 0.110872
R6533 VGND.n773 VGND.n772 0.110872
R6534 VGND.n768 VGND.n767 0.110872
R6535 VGND.n763 VGND.n762 0.110872
R6536 VGND.n758 VGND.n757 0.110872
R6537 VGND.n753 VGND.n752 0.110872
R6538 VGND.n748 VGND.n747 0.110872
R6539 VGND.n743 VGND.n742 0.110872
R6540 VGND.n738 VGND.n737 0.110872
R6541 VGND.n733 VGND.n732 0.110872
R6542 VGND.n728 VGND.n727 0.110872
R6543 VGND.n723 VGND.n722 0.110872
R6544 VGND.n684 VGND.n683 0.110872
R6545 VGND.n1288 VGND.n1287 0.110872
R6546 VGND.n1086 VGND 0.0981562
R6547 VGND.n994 VGND 0.0981562
R6548 VGND.n1055 VGND 0.0981562
R6549 VGND VGND.n143 0.0968542
R6550 VGND VGND.n611 0.0968542
R6551 VGND VGND.n987 0.0968542
R6552 VGND.n1024 VGND 0.0968542
R6553 VGND VGND.n173 0.0968542
R6554 VGND.n15 VGND 0.0968542
R6555 VGND VGND.n2904 0.0968542
R6556 VGND VGND.n60 0.0968542
R6557 VGND.n2933 VGND 0.0968542
R6558 VGND.n44 VGND 0.0968542
R6559 VGND.n2973 VGND 0.0968542
R6560 VGND.n2521 VGND 0.088625
R6561 VGND.n2711 VGND 0.0790114
R6562 VGND VGND.n2710 0.0790114
R6563 VGND VGND.n188 0.0790114
R6564 VGND.n2817 VGND 0.0790114
R6565 VGND VGND.n2816 0.0790114
R6566 VGND.n2811 VGND 0.0790114
R6567 VGND VGND.n2810 0.0790114
R6568 VGND.n2805 VGND 0.0790114
R6569 VGND VGND.n2804 0.0790114
R6570 VGND.n2799 VGND 0.0790114
R6571 VGND VGND.n2798 0.0790114
R6572 VGND.n2793 VGND 0.0790114
R6573 VGND VGND.n2792 0.0790114
R6574 VGND.n2787 VGND 0.0790114
R6575 VGND VGND.n2786 0.0790114
R6576 VGND.n3004 VGND 0.0790114
R6577 VGND.n2713 VGND 0.0790114
R6578 VGND.n2714 VGND 0.0790114
R6579 VGND.n2820 VGND 0.0790114
R6580 VGND VGND.n2819 0.0790114
R6581 VGND.n2814 VGND 0.0790114
R6582 VGND VGND.n2813 0.0790114
R6583 VGND.n2808 VGND 0.0790114
R6584 VGND VGND.n2807 0.0790114
R6585 VGND.n2802 VGND 0.0790114
R6586 VGND VGND.n2801 0.0790114
R6587 VGND.n2796 VGND 0.0790114
R6588 VGND VGND.n2795 0.0790114
R6589 VGND.n2790 VGND 0.0790114
R6590 VGND VGND.n2789 0.0790114
R6591 VGND.n2784 VGND 0.0790114
R6592 VGND.n3002 VGND 0.0790114
R6593 VGND VGND.n2518 0.0790114
R6594 VGND.n2824 VGND 0.0790114
R6595 VGND VGND.n2823 0.0790114
R6596 VGND.n2504 VGND 0.0790114
R6597 VGND VGND.n2503 0.0790114
R6598 VGND VGND.n2502 0.0790114
R6599 VGND VGND.n2501 0.0790114
R6600 VGND VGND.n2500 0.0790114
R6601 VGND VGND.n2499 0.0790114
R6602 VGND VGND.n2498 0.0790114
R6603 VGND VGND.n2497 0.0790114
R6604 VGND VGND.n2496 0.0790114
R6605 VGND VGND.n2495 0.0790114
R6606 VGND VGND.n2494 0.0790114
R6607 VGND VGND.n2493 0.0790114
R6608 VGND VGND.n2492 0.0790114
R6609 VGND.n639 VGND 0.0790114
R6610 VGND.n2827 VGND 0.0790114
R6611 VGND.n375 VGND 0.0790114
R6612 VGND.n2166 VGND 0.0790114
R6613 VGND.n2176 VGND 0.0790114
R6614 VGND.n2192 VGND 0.0790114
R6615 VGND.n2202 VGND 0.0790114
R6616 VGND.n2218 VGND 0.0790114
R6617 VGND.n2228 VGND 0.0790114
R6618 VGND.n2244 VGND 0.0790114
R6619 VGND.n2254 VGND 0.0790114
R6620 VGND.n2275 VGND 0.0790114
R6621 VGND.n2298 VGND 0.0790114
R6622 VGND VGND.n2297 0.0790114
R6623 VGND VGND.n2295 0.0790114
R6624 VGND.n2431 VGND 0.0790114
R6625 VGND.n1434 VGND 0.0790114
R6626 VGND VGND.n1433 0.0790114
R6627 VGND.n2153 VGND 0.0790114
R6628 VGND.n2163 VGND 0.0790114
R6629 VGND.n2179 VGND 0.0790114
R6630 VGND.n2189 VGND 0.0790114
R6631 VGND.n2205 VGND 0.0790114
R6632 VGND.n2215 VGND 0.0790114
R6633 VGND.n2231 VGND 0.0790114
R6634 VGND.n2241 VGND 0.0790114
R6635 VGND.n2257 VGND 0.0790114
R6636 VGND.n2272 VGND 0.0790114
R6637 VGND.n2301 VGND 0.0790114
R6638 VGND.n2302 VGND 0.0790114
R6639 VGND.n2315 VGND 0.0790114
R6640 VGND VGND.n2314 0.0790114
R6641 VGND.n1437 VGND 0.0790114
R6642 VGND.n1497 VGND 0.0790114
R6643 VGND.n2150 VGND 0.0790114
R6644 VGND VGND.n2149 0.0790114
R6645 VGND VGND.n2148 0.0790114
R6646 VGND VGND.n2147 0.0790114
R6647 VGND VGND.n2146 0.0790114
R6648 VGND VGND.n2145 0.0790114
R6649 VGND VGND.n2144 0.0790114
R6650 VGND VGND.n2143 0.0790114
R6651 VGND VGND.n2142 0.0790114
R6652 VGND VGND.n2141 0.0790114
R6653 VGND VGND.n2140 0.0790114
R6654 VGND.n2319 VGND 0.0790114
R6655 VGND VGND.n2318 0.0790114
R6656 VGND.n2126 VGND 0.0790114
R6657 VGND VGND.n1415 0.0790114
R6658 VGND.n1500 VGND 0.0790114
R6659 VGND VGND.n630 0.0790114
R6660 VGND.n1992 VGND 0.0790114
R6661 VGND.n2002 VGND 0.0790114
R6662 VGND.n2018 VGND 0.0790114
R6663 VGND.n2028 VGND 0.0790114
R6664 VGND.n2044 VGND 0.0790114
R6665 VGND.n2054 VGND 0.0790114
R6666 VGND.n2070 VGND 0.0790114
R6667 VGND.n2080 VGND 0.0790114
R6668 VGND.n2101 VGND 0.0790114
R6669 VGND.n2323 VGND 0.0790114
R6670 VGND VGND.n2322 0.0790114
R6671 VGND.n398 VGND 0.0790114
R6672 VGND.n2123 VGND 0.0790114
R6673 VGND VGND.n1413 0.0790114
R6674 VGND VGND.n656 0.0790114
R6675 VGND.n1979 VGND 0.0790114
R6676 VGND.n1989 VGND 0.0790114
R6677 VGND.n2005 VGND 0.0790114
R6678 VGND.n2015 VGND 0.0790114
R6679 VGND.n2031 VGND 0.0790114
R6680 VGND.n2041 VGND 0.0790114
R6681 VGND.n2057 VGND 0.0790114
R6682 VGND.n2067 VGND 0.0790114
R6683 VGND.n2083 VGND 0.0790114
R6684 VGND.n2098 VGND 0.0790114
R6685 VGND.n2326 VGND 0.0790114
R6686 VGND.n2327 VGND 0.0790114
R6687 VGND.n2340 VGND 0.0790114
R6688 VGND VGND.n2339 0.0790114
R6689 VGND.n1410 VGND 0.0790114
R6690 VGND VGND.n1409 0.0790114
R6691 VGND.n1976 VGND 0.0790114
R6692 VGND VGND.n1975 0.0790114
R6693 VGND VGND.n1974 0.0790114
R6694 VGND VGND.n1973 0.0790114
R6695 VGND VGND.n1972 0.0790114
R6696 VGND VGND.n1971 0.0790114
R6697 VGND VGND.n1970 0.0790114
R6698 VGND VGND.n1969 0.0790114
R6699 VGND VGND.n1968 0.0790114
R6700 VGND VGND.n1967 0.0790114
R6701 VGND VGND.n1966 0.0790114
R6702 VGND.n2344 VGND 0.0790114
R6703 VGND VGND.n2343 0.0790114
R6704 VGND.n1952 VGND 0.0790114
R6705 VGND.n1390 VGND 0.0790114
R6706 VGND.n1406 VGND 0.0790114
R6707 VGND VGND.n1405 0.0790114
R6708 VGND.n1818 VGND 0.0790114
R6709 VGND.n1828 VGND 0.0790114
R6710 VGND.n1844 VGND 0.0790114
R6711 VGND.n1854 VGND 0.0790114
R6712 VGND.n1870 VGND 0.0790114
R6713 VGND.n1880 VGND 0.0790114
R6714 VGND.n1896 VGND 0.0790114
R6715 VGND.n1906 VGND 0.0790114
R6716 VGND.n1927 VGND 0.0790114
R6717 VGND.n2348 VGND 0.0790114
R6718 VGND VGND.n2347 0.0790114
R6719 VGND.n454 VGND 0.0790114
R6720 VGND.n1949 VGND 0.0790114
R6721 VGND VGND.n1387 0.0790114
R6722 VGND VGND.n1385 0.0790114
R6723 VGND.n1805 VGND 0.0790114
R6724 VGND.n1815 VGND 0.0790114
R6725 VGND.n1831 VGND 0.0790114
R6726 VGND.n1841 VGND 0.0790114
R6727 VGND.n1857 VGND 0.0790114
R6728 VGND.n1867 VGND 0.0790114
R6729 VGND.n1883 VGND 0.0790114
R6730 VGND.n1893 VGND 0.0790114
R6731 VGND.n1909 VGND 0.0790114
R6732 VGND.n1924 VGND 0.0790114
R6733 VGND.n2351 VGND 0.0790114
R6734 VGND.n2352 VGND 0.0790114
R6735 VGND.n2365 VGND 0.0790114
R6736 VGND VGND.n2364 0.0790114
R6737 VGND VGND.n1369 0.0790114
R6738 VGND VGND.n1368 0.0790114
R6739 VGND.n1802 VGND 0.0790114
R6740 VGND VGND.n1801 0.0790114
R6741 VGND VGND.n1800 0.0790114
R6742 VGND VGND.n1799 0.0790114
R6743 VGND VGND.n1798 0.0790114
R6744 VGND VGND.n1797 0.0790114
R6745 VGND VGND.n1796 0.0790114
R6746 VGND VGND.n1795 0.0790114
R6747 VGND VGND.n1794 0.0790114
R6748 VGND VGND.n1793 0.0790114
R6749 VGND VGND.n1792 0.0790114
R6750 VGND.n2369 VGND 0.0790114
R6751 VGND VGND.n2368 0.0790114
R6752 VGND.n1778 VGND 0.0790114
R6753 VGND.n1529 VGND 0.0790114
R6754 VGND VGND.n1528 0.0790114
R6755 VGND VGND.n1527 0.0790114
R6756 VGND.n1644 VGND 0.0790114
R6757 VGND.n1654 VGND 0.0790114
R6758 VGND.n1670 VGND 0.0790114
R6759 VGND.n1680 VGND 0.0790114
R6760 VGND.n1696 VGND 0.0790114
R6761 VGND.n1706 VGND 0.0790114
R6762 VGND.n1722 VGND 0.0790114
R6763 VGND.n1732 VGND 0.0790114
R6764 VGND.n1753 VGND 0.0790114
R6765 VGND.n2373 VGND 0.0790114
R6766 VGND VGND.n2372 0.0790114
R6767 VGND.n510 VGND 0.0790114
R6768 VGND.n1775 VGND 0.0790114
R6769 VGND.n1532 VGND 0.0790114
R6770 VGND.n1542 VGND 0.0790114
R6771 VGND.n1631 VGND 0.0790114
R6772 VGND.n1641 VGND 0.0790114
R6773 VGND.n1657 VGND 0.0790114
R6774 VGND.n1667 VGND 0.0790114
R6775 VGND.n1683 VGND 0.0790114
R6776 VGND.n1693 VGND 0.0790114
R6777 VGND.n1709 VGND 0.0790114
R6778 VGND.n1719 VGND 0.0790114
R6779 VGND.n1735 VGND 0.0790114
R6780 VGND.n1750 VGND 0.0790114
R6781 VGND.n2376 VGND 0.0790114
R6782 VGND.n2377 VGND 0.0790114
R6783 VGND.n2390 VGND 0.0790114
R6784 VGND VGND.n2389 0.0790114
R6785 VGND VGND.n1299 0.0790114
R6786 VGND.n1545 VGND 0.0790114
R6787 VGND.n1628 VGND 0.0790114
R6788 VGND VGND.n1627 0.0790114
R6789 VGND VGND.n1626 0.0790114
R6790 VGND VGND.n1625 0.0790114
R6791 VGND VGND.n1624 0.0790114
R6792 VGND VGND.n1623 0.0790114
R6793 VGND VGND.n1622 0.0790114
R6794 VGND VGND.n1621 0.0790114
R6795 VGND VGND.n1620 0.0790114
R6796 VGND VGND.n1619 0.0790114
R6797 VGND VGND.n1618 0.0790114
R6798 VGND.n2394 VGND 0.0790114
R6799 VGND VGND.n2393 0.0790114
R6800 VGND.n1604 VGND 0.0790114
R6801 VGND.n896 VGND 0.0790114
R6802 VGND VGND.n895 0.0790114
R6803 VGND VGND.n894 0.0790114
R6804 VGND.n1276 VGND 0.0790114
R6805 VGND VGND.n1275 0.0790114
R6806 VGND.n1268 VGND 0.0790114
R6807 VGND VGND.n1267 0.0790114
R6808 VGND.n1260 VGND 0.0790114
R6809 VGND VGND.n1259 0.0790114
R6810 VGND.n1252 VGND 0.0790114
R6811 VGND VGND.n1251 0.0790114
R6812 VGND.n1244 VGND 0.0790114
R6813 VGND VGND.n1243 0.0790114
R6814 VGND.n2397 VGND 0.0790114
R6815 VGND.n284 VGND 0.0790114
R6816 VGND.n2409 VGND 0.0790114
R6817 VGND.n1120 VGND 0.0790114
R6818 VGND.n1283 VGND 0.0790114
R6819 VGND VGND.n1282 0.0790114
R6820 VGND.n687 VGND 0.0790114
R6821 VGND.n690 VGND 0.0790114
R6822 VGND.n693 VGND 0.0790114
R6823 VGND.n696 VGND 0.0790114
R6824 VGND.n699 VGND 0.0790114
R6825 VGND.n702 VGND 0.0790114
R6826 VGND.n705 VGND 0.0790114
R6827 VGND.n708 VGND 0.0790114
R6828 VGND.n711 VGND 0.0790114
R6829 VGND.n714 VGND 0.0790114
R6830 VGND.n1221 VGND 0.0790114
R6831 VGND.n1236 VGND 0.0790114
R6832 VGND VGND.n1235 0.0790114
R6833 VGND.n1118 VGND 0.0790114
R6834 VGND.n1285 VGND 0.0790114
R6835 VGND.n1280 VGND 0.0790114
R6836 VGND VGND.n1279 0.0790114
R6837 VGND.n1272 VGND 0.0790114
R6838 VGND VGND.n1271 0.0790114
R6839 VGND.n1264 VGND 0.0790114
R6840 VGND VGND.n1263 0.0790114
R6841 VGND.n1256 VGND 0.0790114
R6842 VGND VGND.n1255 0.0790114
R6843 VGND.n1248 VGND 0.0790114
R6844 VGND VGND.n1247 0.0790114
R6845 VGND.n1240 VGND 0.0790114
R6846 VGND VGND.n1239 0.0790114
R6847 VGND VGND.n1238 0.0790114
R6848 VGND.n2412 VGND 0.0790114
R6849 VGND.n3024 VGND.n3023 0.0732323
R6850 VGND.n2655 VGND.n2654 0.0656596
R6851 VGND.n2650 VGND.n2648 0.0656596
R6852 VGND.n2663 VGND.n2662 0.0656596
R6853 VGND.n2646 VGND.n2644 0.0656596
R6854 VGND.n2671 VGND.n2670 0.0656596
R6855 VGND.n2642 VGND.n2640 0.0656596
R6856 VGND.n2679 VGND.n2678 0.0656596
R6857 VGND.n2638 VGND.n2636 0.0656596
R6858 VGND.n2687 VGND.n2686 0.0656596
R6859 VGND.n2634 VGND.n2632 0.0656596
R6860 VGND.n2695 VGND.n2694 0.0656596
R6861 VGND.n2630 VGND.n2628 0.0656596
R6862 VGND.n2703 VGND.n2702 0.0656596
R6863 VGND.n2581 VGND.n2573 0.0656596
R6864 VGND.n2577 VGND.n2572 0.0656596
R6865 VGND.n2565 VGND 0.063
R6866 VGND.n2562 VGND 0.063
R6867 VGND.n2559 VGND 0.063
R6868 VGND.n2556 VGND 0.063
R6869 VGND.n2553 VGND 0.063
R6870 VGND.n2550 VGND 0.063
R6871 VGND.n2547 VGND 0.063
R6872 VGND.n2544 VGND 0.063
R6873 VGND.n2541 VGND 0.063
R6874 VGND.n2538 VGND 0.063
R6875 VGND.n2535 VGND 0.063
R6876 VGND.n2532 VGND 0.063
R6877 VGND.n2529 VGND 0.063
R6878 VGND.n2526 VGND 0.063
R6879 VGND.n2523 VGND 0.063
R6880 VGND.n1108 VGND 0.0603958
R6881 VGND.n1085 VGND 0.0603958
R6882 VGND VGND.n1084 0.0603958
R6883 VGND.n1081 VGND 0.0603958
R6884 VGND.n145 VGND 0.0603958
R6885 VGND VGND.n144 0.0603958
R6886 VGND.n127 VGND 0.0603958
R6887 VGND.n613 VGND 0.0603958
R6888 VGND VGND.n612 0.0603958
R6889 VGND.n595 VGND 0.0603958
R6890 VGND.n989 VGND 0.0603958
R6891 VGND VGND.n988 0.0603958
R6892 VGND.n981 VGND 0.0603958
R6893 VGND.n978 VGND 0.0603958
R6894 VGND.n973 VGND 0.0603958
R6895 VGND.n1023 VGND 0.0603958
R6896 VGND VGND.n1022 0.0603958
R6897 VGND.n1019 VGND 0.0603958
R6898 VGND.n1054 VGND 0.0603958
R6899 VGND VGND.n1053 0.0603958
R6900 VGND.n1050 VGND 0.0603958
R6901 VGND.n175 VGND 0.0603958
R6902 VGND VGND.n174 0.0603958
R6903 VGND.n157 VGND 0.0603958
R6904 VGND VGND.n27 0.0603958
R6905 VGND.n3007 VGND 0.0603958
R6906 VGND.n111 VGND 0.0603958
R6907 VGND VGND.n110 0.0603958
R6908 VGND.n2873 VGND 0.0603958
R6909 VGND VGND.n2872 0.0603958
R6910 VGND.n2906 VGND 0.0603958
R6911 VGND VGND.n2905 0.0603958
R6912 VGND.n2901 VGND 0.0603958
R6913 VGND.n2913 VGND 0.0603958
R6914 VGND.n2914 VGND 0.0603958
R6915 VGND VGND.n2945 0.0603958
R6916 VGND.n2946 VGND 0.0603958
R6917 VGND.n2947 VGND 0.0603958
R6918 VGND VGND.n56 0.0603958
R6919 VGND.n57 VGND 0.0603958
R6920 VGND.n2959 VGND 0.0603958
R6921 VGND VGND.n2985 0.0603958
R6922 VGND.n2986 VGND 0.0603958
R6923 VGND.n2991 VGND 0.0603958
R6924 VGND.n2654 VGND 0.0574853
R6925 VGND.n2650 VGND 0.0574853
R6926 VGND.n2662 VGND 0.0574853
R6927 VGND.n2646 VGND 0.0574853
R6928 VGND.n2670 VGND 0.0574853
R6929 VGND.n2642 VGND 0.0574853
R6930 VGND.n2678 VGND 0.0574853
R6931 VGND.n2638 VGND 0.0574853
R6932 VGND.n2686 VGND 0.0574853
R6933 VGND.n2634 VGND 0.0574853
R6934 VGND.n2694 VGND 0.0574853
R6935 VGND.n2630 VGND 0.0574853
R6936 VGND.n2702 VGND 0.0574853
R6937 VGND.n2581 VGND 0.0574853
R6938 VGND.n2572 VGND 0.0574853
R6939 VGND.n822 VGND 0.0489375
R6940 VGND.n785 VGND 0.0489375
R6941 VGND.n2586 VGND 0.0489375
R6942 VGND.n2583 VGND 0.0489375
R6943 VGND.n2569 VGND 0.0489375
R6944 VGND.n2582 VGND 0.0489375
R6945 VGND.n2621 VGND 0.0489375
R6946 VGND.n2618 VGND 0.0489375
R6947 VGND.n2615 VGND 0.0489375
R6948 VGND.n2612 VGND 0.0489375
R6949 VGND.n2609 VGND 0.0489375
R6950 VGND.n2606 VGND 0.0489375
R6951 VGND.n2603 VGND 0.0489375
R6952 VGND.n2600 VGND 0.0489375
R6953 VGND.n2597 VGND 0.0489375
R6954 VGND.n2594 VGND 0.0489375
R6955 VGND.n2591 VGND 0.0489375
R6956 VGND.n2588 VGND 0.0489375
R6957 VGND.n819 VGND 0.0489375
R6958 VGND.n816 VGND 0.0489375
R6959 VGND.n1137 VGND 0.0489375
R6960 VGND.n807 VGND 0.0489375
R6961 VGND.n805 VGND 0.0489375
R6962 VGND.n1152 VGND 0.0489375
R6963 VGND.n1169 VGND 0.0489375
R6964 VGND.n799 VGND 0.0489375
R6965 VGND.n797 VGND 0.0489375
R6966 VGND.n1184 VGND 0.0489375
R6967 VGND.n1201 VGND 0.0489375
R6968 VGND.n791 VGND 0.0489375
R6969 VGND.n789 VGND 0.0489375
R6970 VGND.n1216 VGND 0.0489375
R6971 VGND VGND.n2575 0.037734
R6972 VGND.n226 VGND 0.037734
R6973 VGND.n2777 VGND 0.037734
R6974 VGND.n2772 VGND 0.037734
R6975 VGND.n2767 VGND 0.037734
R6976 VGND.n2762 VGND 0.037734
R6977 VGND.n2757 VGND 0.037734
R6978 VGND.n2752 VGND 0.037734
R6979 VGND.n2747 VGND 0.037734
R6980 VGND.n2742 VGND 0.037734
R6981 VGND.n2737 VGND 0.037734
R6982 VGND.n2732 VGND 0.037734
R6983 VGND.n2727 VGND 0.037734
R6984 VGND.n2722 VGND 0.037734
R6985 VGND.n2717 VGND 0.037734
R6986 VGND.n231 VGND 0.037734
R6987 VGND VGND.n229 0.037734
R6988 VGND.n2486 VGND 0.037734
R6989 VGND.n2481 VGND 0.037734
R6990 VGND.n2476 VGND 0.037734
R6991 VGND.n2471 VGND 0.037734
R6992 VGND.n2466 VGND 0.037734
R6993 VGND.n2461 VGND 0.037734
R6994 VGND.n2456 VGND 0.037734
R6995 VGND.n2451 VGND 0.037734
R6996 VGND.n2446 VGND 0.037734
R6997 VGND.n2441 VGND 0.037734
R6998 VGND.n2436 VGND 0.037734
R6999 VGND VGND.n247 0.037734
R7000 VGND.n2506 VGND 0.037734
R7001 VGND.n2511 VGND 0.037734
R7002 VGND.n241 VGND 0.037734
R7003 VGND VGND.n239 0.037734
R7004 VGND.n331 VGND 0.037734
R7005 VGND.n2288 VGND 0.037734
R7006 VGND.n2283 VGND 0.037734
R7007 VGND.n2278 VGND 0.037734
R7008 VGND.n339 VGND 0.037734
R7009 VGND.n2247 VGND 0.037734
R7010 VGND.n347 VGND 0.037734
R7011 VGND.n2221 VGND 0.037734
R7012 VGND.n355 VGND 0.037734
R7013 VGND.n2195 VGND 0.037734
R7014 VGND.n363 VGND 0.037734
R7015 VGND.n2169 VGND 0.037734
R7016 VGND.n369 VGND 0.037734
R7017 VGND VGND.n367 0.037734
R7018 VGND.n2829 VGND 0.037734
R7019 VGND VGND.n179 0.037734
R7020 VGND VGND.n2312 0.037734
R7021 VGND.n2305 VGND 0.037734
R7022 VGND.n2265 VGND 0.037734
R7023 VGND.n335 VGND 0.037734
R7024 VGND.n2260 VGND 0.037734
R7025 VGND.n343 VGND 0.037734
R7026 VGND.n2234 VGND 0.037734
R7027 VGND.n351 VGND 0.037734
R7028 VGND.n2208 VGND 0.037734
R7029 VGND.n359 VGND 0.037734
R7030 VGND.n2182 VGND 0.037734
R7031 VGND.n378 VGND 0.037734
R7032 VGND.n2156 VGND 0.037734
R7033 VGND.n1423 VGND 0.037734
R7034 VGND.n1426 VGND 0.037734
R7035 VGND VGND.n1420 0.037734
R7036 VGND.n2128 VGND 0.037734
R7037 VGND.n2133 VGND 0.037734
R7038 VGND.n392 VGND 0.037734
R7039 VGND.n1445 VGND 0.037734
R7040 VGND.n1450 VGND 0.037734
R7041 VGND.n1455 VGND 0.037734
R7042 VGND.n1460 VGND 0.037734
R7043 VGND.n1465 VGND 0.037734
R7044 VGND.n1470 VGND 0.037734
R7045 VGND.n1475 VGND 0.037734
R7046 VGND.n1480 VGND 0.037734
R7047 VGND.n1485 VGND 0.037734
R7048 VGND.n1490 VGND 0.037734
R7049 VGND.n633 VGND 0.037734
R7050 VGND.n1440 VGND 0.037734
R7051 VGND VGND.n637 0.037734
R7052 VGND VGND.n2121 0.037734
R7053 VGND.n2114 VGND 0.037734
R7054 VGND.n2109 VGND 0.037734
R7055 VGND.n2104 VGND 0.037734
R7056 VGND.n406 VGND 0.037734
R7057 VGND.n2073 VGND 0.037734
R7058 VGND.n414 VGND 0.037734
R7059 VGND.n2047 VGND 0.037734
R7060 VGND.n422 VGND 0.037734
R7061 VGND.n2021 VGND 0.037734
R7062 VGND.n430 VGND 0.037734
R7063 VGND.n1995 VGND 0.037734
R7064 VGND.n624 VGND 0.037734
R7065 VGND VGND.n622 0.037734
R7066 VGND.n1502 VGND 0.037734
R7067 VGND VGND.n616 0.037734
R7068 VGND VGND.n2337 0.037734
R7069 VGND.n2330 VGND 0.037734
R7070 VGND.n2091 VGND 0.037734
R7071 VGND.n402 VGND 0.037734
R7072 VGND.n2086 VGND 0.037734
R7073 VGND.n410 VGND 0.037734
R7074 VGND.n2060 VGND 0.037734
R7075 VGND.n418 VGND 0.037734
R7076 VGND.n2034 VGND 0.037734
R7077 VGND.n426 VGND 0.037734
R7078 VGND.n2008 VGND 0.037734
R7079 VGND.n434 VGND 0.037734
R7080 VGND.n1982 VGND 0.037734
R7081 VGND.n646 VGND 0.037734
R7082 VGND.n649 VGND 0.037734
R7083 VGND VGND.n643 0.037734
R7084 VGND.n1954 VGND 0.037734
R7085 VGND.n1959 VGND 0.037734
R7086 VGND.n448 VGND 0.037734
R7087 VGND.n901 VGND 0.037734
R7088 VGND.n906 VGND 0.037734
R7089 VGND.n911 VGND 0.037734
R7090 VGND.n916 VGND 0.037734
R7091 VGND.n921 VGND 0.037734
R7092 VGND.n926 VGND 0.037734
R7093 VGND.n931 VGND 0.037734
R7094 VGND.n936 VGND 0.037734
R7095 VGND.n941 VGND 0.037734
R7096 VGND.n946 VGND 0.037734
R7097 VGND.n951 VGND 0.037734
R7098 VGND.n956 VGND 0.037734
R7099 VGND VGND.n659 0.037734
R7100 VGND VGND.n1947 0.037734
R7101 VGND.n1940 VGND 0.037734
R7102 VGND.n1935 VGND 0.037734
R7103 VGND.n1930 VGND 0.037734
R7104 VGND.n462 VGND 0.037734
R7105 VGND.n1899 VGND 0.037734
R7106 VGND.n470 VGND 0.037734
R7107 VGND.n1873 VGND 0.037734
R7108 VGND.n478 VGND 0.037734
R7109 VGND.n1847 VGND 0.037734
R7110 VGND.n486 VGND 0.037734
R7111 VGND.n1821 VGND 0.037734
R7112 VGND.n665 VGND 0.037734
R7113 VGND.n1398 VGND 0.037734
R7114 VGND.n1393 VGND 0.037734
R7115 VGND VGND.n668 0.037734
R7116 VGND VGND.n2362 0.037734
R7117 VGND.n2355 VGND 0.037734
R7118 VGND.n1917 VGND 0.037734
R7119 VGND.n458 VGND 0.037734
R7120 VGND.n1912 VGND 0.037734
R7121 VGND.n466 VGND 0.037734
R7122 VGND.n1886 VGND 0.037734
R7123 VGND.n474 VGND 0.037734
R7124 VGND.n1860 VGND 0.037734
R7125 VGND.n482 VGND 0.037734
R7126 VGND.n1834 VGND 0.037734
R7127 VGND.n490 VGND 0.037734
R7128 VGND.n1808 VGND 0.037734
R7129 VGND.n1375 VGND 0.037734
R7130 VGND.n1378 VGND 0.037734
R7131 VGND VGND.n1372 0.037734
R7132 VGND.n1780 VGND 0.037734
R7133 VGND.n1785 VGND 0.037734
R7134 VGND.n504 VGND 0.037734
R7135 VGND.n1315 VGND 0.037734
R7136 VGND.n1320 VGND 0.037734
R7137 VGND.n1325 VGND 0.037734
R7138 VGND.n1330 VGND 0.037734
R7139 VGND.n1335 VGND 0.037734
R7140 VGND.n1340 VGND 0.037734
R7141 VGND.n1345 VGND 0.037734
R7142 VGND.n1350 VGND 0.037734
R7143 VGND.n1355 VGND 0.037734
R7144 VGND.n1360 VGND 0.037734
R7145 VGND.n1307 VGND 0.037734
R7146 VGND.n1310 VGND 0.037734
R7147 VGND VGND.n1304 0.037734
R7148 VGND VGND.n1773 0.037734
R7149 VGND.n1766 VGND 0.037734
R7150 VGND.n1761 VGND 0.037734
R7151 VGND.n1756 VGND 0.037734
R7152 VGND.n518 VGND 0.037734
R7153 VGND.n1725 VGND 0.037734
R7154 VGND.n526 VGND 0.037734
R7155 VGND.n1699 VGND 0.037734
R7156 VGND.n534 VGND 0.037734
R7157 VGND.n1673 VGND 0.037734
R7158 VGND.n542 VGND 0.037734
R7159 VGND.n1647 VGND 0.037734
R7160 VGND.n576 VGND 0.037734
R7161 VGND.n1520 VGND 0.037734
R7162 VGND.n1515 VGND 0.037734
R7163 VGND VGND.n572 0.037734
R7164 VGND VGND.n2387 0.037734
R7165 VGND.n2380 VGND 0.037734
R7166 VGND.n1743 VGND 0.037734
R7167 VGND.n514 VGND 0.037734
R7168 VGND.n1738 VGND 0.037734
R7169 VGND.n522 VGND 0.037734
R7170 VGND.n1712 VGND 0.037734
R7171 VGND.n530 VGND 0.037734
R7172 VGND.n1686 VGND 0.037734
R7173 VGND.n538 VGND 0.037734
R7174 VGND.n1660 VGND 0.037734
R7175 VGND.n546 VGND 0.037734
R7176 VGND.n1634 VGND 0.037734
R7177 VGND.n565 VGND 0.037734
R7178 VGND.n1535 VGND 0.037734
R7179 VGND VGND.n568 0.037734
R7180 VGND.n1606 VGND 0.037734
R7181 VGND.n1611 VGND 0.037734
R7182 VGND.n560 VGND 0.037734
R7183 VGND.n1598 VGND 0.037734
R7184 VGND.n1593 VGND 0.037734
R7185 VGND.n1588 VGND 0.037734
R7186 VGND.n1583 VGND 0.037734
R7187 VGND.n1578 VGND 0.037734
R7188 VGND.n1573 VGND 0.037734
R7189 VGND.n1568 VGND 0.037734
R7190 VGND.n1563 VGND 0.037734
R7191 VGND.n1558 VGND 0.037734
R7192 VGND.n1553 VGND 0.037734
R7193 VGND.n1548 VGND 0.037734
R7194 VGND.n673 VGND 0.037734
R7195 VGND VGND.n671 0.037734
R7196 VGND VGND.n2407 0.037734
R7197 VGND.n2400 VGND 0.037734
R7198 VGND.n842 VGND 0.037734
R7199 VGND.n847 VGND 0.037734
R7200 VGND.n852 VGND 0.037734
R7201 VGND.n857 VGND 0.037734
R7202 VGND.n862 VGND 0.037734
R7203 VGND.n867 VGND 0.037734
R7204 VGND.n872 VGND 0.037734
R7205 VGND.n877 VGND 0.037734
R7206 VGND.n882 VGND 0.037734
R7207 VGND.n887 VGND 0.037734
R7208 VGND.n829 VGND 0.037734
R7209 VGND.n837 VGND 0.037734
R7210 VGND.n832 VGND 0.037734
R7211 VGND VGND.n825 0.037734
R7212 VGND VGND.n815 0.037734
R7213 VGND VGND.n1126 0.037734
R7214 VGND.n1129 VGND 0.037734
R7215 VGND VGND.n1136 0.037734
R7216 VGND.n1142 VGND 0.037734
R7217 VGND.n809 VGND 0.037734
R7218 VGND.n1161 VGND 0.037734
R7219 VGND VGND.n1168 0.037734
R7220 VGND.n1174 VGND 0.037734
R7221 VGND.n801 VGND 0.037734
R7222 VGND.n1193 VGND 0.037734
R7223 VGND VGND.n1200 0.037734
R7224 VGND.n1206 VGND 0.037734
R7225 VGND.n793 VGND 0.037734
R7226 VGND.n1225 VGND 0.037734
R7227 VGND VGND.n1232 0.037734
R7228 VGND.n718 VGND 0.037734
R7229 VGND.n777 VGND 0.037734
R7230 VGND.n772 VGND 0.037734
R7231 VGND.n767 VGND 0.037734
R7232 VGND.n762 VGND 0.037734
R7233 VGND.n757 VGND 0.037734
R7234 VGND.n752 VGND 0.037734
R7235 VGND.n747 VGND 0.037734
R7236 VGND.n742 VGND 0.037734
R7237 VGND.n737 VGND 0.037734
R7238 VGND.n732 VGND 0.037734
R7239 VGND.n727 VGND 0.037734
R7240 VGND.n722 VGND 0.037734
R7241 VGND VGND.n684 0.037734
R7242 VGND.n1287 VGND 0.037734
R7243 VGND VGND.n676 0.037734
R7244 VGND.n1112 VGND 0.0343542
R7245 VGND.n1084 VGND 0.0343542
R7246 VGND.n145 VGND 0.0343542
R7247 VGND.n613 VGND 0.0343542
R7248 VGND.n989 VGND 0.0343542
R7249 VGND.n1022 VGND 0.0343542
R7250 VGND.n1053 VGND 0.0343542
R7251 VGND.n175 VGND 0.0343542
R7252 VGND.n3007 VGND 0.0330521
R7253 VGND.n111 VGND 0.0330521
R7254 VGND.n2873 VGND 0.0330521
R7255 VGND.n2906 VGND 0.0330521
R7256 VGND VGND.n2913 0.0330521
R7257 VGND VGND.n2946 0.0330521
R7258 VGND VGND.n57 0.0330521
R7259 VGND VGND.n2986 0.0330521
R7260 VGND.n3006 VGND 0.024
R7261 VGND.n1 VGND 0.024
R7262 VGND.n144 VGND 0.0239375
R7263 VGND.n612 VGND 0.0239375
R7264 VGND.n174 VGND 0.0239375
R7265 VGND.n2905 VGND 0.0239375
R7266 VGND.n2914 VGND 0.0239375
R7267 VGND.n1089 VGND 0.0226354
R7268 VGND VGND.n119 0.0226354
R7269 VGND.n997 VGND 0.0226354
R7270 VGND.n988 VGND 0.0226354
R7271 VGND.n1028 VGND 0.0226354
R7272 VGND VGND.n2919 0.0226354
R7273 VGND.n2957 VGND 0.0226354
R7274 VGND.n2989 VGND 0.0226354
R7275 VGND VGND.n587 0.0213333
R7276 VGND.n993 VGND 0.0213333
R7277 VGND.n1059 VGND 0.0213333
R7278 VGND VGND.n108 0.0213333
R7279 VGND.n110 VGND 0.0213333
R7280 VGND VGND.n2868 0.0213333
R7281 VGND.n2872 VGND 0.0213333
R7282 VGND VGND.n2900 0.0213333
R7283 VGND.n82 VGND 0.0213333
R7284 VGND VGND.n2952 0.0213333
R7285 VGND.n3006 VGND 0.0161667
R7286 VGND.n2576 VGND 0.00980851
R7287 VGND.n3001 VGND 0.00980851
R7288 VGND.n2783 VGND 0.00980851
R7289 VGND VGND.n220 0.00980851
R7290 VGND VGND.n219 0.00980851
R7291 VGND VGND.n214 0.00980851
R7292 VGND VGND.n213 0.00980851
R7293 VGND VGND.n208 0.00980851
R7294 VGND VGND.n207 0.00980851
R7295 VGND VGND.n202 0.00980851
R7296 VGND VGND.n201 0.00980851
R7297 VGND VGND.n196 0.00980851
R7298 VGND VGND.n195 0.00980851
R7299 VGND VGND.n190 0.00980851
R7300 VGND VGND.n189 0.00980851
R7301 VGND.n2715 VGND 0.00980851
R7302 VGND.n235 VGND 0.00980851
R7303 VGND.n2491 VGND 0.00980851
R7304 VGND VGND.n258 0.00980851
R7305 VGND VGND.n257 0.00980851
R7306 VGND VGND.n256 0.00980851
R7307 VGND VGND.n255 0.00980851
R7308 VGND VGND.n254 0.00980851
R7309 VGND VGND.n253 0.00980851
R7310 VGND VGND.n252 0.00980851
R7311 VGND VGND.n251 0.00980851
R7312 VGND VGND.n250 0.00980851
R7313 VGND VGND.n249 0.00980851
R7314 VGND.n248 VGND 0.00980851
R7315 VGND VGND.n2505 0.00980851
R7316 VGND VGND.n186 0.00980851
R7317 VGND VGND.n185 0.00980851
R7318 VGND.n2517 VGND 0.00980851
R7319 VGND.n2430 VGND 0.00980851
R7320 VGND.n2294 VGND 0.00980851
R7321 VGND VGND.n329 0.00980851
R7322 VGND VGND.n328 0.00980851
R7323 VGND.n2276 VGND 0.00980851
R7324 VGND.n2253 VGND 0.00980851
R7325 VGND.n2245 VGND 0.00980851
R7326 VGND.n2227 VGND 0.00980851
R7327 VGND.n2219 VGND 0.00980851
R7328 VGND.n2201 VGND 0.00980851
R7329 VGND.n2193 VGND 0.00980851
R7330 VGND.n2175 VGND 0.00980851
R7331 VGND.n2167 VGND 0.00980851
R7332 VGND.n374 VGND 0.00980851
R7333 VGND VGND.n2828 0.00980851
R7334 VGND.n180 VGND 0.00980851
R7335 VGND.n2313 VGND 0.00980851
R7336 VGND VGND.n324 0.00980851
R7337 VGND.n2303 VGND 0.00980851
R7338 VGND VGND.n327 0.00980851
R7339 VGND.n2271 VGND 0.00980851
R7340 VGND.n2258 VGND 0.00980851
R7341 VGND.n2240 VGND 0.00980851
R7342 VGND.n2232 VGND 0.00980851
R7343 VGND.n2214 VGND 0.00980851
R7344 VGND.n2206 VGND 0.00980851
R7345 VGND.n2188 VGND 0.00980851
R7346 VGND.n2180 VGND 0.00980851
R7347 VGND.n2162 VGND 0.00980851
R7348 VGND.n2154 VGND 0.00980851
R7349 VGND.n1432 VGND 0.00980851
R7350 VGND.n1421 VGND 0.00980851
R7351 VGND VGND.n2127 0.00980851
R7352 VGND VGND.n322 0.00980851
R7353 VGND VGND.n321 0.00980851
R7354 VGND.n2139 VGND 0.00980851
R7355 VGND VGND.n390 0.00980851
R7356 VGND VGND.n389 0.00980851
R7357 VGND VGND.n388 0.00980851
R7358 VGND VGND.n387 0.00980851
R7359 VGND VGND.n386 0.00980851
R7360 VGND VGND.n385 0.00980851
R7361 VGND VGND.n384 0.00980851
R7362 VGND VGND.n383 0.00980851
R7363 VGND VGND.n382 0.00980851
R7364 VGND VGND.n381 0.00980851
R7365 VGND.n1496 VGND 0.00980851
R7366 VGND.n1438 VGND 0.00980851
R7367 VGND.n2122 VGND 0.00980851
R7368 VGND VGND.n399 0.00980851
R7369 VGND VGND.n319 0.00980851
R7370 VGND VGND.n318 0.00980851
R7371 VGND.n2102 VGND 0.00980851
R7372 VGND.n2079 VGND 0.00980851
R7373 VGND.n2071 VGND 0.00980851
R7374 VGND.n2053 VGND 0.00980851
R7375 VGND.n2045 VGND 0.00980851
R7376 VGND.n2027 VGND 0.00980851
R7377 VGND.n2019 VGND 0.00980851
R7378 VGND.n2001 VGND 0.00980851
R7379 VGND.n1993 VGND 0.00980851
R7380 VGND.n629 VGND 0.00980851
R7381 VGND VGND.n1501 0.00980851
R7382 VGND.n617 VGND 0.00980851
R7383 VGND.n2338 VGND 0.00980851
R7384 VGND VGND.n312 0.00980851
R7385 VGND.n2328 VGND 0.00980851
R7386 VGND VGND.n316 0.00980851
R7387 VGND.n2097 VGND 0.00980851
R7388 VGND.n2084 VGND 0.00980851
R7389 VGND.n2066 VGND 0.00980851
R7390 VGND.n2058 VGND 0.00980851
R7391 VGND.n2040 VGND 0.00980851
R7392 VGND.n2032 VGND 0.00980851
R7393 VGND.n2014 VGND 0.00980851
R7394 VGND.n2006 VGND 0.00980851
R7395 VGND.n1988 VGND 0.00980851
R7396 VGND.n1980 VGND 0.00980851
R7397 VGND.n655 VGND 0.00980851
R7398 VGND.n644 VGND 0.00980851
R7399 VGND VGND.n1953 0.00980851
R7400 VGND VGND.n310 0.00980851
R7401 VGND VGND.n309 0.00980851
R7402 VGND.n1965 VGND 0.00980851
R7403 VGND VGND.n446 0.00980851
R7404 VGND VGND.n445 0.00980851
R7405 VGND VGND.n444 0.00980851
R7406 VGND VGND.n443 0.00980851
R7407 VGND VGND.n442 0.00980851
R7408 VGND VGND.n441 0.00980851
R7409 VGND VGND.n440 0.00980851
R7410 VGND VGND.n439 0.00980851
R7411 VGND VGND.n438 0.00980851
R7412 VGND VGND.n437 0.00980851
R7413 VGND VGND.n661 0.00980851
R7414 VGND.n660 VGND 0.00980851
R7415 VGND.n1948 VGND 0.00980851
R7416 VGND VGND.n455 0.00980851
R7417 VGND VGND.n307 0.00980851
R7418 VGND VGND.n306 0.00980851
R7419 VGND.n1928 VGND 0.00980851
R7420 VGND.n1905 VGND 0.00980851
R7421 VGND.n1897 VGND 0.00980851
R7422 VGND.n1879 VGND 0.00980851
R7423 VGND.n1871 VGND 0.00980851
R7424 VGND.n1853 VGND 0.00980851
R7425 VGND.n1845 VGND 0.00980851
R7426 VGND.n1827 VGND 0.00980851
R7427 VGND.n1819 VGND 0.00980851
R7428 VGND.n1404 VGND 0.00980851
R7429 VGND VGND.n663 0.00980851
R7430 VGND.n1391 VGND 0.00980851
R7431 VGND.n2363 VGND 0.00980851
R7432 VGND VGND.n300 0.00980851
R7433 VGND.n2353 VGND 0.00980851
R7434 VGND VGND.n304 0.00980851
R7435 VGND.n1923 VGND 0.00980851
R7436 VGND.n1910 VGND 0.00980851
R7437 VGND.n1892 VGND 0.00980851
R7438 VGND.n1884 VGND 0.00980851
R7439 VGND.n1866 VGND 0.00980851
R7440 VGND.n1858 VGND 0.00980851
R7441 VGND.n1840 VGND 0.00980851
R7442 VGND.n1832 VGND 0.00980851
R7443 VGND.n1814 VGND 0.00980851
R7444 VGND.n1806 VGND 0.00980851
R7445 VGND.n1384 VGND 0.00980851
R7446 VGND.n1373 VGND 0.00980851
R7447 VGND VGND.n1779 0.00980851
R7448 VGND VGND.n298 0.00980851
R7449 VGND VGND.n297 0.00980851
R7450 VGND.n1791 VGND 0.00980851
R7451 VGND VGND.n502 0.00980851
R7452 VGND VGND.n501 0.00980851
R7453 VGND VGND.n500 0.00980851
R7454 VGND VGND.n499 0.00980851
R7455 VGND VGND.n498 0.00980851
R7456 VGND VGND.n497 0.00980851
R7457 VGND VGND.n496 0.00980851
R7458 VGND VGND.n495 0.00980851
R7459 VGND VGND.n494 0.00980851
R7460 VGND VGND.n493 0.00980851
R7461 VGND.n1366 VGND 0.00980851
R7462 VGND.n1305 VGND 0.00980851
R7463 VGND.n1774 VGND 0.00980851
R7464 VGND VGND.n511 0.00980851
R7465 VGND VGND.n295 0.00980851
R7466 VGND VGND.n294 0.00980851
R7467 VGND.n1754 VGND 0.00980851
R7468 VGND.n1731 VGND 0.00980851
R7469 VGND.n1723 VGND 0.00980851
R7470 VGND.n1705 VGND 0.00980851
R7471 VGND.n1697 VGND 0.00980851
R7472 VGND.n1679 VGND 0.00980851
R7473 VGND.n1671 VGND 0.00980851
R7474 VGND.n1653 VGND 0.00980851
R7475 VGND.n1645 VGND 0.00980851
R7476 VGND.n1526 VGND 0.00980851
R7477 VGND VGND.n574 0.00980851
R7478 VGND.n573 VGND 0.00980851
R7479 VGND.n2388 VGND 0.00980851
R7480 VGND VGND.n287 0.00980851
R7481 VGND.n2378 VGND 0.00980851
R7482 VGND VGND.n291 0.00980851
R7483 VGND.n1749 VGND 0.00980851
R7484 VGND.n1736 VGND 0.00980851
R7485 VGND.n1718 VGND 0.00980851
R7486 VGND.n1710 VGND 0.00980851
R7487 VGND.n1692 VGND 0.00980851
R7488 VGND.n1684 VGND 0.00980851
R7489 VGND.n1666 VGND 0.00980851
R7490 VGND.n1658 VGND 0.00980851
R7491 VGND.n1640 VGND 0.00980851
R7492 VGND.n1632 VGND 0.00980851
R7493 VGND.n1541 VGND 0.00980851
R7494 VGND.n1533 VGND 0.00980851
R7495 VGND VGND.n1605 0.00980851
R7496 VGND VGND.n283 0.00980851
R7497 VGND VGND.n282 0.00980851
R7498 VGND.n1617 VGND 0.00980851
R7499 VGND VGND.n558 0.00980851
R7500 VGND VGND.n557 0.00980851
R7501 VGND VGND.n556 0.00980851
R7502 VGND VGND.n555 0.00980851
R7503 VGND VGND.n554 0.00980851
R7504 VGND VGND.n553 0.00980851
R7505 VGND VGND.n552 0.00980851
R7506 VGND VGND.n551 0.00980851
R7507 VGND VGND.n550 0.00980851
R7508 VGND VGND.n549 0.00980851
R7509 VGND.n1546 VGND 0.00980851
R7510 VGND.n1298 VGND 0.00980851
R7511 VGND.n2408 VGND 0.00980851
R7512 VGND VGND.n279 0.00980851
R7513 VGND.n2398 VGND 0.00980851
R7514 VGND VGND.n713 0.00980851
R7515 VGND VGND.n712 0.00980851
R7516 VGND VGND.n707 0.00980851
R7517 VGND VGND.n706 0.00980851
R7518 VGND VGND.n701 0.00980851
R7519 VGND VGND.n700 0.00980851
R7520 VGND VGND.n695 0.00980851
R7521 VGND VGND.n694 0.00980851
R7522 VGND VGND.n689 0.00980851
R7523 VGND VGND.n688 0.00980851
R7524 VGND.n893 VGND 0.00980851
R7525 VGND VGND.n827 0.00980851
R7526 VGND.n826 VGND 0.00980851
R7527 VGND.n1122 VGND 0.00980851
R7528 VGND.n1127 VGND 0.00980851
R7529 VGND VGND.n812 0.00980851
R7530 VGND.n1140 VGND 0.00980851
R7531 VGND.n1148 VGND 0.00980851
R7532 VGND.n1159 VGND 0.00980851
R7533 VGND VGND.n804 0.00980851
R7534 VGND.n1172 VGND 0.00980851
R7535 VGND.n1180 VGND 0.00980851
R7536 VGND.n1191 VGND 0.00980851
R7537 VGND VGND.n796 0.00980851
R7538 VGND.n1204 VGND 0.00980851
R7539 VGND.n1212 VGND 0.00980851
R7540 VGND.n1223 VGND 0.00980851
R7541 VGND VGND.n788 0.00980851
R7542 VGND.n1233 VGND 0.00980851
R7543 VGND.n2413 VGND 0.00980851
R7544 VGND.n783 VGND 0.00980851
R7545 VGND VGND.n716 0.00980851
R7546 VGND VGND.n715 0.00980851
R7547 VGND VGND.n710 0.00980851
R7548 VGND VGND.n709 0.00980851
R7549 VGND VGND.n704 0.00980851
R7550 VGND VGND.n703 0.00980851
R7551 VGND VGND.n698 0.00980851
R7552 VGND VGND.n697 0.00980851
R7553 VGND VGND.n692 0.00980851
R7554 VGND VGND.n691 0.00980851
R7555 VGND VGND.n686 0.00980851
R7556 VGND.n685 VGND 0.00980851
R7557 VGND VGND.n1286 0.00980851
R7558 VGND.n677 VGND 0.00980851
R7559 VGND.n3023 VGND 0.00851991
R7560 VGND.n2654 VGND.n2652 0.00182979
R7561 VGND.n2651 VGND.n2650 0.00182979
R7562 VGND.n2662 VGND.n2660 0.00182979
R7563 VGND.n2647 VGND.n2646 0.00182979
R7564 VGND.n2670 VGND.n2668 0.00182979
R7565 VGND.n2643 VGND.n2642 0.00182979
R7566 VGND.n2678 VGND.n2676 0.00182979
R7567 VGND.n2639 VGND.n2638 0.00182979
R7568 VGND.n2686 VGND.n2684 0.00182979
R7569 VGND.n2635 VGND.n2634 0.00182979
R7570 VGND.n2694 VGND.n2692 0.00182979
R7571 VGND.n2631 VGND.n2630 0.00182979
R7572 VGND.n2702 VGND.n2700 0.00182979
R7573 VGND.n2627 VGND.n2581 0.00182979
R7574 VGND.n2708 VGND.n2572 0.00182979
R7575 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7576 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7577 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7578 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7579 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7580 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7581 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7582 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7583 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7584 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7585 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7586 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7587 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7588 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7589 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7590 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7591 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7592 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7593 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7594 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7595 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7596 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7597 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7598 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7599 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7600 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7601 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7602 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7603 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7604 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7605 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7606 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7607 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7608 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7609 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7610 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7611 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7612 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7613 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7614 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7615 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7616 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7617 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7618 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7619 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7620 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7621 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7622 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7623 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7624 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7625 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7626 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7627 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7628 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7629 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7630 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7631 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7632 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7633 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7634 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7635 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7636 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7637 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7638 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7639 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7640 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7641 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7642 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7643 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7644 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7645 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7646 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7647 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7648 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7649 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7650 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7651 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7652 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7653 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7654 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7655 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7656 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7657 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7658 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7659 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7660 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7661 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7662 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7663 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7664 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7665 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7666 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7667 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7668 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7669 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7670 XThR.Tn[2].n5 XThR.Tn[2].n3 135.249
R7671 XThR.Tn[2].n5 XThR.Tn[2].n4 98.982
R7672 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R7673 XThR.Tn[2].n9 XThR.Tn[2].n8 98.982
R7674 XThR.Tn[2].n7 XThR.Tn[2].n5 36.2672
R7675 XThR.Tn[2].n9 XThR.Tn[2].n7 36.2672
R7676 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7677 XThR.Tn[2].n1 XThR.Tn[2].t4 26.5955
R7678 XThR.Tn[2].n1 XThR.Tn[2].t7 26.5955
R7679 XThR.Tn[2].n0 XThR.Tn[2].t11 26.5955
R7680 XThR.Tn[2].n0 XThR.Tn[2].t10 26.5955
R7681 XThR.Tn[2].n3 XThR.Tn[2].t8 24.9236
R7682 XThR.Tn[2].n3 XThR.Tn[2].t1 24.9236
R7683 XThR.Tn[2].n4 XThR.Tn[2].t3 24.9236
R7684 XThR.Tn[2].n4 XThR.Tn[2].t2 24.9236
R7685 XThR.Tn[2].n6 XThR.Tn[2].t6 24.9236
R7686 XThR.Tn[2].n6 XThR.Tn[2].t9 24.9236
R7687 XThR.Tn[2].n8 XThR.Tn[2].t5 24.9236
R7688 XThR.Tn[2].n8 XThR.Tn[2].t0 24.9236
R7689 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7690 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7691 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7692 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7693 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7694 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7695 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7696 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7697 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7698 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7699 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7700 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7701 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7702 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7703 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7704 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7705 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7706 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7707 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7708 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7709 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7710 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7711 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7712 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7713 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7714 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7715 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7716 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7717 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7718 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7719 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7720 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7721 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7722 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7723 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7724 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7725 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7726 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7727 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7728 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7729 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7730 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7731 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7732 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7733 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7734 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7735 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7736 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7737 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7738 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7739 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7740 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7741 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7742 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7743 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7744 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7745 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7746 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7747 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7748 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7749 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7750 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7751 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7752 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7753 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7754 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7755 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7756 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7757 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7758 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7759 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7760 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7761 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7762 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7763 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7764 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7765 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7766 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7767 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7768 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7769 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7770 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7771 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7772 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7773 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7774 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7775 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7776 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7777 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7778 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7779 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7780 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7781 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7782 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7783 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7784 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7785 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7786 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7787 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7788 VPWR.n2837 VPWR.n2823 2618.82
R7789 VPWR.n2835 VPWR.n2829 2618.82
R7790 VPWR.n2853 VPWR.n2823 1916.47
R7791 VPWR.n2828 VPWR.n2827 1916.47
R7792 VPWR.n2827 VPWR.n2821 1916.47
R7793 VPWR.n2829 VPWR.n2822 1916.47
R7794 VPWR.n2852 VPWR.n2824 1912.94
R7795 VPWR.n2849 VPWR.n2843 1560
R7796 VPWR.n2850 VPWR.n2824 1408.24
R7797 VPWR.n2853 VPWR.n2852 1210.59
R7798 VPWR.n2851 VPWR.n2821 1210.59
R7799 VPWR.n2380 VPWR.t1560 1005.7
R7800 VPWR.t1778 VPWR.n485 1005.7
R7801 VPWR.t1627 VPWR.n2210 1005.7
R7802 VPWR.n639 VPWR.t1735 1005.7
R7803 VPWR.n2184 VPWR.t1461 1005.7
R7804 VPWR.t1568 VPWR.n677 1005.7
R7805 VPWR.t1528 VPWR.n2014 1005.7
R7806 VPWR.n831 VPWR.t1633 1005.7
R7807 VPWR.n1988 VPWR.t1453 1005.7
R7808 VPWR.t1640 VPWR.n869 1005.7
R7809 VPWR.n447 VPWR.t1445 1005.7
R7810 VPWR.t1748 VPWR.n1818 1005.7
R7811 VPWR.t1730 VPWR.n2406 1005.7
R7812 VPWR.n1023 VPWR.t1600 1005.7
R7813 VPWR.t1770 VPWR.n293 1005.7
R7814 VPWR.n1792 VPWR.t1711 1005.7
R7815 VPWR.n2591 VPWR.t1662 1005.7
R7816 VPWR.n1062 VPWR.t1546 1005.7
R7817 VPWR.t1146 VPWR.n2309 983.14
R7818 VPWR.n2310 VPWR.t218 983.14
R7819 VPWR.t778 VPWR.n2319 983.14
R7820 VPWR.n2320 VPWR.t1061 983.14
R7821 VPWR.t1388 VPWR.n2329 983.14
R7822 VPWR.n2330 VPWR.t792 983.14
R7823 VPWR.t352 VPWR.n2339 983.14
R7824 VPWR.n2340 VPWR.t285 983.14
R7825 VPWR.t135 VPWR.n2349 983.14
R7826 VPWR.n2350 VPWR.t896 983.14
R7827 VPWR.t1217 VPWR.n2359 983.14
R7828 VPWR.n2360 VPWR.t1193 983.14
R7829 VPWR.t1211 VPWR.n2369 983.14
R7830 VPWR.n2370 VPWR.t324 983.14
R7831 VPWR.t342 VPWR.n2379 983.14
R7832 VPWR.n542 VPWR.t175 983.14
R7833 VPWR.n541 VPWR.t503 983.14
R7834 VPWR.n537 VPWR.t754 983.14
R7835 VPWR.n533 VPWR.t606 983.14
R7836 VPWR.n529 VPWR.t167 983.14
R7837 VPWR.n525 VPWR.t273 983.14
R7838 VPWR.n521 VPWR.t290 983.14
R7839 VPWR.n517 VPWR.t465 983.14
R7840 VPWR.n513 VPWR.t511 983.14
R7841 VPWR.n509 VPWR.t1370 983.14
R7842 VPWR.n505 VPWR.t121 983.14
R7843 VPWR.n501 VPWR.t853 983.14
R7844 VPWR.n497 VPWR.t92 983.14
R7845 VPWR.n493 VPWR.t433 983.14
R7846 VPWR.n489 VPWR.t181 983.14
R7847 VPWR.n2281 VPWR.t1156 983.14
R7848 VPWR.n2280 VPWR.t226 983.14
R7849 VPWR.n2271 VPWR.t732 983.14
R7850 VPWR.n2270 VPWR.t1017 983.14
R7851 VPWR.n2261 VPWR.t1236 983.14
R7852 VPWR.n2260 VPWR.t241 983.14
R7853 VPWR.n2251 VPWR.t423 983.14
R7854 VPWR.n2250 VPWR.t583 983.14
R7855 VPWR.n2241 VPWR.t1276 983.14
R7856 VPWR.n2240 VPWR.t1303 983.14
R7857 VPWR.n2231 VPWR.t53 983.14
R7858 VPWR.n2230 VPWR.t1836 983.14
R7859 VPWR.n2221 VPWR.t69 983.14
R7860 VPWR.n2220 VPWR.t626 983.14
R7861 VPWR.n2211 VPWR.t528 983.14
R7862 VPWR.t159 VPWR.n582 983.14
R7863 VPWR.t485 VPWR.n586 983.14
R7864 VPWR.t746 VPWR.n590 983.14
R7865 VPWR.t1168 VPWR.n594 983.14
R7866 VPWR.t612 VPWR.n598 983.14
R7867 VPWR.t261 VPWR.n602 983.14
R7868 VPWR.t300 VPWR.n606 983.14
R7869 VPWR.t473 VPWR.n610 983.14
R7870 VPWR.t565 VPWR.n614 983.14
R7871 VPWR.t1376 VPWR.n618 983.14
R7872 VPWR.t131 VPWR.n622 983.14
R7873 VPWR.t1100 VPWR.n626 983.14
R7874 VPWR.t100 VPWR.n630 983.14
R7875 VPWR.t409 VPWR.n634 983.14
R7876 VPWR.t187 VPWR.n638 983.14
R7877 VPWR.t145 VPWR.n2113 983.14
R7878 VPWR.n2114 VPWR.t679 983.14
R7879 VPWR.t766 VPWR.n2123 983.14
R7880 VPWR.n2124 VPWR.t1824 983.14
R7881 VPWR.t1227 VPWR.n2133 983.14
R7882 VPWR.n2134 VPWR.t231 983.14
R7883 VPWR.t1889 VPWR.n2143 983.14
R7884 VPWR.n2144 VPWR.t937 983.14
R7885 VPWR.t370 VPWR.n2153 983.14
R7886 VPWR.n2154 VPWR.t541 983.14
R7887 VPWR.t443 VPWR.n2163 983.14
R7888 VPWR.n2164 VPWR.t955 983.14
R7889 VPWR.t1870 VPWR.n2173 983.14
R7890 VPWR.n2174 VPWR.t1116 983.14
R7891 VPWR.t314 VPWR.n2183 983.14
R7892 VPWR.n734 VPWR.t1144 983.14
R7893 VPWR.n733 VPWR.t216 983.14
R7894 VPWR.n729 VPWR.t780 983.14
R7895 VPWR.n725 VPWR.t1059 983.14
R7896 VPWR.n721 VPWR.t1386 983.14
R7897 VPWR.n717 VPWR.t790 983.14
R7898 VPWR.n713 VPWR.t350 983.14
R7899 VPWR.n709 VPWR.t283 983.14
R7900 VPWR.n705 VPWR.t695 983.14
R7901 VPWR.n701 VPWR.t894 983.14
R7902 VPWR.n697 VPWR.t1322 983.14
R7903 VPWR.n693 VPWR.t1191 983.14
R7904 VPWR.n689 VPWR.t1209 983.14
R7905 VPWR.n685 VPWR.t8 983.14
R7906 VPWR.n681 VPWR.t340 983.14
R7907 VPWR.n2085 VPWR.t827 983.14
R7908 VPWR.n2084 VPWR.t1289 983.14
R7909 VPWR.n2075 VPWR.t774 983.14
R7910 VPWR.n2074 VPWR.t1814 983.14
R7911 VPWR.n2065 VPWR.t1223 983.14
R7912 VPWR.n2064 VPWR.t798 983.14
R7913 VPWR.n2055 VPWR.t358 983.14
R7914 VPWR.n2054 VPWR.t986 983.14
R7915 VPWR.n2045 VPWR.t141 983.14
R7916 VPWR.n2044 VPWR.t902 983.14
R7917 VPWR.n2035 VPWR.t1114 983.14
R7918 VPWR.n2034 VPWR.t1183 983.14
R7919 VPWR.n2025 VPWR.t1213 983.14
R7920 VPWR.n2024 VPWR.t664 983.14
R7921 VPWR.n2015 VPWR.t344 983.14
R7922 VPWR.t458 VPWR.n774 983.14
R7923 VPWR.t224 VPWR.n778 983.14
R7924 VPWR.t734 VPWR.n782 983.14
R7925 VPWR.t1013 VPWR.n786 983.14
R7926 VPWR.t1234 VPWR.n790 983.14
R7927 VPWR.t239 VPWR.n794 983.14
R7928 VPWR.t421 VPWR.n798 983.14
R7929 VPWR.t579 VPWR.n802 983.14
R7930 VPWR.t1274 VPWR.n806 983.14
R7931 VPWR.t1301 VPWR.n810 983.14
R7932 VPWR.t51 VPWR.n814 983.14
R7933 VPWR.t1834 VPWR.n818 983.14
R7934 VPWR.t65 VPWR.n822 983.14
R7935 VPWR.t624 VPWR.n826 983.14
R7936 VPWR.t524 VPWR.n830 983.14
R7937 VPWR.t147 VPWR.n1917 983.14
R7938 VPWR.n1918 VPWR.t681 983.14
R7939 VPWR.t764 VPWR.n1927 983.14
R7940 VPWR.n1928 VPWR.t1021 983.14
R7941 VPWR.t916 VPWR.n1937 983.14
R7942 VPWR.n1938 VPWR.t233 983.14
R7943 VPWR.t1891 VPWR.n1947 983.14
R7944 VPWR.n1948 VPWR.t939 983.14
R7945 VPWR.t493 VPWR.n1957 983.14
R7946 VPWR.n1958 VPWR.t543 983.14
R7947 VPWR.t445 VPWR.n1967 983.14
R7948 VPWR.n1968 VPWR.t857 983.14
R7949 VPWR.t1872 VPWR.n1977 983.14
R7950 VPWR.n1978 VPWR.t1118 983.14
R7951 VPWR.t316 VPWR.n1987 983.14
R7952 VPWR.n926 VPWR.t456 983.14
R7953 VPWR.n925 VPWR.t222 983.14
R7954 VPWR.n921 VPWR.t736 983.14
R7955 VPWR.n917 VPWR.t1011 983.14
R7956 VPWR.n913 VPWR.t1232 983.14
R7957 VPWR.n909 VPWR.t237 983.14
R7958 VPWR.n905 VPWR.t419 983.14
R7959 VPWR.n901 VPWR.t575 983.14
R7960 VPWR.n897 VPWR.t1272 983.14
R7961 VPWR.n893 VPWR.t1299 983.14
R7962 VPWR.n889 VPWR.t49 983.14
R7963 VPWR.n885 VPWR.t1832 983.14
R7964 VPWR.n881 VPWR.t61 983.14
R7965 VPWR.n877 VPWR.t622 983.14
R7966 VPWR.n873 VPWR.t522 983.14
R7967 VPWR.t149 VPWR.n390 983.14
R7968 VPWR.t683 VPWR.n394 983.14
R7969 VPWR.t762 VPWR.n398 983.14
R7970 VPWR.t1025 VPWR.n402 983.14
R7971 VPWR.t918 VPWR.n406 983.14
R7972 VPWR.t235 VPWR.n410 983.14
R7973 VPWR.t1893 VPWR.n414 983.14
R7974 VPWR.t941 VPWR.n418 983.14
R7975 VPWR.t495 VPWR.n422 983.14
R7976 VPWR.t545 VPWR.n426 983.14
R7977 VPWR.t447 VPWR.n430 983.14
R7978 VPWR.t859 VPWR.n434 983.14
R7979 VPWR.t1874 VPWR.n438 983.14
R7980 VPWR.t1120 VPWR.n442 983.14
R7981 VPWR.t320 VPWR.n446 983.14
R7982 VPWR.n1889 VPWR.t157 983.14
R7983 VPWR.n1888 VPWR.t509 983.14
R7984 VPWR.n1879 VPWR.t748 983.14
R7985 VPWR.n1878 VPWR.t1166 983.14
R7986 VPWR.n1869 VPWR.t173 983.14
R7987 VPWR.n1868 VPWR.t257 983.14
R7988 VPWR.n1859 VPWR.t296 983.14
R7989 VPWR.n1858 VPWR.t471 983.14
R7990 VPWR.n1849 VPWR.t641 983.14
R7991 VPWR.n1848 VPWR.t1374 983.14
R7992 VPWR.n1839 VPWR.t127 983.14
R7993 VPWR.n1838 VPWR.t1098 983.14
R7994 VPWR.n1829 VPWR.t98 983.14
R7995 VPWR.n1828 VPWR.t407 983.14
R7996 VPWR.n1819 VPWR.t185 983.14
R7997 VPWR.n2477 VPWR.t161 983.14
R7998 VPWR.n2476 VPWR.t487 983.14
R7999 VPWR.n2467 VPWR.t744 983.14
R8000 VPWR.n2466 VPWR.t1172 983.14
R8001 VPWR.n2457 VPWR.t614 983.14
R8002 VPWR.n2456 VPWR.t263 983.14
R8003 VPWR.n2447 VPWR.t302 983.14
R8004 VPWR.n2446 VPWR.t837 983.14
R8005 VPWR.n2437 VPWR.t567 983.14
R8006 VPWR.n2436 VPWR.t1378 983.14
R8007 VPWR.n2427 VPWR.t133 983.14
R8008 VPWR.n2426 VPWR.t1102 983.14
R8009 VPWR.n2417 VPWR.t102 983.14
R8010 VPWR.n2416 VPWR.t411 983.14
R8011 VPWR.n2407 VPWR.t191 983.14
R8012 VPWR.t1158 VPWR.n966 983.14
R8013 VPWR.t1258 VPWR.n970 983.14
R8014 VPWR.t726 VPWR.n974 983.14
R8015 VPWR.t1055 VPWR.n978 983.14
R8016 VPWR.t477 VPWR.n982 983.14
R8017 VPWR.t247 VPWR.n986 983.14
R8018 VPWR.t429 VPWR.n990 983.14
R8019 VPWR.t587 VPWR.n994 983.14
R8020 VPWR.t689 VPWR.n998 983.14
R8021 VPWR.t1305 VPWR.n1002 983.14
R8022 VPWR.t1316 VPWR.n1006 983.14
R8023 VPWR.t1838 VPWR.n1010 983.14
R8024 VPWR.t1201 VPWR.n1014 983.14
R8025 VPWR.t0 VPWR.n1018 983.14
R8026 VPWR.t336 VPWR.n1022 983.14
R8027 VPWR.n350 VPWR.t177 983.14
R8028 VPWR.n349 VPWR.t505 983.14
R8029 VPWR.n345 VPWR.t752 983.14
R8030 VPWR.n341 VPWR.t608 983.14
R8031 VPWR.n337 VPWR.t169 983.14
R8032 VPWR.n333 VPWR.t253 983.14
R8033 VPWR.n329 VPWR.t292 983.14
R8034 VPWR.n325 VPWR.t469 983.14
R8035 VPWR.n321 VPWR.t637 983.14
R8036 VPWR.n317 VPWR.t1372 983.14
R8037 VPWR.n313 VPWR.t123 983.14
R8038 VPWR.n309 VPWR.t855 983.14
R8039 VPWR.n305 VPWR.t96 983.14
R8040 VPWR.n301 VPWR.t435 983.14
R8041 VPWR.n297 VPWR.t183 983.14
R8042 VPWR.t1681 VPWR.n1468 983.14
R8043 VPWR.t1783 VPWR.n1475 983.14
R8044 VPWR.t1554 VPWR.n1481 983.14
R8045 VPWR.t1656 VPWR.n1492 983.14
R8046 VPWR.n1493 VPWR.t1678 983.14
R8047 VPWR.t1429 VPWR.n1506 983.14
R8048 VPWR.n1507 VPWR.t1551 983.14
R8049 VPWR.t1692 VPWR.n1520 983.14
R8050 VPWR.n1521 VPWR.t1708 983.14
R8051 VPWR.n1536 VPWR.t1448 983.14
R8052 VPWR.n1535 VPWR.t1581 983.14
R8053 VPWR.n1761 VPWR.t1622 983.14
R8054 VPWR.n1760 VPWR.t1458 983.14
R8055 VPWR.n1749 VPWR.t1495 983.14
R8056 VPWR.t1603 VPWR.n1791 983.14
R8057 VPWR.t1609 VPWR.n2506 983.14
R8058 VPWR.n2507 VPWR.t1721 983.14
R8059 VPWR.t1486 VPWR.n2518 983.14
R8060 VPWR.n2519 VPWR.t1594 983.14
R8061 VPWR.t1606 VPWR.n2530 983.14
R8062 VPWR.n2531 VPWR.t1762 983.14
R8063 VPWR.t1483 VPWR.n2542 983.14
R8064 VPWR.n2543 VPWR.t1643 983.14
R8065 VPWR.t1659 VPWR.n2554 983.14
R8066 VPWR.n2555 VPWR.t1789 983.14
R8067 VPWR.t1533 VPWR.n2566 983.14
R8068 VPWR.n2567 VPWR.t1563 983.14
R8069 VPWR.t1413 VPWR.n2578 983.14
R8070 VPWR.n2579 VPWR.t1432 983.14
R8071 VPWR.t1557 VPWR.n2590 983.14
R8072 VPWR.n1594 VPWR.t1492 983.14
R8073 VPWR.n1593 VPWR.t1597 983.14
R8074 VPWR.t1759 VPWR.n1182 983.14
R8075 VPWR.t1477 VPWR.n1185 983.14
R8076 VPWR.n1220 VPWR.t1489 983.14
R8077 VPWR.n1219 VPWR.t1648 983.14
R8078 VPWR.n1216 VPWR.t1756 983.14
R8079 VPWR.n1213 VPWR.t1517 983.14
R8080 VPWR.n1205 VPWR.t1543 983.14
R8081 VPWR.n1202 VPWR.t1670 983.14
R8082 VPWR.n1199 VPWR.t1416 983.14
R8083 VPWR.n1191 VPWR.t1437 983.14
R8084 VPWR.n1188 VPWR.t1675 983.14
R8085 VPWR.n1740 VPWR.t1703 983.14
R8086 VPWR.n1739 VPWR.t1423 983.14
R8087 VPWR.n1308 VPWR.t1242 877.144
R8088 VPWR.n2723 VPWR.t921 877.144
R8089 VPWR.n2843 VPWR.n2822 857.648
R8090 VPWR.n1122 VPWR.t1725 738.074
R8091 VPWR.n99 VPWR.t1465 738.074
R8092 VPWR.n290 VPWR.t1083 738.074
R8093 VPWR.n68 VPWR.t1534 738.074
R8094 VPWR.n346 VPWR.t178 738.074
R8095 VPWR.n98 VPWR.t1610 738.074
R8096 VPWR.n963 VPWR.t1068 738.074
R8097 VPWR.n356 VPWR.t1076 738.074
R8098 VPWR.n357 VPWR.t162 738.074
R8099 VPWR.n318 VPWR.t470 738.074
R8100 VPWR.n75 VPWR.t1644 738.074
R8101 VPWR.n971 VPWR.t1259 738.074
R8102 VPWR.n369 VPWR.t303 738.074
R8103 VPWR.n322 VPWR.t293 738.074
R8104 VPWR.n80 VPWR.t1484 738.074
R8105 VPWR.n932 VPWR.t1080 738.074
R8106 VPWR.n933 VPWR.t158 738.074
R8107 VPWR.n936 VPWR.t510 738.074
R8108 VPWR.n387 VPWR.t1087 738.074
R8109 VPWR.n391 VPWR.t150 738.074
R8110 VPWR.n395 VPWR.t684 738.074
R8111 VPWR.n365 VPWR.t615 738.074
R8112 VPWR.n330 VPWR.t170 738.074
R8113 VPWR.n86 VPWR.t1607 738.074
R8114 VPWR.n937 VPWR.t749 738.074
R8115 VPWR.n403 VPWR.t1026 738.074
R8116 VPWR.n364 VPWR.t1173 738.074
R8117 VPWR.n334 VPWR.t609 738.074
R8118 VPWR.n87 VPWR.t1595 738.074
R8119 VPWR.n481 VPWR.t1095 738.074
R8120 VPWR.n480 VPWR.t1147 738.074
R8121 VPWR.n477 VPWR.t219 738.074
R8122 VPWR.n476 VPWR.t779 738.074
R8123 VPWR.n472 VPWR.t1389 738.074
R8124 VPWR.n469 VPWR.t793 738.074
R8125 VPWR.n468 VPWR.t353 738.074
R8126 VPWR.n465 VPWR.t286 738.074
R8127 VPWR.n464 VPWR.t136 738.074
R8128 VPWR.n461 VPWR.t897 738.074
R8129 VPWR.n460 VPWR.t1218 738.074
R8130 VPWR.n457 VPWR.t1194 738.074
R8131 VPWR.n456 VPWR.t1212 738.074
R8132 VPWR.n453 VPWR.t325 738.074
R8133 VPWR.n452 VPWR.t343 738.074
R8134 VPWR.n473 VPWR.t1062 738.074
R8135 VPWR.n482 VPWR.t1085 738.074
R8136 VPWR.n538 VPWR.t176 738.074
R8137 VPWR.n534 VPWR.t504 738.074
R8138 VPWR.n530 VPWR.t755 738.074
R8139 VPWR.n522 VPWR.t168 738.074
R8140 VPWR.n518 VPWR.t274 738.074
R8141 VPWR.n514 VPWR.t291 738.074
R8142 VPWR.n510 VPWR.t466 738.074
R8143 VPWR.n506 VPWR.t512 738.074
R8144 VPWR.n502 VPWR.t1371 738.074
R8145 VPWR.n498 VPWR.t122 738.074
R8146 VPWR.n494 VPWR.t854 738.074
R8147 VPWR.n490 VPWR.t93 738.074
R8148 VPWR.n486 VPWR.t434 738.074
R8149 VPWR.n483 VPWR.t182 738.074
R8150 VPWR.n526 VPWR.t607 738.074
R8151 VPWR.n548 VPWR.t1070 738.074
R8152 VPWR.n549 VPWR.t1157 738.074
R8153 VPWR.n552 VPWR.t227 738.074
R8154 VPWR.n553 VPWR.t733 738.074
R8155 VPWR.n557 VPWR.t1237 738.074
R8156 VPWR.n560 VPWR.t242 738.074
R8157 VPWR.n561 VPWR.t424 738.074
R8158 VPWR.n564 VPWR.t584 738.074
R8159 VPWR.n565 VPWR.t1277 738.074
R8160 VPWR.n568 VPWR.t1304 738.074
R8161 VPWR.n569 VPWR.t54 738.074
R8162 VPWR.n572 VPWR.t1837 738.074
R8163 VPWR.n573 VPWR.t70 738.074
R8164 VPWR.n576 VPWR.t627 738.074
R8165 VPWR.n577 VPWR.t529 738.074
R8166 VPWR.n556 VPWR.t1018 738.074
R8167 VPWR.n579 VPWR.t1078 738.074
R8168 VPWR.n583 VPWR.t160 738.074
R8169 VPWR.n587 VPWR.t486 738.074
R8170 VPWR.n591 VPWR.t747 738.074
R8171 VPWR.n599 VPWR.t613 738.074
R8172 VPWR.n603 VPWR.t262 738.074
R8173 VPWR.n607 VPWR.t301 738.074
R8174 VPWR.n611 VPWR.t474 738.074
R8175 VPWR.n615 VPWR.t566 738.074
R8176 VPWR.n619 VPWR.t1377 738.074
R8177 VPWR.n623 VPWR.t132 738.074
R8178 VPWR.n627 VPWR.t1101 738.074
R8179 VPWR.n631 VPWR.t101 738.074
R8180 VPWR.n635 VPWR.t410 738.074
R8181 VPWR.n578 VPWR.t188 738.074
R8182 VPWR.n595 VPWR.t1169 738.074
R8183 VPWR.n673 VPWR.t1091 738.074
R8184 VPWR.n672 VPWR.t146 738.074
R8185 VPWR.n669 VPWR.t680 738.074
R8186 VPWR.n668 VPWR.t767 738.074
R8187 VPWR.n664 VPWR.t1228 738.074
R8188 VPWR.n661 VPWR.t232 738.074
R8189 VPWR.n660 VPWR.t1890 738.074
R8190 VPWR.n657 VPWR.t938 738.074
R8191 VPWR.n656 VPWR.t371 738.074
R8192 VPWR.n653 VPWR.t542 738.074
R8193 VPWR.n652 VPWR.t444 738.074
R8194 VPWR.n649 VPWR.t956 738.074
R8195 VPWR.n648 VPWR.t1871 738.074
R8196 VPWR.n645 VPWR.t1117 738.074
R8197 VPWR.n644 VPWR.t315 738.074
R8198 VPWR.n665 VPWR.t1825 738.074
R8199 VPWR.n674 VPWR.t1097 738.074
R8200 VPWR.n730 VPWR.t1145 738.074
R8201 VPWR.n726 VPWR.t217 738.074
R8202 VPWR.n722 VPWR.t781 738.074
R8203 VPWR.n714 VPWR.t1387 738.074
R8204 VPWR.n710 VPWR.t791 738.074
R8205 VPWR.n706 VPWR.t351 738.074
R8206 VPWR.n702 VPWR.t284 738.074
R8207 VPWR.n698 VPWR.t696 738.074
R8208 VPWR.n694 VPWR.t895 738.074
R8209 VPWR.n690 VPWR.t1323 738.074
R8210 VPWR.n686 VPWR.t1192 738.074
R8211 VPWR.n682 VPWR.t1210 738.074
R8212 VPWR.n678 VPWR.t9 738.074
R8213 VPWR.n675 VPWR.t341 738.074
R8214 VPWR.n718 VPWR.t1060 738.074
R8215 VPWR.n740 VPWR.t1093 738.074
R8216 VPWR.n741 VPWR.t828 738.074
R8217 VPWR.n744 VPWR.t1290 738.074
R8218 VPWR.n745 VPWR.t775 738.074
R8219 VPWR.n749 VPWR.t1224 738.074
R8220 VPWR.n752 VPWR.t799 738.074
R8221 VPWR.n753 VPWR.t359 738.074
R8222 VPWR.n756 VPWR.t987 738.074
R8223 VPWR.n757 VPWR.t142 738.074
R8224 VPWR.n760 VPWR.t903 738.074
R8225 VPWR.n761 VPWR.t1115 738.074
R8226 VPWR.n764 VPWR.t1184 738.074
R8227 VPWR.n765 VPWR.t1214 738.074
R8228 VPWR.n768 VPWR.t665 738.074
R8229 VPWR.n769 VPWR.t345 738.074
R8230 VPWR.n748 VPWR.t1815 738.074
R8231 VPWR.n771 VPWR.t1072 738.074
R8232 VPWR.n775 VPWR.t459 738.074
R8233 VPWR.n779 VPWR.t225 738.074
R8234 VPWR.n783 VPWR.t735 738.074
R8235 VPWR.n791 VPWR.t1235 738.074
R8236 VPWR.n795 VPWR.t240 738.074
R8237 VPWR.n799 VPWR.t422 738.074
R8238 VPWR.n803 VPWR.t580 738.074
R8239 VPWR.n807 VPWR.t1275 738.074
R8240 VPWR.n811 VPWR.t1302 738.074
R8241 VPWR.n815 VPWR.t52 738.074
R8242 VPWR.n819 VPWR.t1835 738.074
R8243 VPWR.n823 VPWR.t66 738.074
R8244 VPWR.n827 VPWR.t625 738.074
R8245 VPWR.n770 VPWR.t525 738.074
R8246 VPWR.n787 VPWR.t1014 738.074
R8247 VPWR.n865 VPWR.t1089 738.074
R8248 VPWR.n864 VPWR.t148 738.074
R8249 VPWR.n861 VPWR.t682 738.074
R8250 VPWR.n860 VPWR.t765 738.074
R8251 VPWR.n856 VPWR.t917 738.074
R8252 VPWR.n853 VPWR.t234 738.074
R8253 VPWR.n852 VPWR.t1892 738.074
R8254 VPWR.n849 VPWR.t940 738.074
R8255 VPWR.n848 VPWR.t494 738.074
R8256 VPWR.n845 VPWR.t544 738.074
R8257 VPWR.n844 VPWR.t446 738.074
R8258 VPWR.n841 VPWR.t858 738.074
R8259 VPWR.n840 VPWR.t1873 738.074
R8260 VPWR.n837 VPWR.t1119 738.074
R8261 VPWR.n836 VPWR.t317 738.074
R8262 VPWR.n857 VPWR.t1022 738.074
R8263 VPWR.n866 VPWR.t1074 738.074
R8264 VPWR.n922 VPWR.t457 738.074
R8265 VPWR.n918 VPWR.t223 738.074
R8266 VPWR.n914 VPWR.t737 738.074
R8267 VPWR.n906 VPWR.t1233 738.074
R8268 VPWR.n902 VPWR.t238 738.074
R8269 VPWR.n898 VPWR.t420 738.074
R8270 VPWR.n894 VPWR.t576 738.074
R8271 VPWR.n890 VPWR.t1273 738.074
R8272 VPWR.n886 VPWR.t1300 738.074
R8273 VPWR.n882 VPWR.t50 738.074
R8274 VPWR.n878 VPWR.t1833 738.074
R8275 VPWR.n874 VPWR.t62 738.074
R8276 VPWR.n870 VPWR.t623 738.074
R8277 VPWR.n867 VPWR.t523 738.074
R8278 VPWR.n910 VPWR.t1012 738.074
R8279 VPWR.n940 VPWR.t1167 738.074
R8280 VPWR.n979 VPWR.t1056 738.074
R8281 VPWR.n1179 VPWR.t1478 738.074
R8282 VPWR.n399 VPWR.t763 738.074
R8283 VPWR.n361 VPWR.t745 738.074
R8284 VPWR.n338 VPWR.t753 738.074
R8285 VPWR.n92 VPWR.t1487 738.074
R8286 VPWR.n975 VPWR.t727 738.074
R8287 VPWR.n1183 VPWR.t1760 738.074
R8288 VPWR.n941 VPWR.t174 738.074
R8289 VPWR.n983 VPWR.t478 738.074
R8290 VPWR.n1217 VPWR.t1490 738.074
R8291 VPWR.n407 VPWR.t919 738.074
R8292 VPWR.n415 VPWR.t1894 738.074
R8293 VPWR.n419 VPWR.t942 738.074
R8294 VPWR.n423 VPWR.t496 738.074
R8295 VPWR.n427 VPWR.t546 738.074
R8296 VPWR.n431 VPWR.t448 738.074
R8297 VPWR.n435 VPWR.t860 738.074
R8298 VPWR.n439 VPWR.t1875 738.074
R8299 VPWR.n443 VPWR.t1121 738.074
R8300 VPWR.n386 VPWR.t321 738.074
R8301 VPWR.n411 VPWR.t236 738.074
R8302 VPWR.n368 VPWR.t264 738.074
R8303 VPWR.n326 VPWR.t254 738.074
R8304 VPWR.n81 VPWR.t1763 738.074
R8305 VPWR.n987 VPWR.t248 738.074
R8306 VPWR.n1214 VPWR.t1649 738.074
R8307 VPWR.n944 VPWR.t258 738.074
R8308 VPWR.n948 VPWR.t472 738.074
R8309 VPWR.n949 VPWR.t642 738.074
R8310 VPWR.n952 VPWR.t1375 738.074
R8311 VPWR.n953 VPWR.t128 738.074
R8312 VPWR.n956 VPWR.t1099 738.074
R8313 VPWR.n957 VPWR.t99 738.074
R8314 VPWR.n960 VPWR.t408 738.074
R8315 VPWR.n961 VPWR.t186 738.074
R8316 VPWR.n945 VPWR.t297 738.074
R8317 VPWR.n991 VPWR.t430 738.074
R8318 VPWR.n1206 VPWR.t1757 738.074
R8319 VPWR.n360 VPWR.t488 738.074
R8320 VPWR.n342 VPWR.t506 738.074
R8321 VPWR.n93 VPWR.t1722 738.074
R8322 VPWR.n1180 VPWR.t1598 738.074
R8323 VPWR.n995 VPWR.t588 738.074
R8324 VPWR.n1203 VPWR.t1518 738.074
R8325 VPWR.n372 VPWR.t838 738.074
R8326 VPWR.n376 VPWR.t1379 738.074
R8327 VPWR.n377 VPWR.t134 738.074
R8328 VPWR.n380 VPWR.t1103 738.074
R8329 VPWR.n381 VPWR.t103 738.074
R8330 VPWR.n384 VPWR.t412 738.074
R8331 VPWR.n385 VPWR.t192 738.074
R8332 VPWR.n373 VPWR.t568 738.074
R8333 VPWR.n314 VPWR.t638 738.074
R8334 VPWR.n74 VPWR.t1660 738.074
R8335 VPWR.n1200 VPWR.t1544 738.074
R8336 VPWR.n999 VPWR.t690 738.074
R8337 VPWR.n1003 VPWR.t1306 738.074
R8338 VPWR.n1007 VPWR.t1317 738.074
R8339 VPWR.n1011 VPWR.t1839 738.074
R8340 VPWR.n1015 VPWR.t1202 738.074
R8341 VPWR.n1019 VPWR.t1 738.074
R8342 VPWR.n962 VPWR.t337 738.074
R8343 VPWR.n967 VPWR.t1159 738.074
R8344 VPWR.n1123 VPWR.t1493 738.074
R8345 VPWR.n310 VPWR.t1373 738.074
R8346 VPWR.n69 VPWR.t1790 738.074
R8347 VPWR.n1192 VPWR.t1671 738.074
R8348 VPWR.n1189 VPWR.t1417 738.074
R8349 VPWR.n306 VPWR.t124 738.074
R8350 VPWR.n302 VPWR.t856 738.074
R8351 VPWR.n294 VPWR.t436 738.074
R8352 VPWR.n291 VPWR.t184 738.074
R8353 VPWR.n298 VPWR.t97 738.074
R8354 VPWR.n1058 VPWR.t1676 738.074
R8355 VPWR.n1186 VPWR.t1438 738.074
R8356 VPWR.n63 VPWR.t1564 738.074
R8357 VPWR.n62 VPWR.t1414 738.074
R8358 VPWR.n57 VPWR.t1433 738.074
R8359 VPWR.n56 VPWR.t1558 738.074
R8360 VPWR.n1059 VPWR.t1704 738.074
R8361 VPWR.n1061 VPWR.t1424 738.074
R8362 VPWR.n2856 VPWR.n2821 702.354
R8363 VPWR.n2856 VPWR.n2822 702.354
R8364 VPWR.n2854 VPWR.n2853 702.354
R8365 VPWR.n2854 VPWR.n2821 702.354
R8366 VPWR.n2837 VPWR.n2828 702.354
R8367 VPWR.n2850 VPWR.n2849 702.354
R8368 VPWR.n2835 VPWR.n2828 702.354
R8369 VPWR.n2815 VPWR.t517 651.634
R8370 VPWR.n2831 VPWR.t1081 651.505
R8371 VPWR.n2825 VPWR.t719 651.505
R8372 VPWR.n2862 VPWR.t1801 651.431
R8373 VPWR.n1061 VPWR.t1547 646.071
R8374 VPWR.n1122 VPWR.t1443 646.071
R8375 VPWR.n1059 VPWR.t1696 646.071
R8376 VPWR.n56 VPWR.t1663 646.071
R8377 VPWR.n62 VPWR.t1787 646.071
R8378 VPWR.n99 VPWR.t1572 646.071
R8379 VPWR.n1053 VPWR.t1208 646.071
R8380 VPWR.n1231 VPWR.t455 646.071
R8381 VPWR.n298 VPWR.t1123 646.071
R8382 VPWR.n290 VPWR.t166 646.071
R8383 VPWR.n306 VPWR.t1847 646.071
R8384 VPWR.n68 VPWR.t1526 646.071
R8385 VPWR.n1153 VPWR.t1364 646.071
R8386 VPWR.n346 VPWR.t484 646.071
R8387 VPWR.n98 VPWR.t1701 646.071
R8388 VPWR.n967 VPWR.t1263 646.071
R8389 VPWR.n963 VPWR.t1149 646.071
R8390 VPWR.n999 VPWR.t899 646.071
R8391 VPWR.n373 VPWR.t1913 646.071
R8392 VPWR.n356 VPWR.t1004 646.071
R8393 VPWR.n357 VPWR.t58 646.071
R8394 VPWR.n372 VPWR.t574 646.071
R8395 VPWR.n318 VPWR.t644 646.071
R8396 VPWR.n75 VPWR.t1631 646.071
R8397 VPWR.n971 VPWR.t761 646.071
R8398 VPWR.n369 VPWR.t592 646.071
R8399 VPWR.n322 VPWR.t582 646.071
R8400 VPWR.n80 VPWR.t1503 646.071
R8401 VPWR.n945 VPWR.t586 646.071
R8402 VPWR.n932 VPWR.t1000 646.071
R8403 VPWR.n933 VPWR.t490 646.071
R8404 VPWR.n936 VPWR.t725 646.071
R8405 VPWR.n944 VPWR.t305 646.071
R8406 VPWR.n411 VPWR.t1900 646.071
R8407 VPWR.n387 VPWR.t600 646.071
R8408 VPWR.n391 VPWR.t492 646.071
R8409 VPWR.n395 VPWR.t739 646.071
R8410 VPWR.n407 VPWR.t272 646.071
R8411 VPWR.n365 VPWR.t278 646.071
R8412 VPWR.n330 VPWR.t260 646.071
R8413 VPWR.n86 VPWR.t1744 646.071
R8414 VPWR.n937 VPWR.t1016 646.071
R8415 VPWR.n403 VPWR.t1249 646.071
R8416 VPWR.n364 VPWR.t621 646.071
R8417 VPWR.n334 VPWR.t611 646.071
R8418 VPWR.n87 VPWR.t1589 646.071
R8419 VPWR.n473 VPWR.t1393 646.071
R8420 VPWR.n481 VPWR.t830 646.071
R8421 VPWR.n480 VPWR.t1288 646.071
R8422 VPWR.n477 VPWR.t757 646.071
R8423 VPWR.n476 VPWR.t603 646.071
R8424 VPWR.n472 VPWR.t797 646.071
R8425 VPWR.n469 VPWR.t357 646.071
R8426 VPWR.n468 VPWR.t556 646.071
R8427 VPWR.n465 VPWR.t140 646.071
R8428 VPWR.n464 VPWR.t905 646.071
R8429 VPWR.n461 VPWR.t1222 646.071
R8430 VPWR.n460 VPWR.t1186 646.071
R8431 VPWR.n457 VPWR.t1879 646.071
R8432 VPWR.n456 VPWR.t667 646.071
R8433 VPWR.n453 VPWR.t323 646.071
R8434 VPWR.n452 VPWR.t1561 646.071
R8435 VPWR.n526 VPWR.t172 646.071
R8436 VPWR.n482 VPWR.t164 646.071
R8437 VPWR.n538 VPWR.t508 646.071
R8438 VPWR.n534 VPWR.t731 646.071
R8439 VPWR.n530 VPWR.t1008 646.071
R8440 VPWR.n522 VPWR.t256 646.071
R8441 VPWR.n518 VPWR.t295 646.071
R8442 VPWR.n514 VPWR.t578 646.071
R8443 VPWR.n510 VPWR.t640 646.071
R8444 VPWR.n506 VPWR.t1381 646.071
R8445 VPWR.n502 VPWR.t126 646.071
R8446 VPWR.n498 VPWR.t1105 646.071
R8447 VPWR.n494 VPWR.t64 646.071
R8448 VPWR.n490 VPWR.t414 646.071
R8449 VPWR.n486 VPWR.t519 646.071
R8450 VPWR.n483 VPWR.t1779 646.071
R8451 VPWR.n556 VPWR.t480 646.071
R8452 VPWR.n548 VPWR.t1165 646.071
R8453 VPWR.n549 VPWR.t1261 646.071
R8454 VPWR.n552 VPWR.t769 646.071
R8455 VPWR.n553 VPWR.t1821 646.071
R8456 VPWR.n557 VPWR.t250 646.071
R8457 VPWR.n560 VPWR.t432 646.071
R8458 VPWR.n561 VPWR.t993 646.071
R8459 VPWR.n564 VPWR.t692 646.071
R8460 VPWR.n565 VPWR.t893 646.071
R8461 VPWR.n568 VPWR.t1319 646.071
R8462 VPWR.n569 VPWR.t1190 646.071
R8463 VPWR.n572 VPWR.t1867 646.071
R8464 VPWR.n573 VPWR.t7 646.071
R8465 VPWR.n576 VPWR.t311 646.071
R8466 VPWR.n577 VPWR.t1628 646.071
R8467 VPWR.n595 VPWR.t619 646.071
R8468 VPWR.n579 VPWR.t1002 646.071
R8469 VPWR.n583 VPWR.t1286 646.071
R8470 VPWR.n587 VPWR.t723 646.071
R8471 VPWR.n591 VPWR.t1020 646.071
R8472 VPWR.n599 VPWR.t276 646.071
R8473 VPWR.n603 VPWR.t307 646.071
R8474 VPWR.n607 VPWR.t590 646.071
R8475 VPWR.n611 VPWR.t572 646.071
R8476 VPWR.n615 VPWR.t1911 646.071
R8477 VPWR.n619 VPWR.t1360 646.071
R8478 VPWR.n623 VPWR.t1851 646.071
R8479 VPWR.n627 VPWR.t1204 646.071
R8480 VPWR.n631 VPWR.t1127 646.071
R8481 VPWR.n635 VPWR.t531 646.071
R8482 VPWR.n578 VPWR.t1736 646.071
R8483 VPWR.n665 VPWR.t210 646.071
R8484 VPWR.n673 VPWR.t596 646.071
R8485 VPWR.n672 VPWR.t686 646.071
R8486 VPWR.n669 VPWR.t743 646.071
R8487 VPWR.n668 VPWR.t1171 646.071
R8488 VPWR.n664 VPWR.t268 646.071
R8489 VPWR.n661 VPWR.t1896 646.071
R8490 VPWR.n660 VPWR.t840 646.071
R8491 VPWR.n657 VPWR.t498 646.071
R8492 VPWR.n656 VPWR.t548 646.071
R8493 VPWR.n653 VPWR.t1809 646.071
R8494 VPWR.n652 VPWR.t862 646.071
R8495 VPWR.n649 VPWR.t105 646.071
R8496 VPWR.n648 VPWR.t152 646.071
R8497 VPWR.n645 VPWR.t190 646.071
R8498 VPWR.n644 VPWR.t1462 646.071
R8499 VPWR.n718 VPWR.t1391 646.071
R8500 VPWR.n674 VPWR.t826 646.071
R8501 VPWR.n730 VPWR.t221 646.071
R8502 VPWR.n726 VPWR.t759 646.071
R8503 VPWR.n722 VPWR.t1024 646.071
R8504 VPWR.n714 VPWR.t795 646.071
R8505 VPWR.n710 VPWR.t355 646.071
R8506 VPWR.n706 VPWR.t554 646.071
R8507 VPWR.n702 VPWR.t138 646.071
R8508 VPWR.n698 VPWR.t901 646.071
R8509 VPWR.n694 VPWR.t1220 646.071
R8510 VPWR.n690 VPWR.t1182 646.071
R8511 VPWR.n686 VPWR.t1877 646.071
R8512 VPWR.n682 VPWR.t329 646.071
R8513 VPWR.n678 VPWR.t319 646.071
R8514 VPWR.n675 VPWR.t1569 646.071
R8515 VPWR.n748 VPWR.t1226 646.071
R8516 VPWR.n740 VPWR.t144 646.071
R8517 VPWR.n741 VPWR.t1292 646.071
R8518 VPWR.n744 VPWR.t751 646.071
R8519 VPWR.n745 VPWR.t605 646.071
R8520 VPWR.n749 VPWR.t230 646.071
R8521 VPWR.n752 VPWR.t1888 646.071
R8522 VPWR.n753 VPWR.t468 646.071
R8523 VPWR.n756 VPWR.t369 646.071
R8524 VPWR.n757 VPWR.t540 646.071
R8525 VPWR.n760 VPWR.t442 646.071
R8526 VPWR.n761 VPWR.t954 646.071
R8527 VPWR.n764 VPWR.t95 646.071
R8528 VPWR.n765 VPWR.t669 646.071
R8529 VPWR.n768 VPWR.t180 646.071
R8530 VPWR.n769 VPWR.t1529 646.071
R8531 VPWR.n787 VPWR.t476 646.071
R8532 VPWR.n771 VPWR.t1163 646.071
R8533 VPWR.n775 VPWR.t1257 646.071
R8534 VPWR.n779 VPWR.t771 646.071
R8535 VPWR.n783 VPWR.t1819 646.071
R8536 VPWR.n791 VPWR.t246 646.071
R8537 VPWR.n795 VPWR.t428 646.071
R8538 VPWR.n799 VPWR.t991 646.071
R8539 VPWR.n803 VPWR.t1281 646.071
R8540 VPWR.n807 VPWR.t891 646.071
R8541 VPWR.n811 VPWR.t1315 646.071
R8542 VPWR.n815 VPWR.t1188 646.071
R8543 VPWR.n819 VPWR.t1865 646.071
R8544 VPWR.n823 VPWR.t5 646.071
R8545 VPWR.n827 VPWR.t349 646.071
R8546 VPWR.n770 VPWR.t1634 646.071
R8547 VPWR.n857 VPWR.t212 646.071
R8548 VPWR.n865 VPWR.t598 646.071
R8549 VPWR.n864 VPWR.t688 646.071
R8550 VPWR.n861 VPWR.t741 646.071
R8551 VPWR.n860 VPWR.t1175 646.071
R8552 VPWR.n856 VPWR.t270 646.071
R8553 VPWR.n853 VPWR.t1898 646.071
R8554 VPWR.n852 VPWR.t842 646.071
R8555 VPWR.n849 VPWR.t500 646.071
R8556 VPWR.n848 VPWR.t550 646.071
R8557 VPWR.n845 VPWR.t1811 646.071
R8558 VPWR.n844 VPWR.t864 646.071
R8559 VPWR.n841 VPWR.t107 646.071
R8560 VPWR.n840 VPWR.t154 646.071
R8561 VPWR.n837 VPWR.t194 646.071
R8562 VPWR.n836 VPWR.t1454 646.071
R8563 VPWR.n910 VPWR.t1239 646.071
R8564 VPWR.n866 VPWR.t1161 646.071
R8565 VPWR.n922 VPWR.t1255 646.071
R8566 VPWR.n918 VPWR.t773 646.071
R8567 VPWR.n914 VPWR.t1817 646.071
R8568 VPWR.n906 VPWR.t244 646.071
R8569 VPWR.n902 VPWR.t426 646.071
R8570 VPWR.n898 VPWR.t989 646.071
R8571 VPWR.n894 VPWR.t1279 646.071
R8572 VPWR.n890 VPWR.t889 646.071
R8573 VPWR.n886 VPWR.t56 646.071
R8574 VPWR.n882 VPWR.t1841 646.071
R8575 VPWR.n878 VPWR.t1863 646.071
R8576 VPWR.n874 VPWR.t3 646.071
R8577 VPWR.n870 VPWR.t347 646.071
R8578 VPWR.n867 VPWR.t1641 646.071
R8579 VPWR.n940 VPWR.t617 646.071
R8580 VPWR.n979 VPWR.t482 646.071
R8581 VPWR.n1227 VPWR.t416 646.071
R8582 VPWR.n1179 VPWR.t1473 646.071
R8583 VPWR.n399 VPWR.t1177 646.071
R8584 VPWR.n361 VPWR.t1054 646.071
R8585 VPWR.n338 VPWR.t1010 646.071
R8586 VPWR.n92 VPWR.t1481 646.071
R8587 VPWR.n975 VPWR.t1823 646.071
R8588 VPWR.n1485 VPWR.t1058 646.071
R8589 VPWR.n1183 VPWR.t1752 646.071
R8590 VPWR.n941 VPWR.t266 646.071
R8591 VPWR.n983 VPWR.t252 646.071
R8592 VPWR.n1173 VPWR.t280 646.071
R8593 VPWR.n1217 VPWR.t1620 646.071
R8594 VPWR.n415 VPWR.t844 646.071
R8595 VPWR.n419 VPWR.t502 646.071
R8596 VPWR.n423 VPWR.t552 646.071
R8597 VPWR.n427 VPWR.t1813 646.071
R8598 VPWR.n431 VPWR.t866 646.071
R8599 VPWR.n435 VPWR.t109 646.071
R8600 VPWR.n439 VPWR.t156 646.071
R8601 VPWR.n443 VPWR.t196 646.071
R8602 VPWR.n386 VPWR.t1446 646.071
R8603 VPWR.n368 VPWR.t309 646.071
R8604 VPWR.n326 VPWR.t299 646.071
R8605 VPWR.n81 VPWR.t1468 646.071
R8606 VPWR.n987 VPWR.t1006 646.071
R8607 VPWR.n1169 VPWR.t418 646.071
R8608 VPWR.n1214 VPWR.t1728 646.071
R8609 VPWR.n948 VPWR.t570 646.071
R8610 VPWR.n949 VPWR.t1385 646.071
R8611 VPWR.n952 VPWR.t1358 646.071
R8612 VPWR.n953 VPWR.t1849 646.071
R8613 VPWR.n956 VPWR.t72 646.071
R8614 VPWR.n957 VPWR.t1125 646.071
R8615 VPWR.n960 VPWR.t527 646.071
R8616 VPWR.n961 VPWR.t1749 646.071
R8617 VPWR.n991 VPWR.t936 646.071
R8618 VPWR.n1163 VPWR.t282 646.071
R8619 VPWR.n1206 VPWR.t1768 646.071
R8620 VPWR.n360 VPWR.t721 646.071
R8621 VPWR.n342 VPWR.t729 646.071
R8622 VPWR.n93 VPWR.t1719 646.071
R8623 VPWR.n1479 VPWR.t777 646.071
R8624 VPWR.n1180 VPWR.t1592 646.071
R8625 VPWR.n995 VPWR.t694 646.071
R8626 VPWR.n1159 VPWR.t824 646.071
R8627 VPWR.n1203 VPWR.t1513 646.071
R8628 VPWR.n376 VPWR.t1362 646.071
R8629 VPWR.n377 VPWR.t1853 646.071
R8630 VPWR.n380 VPWR.t1206 646.071
R8631 VPWR.n381 VPWR.t331 646.071
R8632 VPWR.n384 VPWR.t335 646.071
R8633 VPWR.n385 VPWR.t1731 646.071
R8634 VPWR.n314 VPWR.t1383 646.071
R8635 VPWR.n74 VPWR.t1741 646.071
R8636 VPWR.n1149 VPWR.t1915 646.071
R8637 VPWR.n1200 VPWR.t1617 646.071
R8638 VPWR.n1003 VPWR.t1321 646.071
R8639 VPWR.n1007 VPWR.t1196 646.071
R8640 VPWR.n1011 VPWR.t1869 646.071
R8641 VPWR.n1015 VPWR.t327 646.071
R8642 VPWR.n1019 VPWR.t313 646.071
R8643 VPWR.n962 VPWR.t1601 646.071
R8644 VPWR.n1472 VPWR.t60 646.071
R8645 VPWR.n1123 VPWR.t1579 646.071
R8646 VPWR.n310 VPWR.t130 646.071
R8647 VPWR.n69 VPWR.t1508 646.071
R8648 VPWR.n1192 VPWR.t1776 646.071
R8649 VPWR.n1049 VPWR.t114 646.071
R8650 VPWR.n1189 VPWR.t1795 646.071
R8651 VPWR.n302 VPWR.t68 646.071
R8652 VPWR.n294 VPWR.t521 646.071
R8653 VPWR.n291 VPWR.t1771 646.071
R8654 VPWR.n1058 VPWR.t1668 646.071
R8655 VPWR.n1748 VPWR.t333 646.071
R8656 VPWR.n1036 VPWR.t339 646.071
R8657 VPWR.n1032 VPWR.t1712 646.071
R8658 VPWR.n1186 VPWR.t1539 646.071
R8659 VPWR.n63 VPWR.t1654 646.071
R8660 VPWR.n57 VPWR.t1427 646.071
R8661 VPWR.n1230 VPWR.t1521 642.13
R8662 VPWR.n1152 VPWR.t1449 642.13
R8663 VPWR.n1226 VPWR.t1657 642.13
R8664 VPWR.n1484 VPWR.t1555 642.13
R8665 VPWR.n1172 VPWR.t1679 642.13
R8666 VPWR.n1168 VPWR.t1430 642.13
R8667 VPWR.n1162 VPWR.t1552 642.13
R8668 VPWR.n1478 VPWR.t1784 642.13
R8669 VPWR.n1158 VPWR.t1693 642.13
R8670 VPWR.n1148 VPWR.t1709 642.13
R8671 VPWR.n1471 VPWR.t1682 642.13
R8672 VPWR.n1048 VPWR.t1582 642.13
R8673 VPWR.n1747 VPWR.t1459 642.13
R8674 VPWR.n1035 VPWR.t1496 642.13
R8675 VPWR.n1031 VPWR.t1604 642.13
R8676 VPWR.n1052 VPWR.t1623 642.13
R8677 VPWR.n2309 VPWR.t829 629.652
R8678 VPWR.n2310 VPWR.t1287 629.652
R8679 VPWR.n2319 VPWR.t756 629.652
R8680 VPWR.n2320 VPWR.t602 629.652
R8681 VPWR.n2329 VPWR.t1392 629.652
R8682 VPWR.n2330 VPWR.t796 629.652
R8683 VPWR.n2339 VPWR.t356 629.652
R8684 VPWR.n2340 VPWR.t555 629.652
R8685 VPWR.n2349 VPWR.t139 629.652
R8686 VPWR.n2350 VPWR.t904 629.652
R8687 VPWR.n2359 VPWR.t1221 629.652
R8688 VPWR.n2360 VPWR.t1185 629.652
R8689 VPWR.n2369 VPWR.t1878 629.652
R8690 VPWR.n2370 VPWR.t666 629.652
R8691 VPWR.n2379 VPWR.t322 629.652
R8692 VPWR.n542 VPWR.t163 629.652
R8693 VPWR.t507 VPWR.n541 629.652
R8694 VPWR.t730 VPWR.n537 629.652
R8695 VPWR.t1007 VPWR.n533 629.652
R8696 VPWR.t171 VPWR.n529 629.652
R8697 VPWR.t255 VPWR.n525 629.652
R8698 VPWR.t294 VPWR.n521 629.652
R8699 VPWR.t577 VPWR.n517 629.652
R8700 VPWR.t639 VPWR.n513 629.652
R8701 VPWR.t1380 VPWR.n509 629.652
R8702 VPWR.t125 VPWR.n505 629.652
R8703 VPWR.t1104 VPWR.n501 629.652
R8704 VPWR.t63 VPWR.n497 629.652
R8705 VPWR.t413 VPWR.n493 629.652
R8706 VPWR.t518 VPWR.n489 629.652
R8707 VPWR.n2281 VPWR.t1164 629.652
R8708 VPWR.t1260 VPWR.n2280 629.652
R8709 VPWR.n2271 VPWR.t768 629.652
R8710 VPWR.t1820 VPWR.n2270 629.652
R8711 VPWR.n2261 VPWR.t479 629.652
R8712 VPWR.t249 VPWR.n2260 629.652
R8713 VPWR.n2251 VPWR.t431 629.652
R8714 VPWR.t992 VPWR.n2250 629.652
R8715 VPWR.n2241 VPWR.t691 629.652
R8716 VPWR.t892 VPWR.n2240 629.652
R8717 VPWR.n2231 VPWR.t1318 629.652
R8718 VPWR.t1189 VPWR.n2230 629.652
R8719 VPWR.n2221 VPWR.t1866 629.652
R8720 VPWR.t6 VPWR.n2220 629.652
R8721 VPWR.n2211 VPWR.t310 629.652
R8722 VPWR.n582 VPWR.t1001 629.652
R8723 VPWR.n586 VPWR.t1285 629.652
R8724 VPWR.n590 VPWR.t722 629.652
R8725 VPWR.n594 VPWR.t1019 629.652
R8726 VPWR.n598 VPWR.t618 629.652
R8727 VPWR.n602 VPWR.t275 629.652
R8728 VPWR.n606 VPWR.t306 629.652
R8729 VPWR.n610 VPWR.t589 629.652
R8730 VPWR.n614 VPWR.t571 629.652
R8731 VPWR.n618 VPWR.t1910 629.652
R8732 VPWR.n622 VPWR.t1359 629.652
R8733 VPWR.n626 VPWR.t1850 629.652
R8734 VPWR.n630 VPWR.t1203 629.652
R8735 VPWR.n634 VPWR.t1126 629.652
R8736 VPWR.n638 VPWR.t530 629.652
R8737 VPWR.n2113 VPWR.t595 629.652
R8738 VPWR.n2114 VPWR.t685 629.652
R8739 VPWR.n2123 VPWR.t742 629.652
R8740 VPWR.n2124 VPWR.t1170 629.652
R8741 VPWR.n2133 VPWR.t209 629.652
R8742 VPWR.n2134 VPWR.t267 629.652
R8743 VPWR.n2143 VPWR.t1895 629.652
R8744 VPWR.n2144 VPWR.t839 629.652
R8745 VPWR.n2153 VPWR.t497 629.652
R8746 VPWR.n2154 VPWR.t547 629.652
R8747 VPWR.n2163 VPWR.t1808 629.652
R8748 VPWR.n2164 VPWR.t861 629.652
R8749 VPWR.n2173 VPWR.t104 629.652
R8750 VPWR.n2174 VPWR.t151 629.652
R8751 VPWR.n2183 VPWR.t189 629.652
R8752 VPWR.n734 VPWR.t825 629.652
R8753 VPWR.t220 VPWR.n733 629.652
R8754 VPWR.t758 VPWR.n729 629.652
R8755 VPWR.t1023 VPWR.n725 629.652
R8756 VPWR.t1390 VPWR.n721 629.652
R8757 VPWR.t794 VPWR.n717 629.652
R8758 VPWR.t354 VPWR.n713 629.652
R8759 VPWR.t553 VPWR.n709 629.652
R8760 VPWR.t137 VPWR.n705 629.652
R8761 VPWR.t900 VPWR.n701 629.652
R8762 VPWR.t1219 VPWR.n697 629.652
R8763 VPWR.t1181 VPWR.n693 629.652
R8764 VPWR.t1876 VPWR.n689 629.652
R8765 VPWR.t328 VPWR.n685 629.652
R8766 VPWR.t318 VPWR.n681 629.652
R8767 VPWR.n2085 VPWR.t143 629.652
R8768 VPWR.t1291 VPWR.n2084 629.652
R8769 VPWR.n2075 VPWR.t750 629.652
R8770 VPWR.t604 VPWR.n2074 629.652
R8771 VPWR.n2065 VPWR.t1225 629.652
R8772 VPWR.t229 VPWR.n2064 629.652
R8773 VPWR.n2055 VPWR.t1887 629.652
R8774 VPWR.t467 VPWR.n2054 629.652
R8775 VPWR.n2045 VPWR.t368 629.652
R8776 VPWR.t539 VPWR.n2044 629.652
R8777 VPWR.n2035 VPWR.t441 629.652
R8778 VPWR.t953 VPWR.n2034 629.652
R8779 VPWR.n2025 VPWR.t94 629.652
R8780 VPWR.t668 VPWR.n2024 629.652
R8781 VPWR.n2015 VPWR.t179 629.652
R8782 VPWR.n774 VPWR.t1162 629.652
R8783 VPWR.n778 VPWR.t1256 629.652
R8784 VPWR.n782 VPWR.t770 629.652
R8785 VPWR.n786 VPWR.t1818 629.652
R8786 VPWR.n790 VPWR.t475 629.652
R8787 VPWR.n794 VPWR.t245 629.652
R8788 VPWR.n798 VPWR.t427 629.652
R8789 VPWR.n802 VPWR.t990 629.652
R8790 VPWR.n806 VPWR.t1280 629.652
R8791 VPWR.n810 VPWR.t890 629.652
R8792 VPWR.n814 VPWR.t1314 629.652
R8793 VPWR.n818 VPWR.t1187 629.652
R8794 VPWR.n822 VPWR.t1864 629.652
R8795 VPWR.n826 VPWR.t4 629.652
R8796 VPWR.n830 VPWR.t348 629.652
R8797 VPWR.n1917 VPWR.t597 629.652
R8798 VPWR.n1918 VPWR.t687 629.652
R8799 VPWR.n1927 VPWR.t740 629.652
R8800 VPWR.n1928 VPWR.t1174 629.652
R8801 VPWR.n1937 VPWR.t211 629.652
R8802 VPWR.n1938 VPWR.t269 629.652
R8803 VPWR.n1947 VPWR.t1897 629.652
R8804 VPWR.n1948 VPWR.t841 629.652
R8805 VPWR.n1957 VPWR.t499 629.652
R8806 VPWR.n1958 VPWR.t549 629.652
R8807 VPWR.n1967 VPWR.t1810 629.652
R8808 VPWR.n1968 VPWR.t863 629.652
R8809 VPWR.n1977 VPWR.t106 629.652
R8810 VPWR.n1978 VPWR.t153 629.652
R8811 VPWR.n1987 VPWR.t193 629.652
R8812 VPWR.n926 VPWR.t1160 629.652
R8813 VPWR.t1254 VPWR.n925 629.652
R8814 VPWR.t772 VPWR.n921 629.652
R8815 VPWR.t1816 VPWR.n917 629.652
R8816 VPWR.t1238 VPWR.n913 629.652
R8817 VPWR.t243 VPWR.n909 629.652
R8818 VPWR.t425 VPWR.n905 629.652
R8819 VPWR.t988 VPWR.n901 629.652
R8820 VPWR.t1278 VPWR.n897 629.652
R8821 VPWR.t888 VPWR.n893 629.652
R8822 VPWR.t55 VPWR.n889 629.652
R8823 VPWR.t1840 VPWR.n885 629.652
R8824 VPWR.t1862 VPWR.n881 629.652
R8825 VPWR.t2 VPWR.n877 629.652
R8826 VPWR.t346 VPWR.n873 629.652
R8827 VPWR.n390 VPWR.t599 629.652
R8828 VPWR.n394 VPWR.t491 629.652
R8829 VPWR.n398 VPWR.t738 629.652
R8830 VPWR.n402 VPWR.t1176 629.652
R8831 VPWR.n406 VPWR.t1248 629.652
R8832 VPWR.n410 VPWR.t271 629.652
R8833 VPWR.n414 VPWR.t1899 629.652
R8834 VPWR.n418 VPWR.t843 629.652
R8835 VPWR.n422 VPWR.t501 629.652
R8836 VPWR.n426 VPWR.t551 629.652
R8837 VPWR.n430 VPWR.t1812 629.652
R8838 VPWR.n434 VPWR.t865 629.652
R8839 VPWR.n438 VPWR.t108 629.652
R8840 VPWR.n442 VPWR.t155 629.652
R8841 VPWR.n446 VPWR.t195 629.652
R8842 VPWR.n1889 VPWR.t999 629.652
R8843 VPWR.t489 VPWR.n1888 629.652
R8844 VPWR.n1879 VPWR.t724 629.652
R8845 VPWR.t1015 VPWR.n1878 629.652
R8846 VPWR.n1869 VPWR.t616 629.652
R8847 VPWR.t265 VPWR.n1868 629.652
R8848 VPWR.n1859 VPWR.t304 629.652
R8849 VPWR.t585 VPWR.n1858 629.652
R8850 VPWR.n1849 VPWR.t569 629.652
R8851 VPWR.t1384 VPWR.n1848 629.652
R8852 VPWR.n1839 VPWR.t1357 629.652
R8853 VPWR.t1848 VPWR.n1838 629.652
R8854 VPWR.n1829 VPWR.t71 629.652
R8855 VPWR.t1124 VPWR.n1828 629.652
R8856 VPWR.n1819 VPWR.t526 629.652
R8857 VPWR.n2477 VPWR.t1003 629.652
R8858 VPWR.t57 VPWR.n2476 629.652
R8859 VPWR.n2467 VPWR.t720 629.652
R8860 VPWR.t1053 VPWR.n2466 629.652
R8861 VPWR.n2457 VPWR.t620 629.652
R8862 VPWR.t277 VPWR.n2456 629.652
R8863 VPWR.n2447 VPWR.t308 629.652
R8864 VPWR.t591 VPWR.n2446 629.652
R8865 VPWR.n2437 VPWR.t573 629.652
R8866 VPWR.t1912 VPWR.n2436 629.652
R8867 VPWR.n2427 VPWR.t1361 629.652
R8868 VPWR.t1852 VPWR.n2426 629.652
R8869 VPWR.n2417 VPWR.t1205 629.652
R8870 VPWR.t330 VPWR.n2416 629.652
R8871 VPWR.n2407 VPWR.t334 629.652
R8872 VPWR.n966 VPWR.t1148 629.652
R8873 VPWR.n970 VPWR.t1262 629.652
R8874 VPWR.n974 VPWR.t760 629.652
R8875 VPWR.n978 VPWR.t1822 629.652
R8876 VPWR.n982 VPWR.t481 629.652
R8877 VPWR.n986 VPWR.t251 629.652
R8878 VPWR.n990 VPWR.t1005 629.652
R8879 VPWR.n994 VPWR.t935 629.652
R8880 VPWR.n998 VPWR.t693 629.652
R8881 VPWR.n1002 VPWR.t898 629.652
R8882 VPWR.n1006 VPWR.t1320 629.652
R8883 VPWR.n1010 VPWR.t1195 629.652
R8884 VPWR.n1014 VPWR.t1868 629.652
R8885 VPWR.n1018 VPWR.t326 629.652
R8886 VPWR.n1022 VPWR.t312 629.652
R8887 VPWR.n350 VPWR.t165 629.652
R8888 VPWR.t483 VPWR.n349 629.652
R8889 VPWR.t728 VPWR.n345 629.652
R8890 VPWR.t1009 VPWR.n341 629.652
R8891 VPWR.t610 VPWR.n337 629.652
R8892 VPWR.t259 VPWR.n333 629.652
R8893 VPWR.t298 VPWR.n329 629.652
R8894 VPWR.t581 VPWR.n325 629.652
R8895 VPWR.t643 VPWR.n321 629.652
R8896 VPWR.t1382 VPWR.n317 629.652
R8897 VPWR.t129 VPWR.n313 629.652
R8898 VPWR.t1846 VPWR.n309 629.652
R8899 VPWR.t67 VPWR.n305 629.652
R8900 VPWR.t1122 VPWR.n301 629.652
R8901 VPWR.t520 VPWR.n297 629.652
R8902 VPWR.n1468 VPWR.t454 629.652
R8903 VPWR.n1475 VPWR.t59 629.652
R8904 VPWR.n1481 VPWR.t776 629.652
R8905 VPWR.n1492 VPWR.t1057 629.652
R8906 VPWR.n1493 VPWR.t415 629.652
R8907 VPWR.n1506 VPWR.t279 629.652
R8908 VPWR.n1507 VPWR.t417 629.652
R8909 VPWR.n1520 VPWR.t281 629.652
R8910 VPWR.n1521 VPWR.t823 629.652
R8911 VPWR.n1536 VPWR.t1914 629.652
R8912 VPWR.t1363 VPWR.n1535 629.652
R8913 VPWR.n1761 VPWR.t113 629.652
R8914 VPWR.t1207 VPWR.n1760 629.652
R8915 VPWR.n1749 VPWR.t332 629.652
R8916 VPWR.n1791 VPWR.t338 629.652
R8917 VPWR.n2506 VPWR.t1571 629.652
R8918 VPWR.n2507 VPWR.t1700 629.652
R8919 VPWR.n2518 VPWR.t1718 629.652
R8920 VPWR.n2519 VPWR.t1480 629.652
R8921 VPWR.n2530 VPWR.t1588 629.652
R8922 VPWR.n2531 VPWR.t1743 629.652
R8923 VPWR.n2542 VPWR.t1467 629.652
R8924 VPWR.n2543 VPWR.t1502 629.652
R8925 VPWR.n2554 VPWR.t1630 629.652
R8926 VPWR.n2555 VPWR.t1740 629.652
R8927 VPWR.n2566 VPWR.t1507 629.652
R8928 VPWR.n2567 VPWR.t1525 629.652
R8929 VPWR.n2578 VPWR.t1653 629.652
R8930 VPWR.n2579 VPWR.t1786 629.652
R8931 VPWR.n2590 VPWR.t1426 629.652
R8932 VPWR.n1594 VPWR.t1442 629.652
R8933 VPWR.t1578 VPWR.n1593 629.652
R8934 VPWR.n1182 VPWR.t1591 629.652
R8935 VPWR.n1185 VPWR.t1751 629.652
R8936 VPWR.n1220 VPWR.t1472 629.652
R8937 VPWR.t1619 VPWR.n1219 629.652
R8938 VPWR.t1727 VPWR.n1216 629.652
R8939 VPWR.t1767 VPWR.n1213 629.652
R8940 VPWR.t1512 VPWR.n1205 629.652
R8941 VPWR.t1616 VPWR.n1202 629.652
R8942 VPWR.t1775 VPWR.n1199 629.652
R8943 VPWR.t1794 VPWR.n1191 629.652
R8944 VPWR.t1538 VPWR.n1188 629.652
R8945 VPWR.n1740 VPWR.t1667 629.652
R8946 VPWR.t1695 VPWR.n1739 629.652
R8947 VPWR.n2836 VPWR.t718 531.804
R8948 VPWR.n2855 VPWR.t718 531.804
R8949 VPWR.n2851 VPWR.n2850 504.707
R8950 VPWR.t829 VPWR.t376 486.048
R8951 VPWR.t1287 VPWR.t453 486.048
R8952 VPWR.t1856 VPWR.t756 486.048
R8953 VPWR.t602 VPWR.t1855 486.048
R8954 VPWR.t375 VPWR.t1392 486.048
R8955 VPWR.t796 VPWR.t451 486.048
R8956 VPWR.t450 VPWR.t356 486.048
R8957 VPWR.t555 VPWR.t374 486.048
R8958 VPWR.t1216 VPWR.t139 486.048
R8959 VPWR.t904 VPWR.t452 486.048
R8960 VPWR.t1854 VPWR.t1221 486.048
R8961 VPWR.t1185 VPWR.t377 486.048
R8962 VPWR.t449 VPWR.t1878 486.048
R8963 VPWR.t666 VPWR.t1858 486.048
R8964 VPWR.t1857 VPWR.t322 486.048
R8965 VPWR.t1560 VPWR.t1215 486.048
R8966 VPWR.t163 VPWR.t978 486.048
R8967 VPWR.t1365 VPWR.t507 486.048
R8968 VPWR.t949 VPWR.t730 486.048
R8969 VPWR.t981 VPWR.t1007 486.048
R8970 VPWR.t1369 VPWR.t171 486.048
R8971 VPWR.t976 VPWR.t255 486.048
R8972 VPWR.t975 VPWR.t294 486.048
R8973 VPWR.t1368 VPWR.t577 486.048
R8974 VPWR.t1367 VPWR.t639 486.048
R8975 VPWR.t977 VPWR.t1380 486.048
R8976 VPWR.t980 VPWR.t125 486.048
R8977 VPWR.t979 VPWR.t1104 486.048
R8978 VPWR.t974 VPWR.t63 486.048
R8979 VPWR.t973 VPWR.t413 486.048
R8980 VPWR.t950 VPWR.t518 486.048
R8981 VPWR.t1366 VPWR.t1778 486.048
R8982 VPWR.t1164 VPWR.t1807 486.048
R8983 VPWR.t1802 VPWR.t1260 486.048
R8984 VPWR.t768 VPWR.t1345 486.048
R8985 VPWR.t1344 VPWR.t1820 486.048
R8986 VPWR.t479 VPWR.t1806 486.048
R8987 VPWR.t1350 VPWR.t249 486.048
R8988 VPWR.t431 VPWR.t1349 486.048
R8989 VPWR.t1805 VPWR.t992 486.048
R8990 VPWR.t691 VPWR.t1804 486.048
R8991 VPWR.t1351 VPWR.t892 486.048
R8992 VPWR.t1318 VPWR.t1343 486.048
R8993 VPWR.t1342 VPWR.t1189 486.048
R8994 VPWR.t1866 VPWR.t1348 486.048
R8995 VPWR.t1347 VPWR.t6 486.048
R8996 VPWR.t310 VPWR.t1346 486.048
R8997 VPWR.t1803 VPWR.t1627 486.048
R8998 VPWR.t1001 VPWR.t944 486.048
R8999 VPWR.t1285 VPWR.t1049 486.048
R9000 VPWR.t722 VPWR.t948 486.048
R9001 VPWR.t1019 VPWR.t947 486.048
R9002 VPWR.t618 VPWR.t943 486.048
R9003 VPWR.t275 VPWR.t1047 486.048
R9004 VPWR.t306 VPWR.t1046 486.048
R9005 VPWR.t589 VPWR.t1052 486.048
R9006 VPWR.t571 VPWR.t1051 486.048
R9007 VPWR.t1910 VPWR.t1048 486.048
R9008 VPWR.t1359 VPWR.t946 486.048
R9009 VPWR.t1850 VPWR.t945 486.048
R9010 VPWR.t1203 VPWR.t1045 486.048
R9011 VPWR.t1126 VPWR.t1044 486.048
R9012 VPWR.t530 VPWR.t513 486.048
R9013 VPWR.t1735 VPWR.t1050 486.048
R9014 VPWR.t595 VPWR.t199 486.048
R9015 VPWR.t685 VPWR.t1178 486.048
R9016 VPWR.t594 VPWR.t742 486.048
R9017 VPWR.t1170 VPWR.t593 486.048
R9018 VPWR.t198 VPWR.t209 486.048
R9019 VPWR.t267 VPWR.t1245 486.048
R9020 VPWR.t1244 VPWR.t1895 486.048
R9021 VPWR.t839 VPWR.t197 486.048
R9022 VPWR.t1180 VPWR.t497 486.048
R9023 VPWR.t547 VPWR.t1246 486.048
R9024 VPWR.t671 VPWR.t1808 486.048
R9025 VPWR.t861 VPWR.t670 486.048
R9026 VPWR.t1243 VPWR.t104 486.048
R9027 VPWR.t151 VPWR.t673 486.048
R9028 VPWR.t672 VPWR.t189 486.048
R9029 VPWR.t1461 VPWR.t1179 486.048
R9030 VPWR.t825 VPWR.t705 486.048
R9031 VPWR.t46 VPWR.t220 486.048
R9032 VPWR.t907 VPWR.t758 486.048
R9033 VPWR.t906 VPWR.t1023 486.048
R9034 VPWR.t704 VPWR.t1390 486.048
R9035 VPWR.t1199 VPWR.t794 486.048
R9036 VPWR.t1198 VPWR.t354 486.048
R9037 VPWR.t289 VPWR.t553 486.048
R9038 VPWR.t48 VPWR.t137 486.048
R9039 VPWR.t1200 VPWR.t900 486.048
R9040 VPWR.t707 VPWR.t1219 486.048
R9041 VPWR.t706 VPWR.t1181 486.048
R9042 VPWR.t1197 VPWR.t1876 486.048
R9043 VPWR.t909 VPWR.t328 486.048
R9044 VPWR.t908 VPWR.t318 486.048
R9045 VPWR.t47 VPWR.t1568 486.048
R9046 VPWR.t143 VPWR.t1883 486.048
R9047 VPWR.t386 VPWR.t1291 486.048
R9048 VPWR.t750 VPWR.t379 486.048
R9049 VPWR.t1886 VPWR.t604 486.048
R9050 VPWR.t1225 VPWR.t1882 486.048
R9051 VPWR.t384 VPWR.t229 486.048
R9052 VPWR.t1887 VPWR.t383 486.048
R9053 VPWR.t1881 VPWR.t467 486.048
R9054 VPWR.t368 VPWR.t1880 486.048
R9055 VPWR.t385 VPWR.t539 486.048
R9056 VPWR.t441 VPWR.t1885 486.048
R9057 VPWR.t1884 VPWR.t953 486.048
R9058 VPWR.t94 VPWR.t382 486.048
R9059 VPWR.t381 VPWR.t668 486.048
R9060 VPWR.t179 VPWR.t380 486.048
R9061 VPWR.t378 VPWR.t1528 486.048
R9062 VPWR.t1162 VPWR.t1339 486.048
R9063 VPWR.t1256 VPWR.t1334 486.048
R9064 VPWR.t770 VPWR.t1030 486.048
R9065 VPWR.t1818 VPWR.t1029 486.048
R9066 VPWR.t475 VPWR.t1338 486.048
R9067 VPWR.t245 VPWR.t1035 486.048
R9068 VPWR.t427 VPWR.t1034 486.048
R9069 VPWR.t990 VPWR.t1337 486.048
R9070 VPWR.t1280 VPWR.t1336 486.048
R9071 VPWR.t890 VPWR.t1036 486.048
R9072 VPWR.t1314 VPWR.t1028 486.048
R9073 VPWR.t1187 VPWR.t1027 486.048
R9074 VPWR.t1864 VPWR.t1033 486.048
R9075 VPWR.t4 VPWR.t1032 486.048
R9076 VPWR.t348 VPWR.t1031 486.048
R9077 VPWR.t1633 VPWR.t1335 486.048
R9078 VPWR.t597 VPWR.t363 486.048
R9079 VPWR.t687 VPWR.t1826 486.048
R9080 VPWR.t532 VPWR.t740 486.048
R9081 VPWR.t1174 VPWR.t366 486.048
R9082 VPWR.t362 VPWR.t211 486.048
R9083 VPWR.t269 VPWR.t537 486.048
R9084 VPWR.t536 VPWR.t1897 486.048
R9085 VPWR.t841 VPWR.t361 486.048
R9086 VPWR.t360 VPWR.t499 486.048
R9087 VPWR.t549 VPWR.t538 486.048
R9088 VPWR.t365 VPWR.t1810 486.048
R9089 VPWR.t863 VPWR.t364 486.048
R9090 VPWR.t535 VPWR.t106 486.048
R9091 VPWR.t153 VPWR.t534 486.048
R9092 VPWR.t533 VPWR.t193 486.048
R9093 VPWR.t1453 VPWR.t1827 486.048
R9094 VPWR.t1160 VPWR.t120 486.048
R9095 VPWR.t115 VPWR.t1254 486.048
R9096 VPWR.t871 VPWR.t772 486.048
R9097 VPWR.t1231 VPWR.t1816 486.048
R9098 VPWR.t119 VPWR.t1238 486.048
R9099 VPWR.t876 VPWR.t243 486.048
R9100 VPWR.t875 VPWR.t425 486.048
R9101 VPWR.t118 VPWR.t988 486.048
R9102 VPWR.t117 VPWR.t1278 486.048
R9103 VPWR.t877 VPWR.t888 486.048
R9104 VPWR.t1230 VPWR.t55 486.048
R9105 VPWR.t1229 VPWR.t1840 486.048
R9106 VPWR.t874 VPWR.t1862 486.048
R9107 VPWR.t873 VPWR.t2 486.048
R9108 VPWR.t872 VPWR.t346 486.048
R9109 VPWR.t116 VPWR.t1640 486.048
R9110 VPWR.t599 VPWR.t678 486.048
R9111 VPWR.t491 VPWR.t1247 486.048
R9112 VPWR.t738 VPWR.t632 486.048
R9113 VPWR.t1176 VPWR.t631 486.048
R9114 VPWR.t1248 VPWR.t677 486.048
R9115 VPWR.t271 VPWR.t207 486.048
R9116 VPWR.t1899 VPWR.t206 486.048
R9117 VPWR.t843 VPWR.t676 486.048
R9118 VPWR.t501 VPWR.t675 486.048
R9119 VPWR.t551 VPWR.t208 486.048
R9120 VPWR.t1812 VPWR.t630 486.048
R9121 VPWR.t865 VPWR.t629 486.048
R9122 VPWR.t108 VPWR.t205 486.048
R9123 VPWR.t155 VPWR.t204 486.048
R9124 VPWR.t195 VPWR.t203 486.048
R9125 VPWR.t1445 VPWR.t674 486.048
R9126 VPWR.t999 VPWR.t21 486.048
R9127 VPWR.t1330 VPWR.t489 486.048
R9128 VPWR.t724 VPWR.t1333 486.048
R9129 VPWR.t24 VPWR.t1015 486.048
R9130 VPWR.t616 VPWR.t20 486.048
R9131 VPWR.t1328 VPWR.t265 486.048
R9132 VPWR.t304 VPWR.t1153 486.048
R9133 VPWR.t19 VPWR.t585 486.048
R9134 VPWR.t569 VPWR.t1332 486.048
R9135 VPWR.t1329 VPWR.t1384 486.048
R9136 VPWR.t1357 VPWR.t23 486.048
R9137 VPWR.t22 VPWR.t1848 486.048
R9138 VPWR.t71 VPWR.t1152 486.048
R9139 VPWR.t1151 VPWR.t1124 486.048
R9140 VPWR.t526 VPWR.t1150 486.048
R9141 VPWR.t1331 VPWR.t1748 486.048
R9142 VPWR.t1003 VPWR.t1356 486.048
R9143 VPWR.t1861 VPWR.t57 486.048
R9144 VPWR.t720 VPWR.t816 486.048
R9145 VPWR.t202 VPWR.t1053 486.048
R9146 VPWR.t620 VPWR.t1355 486.048
R9147 VPWR.t1859 VPWR.t277 486.048
R9148 VPWR.t308 VPWR.t820 486.048
R9149 VPWR.t1354 VPWR.t591 486.048
R9150 VPWR.t573 VPWR.t1353 486.048
R9151 VPWR.t1860 VPWR.t1912 486.048
R9152 VPWR.t1361 VPWR.t201 486.048
R9153 VPWR.t200 VPWR.t1852 486.048
R9154 VPWR.t1205 VPWR.t819 486.048
R9155 VPWR.t818 VPWR.t330 486.048
R9156 VPWR.t334 VPWR.t817 486.048
R9157 VPWR.t1352 VPWR.t1730 486.048
R9158 VPWR.t1148 VPWR.t697 486.048
R9159 VPWR.t1262 VPWR.t215 486.048
R9160 VPWR.t760 VPWR.t701 486.048
R9161 VPWR.t1822 VPWR.t700 486.048
R9162 VPWR.t481 VPWR.t636 486.048
R9163 VPWR.t251 VPWR.t213 486.048
R9164 VPWR.t1005 VPWR.t985 486.048
R9165 VPWR.t935 VPWR.t635 486.048
R9166 VPWR.t693 VPWR.t634 486.048
R9167 VPWR.t898 VPWR.t214 486.048
R9168 VPWR.t1320 VPWR.t699 486.048
R9169 VPWR.t1195 VPWR.t698 486.048
R9170 VPWR.t1868 VPWR.t984 486.048
R9171 VPWR.t326 VPWR.t983 486.048
R9172 VPWR.t312 VPWR.t982 486.048
R9173 VPWR.t1600 VPWR.t633 486.048
R9174 VPWR.t165 VPWR.t711 486.048
R9175 VPWR.t1042 VPWR.t483 486.048
R9176 VPWR.t662 VPWR.t728 486.048
R9177 VPWR.t661 VPWR.t1009 486.048
R9178 VPWR.t710 VPWR.t610 486.048
R9179 VPWR.t1040 VPWR.t259 486.048
R9180 VPWR.t1039 VPWR.t298 486.048
R9181 VPWR.t709 VPWR.t581 486.048
R9182 VPWR.t708 VPWR.t643 486.048
R9183 VPWR.t1041 VPWR.t1382 486.048
R9184 VPWR.t713 VPWR.t129 486.048
R9185 VPWR.t712 VPWR.t1846 486.048
R9186 VPWR.t1038 VPWR.t67 486.048
R9187 VPWR.t1037 VPWR.t1122 486.048
R9188 VPWR.t663 VPWR.t520 486.048
R9189 VPWR.t1043 VPWR.t1770 486.048
R9190 VPWR.t454 VPWR.t1505 486.048
R9191 VPWR.t59 VPWR.t1636 486.048
R9192 VPWR.t776 VPWR.t1765 486.048
R9193 VPWR.t1057 VPWR.t1421 486.048
R9194 VPWR.t415 VPWR.t1531 486.048
R9195 VPWR.t1686 VPWR.t279 486.048
R9196 VPWR.t417 VPWR.t1688 486.048
R9197 VPWR.t1536 VPWR.t281 486.048
R9198 VPWR.t823 VPWR.t1566 486.048
R9199 VPWR.t1684 VPWR.t1914 486.048
R9200 VPWR.t1435 VPWR.t1363 486.048
R9201 VPWR.t1451 VPWR.t113 486.048
R9202 VPWR.t1698 VPWR.t1207 486.048
R9203 VPWR.t332 VPWR.t1716 486.048
R9204 VPWR.t1754 VPWR.t338 486.048
R9205 VPWR.t1711 VPWR.t1586 486.048
R9206 VPWR.t1571 VPWR.t1440 486.048
R9207 VPWR.t1700 VPWR.t1576 486.048
R9208 VPWR.t1706 VPWR.t1718 486.048
R9209 VPWR.t1480 VPWR.t1746 486.048
R9210 VPWR.t1470 VPWR.t1588 486.048
R9211 VPWR.t1743 VPWR.t1614 486.048
R9212 VPWR.t1638 VPWR.t1467 486.048
R9213 VPWR.t1502 VPWR.t1475 486.048
R9214 VPWR.t1510 VPWR.t1630 486.048
R9215 VPWR.t1740 VPWR.t1612 486.048
R9216 VPWR.t1773 VPWR.t1507 486.048
R9217 VPWR.t1525 VPWR.t1792 486.048
R9218 VPWR.t1646 VPWR.t1653 486.048
R9219 VPWR.t1786 VPWR.t1665 486.048
R9220 VPWR.t1690 VPWR.t1426 486.048
R9221 VPWR.t1662 VPWR.t1541 486.048
R9222 VPWR.t1442 VPWR.t1714 486.048
R9223 VPWR.t1456 VPWR.t1578 486.048
R9224 VPWR.t1591 VPWR.t1584 486.048
R9225 VPWR.t1751 VPWR.t1625 486.048
R9226 VPWR.t1472 VPWR.t1733 486.048
R9227 VPWR.t1500 VPWR.t1619 486.048
R9228 VPWR.t1515 VPWR.t1727 486.048
R9229 VPWR.t1738 VPWR.t1767 486.048
R9230 VPWR.t1781 VPWR.t1512 486.048
R9231 VPWR.t1498 VPWR.t1616 486.048
R9232 VPWR.t1651 VPWR.t1775 486.048
R9233 VPWR.t1673 VPWR.t1794 486.048
R9234 VPWR.t1523 VPWR.t1538 486.048
R9235 VPWR.t1549 VPWR.t1667 486.048
R9236 VPWR.t1574 VPWR.t1695 486.048
R9237 VPWR.t1546 VPWR.t1419 486.048
R9238 VPWR.t376 VPWR.t1094 463.954
R9239 VPWR.t453 VPWR.t1146 463.954
R9240 VPWR.t218 VPWR.t1856 463.954
R9241 VPWR.t1855 VPWR.t778 463.954
R9242 VPWR.t1061 VPWR.t375 463.954
R9243 VPWR.t451 VPWR.t1388 463.954
R9244 VPWR.t792 VPWR.t450 463.954
R9245 VPWR.t374 VPWR.t352 463.954
R9246 VPWR.t285 VPWR.t1216 463.954
R9247 VPWR.t452 VPWR.t135 463.954
R9248 VPWR.t896 VPWR.t1854 463.954
R9249 VPWR.t377 VPWR.t1217 463.954
R9250 VPWR.t1193 VPWR.t449 463.954
R9251 VPWR.t1858 VPWR.t1211 463.954
R9252 VPWR.t324 VPWR.t1857 463.954
R9253 VPWR.t1215 VPWR.t342 463.954
R9254 VPWR.t978 VPWR.t1084 463.954
R9255 VPWR.t175 VPWR.t1365 463.954
R9256 VPWR.t503 VPWR.t949 463.954
R9257 VPWR.t754 VPWR.t981 463.954
R9258 VPWR.t606 VPWR.t1369 463.954
R9259 VPWR.t167 VPWR.t976 463.954
R9260 VPWR.t273 VPWR.t975 463.954
R9261 VPWR.t290 VPWR.t1368 463.954
R9262 VPWR.t465 VPWR.t1367 463.954
R9263 VPWR.t511 VPWR.t977 463.954
R9264 VPWR.t1370 VPWR.t980 463.954
R9265 VPWR.t121 VPWR.t979 463.954
R9266 VPWR.t853 VPWR.t974 463.954
R9267 VPWR.t92 VPWR.t973 463.954
R9268 VPWR.t433 VPWR.t950 463.954
R9269 VPWR.t181 VPWR.t1366 463.954
R9270 VPWR.t1807 VPWR.t1069 463.954
R9271 VPWR.t1156 VPWR.t1802 463.954
R9272 VPWR.t1345 VPWR.t226 463.954
R9273 VPWR.t732 VPWR.t1344 463.954
R9274 VPWR.t1806 VPWR.t1017 463.954
R9275 VPWR.t1236 VPWR.t1350 463.954
R9276 VPWR.t1349 VPWR.t241 463.954
R9277 VPWR.t423 VPWR.t1805 463.954
R9278 VPWR.t1804 VPWR.t583 463.954
R9279 VPWR.t1276 VPWR.t1351 463.954
R9280 VPWR.t1343 VPWR.t1303 463.954
R9281 VPWR.t53 VPWR.t1342 463.954
R9282 VPWR.t1348 VPWR.t1836 463.954
R9283 VPWR.t69 VPWR.t1347 463.954
R9284 VPWR.t1346 VPWR.t626 463.954
R9285 VPWR.t528 VPWR.t1803 463.954
R9286 VPWR.t944 VPWR.t1077 463.954
R9287 VPWR.t1049 VPWR.t159 463.954
R9288 VPWR.t948 VPWR.t485 463.954
R9289 VPWR.t947 VPWR.t746 463.954
R9290 VPWR.t943 VPWR.t1168 463.954
R9291 VPWR.t1047 VPWR.t612 463.954
R9292 VPWR.t1046 VPWR.t261 463.954
R9293 VPWR.t1052 VPWR.t300 463.954
R9294 VPWR.t1051 VPWR.t473 463.954
R9295 VPWR.t1048 VPWR.t565 463.954
R9296 VPWR.t946 VPWR.t1376 463.954
R9297 VPWR.t945 VPWR.t131 463.954
R9298 VPWR.t1045 VPWR.t1100 463.954
R9299 VPWR.t1044 VPWR.t100 463.954
R9300 VPWR.t513 VPWR.t409 463.954
R9301 VPWR.t1050 VPWR.t187 463.954
R9302 VPWR.t199 VPWR.t1090 463.954
R9303 VPWR.t1178 VPWR.t145 463.954
R9304 VPWR.t679 VPWR.t594 463.954
R9305 VPWR.t593 VPWR.t766 463.954
R9306 VPWR.t1824 VPWR.t198 463.954
R9307 VPWR.t1245 VPWR.t1227 463.954
R9308 VPWR.t231 VPWR.t1244 463.954
R9309 VPWR.t197 VPWR.t1889 463.954
R9310 VPWR.t937 VPWR.t1180 463.954
R9311 VPWR.t1246 VPWR.t370 463.954
R9312 VPWR.t541 VPWR.t671 463.954
R9313 VPWR.t670 VPWR.t443 463.954
R9314 VPWR.t955 VPWR.t1243 463.954
R9315 VPWR.t673 VPWR.t1870 463.954
R9316 VPWR.t1116 VPWR.t672 463.954
R9317 VPWR.t1179 VPWR.t314 463.954
R9318 VPWR.t705 VPWR.t1096 463.954
R9319 VPWR.t1144 VPWR.t46 463.954
R9320 VPWR.t216 VPWR.t907 463.954
R9321 VPWR.t780 VPWR.t906 463.954
R9322 VPWR.t1059 VPWR.t704 463.954
R9323 VPWR.t1386 VPWR.t1199 463.954
R9324 VPWR.t790 VPWR.t1198 463.954
R9325 VPWR.t350 VPWR.t289 463.954
R9326 VPWR.t283 VPWR.t48 463.954
R9327 VPWR.t695 VPWR.t1200 463.954
R9328 VPWR.t894 VPWR.t707 463.954
R9329 VPWR.t1322 VPWR.t706 463.954
R9330 VPWR.t1191 VPWR.t1197 463.954
R9331 VPWR.t1209 VPWR.t909 463.954
R9332 VPWR.t8 VPWR.t908 463.954
R9333 VPWR.t340 VPWR.t47 463.954
R9334 VPWR.t1883 VPWR.t1092 463.954
R9335 VPWR.t827 VPWR.t386 463.954
R9336 VPWR.t379 VPWR.t1289 463.954
R9337 VPWR.t774 VPWR.t1886 463.954
R9338 VPWR.t1882 VPWR.t1814 463.954
R9339 VPWR.t1223 VPWR.t384 463.954
R9340 VPWR.t383 VPWR.t798 463.954
R9341 VPWR.t358 VPWR.t1881 463.954
R9342 VPWR.t1880 VPWR.t986 463.954
R9343 VPWR.t141 VPWR.t385 463.954
R9344 VPWR.t1885 VPWR.t902 463.954
R9345 VPWR.t1114 VPWR.t1884 463.954
R9346 VPWR.t382 VPWR.t1183 463.954
R9347 VPWR.t1213 VPWR.t381 463.954
R9348 VPWR.t380 VPWR.t664 463.954
R9349 VPWR.t344 VPWR.t378 463.954
R9350 VPWR.t1339 VPWR.t1071 463.954
R9351 VPWR.t1334 VPWR.t458 463.954
R9352 VPWR.t1030 VPWR.t224 463.954
R9353 VPWR.t1029 VPWR.t734 463.954
R9354 VPWR.t1338 VPWR.t1013 463.954
R9355 VPWR.t1035 VPWR.t1234 463.954
R9356 VPWR.t1034 VPWR.t239 463.954
R9357 VPWR.t1337 VPWR.t421 463.954
R9358 VPWR.t1336 VPWR.t579 463.954
R9359 VPWR.t1036 VPWR.t1274 463.954
R9360 VPWR.t1028 VPWR.t1301 463.954
R9361 VPWR.t1027 VPWR.t51 463.954
R9362 VPWR.t1033 VPWR.t1834 463.954
R9363 VPWR.t1032 VPWR.t65 463.954
R9364 VPWR.t1031 VPWR.t624 463.954
R9365 VPWR.t1335 VPWR.t524 463.954
R9366 VPWR.t363 VPWR.t1088 463.954
R9367 VPWR.t1826 VPWR.t147 463.954
R9368 VPWR.t681 VPWR.t532 463.954
R9369 VPWR.t366 VPWR.t764 463.954
R9370 VPWR.t1021 VPWR.t362 463.954
R9371 VPWR.t537 VPWR.t916 463.954
R9372 VPWR.t233 VPWR.t536 463.954
R9373 VPWR.t361 VPWR.t1891 463.954
R9374 VPWR.t939 VPWR.t360 463.954
R9375 VPWR.t538 VPWR.t493 463.954
R9376 VPWR.t543 VPWR.t365 463.954
R9377 VPWR.t364 VPWR.t445 463.954
R9378 VPWR.t857 VPWR.t535 463.954
R9379 VPWR.t534 VPWR.t1872 463.954
R9380 VPWR.t1118 VPWR.t533 463.954
R9381 VPWR.t1827 VPWR.t316 463.954
R9382 VPWR.t120 VPWR.t1073 463.954
R9383 VPWR.t456 VPWR.t115 463.954
R9384 VPWR.t222 VPWR.t871 463.954
R9385 VPWR.t736 VPWR.t1231 463.954
R9386 VPWR.t1011 VPWR.t119 463.954
R9387 VPWR.t1232 VPWR.t876 463.954
R9388 VPWR.t237 VPWR.t875 463.954
R9389 VPWR.t419 VPWR.t118 463.954
R9390 VPWR.t575 VPWR.t117 463.954
R9391 VPWR.t1272 VPWR.t877 463.954
R9392 VPWR.t1299 VPWR.t1230 463.954
R9393 VPWR.t49 VPWR.t1229 463.954
R9394 VPWR.t1832 VPWR.t874 463.954
R9395 VPWR.t61 VPWR.t873 463.954
R9396 VPWR.t622 VPWR.t872 463.954
R9397 VPWR.t522 VPWR.t116 463.954
R9398 VPWR.t678 VPWR.t1086 463.954
R9399 VPWR.t1247 VPWR.t149 463.954
R9400 VPWR.t632 VPWR.t683 463.954
R9401 VPWR.t631 VPWR.t762 463.954
R9402 VPWR.t677 VPWR.t1025 463.954
R9403 VPWR.t207 VPWR.t918 463.954
R9404 VPWR.t206 VPWR.t235 463.954
R9405 VPWR.t676 VPWR.t1893 463.954
R9406 VPWR.t675 VPWR.t941 463.954
R9407 VPWR.t208 VPWR.t495 463.954
R9408 VPWR.t630 VPWR.t545 463.954
R9409 VPWR.t629 VPWR.t447 463.954
R9410 VPWR.t205 VPWR.t859 463.954
R9411 VPWR.t204 VPWR.t1874 463.954
R9412 VPWR.t203 VPWR.t1120 463.954
R9413 VPWR.t674 VPWR.t320 463.954
R9414 VPWR.t21 VPWR.t1079 463.954
R9415 VPWR.t157 VPWR.t1330 463.954
R9416 VPWR.t1333 VPWR.t509 463.954
R9417 VPWR.t748 VPWR.t24 463.954
R9418 VPWR.t20 VPWR.t1166 463.954
R9419 VPWR.t173 VPWR.t1328 463.954
R9420 VPWR.t1153 VPWR.t257 463.954
R9421 VPWR.t296 VPWR.t19 463.954
R9422 VPWR.t1332 VPWR.t471 463.954
R9423 VPWR.t641 VPWR.t1329 463.954
R9424 VPWR.t23 VPWR.t1374 463.954
R9425 VPWR.t127 VPWR.t22 463.954
R9426 VPWR.t1152 VPWR.t1098 463.954
R9427 VPWR.t98 VPWR.t1151 463.954
R9428 VPWR.t1150 VPWR.t407 463.954
R9429 VPWR.t185 VPWR.t1331 463.954
R9430 VPWR.t1356 VPWR.t1075 463.954
R9431 VPWR.t161 VPWR.t1861 463.954
R9432 VPWR.t816 VPWR.t487 463.954
R9433 VPWR.t744 VPWR.t202 463.954
R9434 VPWR.t1355 VPWR.t1172 463.954
R9435 VPWR.t614 VPWR.t1859 463.954
R9436 VPWR.t820 VPWR.t263 463.954
R9437 VPWR.t302 VPWR.t1354 463.954
R9438 VPWR.t1353 VPWR.t837 463.954
R9439 VPWR.t567 VPWR.t1860 463.954
R9440 VPWR.t201 VPWR.t1378 463.954
R9441 VPWR.t133 VPWR.t200 463.954
R9442 VPWR.t819 VPWR.t1102 463.954
R9443 VPWR.t102 VPWR.t818 463.954
R9444 VPWR.t817 VPWR.t411 463.954
R9445 VPWR.t191 VPWR.t1352 463.954
R9446 VPWR.t697 VPWR.t1067 463.954
R9447 VPWR.t215 VPWR.t1158 463.954
R9448 VPWR.t701 VPWR.t1258 463.954
R9449 VPWR.t700 VPWR.t726 463.954
R9450 VPWR.t636 VPWR.t1055 463.954
R9451 VPWR.t213 VPWR.t477 463.954
R9452 VPWR.t985 VPWR.t247 463.954
R9453 VPWR.t635 VPWR.t429 463.954
R9454 VPWR.t634 VPWR.t587 463.954
R9455 VPWR.t214 VPWR.t689 463.954
R9456 VPWR.t699 VPWR.t1305 463.954
R9457 VPWR.t698 VPWR.t1316 463.954
R9458 VPWR.t984 VPWR.t1838 463.954
R9459 VPWR.t983 VPWR.t1201 463.954
R9460 VPWR.t982 VPWR.t0 463.954
R9461 VPWR.t633 VPWR.t336 463.954
R9462 VPWR.t711 VPWR.t1082 463.954
R9463 VPWR.t177 VPWR.t1042 463.954
R9464 VPWR.t505 VPWR.t662 463.954
R9465 VPWR.t752 VPWR.t661 463.954
R9466 VPWR.t608 VPWR.t710 463.954
R9467 VPWR.t169 VPWR.t1040 463.954
R9468 VPWR.t253 VPWR.t1039 463.954
R9469 VPWR.t292 VPWR.t709 463.954
R9470 VPWR.t469 VPWR.t708 463.954
R9471 VPWR.t637 VPWR.t1041 463.954
R9472 VPWR.t1372 VPWR.t713 463.954
R9473 VPWR.t123 VPWR.t712 463.954
R9474 VPWR.t855 VPWR.t1038 463.954
R9475 VPWR.t96 VPWR.t1037 463.954
R9476 VPWR.t435 VPWR.t663 463.954
R9477 VPWR.t183 VPWR.t1043 463.954
R9478 VPWR.t1505 VPWR.t1520 463.954
R9479 VPWR.t1636 VPWR.t1681 463.954
R9480 VPWR.t1765 VPWR.t1783 463.954
R9481 VPWR.t1421 VPWR.t1554 463.954
R9482 VPWR.t1531 VPWR.t1656 463.954
R9483 VPWR.t1678 VPWR.t1686 463.954
R9484 VPWR.t1688 VPWR.t1429 463.954
R9485 VPWR.t1551 VPWR.t1536 463.954
R9486 VPWR.t1566 VPWR.t1692 463.954
R9487 VPWR.t1708 VPWR.t1684 463.954
R9488 VPWR.t1448 VPWR.t1435 463.954
R9489 VPWR.t1581 VPWR.t1451 463.954
R9490 VPWR.t1622 VPWR.t1698 463.954
R9491 VPWR.t1716 VPWR.t1458 463.954
R9492 VPWR.t1495 VPWR.t1754 463.954
R9493 VPWR.t1586 VPWR.t1603 463.954
R9494 VPWR.t1440 VPWR.t1464 463.954
R9495 VPWR.t1576 VPWR.t1609 463.954
R9496 VPWR.t1721 VPWR.t1706 463.954
R9497 VPWR.t1746 VPWR.t1486 463.954
R9498 VPWR.t1594 VPWR.t1470 463.954
R9499 VPWR.t1614 VPWR.t1606 463.954
R9500 VPWR.t1762 VPWR.t1638 463.954
R9501 VPWR.t1475 VPWR.t1483 463.954
R9502 VPWR.t1643 VPWR.t1510 463.954
R9503 VPWR.t1612 VPWR.t1659 463.954
R9504 VPWR.t1789 VPWR.t1773 463.954
R9505 VPWR.t1792 VPWR.t1533 463.954
R9506 VPWR.t1563 VPWR.t1646 463.954
R9507 VPWR.t1665 VPWR.t1413 463.954
R9508 VPWR.t1432 VPWR.t1690 463.954
R9509 VPWR.t1541 VPWR.t1557 463.954
R9510 VPWR.t1714 VPWR.t1724 463.954
R9511 VPWR.t1492 VPWR.t1456 463.954
R9512 VPWR.t1584 VPWR.t1597 463.954
R9513 VPWR.t1625 VPWR.t1759 463.954
R9514 VPWR.t1733 VPWR.t1477 463.954
R9515 VPWR.t1489 VPWR.t1500 463.954
R9516 VPWR.t1648 VPWR.t1515 463.954
R9517 VPWR.t1756 VPWR.t1738 463.954
R9518 VPWR.t1517 VPWR.t1781 463.954
R9519 VPWR.t1543 VPWR.t1498 463.954
R9520 VPWR.t1670 VPWR.t1651 463.954
R9521 VPWR.t1416 VPWR.t1673 463.954
R9522 VPWR.t1437 VPWR.t1523 463.954
R9523 VPWR.t1675 VPWR.t1549 463.954
R9524 VPWR.t1703 VPWR.t1574 463.954
R9525 VPWR.t1419 VPWR.t1423 463.954
R9526 VPWR.n2626 VPWR.t804 428.822
R9527 VPWR.n1595 VPWR.n1594 376.045
R9528 VPWR.n2506 VPWR.n2505 376.045
R9529 VPWR.n1468 VPWR.n1467 376.045
R9530 VPWR.n351 VPWR.n350 376.045
R9531 VPWR.n2568 VPWR.n2567 376.045
R9532 VPWR.n1535 VPWR.n1534 376.045
R9533 VPWR.n349 VPWR.n348 376.045
R9534 VPWR.n2508 VPWR.n2507 376.045
R9535 VPWR.n966 VPWR.n965 376.045
R9536 VPWR.n2478 VPWR.n2477 376.045
R9537 VPWR.n2476 VPWR.n2475 376.045
R9538 VPWR.n321 VPWR.n320 376.045
R9539 VPWR.n2554 VPWR.n2553 376.045
R9540 VPWR.n974 VPWR.n973 376.045
R9541 VPWR.n2446 VPWR.n2445 376.045
R9542 VPWR.n325 VPWR.n324 376.045
R9543 VPWR.n2544 VPWR.n2543 376.045
R9544 VPWR.n1890 VPWR.n1889 376.045
R9545 VPWR.n1888 VPWR.n1887 376.045
R9546 VPWR.n1880 VPWR.n1879 376.045
R9547 VPWR.n390 VPWR.n389 376.045
R9548 VPWR.n394 VPWR.n393 376.045
R9549 VPWR.n398 VPWR.n397 376.045
R9550 VPWR.n2456 VPWR.n2455 376.045
R9551 VPWR.n333 VPWR.n332 376.045
R9552 VPWR.n2532 VPWR.n2531 376.045
R9553 VPWR.n1878 VPWR.n1877 376.045
R9554 VPWR.n406 VPWR.n405 376.045
R9555 VPWR.n2458 VPWR.n2457 376.045
R9556 VPWR.n337 VPWR.n336 376.045
R9557 VPWR.n2530 VPWR.n2529 376.045
R9558 VPWR.n2309 VPWR.n2308 376.045
R9559 VPWR.n2311 VPWR.n2310 376.045
R9560 VPWR.n2319 VPWR.n2318 376.045
R9561 VPWR.n2321 VPWR.n2320 376.045
R9562 VPWR.n2331 VPWR.n2330 376.045
R9563 VPWR.n2339 VPWR.n2338 376.045
R9564 VPWR.n2341 VPWR.n2340 376.045
R9565 VPWR.n2349 VPWR.n2348 376.045
R9566 VPWR.n2351 VPWR.n2350 376.045
R9567 VPWR.n2359 VPWR.n2358 376.045
R9568 VPWR.n2361 VPWR.n2360 376.045
R9569 VPWR.n2369 VPWR.n2368 376.045
R9570 VPWR.n2371 VPWR.n2370 376.045
R9571 VPWR.n2379 VPWR.n2378 376.045
R9572 VPWR.n2329 VPWR.n2328 376.045
R9573 VPWR.n543 VPWR.n542 376.045
R9574 VPWR.n541 VPWR.n540 376.045
R9575 VPWR.n537 VPWR.n536 376.045
R9576 VPWR.n533 VPWR.n532 376.045
R9577 VPWR.n525 VPWR.n524 376.045
R9578 VPWR.n521 VPWR.n520 376.045
R9579 VPWR.n517 VPWR.n516 376.045
R9580 VPWR.n513 VPWR.n512 376.045
R9581 VPWR.n509 VPWR.n508 376.045
R9582 VPWR.n505 VPWR.n504 376.045
R9583 VPWR.n501 VPWR.n500 376.045
R9584 VPWR.n497 VPWR.n496 376.045
R9585 VPWR.n493 VPWR.n492 376.045
R9586 VPWR.n489 VPWR.n488 376.045
R9587 VPWR.n529 VPWR.n528 376.045
R9588 VPWR.n2282 VPWR.n2281 376.045
R9589 VPWR.n2280 VPWR.n2279 376.045
R9590 VPWR.n2272 VPWR.n2271 376.045
R9591 VPWR.n2270 VPWR.n2269 376.045
R9592 VPWR.n2260 VPWR.n2259 376.045
R9593 VPWR.n2252 VPWR.n2251 376.045
R9594 VPWR.n2250 VPWR.n2249 376.045
R9595 VPWR.n2242 VPWR.n2241 376.045
R9596 VPWR.n2240 VPWR.n2239 376.045
R9597 VPWR.n2232 VPWR.n2231 376.045
R9598 VPWR.n2230 VPWR.n2229 376.045
R9599 VPWR.n2222 VPWR.n2221 376.045
R9600 VPWR.n2220 VPWR.n2219 376.045
R9601 VPWR.n2212 VPWR.n2211 376.045
R9602 VPWR.n2262 VPWR.n2261 376.045
R9603 VPWR.n582 VPWR.n581 376.045
R9604 VPWR.n586 VPWR.n585 376.045
R9605 VPWR.n590 VPWR.n589 376.045
R9606 VPWR.n594 VPWR.n593 376.045
R9607 VPWR.n602 VPWR.n601 376.045
R9608 VPWR.n606 VPWR.n605 376.045
R9609 VPWR.n610 VPWR.n609 376.045
R9610 VPWR.n614 VPWR.n613 376.045
R9611 VPWR.n618 VPWR.n617 376.045
R9612 VPWR.n622 VPWR.n621 376.045
R9613 VPWR.n626 VPWR.n625 376.045
R9614 VPWR.n630 VPWR.n629 376.045
R9615 VPWR.n634 VPWR.n633 376.045
R9616 VPWR.n638 VPWR.n637 376.045
R9617 VPWR.n598 VPWR.n597 376.045
R9618 VPWR.n2113 VPWR.n2112 376.045
R9619 VPWR.n2115 VPWR.n2114 376.045
R9620 VPWR.n2123 VPWR.n2122 376.045
R9621 VPWR.n2125 VPWR.n2124 376.045
R9622 VPWR.n2135 VPWR.n2134 376.045
R9623 VPWR.n2143 VPWR.n2142 376.045
R9624 VPWR.n2145 VPWR.n2144 376.045
R9625 VPWR.n2153 VPWR.n2152 376.045
R9626 VPWR.n2155 VPWR.n2154 376.045
R9627 VPWR.n2163 VPWR.n2162 376.045
R9628 VPWR.n2165 VPWR.n2164 376.045
R9629 VPWR.n2173 VPWR.n2172 376.045
R9630 VPWR.n2175 VPWR.n2174 376.045
R9631 VPWR.n2183 VPWR.n2182 376.045
R9632 VPWR.n2133 VPWR.n2132 376.045
R9633 VPWR.n735 VPWR.n734 376.045
R9634 VPWR.n733 VPWR.n732 376.045
R9635 VPWR.n729 VPWR.n728 376.045
R9636 VPWR.n725 VPWR.n724 376.045
R9637 VPWR.n717 VPWR.n716 376.045
R9638 VPWR.n713 VPWR.n712 376.045
R9639 VPWR.n709 VPWR.n708 376.045
R9640 VPWR.n705 VPWR.n704 376.045
R9641 VPWR.n701 VPWR.n700 376.045
R9642 VPWR.n697 VPWR.n696 376.045
R9643 VPWR.n693 VPWR.n692 376.045
R9644 VPWR.n689 VPWR.n688 376.045
R9645 VPWR.n685 VPWR.n684 376.045
R9646 VPWR.n681 VPWR.n680 376.045
R9647 VPWR.n721 VPWR.n720 376.045
R9648 VPWR.n2086 VPWR.n2085 376.045
R9649 VPWR.n2084 VPWR.n2083 376.045
R9650 VPWR.n2076 VPWR.n2075 376.045
R9651 VPWR.n2074 VPWR.n2073 376.045
R9652 VPWR.n2064 VPWR.n2063 376.045
R9653 VPWR.n2056 VPWR.n2055 376.045
R9654 VPWR.n2054 VPWR.n2053 376.045
R9655 VPWR.n2046 VPWR.n2045 376.045
R9656 VPWR.n2044 VPWR.n2043 376.045
R9657 VPWR.n2036 VPWR.n2035 376.045
R9658 VPWR.n2034 VPWR.n2033 376.045
R9659 VPWR.n2026 VPWR.n2025 376.045
R9660 VPWR.n2024 VPWR.n2023 376.045
R9661 VPWR.n2016 VPWR.n2015 376.045
R9662 VPWR.n2066 VPWR.n2065 376.045
R9663 VPWR.n774 VPWR.n773 376.045
R9664 VPWR.n778 VPWR.n777 376.045
R9665 VPWR.n782 VPWR.n781 376.045
R9666 VPWR.n786 VPWR.n785 376.045
R9667 VPWR.n794 VPWR.n793 376.045
R9668 VPWR.n798 VPWR.n797 376.045
R9669 VPWR.n802 VPWR.n801 376.045
R9670 VPWR.n806 VPWR.n805 376.045
R9671 VPWR.n810 VPWR.n809 376.045
R9672 VPWR.n814 VPWR.n813 376.045
R9673 VPWR.n818 VPWR.n817 376.045
R9674 VPWR.n822 VPWR.n821 376.045
R9675 VPWR.n826 VPWR.n825 376.045
R9676 VPWR.n830 VPWR.n829 376.045
R9677 VPWR.n790 VPWR.n789 376.045
R9678 VPWR.n1917 VPWR.n1916 376.045
R9679 VPWR.n1919 VPWR.n1918 376.045
R9680 VPWR.n1927 VPWR.n1926 376.045
R9681 VPWR.n1929 VPWR.n1928 376.045
R9682 VPWR.n1939 VPWR.n1938 376.045
R9683 VPWR.n1947 VPWR.n1946 376.045
R9684 VPWR.n1949 VPWR.n1948 376.045
R9685 VPWR.n1957 VPWR.n1956 376.045
R9686 VPWR.n1959 VPWR.n1958 376.045
R9687 VPWR.n1967 VPWR.n1966 376.045
R9688 VPWR.n1969 VPWR.n1968 376.045
R9689 VPWR.n1977 VPWR.n1976 376.045
R9690 VPWR.n1979 VPWR.n1978 376.045
R9691 VPWR.n1987 VPWR.n1986 376.045
R9692 VPWR.n1937 VPWR.n1936 376.045
R9693 VPWR.n927 VPWR.n926 376.045
R9694 VPWR.n925 VPWR.n924 376.045
R9695 VPWR.n921 VPWR.n920 376.045
R9696 VPWR.n917 VPWR.n916 376.045
R9697 VPWR.n909 VPWR.n908 376.045
R9698 VPWR.n905 VPWR.n904 376.045
R9699 VPWR.n901 VPWR.n900 376.045
R9700 VPWR.n897 VPWR.n896 376.045
R9701 VPWR.n893 VPWR.n892 376.045
R9702 VPWR.n889 VPWR.n888 376.045
R9703 VPWR.n885 VPWR.n884 376.045
R9704 VPWR.n881 VPWR.n880 376.045
R9705 VPWR.n877 VPWR.n876 376.045
R9706 VPWR.n873 VPWR.n872 376.045
R9707 VPWR.n913 VPWR.n912 376.045
R9708 VPWR.n1870 VPWR.n1869 376.045
R9709 VPWR.n982 VPWR.n981 376.045
R9710 VPWR.n1494 VPWR.n1493 376.045
R9711 VPWR.n1221 VPWR.n1220 376.045
R9712 VPWR.n402 VPWR.n401 376.045
R9713 VPWR.n2466 VPWR.n2465 376.045
R9714 VPWR.n341 VPWR.n340 376.045
R9715 VPWR.n2520 VPWR.n2519 376.045
R9716 VPWR.n978 VPWR.n977 376.045
R9717 VPWR.n1492 VPWR.n1491 376.045
R9718 VPWR.n1185 VPWR.n1184 376.045
R9719 VPWR.n1868 VPWR.n1867 376.045
R9720 VPWR.n986 VPWR.n985 376.045
R9721 VPWR.n1506 VPWR.n1505 376.045
R9722 VPWR.n1219 VPWR.n1218 376.045
R9723 VPWR.n410 VPWR.n409 376.045
R9724 VPWR.n418 VPWR.n417 376.045
R9725 VPWR.n422 VPWR.n421 376.045
R9726 VPWR.n426 VPWR.n425 376.045
R9727 VPWR.n430 VPWR.n429 376.045
R9728 VPWR.n434 VPWR.n433 376.045
R9729 VPWR.n438 VPWR.n437 376.045
R9730 VPWR.n442 VPWR.n441 376.045
R9731 VPWR.n446 VPWR.n445 376.045
R9732 VPWR.n414 VPWR.n413 376.045
R9733 VPWR.n2448 VPWR.n2447 376.045
R9734 VPWR.n329 VPWR.n328 376.045
R9735 VPWR.n2542 VPWR.n2541 376.045
R9736 VPWR.n990 VPWR.n989 376.045
R9737 VPWR.n1508 VPWR.n1507 376.045
R9738 VPWR.n1216 VPWR.n1215 376.045
R9739 VPWR.n1860 VPWR.n1859 376.045
R9740 VPWR.n1850 VPWR.n1849 376.045
R9741 VPWR.n1848 VPWR.n1847 376.045
R9742 VPWR.n1840 VPWR.n1839 376.045
R9743 VPWR.n1838 VPWR.n1837 376.045
R9744 VPWR.n1830 VPWR.n1829 376.045
R9745 VPWR.n1828 VPWR.n1827 376.045
R9746 VPWR.n1820 VPWR.n1819 376.045
R9747 VPWR.n1858 VPWR.n1857 376.045
R9748 VPWR.n994 VPWR.n993 376.045
R9749 VPWR.n1520 VPWR.n1519 376.045
R9750 VPWR.n1213 VPWR.n1212 376.045
R9751 VPWR.n2468 VPWR.n2467 376.045
R9752 VPWR.n345 VPWR.n344 376.045
R9753 VPWR.n2518 VPWR.n2517 376.045
R9754 VPWR.n1481 VPWR.n1480 376.045
R9755 VPWR.n1182 VPWR.n1181 376.045
R9756 VPWR.n998 VPWR.n997 376.045
R9757 VPWR.n1522 VPWR.n1521 376.045
R9758 VPWR.n1205 VPWR.n1204 376.045
R9759 VPWR.n2438 VPWR.n2437 376.045
R9760 VPWR.n2428 VPWR.n2427 376.045
R9761 VPWR.n2426 VPWR.n2425 376.045
R9762 VPWR.n2418 VPWR.n2417 376.045
R9763 VPWR.n2416 VPWR.n2415 376.045
R9764 VPWR.n2408 VPWR.n2407 376.045
R9765 VPWR.n2436 VPWR.n2435 376.045
R9766 VPWR.n317 VPWR.n316 376.045
R9767 VPWR.n2556 VPWR.n2555 376.045
R9768 VPWR.n1537 VPWR.n1536 376.045
R9769 VPWR.n1202 VPWR.n1201 376.045
R9770 VPWR.n1002 VPWR.n1001 376.045
R9771 VPWR.n1006 VPWR.n1005 376.045
R9772 VPWR.n1010 VPWR.n1009 376.045
R9773 VPWR.n1014 VPWR.n1013 376.045
R9774 VPWR.n1018 VPWR.n1017 376.045
R9775 VPWR.n1022 VPWR.n1021 376.045
R9776 VPWR.n970 VPWR.n969 376.045
R9777 VPWR.n1475 VPWR.n1474 376.045
R9778 VPWR.n1593 VPWR.n1592 376.045
R9779 VPWR.n313 VPWR.n312 376.045
R9780 VPWR.n2566 VPWR.n2565 376.045
R9781 VPWR.n1199 VPWR.n1198 376.045
R9782 VPWR.n1762 VPWR.n1761 376.045
R9783 VPWR.n1191 VPWR.n1190 376.045
R9784 VPWR.n309 VPWR.n308 376.045
R9785 VPWR.n305 VPWR.n304 376.045
R9786 VPWR.n297 VPWR.n296 376.045
R9787 VPWR.n301 VPWR.n300 376.045
R9788 VPWR.n1741 VPWR.n1740 376.045
R9789 VPWR.n1750 VPWR.n1749 376.045
R9790 VPWR.n1791 VPWR.n1790 376.045
R9791 VPWR.n1760 VPWR.n1759 376.045
R9792 VPWR.n1188 VPWR.n1187 376.045
R9793 VPWR.n2578 VPWR.n2577 376.045
R9794 VPWR.n2580 VPWR.n2579 376.045
R9795 VPWR.n2590 VPWR.n2589 376.045
R9796 VPWR.n1739 VPWR.n1738 376.045
R9797 VPWR.n1339 VPWR.t648 342.841
R9798 VPWR.n1378 VPWR.t1265 342.841
R9799 VPWR.n1415 VPWR.t657 342.841
R9800 VPWR.n2693 VPWR.t1143 342.841
R9801 VPWR.n2656 VPWR.t964 342.841
R9802 VPWR.n2599 VPWR.t805 342.841
R9803 VPWR.n1339 VPWR.t403 342.839
R9804 VPWR.n1378 VPWR.t934 342.839
R9805 VPWR.n1415 VPWR.t390 342.839
R9806 VPWR.n2693 VPWR.t1904 342.839
R9807 VPWR.n2656 VPWR.t1400 342.839
R9808 VPWR.n2599 VPWR.t1135 342.839
R9809 VPWR.n2842 VPWR.n2824 339.212
R9810 VPWR.n1306 VPWR.t440 338.488
R9811 VPWR.n2729 VPWR.t1113 338.488
R9812 VPWR.n1315 VPWR.n1314 327.377
R9813 VPWR.n1308 VPWR.n1307 327.377
R9814 VPWR.n1322 VPWR.n1321 327.377
R9815 VPWR.n1352 VPWR.n1350 327.377
R9816 VPWR.n1345 VPWR.n1343 327.377
R9817 VPWR.n1360 VPWR.n1358 327.377
R9818 VPWR.n1391 VPWR.n1389 327.377
R9819 VPWR.n1384 VPWR.n1382 327.377
R9820 VPWR.n1399 VPWR.n1397 327.377
R9821 VPWR.n1428 VPWR.n1426 327.377
R9822 VPWR.n1421 VPWR.n1419 327.377
R9823 VPWR.n1436 VPWR.n1434 327.377
R9824 VPWR.n1324 VPWR.n1323 327.375
R9825 VPWR.n1352 VPWR.n1351 327.375
R9826 VPWR.n1345 VPWR.n1344 327.375
R9827 VPWR.n1360 VPWR.n1359 327.375
R9828 VPWR.n1391 VPWR.n1390 327.375
R9829 VPWR.n1384 VPWR.n1383 327.375
R9830 VPWR.n1399 VPWR.n1398 327.375
R9831 VPWR.n1428 VPWR.n1427 327.375
R9832 VPWR.n1421 VPWR.n1420 327.375
R9833 VPWR.n1436 VPWR.n1435 327.375
R9834 VPWR.n1 VPWR 325.546
R9835 VPWR.n2667 VPWR.t1142 322.262
R9836 VPWR.n2630 VPWR.t963 322.262
R9837 VPWR.n2805 VPWR.n2804 321.642
R9838 VPWR.n2722 VPWR.n2712 320.976
R9839 VPWR.n2716 VPWR.n2715 320.976
R9840 VPWR.n2710 VPWR.n2709 320.976
R9841 VPWR.n2680 VPWR.n2679 320.976
R9842 VPWR.n2686 VPWR.n2675 320.976
R9843 VPWR.n2672 VPWR.n2671 320.976
R9844 VPWR.n2643 VPWR.n2642 320.976
R9845 VPWR.n2649 VPWR.n2638 320.976
R9846 VPWR.n2635 VPWR.n2634 320.976
R9847 VPWR.n2610 VPWR.n2606 320.976
R9848 VPWR.n2614 VPWR.n2613 320.976
R9849 VPWR.n2620 VPWR.n2602 320.976
R9850 VPWR.n2727 VPWR.n2708 320.976
R9851 VPWR.n2680 VPWR.n2678 320.976
R9852 VPWR.n2686 VPWR.n2674 320.976
R9853 VPWR.n2672 VPWR.n2670 320.976
R9854 VPWR.n2643 VPWR.n2641 320.976
R9855 VPWR.n2649 VPWR.n2637 320.976
R9856 VPWR.n2635 VPWR.n2633 320.976
R9857 VPWR.n2610 VPWR.n2605 320.976
R9858 VPWR.n2614 VPWR.n2612 320.976
R9859 VPWR.n2620 VPWR.n2601 320.976
R9860 VPWR.n2801 VPWR 319.627
R9861 VPWR.n6 VPWR.n5 316.245
R9862 VPWR.n1241 VPWR.n1239 316.245
R9863 VPWR.n1264 VPWR.n1262 316.245
R9864 VPWR.n1288 VPWR.n1286 316.245
R9865 VPWR.n2784 VPWR.n2783 316.245
R9866 VPWR.n2764 VPWR.n2763 316.245
R9867 VPWR.n2745 VPWR.n2744 316.245
R9868 VPWR.n1241 VPWR.n1240 316.245
R9869 VPWR.n1264 VPWR.n1263 316.245
R9870 VPWR.n1288 VPWR.n1287 316.245
R9871 VPWR.n2784 VPWR.n2782 316.245
R9872 VPWR.n2764 VPWR.n2762 316.245
R9873 VPWR.n2745 VPWR.n2743 316.245
R9874 VPWR.n2630 VPWR.t514 313.87
R9875 VPWR.n10 VPWR.n4 310.502
R9876 VPWR.n1246 VPWR.n1238 310.502
R9877 VPWR.n1269 VPWR.n1261 310.502
R9878 VPWR.n1293 VPWR.n1285 310.502
R9879 VPWR.n2803 VPWR.n2802 310.502
R9880 VPWR.n2788 VPWR.n2787 310.502
R9881 VPWR.n2768 VPWR.n2767 310.502
R9882 VPWR.n2749 VPWR.n2748 310.502
R9883 VPWR.n1246 VPWR.n1245 310.5
R9884 VPWR.n1269 VPWR.n1268 310.5
R9885 VPWR.n1293 VPWR.n1292 310.5
R9886 VPWR.n2788 VPWR.n2786 310.5
R9887 VPWR.n2768 VPWR.n2766 310.5
R9888 VPWR.n2749 VPWR.n2747 310.5
R9889 VPWR.n2834 VPWR.n2833 279.341
R9890 VPWR.n2839 VPWR.n2838 279.341
R9891 VPWR.n1412 VPWR.t367 255.905
R9892 VPWR.n2663 VPWR.t515 255.905
R9893 VPWR.n1275 VPWR.t562 255.904
R9894 VPWR.n1412 VPWR.t1284 255.904
R9895 VPWR.n2774 VPWR.t1408 255.904
R9896 VPWR.n2663 VPWR.t628 255.904
R9897 VPWR.n1303 VPWR.t1253 254.019
R9898 VPWR.n2735 VPWR.t997 254.019
R9899 VPWR.n1335 VPWR.t1251 252.948
R9900 VPWR.n2737 VPWR.t995 252.948
R9901 VPWR.n1373 VPWR.t714 250.722
R9902 VPWR.n2700 VPWR.t1283 250.722
R9903 VPWR.n1310 VPWR.t836 249.901
R9904 VPWR.n1346 VPWR.t847 249.901
R9905 VPWR.n1385 VPWR.t75 249.901
R9906 VPWR.n1422 VPWR.t849 249.901
R9907 VPWR.n2714 VPWR.t1924 249.901
R9908 VPWR.n2677 VPWR.t878 249.901
R9909 VPWR.n2640 VPWR.t85 249.901
R9910 VPWR.n2607 VPWR.t1844 249.901
R9911 VPWR.n1346 VPWR.t1313 249.901
R9912 VPWR.n1385 VPWR.t45 249.901
R9913 VPWR.n1422 VPWR.t601 249.901
R9914 VPWR.n2677 VPWR.t87 249.901
R9915 VPWR.n2640 VPWR.t1845 249.901
R9916 VPWR.n2607 VPWR.t924 249.901
R9917 VPWR.n1253 VPWR.t1154 249.363
R9918 VPWR.n1338 VPWR.t717 249.363
R9919 VPWR.n2811 VPWR.t26 249.363
R9920 VPWR.n2795 VPWR.t1916 249.363
R9921 VPWR.n2698 VPWR.t564 249.363
R9922 VPWR.n17 VPWR.t464 249.362
R9923 VPWR.n1253 VPWR.t715 249.362
R9924 VPWR.n2795 VPWR.t32 249.362
R9925 VPWR.t557 VPWR.t463 248.599
R9926 VPWR.t437 VPWR.t784 248.599
R9927 VPWR.t784 VPWR.t788 248.599
R9928 VPWR.t788 VPWR.t1295 248.599
R9929 VPWR.t1295 VPWR.t1240 248.599
R9930 VPWR.t1240 VPWR.t831 248.599
R9931 VPWR.t831 VPWR.t846 248.599
R9932 VPWR.t846 VPWR.t851 248.599
R9933 VPWR.t1309 VPWR.t1311 248.599
R9934 VPWR.t1311 VPWR.t835 248.599
R9935 VPWR.t81 VPWR.t887 248.599
R9936 VPWR.t912 VPWR.t81 248.599
R9937 VPWR.t1325 VPWR.t912 248.599
R9938 VPWR.t1110 VPWR.t1325 248.599
R9939 VPWR.t869 VPWR.t1110 248.599
R9940 VPWR.t1065 VPWR.t869 248.599
R9941 VPWR.t1063 VPWR.t1065 248.599
R9942 VPWR.t1409 VPWR.t25 248.599
R9943 VPWR.t14 VPWR.t1923 248.599
R9944 VPWR.t1919 VPWR.t14 248.599
R9945 VPWR.n15 VPWR.t558 247.394
R9946 VPWR.n1251 VPWR.t560 247.394
R9947 VPWR.n2809 VPWR.t1410 247.394
R9948 VPWR.n2793 VPWR.t1404 247.394
R9949 VPWR.n1251 VPWR.t559 247.394
R9950 VPWR.n2793 VPWR.t1406 247.394
R9951 VPWR.n1304 VPWR.t36 244.737
R9952 VPWR.n2730 VPWR.t1831 244.737
R9953 VPWR.n1374 VPWR.t1909 243.886
R9954 VPWR.n2701 VPWR.t461 243.886
R9955 VPWR.n1277 VPWR.t462 243.512
R9956 VPWR.n1300 VPWR.t1155 243.512
R9957 VPWR.n1303 VPWR.t650 243.512
R9958 VPWR.n2776 VPWR.t28 243.512
R9959 VPWR.n2756 VPWR.t1917 243.512
R9960 VPWR.n2735 VPWR.t822 243.512
R9961 VPWR.n1300 VPWR.t716 243.512
R9962 VPWR.n2756 VPWR.t30 243.512
R9963 VPWR.n1329 VPWR.t1252 238.339
R9964 VPWR.n2705 VPWR.t996 238.339
R9965 VPWR.n2855 VPWR.t516 237.99
R9966 VPWR.n2667 VPWR.t563 234.982
R9967 VPWR.t1307 VPWR.t1309 228.101
R9968 VPWR.t928 VPWR.t1919 228.101
R9969 VPWR.n2801 VPWR 224.923
R9970 VPWR.n1 VPWR 219.004
R9971 VPWR.n1444 VPWR.n1443 214.613
R9972 VPWR.n1444 VPWR.n1442 214.613
R9973 VPWR.n1236 VPWR.n1235 214.326
R9974 VPWR.n1259 VPWR.n1258 214.326
R9975 VPWR.n1283 VPWR.n1282 214.326
R9976 VPWR.n1368 VPWR.n1367 214.326
R9977 VPWR.n1407 VPWR.n1406 214.326
R9978 VPWR.n1236 VPWR.n1234 214.326
R9979 VPWR.n1259 VPWR.n1257 214.326
R9980 VPWR.n1283 VPWR.n1281 214.326
R9981 VPWR.n1368 VPWR.n1366 214.326
R9982 VPWR.n1407 VPWR.n1405 214.326
R9983 VPWR.n2 VPWR.n1 213.119
R9984 VPWR.n2808 VPWR.n2801 213.119
R9985 VPWR VPWR.t557 207.166
R9986 VPWR.n2840 VPWR.n2839 204.424
R9987 VPWR.n2830 VPWR.n2817 204.424
R9988 VPWR.n2833 VPWR.n2820 204.424
R9989 VPWR.n2844 VPWR.n2841 204.048
R9990 VPWR VPWR.t1063 201.246
R9991 VPWR.t835 VPWR 189.409
R9992 VPWR.n2741 VPWR 184.63
R9993 VPWR.n1329 VPWR 182.952
R9994 VPWR.n2760 VPWR 182.952
R9995 VPWR.n2780 VPWR 181.273
R9996 VPWR.t514 VPWR 177.916
R9997 VPWR.n2848 VPWR.n2847 166.4
R9998 VPWR.n1770 VPWR.n1768 161.365
R9999 VPWR.n1041 VPWR.n1039 161.365
R10000 VPWR.n1545 VPWR.n1543 161.365
R10001 VPWR.n1550 VPWR.n1548 161.365
R10002 VPWR.n1555 VPWR.n1553 161.365
R10003 VPWR.n1560 VPWR.n1558 161.365
R10004 VPWR.n1565 VPWR.n1563 161.365
R10005 VPWR.n1570 VPWR.n1568 161.365
R10006 VPWR.n1575 VPWR.n1573 161.365
R10007 VPWR.n1580 VPWR.n1578 161.365
R10008 VPWR.n1135 VPWR.n1133 161.365
R10009 VPWR.n1460 VPWR.n1458 161.365
R10010 VPWR.n1455 VPWR.n1453 161.365
R10011 VPWR.n1775 VPWR.n1773 161.365
R10012 VPWR.n1783 VPWR.n1781 161.365
R10013 VPWR.n1779 VPWR.n1777 161.365
R10014 VPWR VPWR.n53 161.363
R10015 VPWR VPWR.n51 161.363
R10016 VPWR VPWR.n49 161.363
R10017 VPWR VPWR.n47 161.363
R10018 VPWR VPWR.n45 161.363
R10019 VPWR VPWR.n43 161.363
R10020 VPWR VPWR.n41 161.363
R10021 VPWR VPWR.n39 161.363
R10022 VPWR VPWR.n37 161.363
R10023 VPWR VPWR.n35 161.363
R10024 VPWR VPWR.n33 161.363
R10025 VPWR VPWR.n31 161.363
R10026 VPWR VPWR.n29 161.363
R10027 VPWR VPWR.n27 161.363
R10028 VPWR VPWR.n25 161.363
R10029 VPWR VPWR.n23 161.363
R10030 VPWR.n1115 VPWR.n1114 161.303
R10031 VPWR.n107 VPWR.n106 161.303
R10032 VPWR.n1120 VPWR.n1119 161.3
R10033 VPWR.n1599 VPWR.n1598 161.3
R10034 VPWR.n1602 VPWR.n1601 161.3
R10035 VPWR.n1111 VPWR.n1110 161.3
R10036 VPWR.n1126 VPWR.n1125 161.3
R10037 VPWR.n1107 VPWR.n1106 161.3
R10038 VPWR.n1612 VPWR.n1611 161.3
R10039 VPWR.n1615 VPWR.n1614 161.3
R10040 VPWR.n1618 VPWR.n1617 161.3
R10041 VPWR.n1623 VPWR.n1622 161.3
R10042 VPWR.n1626 VPWR.n1625 161.3
R10043 VPWR.n1629 VPWR.n1628 161.3
R10044 VPWR.n1101 VPWR.n1100 161.3
R10045 VPWR.n1177 VPWR.n1176 161.3
R10046 VPWR.n1097 VPWR.n1096 161.3
R10047 VPWR.n1639 VPWR.n1638 161.3
R10048 VPWR.n1642 VPWR.n1641 161.3
R10049 VPWR.n1645 VPWR.n1644 161.3
R10050 VPWR.n1650 VPWR.n1649 161.3
R10051 VPWR.n1653 VPWR.n1652 161.3
R10052 VPWR.n1656 VPWR.n1655 161.3
R10053 VPWR.n1091 VPWR.n1090 161.3
R10054 VPWR.n1209 VPWR.n1208 161.3
R10055 VPWR.n1087 VPWR.n1086 161.3
R10056 VPWR.n1666 VPWR.n1665 161.3
R10057 VPWR.n1669 VPWR.n1668 161.3
R10058 VPWR.n1672 VPWR.n1671 161.3
R10059 VPWR.n1677 VPWR.n1676 161.3
R10060 VPWR.n1680 VPWR.n1679 161.3
R10061 VPWR.n1683 VPWR.n1682 161.3
R10062 VPWR.n1081 VPWR.n1080 161.3
R10063 VPWR.n1195 VPWR.n1194 161.3
R10064 VPWR.n1077 VPWR.n1076 161.3
R10065 VPWR.n1693 VPWR.n1692 161.3
R10066 VPWR.n1696 VPWR.n1695 161.3
R10067 VPWR.n1699 VPWR.n1698 161.3
R10068 VPWR.n1704 VPWR.n1703 161.3
R10069 VPWR.n1707 VPWR.n1706 161.3
R10070 VPWR.n1710 VPWR.n1709 161.3
R10071 VPWR.n1070 VPWR.n1069 161.3
R10072 VPWR.n1719 VPWR.n1718 161.3
R10073 VPWR.n1722 VPWR.n1721 161.3
R10074 VPWR.n1717 VPWR.n1716 161.3
R10075 VPWR.n1734 VPWR.n1733 161.3
R10076 VPWR.n1117 VPWR.n1116 161.3
R10077 VPWR.n1731 VPWR.n1730 161.3
R10078 VPWR.n1065 VPWR.n1064 161.3
R10079 VPWR.n126 VPWR.n125 161.3
R10080 VPWR.n117 VPWR.n116 161.3
R10081 VPWR.n120 VPWR.n119 161.3
R10082 VPWR.n115 VPWR.n114 161.3
R10083 VPWR.n138 VPWR.n137 161.3
R10084 VPWR.n128 VPWR.n127 161.3
R10085 VPWR.n109 VPWR.n108 161.3
R10086 VPWR.n105 VPWR.n104 161.3
R10087 VPWR.n288 VPWR.n287 161.3
R10088 VPWR.n285 VPWR.n284 161.3
R10089 VPWR.n101 VPWR.n100 161.3
R10090 VPWR.n272 VPWR.n271 161.3
R10091 VPWR.n275 VPWR.n274 161.3
R10092 VPWR.n270 VPWR.n269 161.3
R10093 VPWR.n260 VPWR.n259 161.3
R10094 VPWR.n263 VPWR.n262 161.3
R10095 VPWR.n258 VPWR.n257 161.3
R10096 VPWR.n248 VPWR.n247 161.3
R10097 VPWR.n251 VPWR.n250 161.3
R10098 VPWR.n246 VPWR.n245 161.3
R10099 VPWR.n236 VPWR.n235 161.3
R10100 VPWR.n239 VPWR.n238 161.3
R10101 VPWR.n234 VPWR.n233 161.3
R10102 VPWR.n224 VPWR.n223 161.3
R10103 VPWR.n227 VPWR.n226 161.3
R10104 VPWR.n222 VPWR.n221 161.3
R10105 VPWR.n212 VPWR.n211 161.3
R10106 VPWR.n215 VPWR.n214 161.3
R10107 VPWR.n210 VPWR.n209 161.3
R10108 VPWR.n200 VPWR.n199 161.3
R10109 VPWR.n203 VPWR.n202 161.3
R10110 VPWR.n198 VPWR.n197 161.3
R10111 VPWR.n188 VPWR.n187 161.3
R10112 VPWR.n191 VPWR.n190 161.3
R10113 VPWR.n186 VPWR.n185 161.3
R10114 VPWR.n176 VPWR.n175 161.3
R10115 VPWR.n179 VPWR.n178 161.3
R10116 VPWR.n174 VPWR.n173 161.3
R10117 VPWR.n164 VPWR.n163 161.3
R10118 VPWR.n167 VPWR.n166 161.3
R10119 VPWR.n162 VPWR.n161 161.3
R10120 VPWR.n152 VPWR.n151 161.3
R10121 VPWR.n155 VPWR.n154 161.3
R10122 VPWR.n150 VPWR.n149 161.3
R10123 VPWR.n140 VPWR.n139 161.3
R10124 VPWR.n143 VPWR.n142 161.3
R10125 VPWR.n131 VPWR.n130 161.3
R10126 VPWR.n1601 VPWR.t1455 161.202
R10127 VPWR.n1106 VPWR.t1583 161.202
R10128 VPWR.n1617 VPWR.t1624 161.202
R10129 VPWR.n1628 VPWR.t1732 161.202
R10130 VPWR.n1096 VPWR.t1499 161.202
R10131 VPWR.n1644 VPWR.t1514 161.202
R10132 VPWR.n1655 VPWR.t1737 161.202
R10133 VPWR.n1086 VPWR.t1780 161.202
R10134 VPWR.n1671 VPWR.t1497 161.202
R10135 VPWR.n1682 VPWR.t1650 161.202
R10136 VPWR.n1076 VPWR.t1672 161.202
R10137 VPWR.n1698 VPWR.t1522 161.202
R10138 VPWR.n1709 VPWR.t1548 161.202
R10139 VPWR.n1721 VPWR.t1573 161.202
R10140 VPWR.n1116 VPWR.t1713 161.202
R10141 VPWR.n1730 VPWR.t1418 161.202
R10142 VPWR.n119 VPWR.t1540 161.202
R10143 VPWR.n108 VPWR.t1439 161.202
R10144 VPWR.n284 VPWR.t1575 161.202
R10145 VPWR.n274 VPWR.t1705 161.202
R10146 VPWR.n262 VPWR.t1745 161.202
R10147 VPWR.n250 VPWR.t1469 161.202
R10148 VPWR.n238 VPWR.t1613 161.202
R10149 VPWR.n226 VPWR.t1637 161.202
R10150 VPWR.n214 VPWR.t1474 161.202
R10151 VPWR.n202 VPWR.t1509 161.202
R10152 VPWR.n190 VPWR.t1611 161.202
R10153 VPWR.n178 VPWR.t1772 161.202
R10154 VPWR.n166 VPWR.t1791 161.202
R10155 VPWR.n154 VPWR.t1645 161.202
R10156 VPWR.n1768 VPWR.t1697 161.202
R10157 VPWR.n1039 VPWR.t1450 161.202
R10158 VPWR.n1543 VPWR.t1434 161.202
R10159 VPWR.n1548 VPWR.t1683 161.202
R10160 VPWR.n1553 VPWR.t1565 161.202
R10161 VPWR.n1558 VPWR.t1535 161.202
R10162 VPWR.n1563 VPWR.t1687 161.202
R10163 VPWR.n1568 VPWR.t1685 161.202
R10164 VPWR.n1573 VPWR.t1530 161.202
R10165 VPWR.n1578 VPWR.t1420 161.202
R10166 VPWR.n1133 VPWR.t1764 161.202
R10167 VPWR.n1458 VPWR.t1635 161.202
R10168 VPWR.n1453 VPWR.t1504 161.202
R10169 VPWR.n1773 VPWR.t1715 161.202
R10170 VPWR.n1781 VPWR.t1753 161.202
R10171 VPWR.n1777 VPWR.t1585 161.202
R10172 VPWR.n142 VPWR.t1664 161.202
R10173 VPWR.n130 VPWR.t1689 161.202
R10174 VPWR.n1119 VPWR.t1441 161.106
R10175 VPWR.n1110 VPWR.t1577 161.106
R10176 VPWR.n1611 VPWR.t1590 161.106
R10177 VPWR.n1622 VPWR.t1750 161.106
R10178 VPWR.n1100 VPWR.t1471 161.106
R10179 VPWR.n1638 VPWR.t1618 161.106
R10180 VPWR.n1649 VPWR.t1726 161.106
R10181 VPWR.n1090 VPWR.t1766 161.106
R10182 VPWR.n1665 VPWR.t1511 161.106
R10183 VPWR.n1676 VPWR.t1615 161.106
R10184 VPWR.n1080 VPWR.t1774 161.106
R10185 VPWR.n1692 VPWR.t1793 161.106
R10186 VPWR.n1703 VPWR.t1537 161.106
R10187 VPWR.n1069 VPWR.t1666 161.106
R10188 VPWR.n1716 VPWR.t1694 161.106
R10189 VPWR.n1064 VPWR.t1545 161.106
R10190 VPWR.n125 VPWR.t1425 161.106
R10191 VPWR.n114 VPWR.t1661 161.106
R10192 VPWR.n137 VPWR.t1785 161.106
R10193 VPWR.n104 VPWR.t1570 161.106
R10194 VPWR.n100 VPWR.t1699 161.106
R10195 VPWR.n269 VPWR.t1717 161.106
R10196 VPWR.n257 VPWR.t1479 161.106
R10197 VPWR.n245 VPWR.t1587 161.106
R10198 VPWR.n233 VPWR.t1742 161.106
R10199 VPWR.n221 VPWR.t1466 161.106
R10200 VPWR.n209 VPWR.t1501 161.106
R10201 VPWR.n197 VPWR.t1629 161.106
R10202 VPWR.n185 VPWR.t1739 161.106
R10203 VPWR.n173 VPWR.t1506 161.106
R10204 VPWR.n161 VPWR.t1524 161.106
R10205 VPWR.n149 VPWR.t1652 161.106
R10206 VPWR.n53 VPWR.t1769 161.106
R10207 VPWR.n51 VPWR.t1729 161.106
R10208 VPWR.n49 VPWR.t1444 161.106
R10209 VPWR.n47 VPWR.t1559 161.106
R10210 VPWR.n45 VPWR.t1777 161.106
R10211 VPWR.n43 VPWR.t1626 161.106
R10212 VPWR.n41 VPWR.t1734 161.106
R10213 VPWR.n39 VPWR.t1460 161.106
R10214 VPWR.n37 VPWR.t1567 161.106
R10215 VPWR.n35 VPWR.t1527 161.106
R10216 VPWR.n33 VPWR.t1632 161.106
R10217 VPWR.n31 VPWR.t1452 161.106
R10218 VPWR.n29 VPWR.t1639 161.106
R10219 VPWR.n27 VPWR.t1747 161.106
R10220 VPWR.n25 VPWR.t1599 161.106
R10221 VPWR.n23 VPWR.t1710 161.106
R10222 VPWR.n1598 VPWR.t1491 159.978
R10223 VPWR.n1125 VPWR.t1596 159.978
R10224 VPWR.n1614 VPWR.t1758 159.978
R10225 VPWR.n1625 VPWR.t1476 159.978
R10226 VPWR.n1176 VPWR.t1488 159.978
R10227 VPWR.n1641 VPWR.t1647 159.978
R10228 VPWR.n1652 VPWR.t1755 159.978
R10229 VPWR.n1208 VPWR.t1516 159.978
R10230 VPWR.n1668 VPWR.t1542 159.978
R10231 VPWR.n1679 VPWR.t1669 159.978
R10232 VPWR.n1194 VPWR.t1415 159.978
R10233 VPWR.n1695 VPWR.t1436 159.978
R10234 VPWR.n1706 VPWR.t1674 159.978
R10235 VPWR.n1718 VPWR.t1702 159.978
R10236 VPWR.n1733 VPWR.t1422 159.978
R10237 VPWR.n1114 VPWR.t1723 159.978
R10238 VPWR.n116 VPWR.t1556 159.978
R10239 VPWR.n127 VPWR.t1431 159.978
R10240 VPWR.n106 VPWR.t1463 159.978
R10241 VPWR.n287 VPWR.t1608 159.978
R10242 VPWR.n271 VPWR.t1720 159.978
R10243 VPWR.n259 VPWR.t1485 159.978
R10244 VPWR.n247 VPWR.t1593 159.978
R10245 VPWR.n235 VPWR.t1605 159.978
R10246 VPWR.n223 VPWR.t1761 159.978
R10247 VPWR.n211 VPWR.t1482 159.978
R10248 VPWR.n199 VPWR.t1642 159.978
R10249 VPWR.n187 VPWR.t1658 159.978
R10250 VPWR.n175 VPWR.t1788 159.978
R10251 VPWR.n163 VPWR.t1532 159.978
R10252 VPWR.n151 VPWR.t1562 159.978
R10253 VPWR.n1228 VPWR.t1519 159.978
R10254 VPWR.n1150 VPWR.t1447 159.978
R10255 VPWR.n1224 VPWR.t1655 159.978
R10256 VPWR.n1482 VPWR.t1553 159.978
R10257 VPWR.n1170 VPWR.t1677 159.978
R10258 VPWR.n1166 VPWR.t1428 159.978
R10259 VPWR.n1160 VPWR.t1550 159.978
R10260 VPWR.n1476 VPWR.t1782 159.978
R10261 VPWR.n1156 VPWR.t1691 159.978
R10262 VPWR.n1146 VPWR.t1707 159.978
R10263 VPWR.n1469 VPWR.t1680 159.978
R10264 VPWR.n1046 VPWR.t1580 159.978
R10265 VPWR.n1745 VPWR.t1457 159.978
R10266 VPWR.n1033 VPWR.t1494 159.978
R10267 VPWR.n1029 VPWR.t1602 159.978
R10268 VPWR.n1050 VPWR.t1621 159.978
R10269 VPWR.n139 VPWR.t1412 159.978
R10270 VPWR.n1229 VPWR.n1228 152
R10271 VPWR.n1151 VPWR.n1150 152
R10272 VPWR.n1225 VPWR.n1224 152
R10273 VPWR.n1483 VPWR.n1482 152
R10274 VPWR.n1171 VPWR.n1170 152
R10275 VPWR.n1167 VPWR.n1166 152
R10276 VPWR.n1161 VPWR.n1160 152
R10277 VPWR.n1477 VPWR.n1476 152
R10278 VPWR.n1157 VPWR.n1156 152
R10279 VPWR.n1147 VPWR.n1146 152
R10280 VPWR.n1470 VPWR.n1469 152
R10281 VPWR.n1047 VPWR.n1046 152
R10282 VPWR.n1746 VPWR.n1745 152
R10283 VPWR.n1034 VPWR.n1033 152
R10284 VPWR.n1030 VPWR.n1029 152
R10285 VPWR.n1051 VPWR.n1050 152
R10286 VPWR.n2845 VPWR.n2844 150.213
R10287 VPWR.n1601 VPWR.t2063 145.137
R10288 VPWR.n1106 VPWR.t2014 145.137
R10289 VPWR.n1617 VPWR.t2000 145.137
R10290 VPWR.n1628 VPWR.t1962 145.137
R10291 VPWR.n1096 VPWR.t2049 145.137
R10292 VPWR.n1644 VPWR.t2042 145.137
R10293 VPWR.n1655 VPWR.t1959 145.137
R10294 VPWR.n1086 VPWR.t1945 145.137
R10295 VPWR.n1671 VPWR.t2050 145.137
R10296 VPWR.n1682 VPWR.t1993 145.137
R10297 VPWR.n1076 VPWR.t1988 145.137
R10298 VPWR.n1698 VPWR.t2040 145.137
R10299 VPWR.n1709 VPWR.t2033 145.137
R10300 VPWR.n1721 VPWR.t2019 145.137
R10301 VPWR.n1116 VPWR.t1969 145.137
R10302 VPWR.n1730 VPWR.t1937 145.137
R10303 VPWR.n119 VPWR.t2048 145.137
R10304 VPWR.n108 VPWR.t1934 145.137
R10305 VPWR.n284 VPWR.t2030 145.137
R10306 VPWR.n274 VPWR.t1983 145.137
R10307 VPWR.n262 VPWR.t1971 145.137
R10308 VPWR.n250 VPWR.t1930 145.137
R10309 VPWR.n238 VPWR.t2016 145.137
R10310 VPWR.n226 VPWR.t2008 145.137
R10311 VPWR.n214 VPWR.t1928 145.137
R10312 VPWR.n202 VPWR.t2057 145.137
R10313 VPWR.n190 VPWR.t2017 145.137
R10314 VPWR.n178 VPWR.t1961 145.137
R10315 VPWR.n166 VPWR.t1952 145.137
R10316 VPWR.n154 VPWR.t2007 145.137
R10317 VPWR.n1768 VPWR.t1976 145.137
R10318 VPWR.n1039 VPWR.t2065 145.137
R10319 VPWR.n1543 VPWR.t1929 145.137
R10320 VPWR.n1548 VPWR.t1986 145.137
R10321 VPWR.n1553 VPWR.t2025 145.137
R10322 VPWR.n1558 VPWR.t2037 145.137
R10323 VPWR.n1563 VPWR.t1979 145.137
R10324 VPWR.n1568 VPWR.t1985 145.137
R10325 VPWR.n1573 VPWR.t2039 145.137
R10326 VPWR.n1578 VPWR.t1936 145.137
R10327 VPWR.n1133 VPWR.t1950 145.137
R10328 VPWR.n1458 VPWR.t1996 145.137
R10329 VPWR.n1453 VPWR.t2045 145.137
R10330 VPWR.n1773 VPWR.t1968 145.137
R10331 VPWR.n1781 VPWR.t1953 145.137
R10332 VPWR.n1777 VPWR.t2013 145.137
R10333 VPWR.n142 VPWR.t1999 145.137
R10334 VPWR.n130 VPWR.t1990 145.137
R10335 VPWR.n1119 VPWR.t2067 145.038
R10336 VPWR.n1110 VPWR.t2018 145.038
R10337 VPWR.n1611 VPWR.t2010 145.038
R10338 VPWR.n1622 VPWR.t1955 145.038
R10339 VPWR.n1100 VPWR.t2059 145.038
R10340 VPWR.n1638 VPWR.t2002 145.038
R10341 VPWR.n1649 VPWR.t1964 145.038
R10342 VPWR.n1090 VPWR.t1949 145.038
R10343 VPWR.n1665 VPWR.t2043 145.038
R10344 VPWR.n1676 VPWR.t2003 145.038
R10345 VPWR.n1080 VPWR.t1947 145.038
R10346 VPWR.n1692 VPWR.t1939 145.038
R10347 VPWR.n1703 VPWR.t2036 145.038
R10348 VPWR.n1069 VPWR.t1989 145.038
R10349 VPWR.n1716 VPWR.t1977 145.038
R10350 VPWR.n1064 VPWR.t2034 145.038
R10351 VPWR.n125 VPWR.t1940 145.038
R10352 VPWR.n114 VPWR.t2001 145.038
R10353 VPWR.n137 VPWR.t1954 145.038
R10354 VPWR.n104 VPWR.t2032 145.038
R10355 VPWR.n100 VPWR.t1987 145.038
R10356 VPWR.n269 VPWR.t1980 145.038
R10357 VPWR.n257 VPWR.t2068 145.038
R10358 VPWR.n245 VPWR.t2027 145.038
R10359 VPWR.n233 VPWR.t1972 145.038
R10360 VPWR.n221 VPWR.t1931 145.038
R10361 VPWR.n209 VPWR.t2060 145.038
R10362 VPWR.n197 VPWR.t2009 145.038
R10363 VPWR.n185 VPWR.t1973 145.038
R10364 VPWR.n173 VPWR.t2058 145.038
R10365 VPWR.n161 VPWR.t2052 145.038
R10366 VPWR.n149 VPWR.t2004 145.038
R10367 VPWR.n53 VPWR.t2053 145.038
R10368 VPWR.n51 VPWR.t1963 145.038
R10369 VPWR.n49 VPWR.t2066 145.038
R10370 VPWR.n47 VPWR.t2026 145.038
R10371 VPWR.n45 VPWR.t1946 145.038
R10372 VPWR.n43 VPWR.t2051 145.038
R10373 VPWR.n41 VPWR.t2069 145.038
R10374 VPWR.n39 VPWR.t2028 145.038
R10375 VPWR.n37 VPWR.t2022 145.038
R10376 VPWR.n35 VPWR.t1943 145.038
R10377 VPWR.n33 VPWR.t1997 145.038
R10378 VPWR.n31 VPWR.t2064 145.038
R10379 VPWR.n29 VPWR.t1995 145.038
R10380 VPWR.n27 VPWR.t1956 145.038
R10381 VPWR.n25 VPWR.t2021 145.038
R10382 VPWR.n23 VPWR.t1970 145.038
R10383 VPWR.n1598 VPWR.t1966 143.911
R10384 VPWR.n1125 VPWR.t2062 143.911
R10385 VPWR.n1614 VPWR.t2047 143.911
R10386 VPWR.n1625 VPWR.t1965 143.911
R10387 VPWR.n1176 VPWR.t1958 143.911
R10388 VPWR.n1641 VPWR.t1944 143.911
R10389 VPWR.n1652 VPWR.t2005 143.911
R10390 VPWR.n1208 VPWR.t1992 143.911
R10391 VPWR.n1668 VPWR.t1941 143.911
R10392 VPWR.n1679 VPWR.t2038 143.911
R10393 VPWR.n1194 VPWR.t2031 143.911
R10394 VPWR.n1695 VPWR.t1978 143.911
R10395 VPWR.n1706 VPWR.t1935 143.911
R10396 VPWR.n1718 VPWR.t2024 143.911
R10397 VPWR.n1733 VPWR.t1984 143.911
R10398 VPWR.n1114 VPWR.t2012 143.911
R10399 VPWR.n116 VPWR.t1951 143.911
R10400 VPWR.n127 VPWR.t1991 143.911
R10401 VPWR.n106 VPWR.t1981 143.911
R10402 VPWR.n287 VPWR.t1933 143.911
R10403 VPWR.n271 VPWR.t2029 143.911
R10404 VPWR.n259 VPWR.t2015 143.911
R10405 VPWR.n247 VPWR.t1932 143.911
R10406 VPWR.n235 VPWR.t1926 143.911
R10407 VPWR.n223 VPWR.t2056 143.911
R10408 VPWR.n211 VPWR.t1974 143.911
R10409 VPWR.n199 VPWR.t1960 143.911
R10410 VPWR.n187 VPWR.t2054 143.911
R10411 VPWR.n175 VPWR.t2006 143.911
R10412 VPWR.n163 VPWR.t1998 143.911
R10413 VPWR.n151 VPWR.t1942 143.911
R10414 VPWR.n1228 VPWR.t1948 143.911
R10415 VPWR.n1150 VPWR.t1975 143.911
R10416 VPWR.n1224 VPWR.t2041 143.911
R10417 VPWR.n1482 VPWR.t1982 143.911
R10418 VPWR.n1170 VPWR.t2035 143.911
R10419 VPWR.n1166 VPWR.t2023 143.911
R10420 VPWR.n1160 VPWR.t1938 143.911
R10421 VPWR.n1476 VPWR.t1994 143.911
R10422 VPWR.n1156 VPWR.t1927 143.911
R10423 VPWR.n1146 VPWR.t2020 143.911
R10424 VPWR.n1469 VPWR.t2044 143.911
R10425 VPWR.n1046 VPWR.t1967 143.911
R10426 VPWR.n1745 VPWR.t2011 143.911
R10427 VPWR.n1033 VPWR.t1957 143.911
R10428 VPWR.n1029 VPWR.t2061 143.911
R10429 VPWR.n1050 VPWR.t2055 143.911
R10430 VPWR.n139 VPWR.t2046 143.911
R10431 VPWR.t1293 VPWR.t1307 140.989
R10432 VPWR.t922 VPWR.t16 140.989
R10433 VPWR.t88 VPWR.t922 140.989
R10434 VPWR.t884 VPWR.t88 140.989
R10435 VPWR.t659 VPWR.t884 140.989
R10436 VPWR.t405 VPWR.t659 140.989
R10437 VPWR.t1132 VPWR.t405 140.989
R10438 VPWR.t1128 VPWR.t1132 140.989
R10439 VPWR.t1403 VPWR.t31 140.989
R10440 VPWR.t1918 VPWR.t911 140.989
R10441 VPWR.t10 VPWR.t1918 140.989
R10442 VPWR.t91 VPWR.t10 140.989
R10443 VPWR.t957 VPWR.t91 140.989
R10444 VPWR.t969 VPWR.t957 140.989
R10445 VPWR.t961 VPWR.t969 140.989
R10446 VPWR.t965 VPWR.t961 140.989
R10447 VPWR.t1324 VPWR.t879 140.989
R10448 VPWR.t927 VPWR.t1324 140.989
R10449 VPWR.t13 VPWR.t927 140.989
R10450 VPWR.t808 VPWR.t13 140.989
R10451 VPWR.t806 VPWR.t808 140.989
R10452 VPWR.t812 VPWR.t806 140.989
R10453 VPWR.t800 VPWR.t812 140.989
R10454 VPWR.t1108 VPWR.t928 140.989
R10455 VPWR.t17 VPWR.t86 140.989
R10456 VPWR.t1828 VPWR.t17 140.989
R10457 VPWR.t930 VPWR.t1828 140.989
R10458 VPWR.t1130 VPWR.t930 140.989
R10459 VPWR.t782 VPWR.t1130 140.989
R10460 VPWR.t372 VPWR.t782 140.989
R10461 VPWR.t1142 VPWR.t372 140.989
R10462 VPWR.t880 VPWR.t84 140.989
R10463 VPWR.t1326 VPWR.t880 140.989
R10464 VPWR.t82 VPWR.t1326 140.989
R10465 VPWR.t967 VPWR.t82 140.989
R10466 VPWR.t959 VPWR.t967 140.989
R10467 VPWR.t971 VPWR.t959 140.989
R10468 VPWR.t963 VPWR.t971 140.989
R10469 VPWR.t89 VPWR.t923 140.989
R10470 VPWR.t885 VPWR.t89 140.989
R10471 VPWR.t925 VPWR.t885 140.989
R10472 VPWR.t810 VPWR.t925 140.989
R10473 VPWR.t814 VPWR.t810 140.989
R10474 VPWR.t802 VPWR.t814 140.989
R10475 VPWR.t804 VPWR.t802 140.989
R10476 VPWR VPWR.n1442 133.312
R10477 VPWR.n2841 VPWR.n2840 129.13
R10478 VPWR.n2858 VPWR.n2819 129.13
R10479 VPWR.n2780 VPWR 127.562
R10480 VPWR.n2760 VPWR 127.562
R10481 VPWR.n2741 VPWR 127.562
R10482 VPWR VPWR.t1830 125.883
R10483 VPWR.n2705 VPWR 125.883
R10484 VPWR.t1405 VPWR.t29 120.849
R10485 VPWR.t649 VPWR.t1250 117.492
R10486 VPWR.t821 VPWR.t994 117.492
R10487 VPWR.t460 VPWR 115.814
R10488 VPWR VPWR.t1128 114.135
R10489 VPWR VPWR.t965 114.135
R10490 VPWR VPWR.t800 114.135
R10491 VPWR.n2859 VPWR.n2817 111.059
R10492 VPWR.t228 VPWR 107.421
R10493 VPWR.n1330 VPWR.n1329 106.561
R10494 VPWR.n2781 VPWR.n2780 106.561
R10495 VPWR.n2761 VPWR.n2760 106.561
R10496 VPWR.n2742 VPWR.n2741 106.561
R10497 VPWR.n2706 VPWR.n2705 106.561
R10498 VPWR.n2668 VPWR.n2667 106.561
R10499 VPWR.n2631 VPWR.n2630 106.561
R10500 VPWR VPWR.t1409 106.543
R10501 VPWR VPWR.n1234 104.8
R10502 VPWR VPWR.n1257 104.8
R10503 VPWR VPWR.n1281 104.8
R10504 VPWR VPWR.n1366 104.8
R10505 VPWR VPWR.n1405 104.8
R10506 VPWR.n1443 VPWR 100.883
R10507 VPWR VPWR.t437 100.624
R10508 VPWR.t1800 VPWR.t516 97.9386
R10509 VPWR.n2859 VPWR.n2858 93.3652
R10510 VPWR.n1231 VPWR.n1230 91.8492
R10511 VPWR.n1153 VPWR.n1152 91.8492
R10512 VPWR.n1227 VPWR.n1226 91.8492
R10513 VPWR.n1485 VPWR.n1484 91.8492
R10514 VPWR.n1173 VPWR.n1172 91.8492
R10515 VPWR.n1169 VPWR.n1168 91.8492
R10516 VPWR.n1163 VPWR.n1162 91.8492
R10517 VPWR.n1479 VPWR.n1478 91.8492
R10518 VPWR.n1159 VPWR.n1158 91.8492
R10519 VPWR.n1149 VPWR.n1148 91.8492
R10520 VPWR.n1472 VPWR.n1471 91.8492
R10521 VPWR.n1049 VPWR.n1048 91.8492
R10522 VPWR.n1748 VPWR.n1747 91.8492
R10523 VPWR.n1036 VPWR.n1035 91.8492
R10524 VPWR.n1032 VPWR.n1031 91.8492
R10525 VPWR.n1053 VPWR.n1052 91.8492
R10526 VPWR.n2847 VPWR.n2820 91.4829
R10527 VPWR.t1800 VPWR.n2842 90.0872
R10528 VPWR.t1923 VPWR 88.7855
R10529 VPWR.n1235 VPWR 79.407
R10530 VPWR.n1258 VPWR 79.407
R10531 VPWR.n1282 VPWR 79.407
R10532 VPWR.n1367 VPWR 79.407
R10533 VPWR.n1406 VPWR 79.407
R10534 VPWR.t563 VPWR.t1282 78.8874
R10535 VPWR.n2840 VPWR.n2818 74.9181
R10536 VPWR.n2858 VPWR.n2818 74.9181
R10537 VPWR.n2858 VPWR.n2857 74.9181
R10538 VPWR.n2857 VPWR.n2820 74.9181
R10539 VPWR.t35 VPWR.t439 70.4952
R10540 VPWR.t439 VPWR.t39 70.4952
R10541 VPWR.t39 VPWR.t786 70.4952
R10542 VPWR.t786 VPWR.t1798 70.4952
R10543 VPWR.t1798 VPWR.t1297 70.4952
R10544 VPWR.t1297 VPWR.t1241 70.4952
R10545 VPWR.t1241 VPWR.t1293 70.4952
R10546 VPWR.t920 VPWR.t1108 70.4952
R10547 VPWR.t867 VPWR.t920 70.4952
R10548 VPWR.t11 VPWR.t867 70.4952
R10549 VPWR.t1106 VPWR.t11 70.4952
R10550 VPWR.t882 VPWR.t1106 70.4952
R10551 VPWR.t1112 VPWR.t882 70.4952
R10552 VPWR.t1830 VPWR.t1112 70.4952
R10553 VPWR VPWR.t35 68.8168
R10554 VPWR.t1411 VPWR.t1407 68.8168
R10555 VPWR.t1282 VPWR.t460 62.103
R10556 VPWR VPWR.t1403 60.4245
R10557 VPWR.n2849 VPWR.n2842 59.762
R10558 VPWR.n2845 VPWR.n2819 53.8358
R10559 VPWR.t1407 VPWR.t27 52.0323
R10560 VPWR.t998 VPWR 50.3539
R10561 VPWR VPWR.t1411 50.3539
R10562 VPWR VPWR.t1405 50.3539
R10563 VPWR.t86 VPWR 50.3539
R10564 VPWR.t84 VPWR 50.3539
R10565 VPWR.t923 VPWR 50.3539
R10566 VPWR.n2854 VPWR.n2818 46.2505
R10567 VPWR.n2855 VPWR.n2854 46.2505
R10568 VPWR.n2835 VPWR.n2834 46.2505
R10569 VPWR.n2836 VPWR.n2835 46.2505
R10570 VPWR.n2838 VPWR.n2837 46.2505
R10571 VPWR.n2837 VPWR.n2836 46.2505
R10572 VPWR.n2844 VPWR.n2824 46.2505
R10573 VPWR.n2857 VPWR.n2856 46.2505
R10574 VPWR.n2856 VPWR.n2855 46.2505
R10575 VPWR.n2849 VPWR.n2848 46.2505
R10576 VPWR.n2846 VPWR.n2845 45.9299
R10577 VPWR.n2832 VPWR.n2830 44.8005
R10578 VPWR.n2830 VPWR.n2826 44.8005
R10579 VPWR.n2847 VPWR.n2843 37.0005
R10580 VPWR.n2843 VPWR.t516 37.0005
R10581 VPWR.n1230 VPWR.n1229 34.7473
R10582 VPWR.n1152 VPWR.n1151 34.7473
R10583 VPWR.n1226 VPWR.n1225 34.7473
R10584 VPWR.n1484 VPWR.n1483 34.7473
R10585 VPWR.n1172 VPWR.n1171 34.7473
R10586 VPWR.n1168 VPWR.n1167 34.7473
R10587 VPWR.n1162 VPWR.n1161 34.7473
R10588 VPWR.n1478 VPWR.n1477 34.7473
R10589 VPWR.n1158 VPWR.n1157 34.7473
R10590 VPWR.n1148 VPWR.n1147 34.7473
R10591 VPWR.n1471 VPWR.n1470 34.7473
R10592 VPWR.n1048 VPWR.n1047 34.7473
R10593 VPWR.n1747 VPWR.n1746 34.7473
R10594 VPWR.n1035 VPWR.n1034 34.7473
R10595 VPWR.n1031 VPWR.n1030 34.7473
R10596 VPWR.n1052 VPWR.n1051 34.7473
R10597 VPWR.n1299 VPWR.n1298 34.6358
R10598 VPWR.n1357 VPWR.n1341 34.6358
R10599 VPWR.n1362 VPWR.n1361 34.6358
R10600 VPWR.n1396 VPWR.n1380 34.6358
R10601 VPWR.n1401 VPWR.n1400 34.6358
R10602 VPWR.n1411 VPWR.n1377 34.6358
R10603 VPWR.n1433 VPWR.n1417 34.6358
R10604 VPWR.n1438 VPWR.n1437 34.6358
R10605 VPWR.n2755 VPWR.n2754 34.6358
R10606 VPWR.n2721 VPWR.n2713 34.6358
R10607 VPWR.n2728 VPWR.n2727 34.6358
R10608 VPWR.n2685 VPWR.n2676 34.6358
R10609 VPWR.n2688 VPWR.n2687 34.6358
R10610 VPWR.n2692 VPWR.n2691 34.6358
R10611 VPWR.n2648 VPWR.n2639 34.6358
R10612 VPWR.n2651 VPWR.n2650 34.6358
R10613 VPWR.n2655 VPWR.n2654 34.6358
R10614 VPWR.n2662 VPWR.n2661 34.6358
R10615 VPWR.n2615 VPWR.n2611 34.6358
R10616 VPWR.n2619 VPWR.n2603 34.6358
R10617 VPWR.n2622 VPWR.n2621 34.6358
R10618 VPWR.n1316 VPWR.n1315 32.0005
R10619 VPWR.n1353 VPWR.n1352 32.0005
R10620 VPWR.n1392 VPWR.n1391 32.0005
R10621 VPWR.n1429 VPWR.n1428 32.0005
R10622 VPWR.n2717 VPWR.n2716 30.8711
R10623 VPWR.n2681 VPWR.n2680 30.8711
R10624 VPWR.n2644 VPWR.n2643 30.8711
R10625 VPWR.n2610 VPWR.n2609 30.8711
R10626 VPWR.n2834 VPWR.n2832 30.1181
R10627 VPWR.n2838 VPWR.n2826 30.1181
R10628 VPWR.n2848 VPWR.n2846 28.9887
R10629 VPWR.n1325 VPWR.n1324 28.2358
R10630 VPWR.n5 VPWR.t789 26.5955
R10631 VPWR.n5 VPWR.t1296 26.5955
R10632 VPWR.n4 VPWR.t438 26.5955
R10633 VPWR.n4 VPWR.t785 26.5955
R10634 VPWR.n1240 VPWR.t401 26.5955
R10635 VPWR.n1240 VPWR.t400 26.5955
R10636 VPWR.n1239 VPWR.t647 26.5955
R10637 VPWR.n1239 VPWR.t951 26.5955
R10638 VPWR.n1245 VPWR.t396 26.5955
R10639 VPWR.n1245 VPWR.t402 26.5955
R10640 VPWR.n1238 VPWR.t702 26.5955
R10641 VPWR.n1238 VPWR.t646 26.5955
R10642 VPWR.n1263 VPWR.t1340 26.5955
R10643 VPWR.n1263 VPWR.t1341 26.5955
R10644 VPWR.n1262 VPWR.t1266 26.5955
R10645 VPWR.n1262 VPWR.t1264 26.5955
R10646 VPWR.n1268 VPWR.t933 26.5955
R10647 VPWR.n1268 VPWR.t1402 26.5955
R10648 VPWR.n1261 VPWR.t1269 26.5955
R10649 VPWR.n1261 VPWR.t1267 26.5955
R10650 VPWR.n1287 VPWR.t388 26.5955
R10651 VPWR.n1287 VPWR.t395 26.5955
R10652 VPWR.n1286 VPWR.t655 26.5955
R10653 VPWR.n1286 VPWR.t654 26.5955
R10654 VPWR.n1292 VPWR.t392 26.5955
R10655 VPWR.n1292 VPWR.t389 26.5955
R10656 VPWR.n1285 VPWR.t658 26.5955
R10657 VPWR.n1285 VPWR.t656 26.5955
R10658 VPWR.n1314 VPWR.t1310 26.5955
R10659 VPWR.n1314 VPWR.t1312 26.5955
R10660 VPWR.n1307 VPWR.t1294 26.5955
R10661 VPWR.n1307 VPWR.t1308 26.5955
R10662 VPWR.n1321 VPWR.t787 26.5955
R10663 VPWR.n1321 VPWR.t1298 26.5955
R10664 VPWR.n1323 VPWR.t40 26.5955
R10665 VPWR.n1323 VPWR.t1799 26.5955
R10666 VPWR.n1351 VPWR.t850 26.5955
R10667 VPWR.n1351 VPWR.t1796 26.5955
R10668 VPWR.n1350 VPWR.t110 26.5955
R10669 VPWR.n1350 VPWR.t832 26.5955
R10670 VPWR.n1344 VPWR.t404 26.5955
R10671 VPWR.n1344 VPWR.t845 26.5955
R10672 VPWR.n1343 VPWR.t703 26.5955
R10673 VPWR.n1343 VPWR.t78 26.5955
R10674 VPWR.n1359 VPWR.t399 26.5955
R10675 VPWR.n1359 VPWR.t398 26.5955
R10676 VPWR.n1358 VPWR.t952 26.5955
R10677 VPWR.n1358 VPWR.t645 26.5955
R10678 VPWR.n1390 VPWR.t76 26.5955
R10679 VPWR.n1390 VPWR.t112 26.5955
R10680 VPWR.n1389 VPWR.t852 26.5955
R10681 VPWR.n1389 VPWR.t1797 26.5955
R10682 VPWR.n1383 VPWR.t288 26.5955
R10683 VPWR.n1383 VPWR.t73 26.5955
R10684 VPWR.n1382 VPWR.t1270 26.5955
R10685 VPWR.n1382 VPWR.t848 26.5955
R10686 VPWR.n1398 VPWR.t287 26.5955
R10687 VPWR.n1398 VPWR.t932 26.5955
R10688 VPWR.n1397 VPWR.t1271 26.5955
R10689 VPWR.n1397 VPWR.t1268 26.5955
R10690 VPWR.n1427 VPWR.t34 26.5955
R10691 VPWR.n1427 VPWR.t41 26.5955
R10692 VPWR.n1426 VPWR.t111 26.5955
R10693 VPWR.n1426 VPWR.t833 26.5955
R10694 VPWR.n1420 VPWR.t391 26.5955
R10695 VPWR.n1420 VPWR.t834 26.5955
R10696 VPWR.n1419 VPWR.t652 26.5955
R10697 VPWR.n1419 VPWR.t80 26.5955
R10698 VPWR.n1435 VPWR.t394 26.5955
R10699 VPWR.n1435 VPWR.t393 26.5955
R10700 VPWR.n1434 VPWR.t653 26.5955
R10701 VPWR.n1434 VPWR.t651 26.5955
R10702 VPWR.n2802 VPWR.t1066 26.5955
R10703 VPWR.n2802 VPWR.t1064 26.5955
R10704 VPWR.n2804 VPWR.t1111 26.5955
R10705 VPWR.n2804 VPWR.t870 26.5955
R10706 VPWR.n2782 VPWR.t1908 26.5955
R10707 VPWR.n2782 VPWR.t1905 26.5955
R10708 VPWR.n2783 VPWR.t660 26.5955
R10709 VPWR.n2783 VPWR.t406 26.5955
R10710 VPWR.n2786 VPWR.t1901 26.5955
R10711 VPWR.n2786 VPWR.t1902 26.5955
R10712 VPWR.n2787 VPWR.t1133 26.5955
R10713 VPWR.n2787 VPWR.t1129 26.5955
R10714 VPWR.n2762 VPWR.t1396 26.5955
R10715 VPWR.n2762 VPWR.t1401 26.5955
R10716 VPWR.n2763 VPWR.t958 26.5955
R10717 VPWR.n2763 VPWR.t970 26.5955
R10718 VPWR.n2766 VPWR.t1397 26.5955
R10719 VPWR.n2766 VPWR.t1398 26.5955
R10720 VPWR.n2767 VPWR.t962 26.5955
R10721 VPWR.n2767 VPWR.t966 26.5955
R10722 VPWR.n2743 VPWR.t1139 26.5955
R10723 VPWR.n2743 VPWR.t1136 26.5955
R10724 VPWR.n2744 VPWR.t809 26.5955
R10725 VPWR.n2744 VPWR.t807 26.5955
R10726 VPWR.n2747 VPWR.t1140 26.5955
R10727 VPWR.n2747 VPWR.t1141 26.5955
R10728 VPWR.n2748 VPWR.t813 26.5955
R10729 VPWR.n2748 VPWR.t801 26.5955
R10730 VPWR.n2708 VPWR.t12 26.5955
R10731 VPWR.n2708 VPWR.t883 26.5955
R10732 VPWR.n2712 VPWR.t929 26.5955
R10733 VPWR.n2712 VPWR.t1109 26.5955
R10734 VPWR.n2715 VPWR.t15 26.5955
R10735 VPWR.n2715 VPWR.t1920 26.5955
R10736 VPWR.n2709 VPWR.t868 26.5955
R10737 VPWR.n2709 VPWR.t1107 26.5955
R10738 VPWR.n2679 VPWR.t18 26.5955
R10739 VPWR.n2679 VPWR.t1921 26.5955
R10740 VPWR.n2678 VPWR.t914 26.5955
R10741 VPWR.n2678 VPWR.t1829 26.5955
R10742 VPWR.n2675 VPWR.t931 26.5955
R10743 VPWR.n2675 VPWR.t1131 26.5955
R10744 VPWR.n2674 VPWR.t1925 26.5955
R10745 VPWR.n2674 VPWR.t1906 26.5955
R10746 VPWR.n2671 VPWR.t783 26.5955
R10747 VPWR.n2671 VPWR.t373 26.5955
R10748 VPWR.n2670 VPWR.t1903 26.5955
R10749 VPWR.n2670 VPWR.t1907 26.5955
R10750 VPWR.n2642 VPWR.t913 26.5955
R10751 VPWR.n2642 VPWR.t1327 26.5955
R10752 VPWR.n2641 VPWR.t881 26.5955
R10753 VPWR.n2641 VPWR.t1842 26.5955
R10754 VPWR.n2638 VPWR.t1922 26.5955
R10755 VPWR.n2638 VPWR.t968 26.5955
R10756 VPWR.n2637 VPWR.t83 26.5955
R10757 VPWR.n2637 VPWR.t1394 26.5955
R10758 VPWR.n2634 VPWR.t960 26.5955
R10759 VPWR.n2634 VPWR.t972 26.5955
R10760 VPWR.n2633 VPWR.t1399 26.5955
R10761 VPWR.n2633 VPWR.t1395 26.5955
R10762 VPWR.n2606 VPWR.t915 26.5955
R10763 VPWR.n2606 VPWR.t910 26.5955
R10764 VPWR.n2605 VPWR.t90 26.5955
R10765 VPWR.n2605 VPWR.t886 26.5955
R10766 VPWR.n2613 VPWR.t926 26.5955
R10767 VPWR.n2613 VPWR.t811 26.5955
R10768 VPWR.n2612 VPWR.t1843 26.5955
R10769 VPWR.n2612 VPWR.t1137 26.5955
R10770 VPWR.n2602 VPWR.t815 26.5955
R10771 VPWR.n2602 VPWR.t803 26.5955
R10772 VPWR.n2601 VPWR.t1134 26.5955
R10773 VPWR.n2601 VPWR.t1138 26.5955
R10774 VPWR.n17 VPWR.n16 25.977
R10775 VPWR.n1253 VPWR.n1252 25.977
R10776 VPWR.n1313 VPWR.n1310 25.977
R10777 VPWR.n1349 VPWR.n1346 25.977
R10778 VPWR.n1372 VPWR.n1338 25.977
R10779 VPWR.n1388 VPWR.n1385 25.977
R10780 VPWR.n1425 VPWR.n1422 25.977
R10781 VPWR.n2811 VPWR.n2810 25.977
R10782 VPWR.n2795 VPWR.n2794 25.977
R10783 VPWR.n2717 VPWR.n2714 25.977
R10784 VPWR.n2681 VPWR.n2677 25.977
R10785 VPWR.n2699 VPWR.n2698 25.977
R10786 VPWR.n2644 VPWR.n2640 25.977
R10787 VPWR.n2609 VPWR.n2607 25.977
R10788 VPWR.n1335 VPWR.n1334 25.224
R10789 VPWR.n2737 VPWR.n2736 25.224
R10790 VPWR.n2722 VPWR.n2721 24.8476
R10791 VPWR.n2686 VPWR.n2685 24.8476
R10792 VPWR.n2649 VPWR.n2648 24.8476
R10793 VPWR.n2615 VPWR.n2614 24.8476
R10794 VPWR.n16 VPWR.n15 24.4711
R10795 VPWR.n1252 VPWR.n1251 24.4711
R10796 VPWR.n1315 VPWR.n1313 24.4711
R10797 VPWR.n1352 VPWR.n1349 24.4711
R10798 VPWR.n1391 VPWR.n1388 24.4711
R10799 VPWR.n1428 VPWR.n1425 24.4711
R10800 VPWR.n2810 VPWR.n2809 24.4711
R10801 VPWR.n2794 VPWR.n2793 24.4711
R10802 VPWR.n11 VPWR.n2 23.7181
R10803 VPWR.n1247 VPWR.n1236 23.7181
R10804 VPWR.n1270 VPWR.n1259 23.7181
R10805 VPWR.n1274 VPWR.n1259 23.7181
R10806 VPWR.n1294 VPWR.n1283 23.7181
R10807 VPWR.n1298 VPWR.n1283 23.7181
R10808 VPWR.n1330 VPWR.n1328 23.7181
R10809 VPWR.n1368 VPWR.n1365 23.7181
R10810 VPWR.n1407 VPWR.n1404 23.7181
R10811 VPWR.n1407 VPWR.n1377 23.7181
R10812 VPWR.n1444 VPWR.n1441 23.7181
R10813 VPWR.n2808 VPWR.n2807 23.7181
R10814 VPWR.n2789 VPWR.n2781 23.7181
R10815 VPWR.n2769 VPWR.n2761 23.7181
R10816 VPWR.n2773 VPWR.n2761 23.7181
R10817 VPWR.n2750 VPWR.n2742 23.7181
R10818 VPWR.n2754 VPWR.n2742 23.7181
R10819 VPWR.n2731 VPWR.n2706 23.7181
R10820 VPWR.n2694 VPWR.n2668 23.7181
R10821 VPWR.n2657 VPWR.n2631 23.7181
R10822 VPWR.n2661 VPWR.n2631 23.7181
R10823 VPWR.n2626 VPWR.n2625 23.7181
R10824 VPWR.t1252 VPWR.t649 23.4987
R10825 VPWR.t996 VPWR.t821 23.4987
R10826 VPWR.n2852 VPWR.n2841 23.1255
R10827 VPWR.n2852 VPWR.t1800 23.1255
R10828 VPWR.n2851 VPWR.n2819 23.1255
R10829 VPWR.t1800 VPWR.n2851 23.1255
R10830 VPWR.n11 VPWR.n10 22.9652
R10831 VPWR.n1247 VPWR.n1246 22.9652
R10832 VPWR.n1270 VPWR.n1269 22.9652
R10833 VPWR.n1294 VPWR.n1293 22.9652
R10834 VPWR.n2807 VPWR.n2803 22.9652
R10835 VPWR.n2789 VPWR.n2788 22.9652
R10836 VPWR.n2769 VPWR.n2768 22.9652
R10837 VPWR.n2750 VPWR.n2749 22.9652
R10838 VPWR.n1320 VPWR.n1308 22.2123
R10839 VPWR.n2724 VPWR.n2723 22.2123
R10840 VPWR.n10 VPWR.n3 21.4593
R10841 VPWR.n1246 VPWR.n1237 21.4593
R10842 VPWR.n1269 VPWR.n1260 21.4593
R10843 VPWR.n1293 VPWR.n1284 21.4593
R10844 VPWR.n1442 VPWR.t79 20.5957
R10845 VPWR.n1443 VPWR.t33 20.5957
R10846 VPWR.n1277 VPWR.n1276 19.9534
R10847 VPWR.n1300 VPWR.n1299 19.9534
R10848 VPWR.n1334 VPWR.n1303 19.9534
R10849 VPWR.n2776 VPWR.n2775 19.9534
R10850 VPWR.n2756 VPWR.n2755 19.9534
R10851 VPWR.n2736 VPWR.n2735 19.9534
R10852 VPWR.n2724 VPWR.n2710 18.824
R10853 VPWR.n2688 VPWR.n2672 18.824
R10854 VPWR.n2651 VPWR.n2635 18.824
R10855 VPWR.n2620 VPWR.n2619 18.824
R10856 VPWR.n1316 VPWR.n1308 18.4476
R10857 VPWR.n1353 VPWR.n1345 18.4476
R10858 VPWR.n1373 VPWR.n1372 18.4476
R10859 VPWR.n1392 VPWR.n1384 18.4476
R10860 VPWR.n1429 VPWR.n1421 18.4476
R10861 VPWR.n2700 VPWR.n2699 18.4476
R10862 VPWR.n1413 VPWR.n1412 17.5829
R10863 VPWR.n2664 VPWR.n2663 17.5829
R10864 VPWR.n6 VPWR.n3 16.9417
R10865 VPWR.n1241 VPWR.n1237 16.9417
R10866 VPWR.n1264 VPWR.n1260 16.9417
R10867 VPWR.n1288 VPWR.n1284 16.9417
R10868 VPWR.n2730 VPWR.n2729 16.5652
R10869 VPWR.n1306 VPWR.n1304 16.1887
R10870 VPWR.n1374 VPWR.n1373 16.1887
R10871 VPWR.n2701 VPWR.n2700 16.1887
R10872 VPWR.n1235 VPWR.t43 16.0935
R10873 VPWR.n1258 VPWR.t561 16.0935
R10874 VPWR.n1282 VPWR.t387 16.0935
R10875 VPWR.n1367 VPWR.t397 16.0935
R10876 VPWR.n1406 VPWR.t44 16.0935
R10877 VPWR.n1234 VPWR.t38 16.0935
R10878 VPWR.n1257 VPWR.t42 16.0935
R10879 VPWR.n1281 VPWR.t37 16.0935
R10880 VPWR.n1366 VPWR.t77 16.0935
R10881 VPWR.n1405 VPWR.t74 16.0935
R10882 VPWR.n1325 VPWR.n1306 15.8123
R10883 VPWR.n2727 VPWR.n2710 15.8123
R10884 VPWR.n2729 VPWR.n2728 15.8123
R10885 VPWR.n2691 VPWR.n2672 15.8123
R10886 VPWR.n2654 VPWR.n2635 15.8123
R10887 VPWR.n2621 VPWR.n2620 15.8123
R10888 VPWR.n1330 VPWR.n1303 13.5534
R10889 VPWR.n2735 VPWR.n2706 13.5534
R10890 VPWR.n2839 VPWR.n2823 13.2148
R10891 VPWR.n2823 VPWR.t718 13.2148
R10892 VPWR.n2827 VPWR.n2817 13.2148
R10893 VPWR.n2827 VPWR.t718 13.2148
R10894 VPWR.n2833 VPWR.n2829 13.2148
R10895 VPWR.n2829 VPWR.t718 13.2148
R10896 VPWR.n15 VPWR.n2 12.8005
R10897 VPWR.n1251 VPWR.n1236 12.8005
R10898 VPWR.n1368 VPWR.n1338 12.8005
R10899 VPWR.n2809 VPWR.n2808 12.8005
R10900 VPWR.n2793 VPWR.n2781 12.8005
R10901 VPWR.n2698 VPWR.n2668 12.8005
R10902 VPWR.n1322 VPWR.n1320 12.424
R10903 VPWR.n1360 VPWR.n1357 12.424
R10904 VPWR.n1399 VPWR.n1396 12.424
R10905 VPWR.n1436 VPWR.n1433 12.424
R10906 VPWR.n1276 VPWR.n1275 10.5417
R10907 VPWR.n1412 VPWR.n1411 10.5417
R10908 VPWR.n2775 VPWR.n2774 10.5417
R10909 VPWR.n2663 VPWR.n2662 10.5417
R10910 VPWR.n2687 VPWR.n2686 9.78874
R10911 VPWR.n2650 VPWR.n2649 9.78874
R10912 VPWR.n2614 VPWR.n2603 9.78874
R10913 VPWR.n1361 VPWR.n1360 9.41227
R10914 VPWR.n1365 VPWR.n1339 9.41227
R10915 VPWR.n1400 VPWR.n1399 9.41227
R10916 VPWR.n1404 VPWR.n1378 9.41227
R10917 VPWR.n1437 VPWR.n1436 9.41227
R10918 VPWR.n1441 VPWR.n1415 9.41227
R10919 VPWR.n2694 VPWR.n2693 9.41227
R10920 VPWR.n2657 VPWR.n2656 9.41227
R10921 VPWR.n2625 VPWR.n2599 9.41227
R10922 VPWR.n1229 VPWR 9.37021
R10923 VPWR.n1151 VPWR 9.37021
R10924 VPWR.n1225 VPWR 9.37021
R10925 VPWR.n1483 VPWR 9.37021
R10926 VPWR.n1171 VPWR 9.37021
R10927 VPWR.n1167 VPWR 9.37021
R10928 VPWR.n1161 VPWR 9.37021
R10929 VPWR.n1477 VPWR 9.37021
R10930 VPWR.n1157 VPWR 9.37021
R10931 VPWR.n1147 VPWR 9.37021
R10932 VPWR.n1470 VPWR 9.37021
R10933 VPWR.n1047 VPWR 9.37021
R10934 VPWR.n1746 VPWR 9.37021
R10935 VPWR.n1034 VPWR 9.37021
R10936 VPWR.n1030 VPWR 9.37021
R10937 VPWR.n1051 VPWR 9.37021
R10938 VPWR.n1467 VPWR.n1466 9.33404
R10939 VPWR.n352 VPWR.n351 9.33404
R10940 VPWR.n1534 VPWR.n1533 9.33404
R10941 VPWR.n348 VPWR.n347 9.33404
R10942 VPWR.n965 VPWR.n964 9.33404
R10943 VPWR.n2479 VPWR.n2478 9.33404
R10944 VPWR.n2475 VPWR.n2474 9.33404
R10945 VPWR.n320 VPWR.n319 9.33404
R10946 VPWR.n973 VPWR.n972 9.33404
R10947 VPWR.n2445 VPWR.n2444 9.33404
R10948 VPWR.n324 VPWR.n323 9.33404
R10949 VPWR.n1891 VPWR.n1890 9.33404
R10950 VPWR.n1887 VPWR.n1886 9.33404
R10951 VPWR.n1881 VPWR.n1880 9.33404
R10952 VPWR.n389 VPWR.n388 9.33404
R10953 VPWR.n393 VPWR.n392 9.33404
R10954 VPWR.n397 VPWR.n396 9.33404
R10955 VPWR.n2455 VPWR.n2454 9.33404
R10956 VPWR.n332 VPWR.n331 9.33404
R10957 VPWR.n1877 VPWR.n1876 9.33404
R10958 VPWR.n405 VPWR.n404 9.33404
R10959 VPWR.n2459 VPWR.n2458 9.33404
R10960 VPWR.n336 VPWR.n335 9.33404
R10961 VPWR.n2308 VPWR.n2307 9.33404
R10962 VPWR.n2312 VPWR.n2311 9.33404
R10963 VPWR.n2318 VPWR.n2317 9.33404
R10964 VPWR.n2322 VPWR.n2321 9.33404
R10965 VPWR.n2332 VPWR.n2331 9.33404
R10966 VPWR.n2338 VPWR.n2337 9.33404
R10967 VPWR.n2342 VPWR.n2341 9.33404
R10968 VPWR.n2348 VPWR.n2347 9.33404
R10969 VPWR.n2352 VPWR.n2351 9.33404
R10970 VPWR.n2358 VPWR.n2357 9.33404
R10971 VPWR.n2362 VPWR.n2361 9.33404
R10972 VPWR.n2368 VPWR.n2367 9.33404
R10973 VPWR.n2372 VPWR.n2371 9.33404
R10974 VPWR.n2378 VPWR.n2377 9.33404
R10975 VPWR.n2381 VPWR.n2380 9.33404
R10976 VPWR.n2328 VPWR.n2327 9.33404
R10977 VPWR.n544 VPWR.n543 9.33404
R10978 VPWR.n540 VPWR.n539 9.33404
R10979 VPWR.n536 VPWR.n535 9.33404
R10980 VPWR.n532 VPWR.n531 9.33404
R10981 VPWR.n524 VPWR.n523 9.33404
R10982 VPWR.n520 VPWR.n519 9.33404
R10983 VPWR.n516 VPWR.n515 9.33404
R10984 VPWR.n512 VPWR.n511 9.33404
R10985 VPWR.n508 VPWR.n507 9.33404
R10986 VPWR.n504 VPWR.n503 9.33404
R10987 VPWR.n500 VPWR.n499 9.33404
R10988 VPWR.n496 VPWR.n495 9.33404
R10989 VPWR.n492 VPWR.n491 9.33404
R10990 VPWR.n488 VPWR.n487 9.33404
R10991 VPWR.n485 VPWR.n484 9.33404
R10992 VPWR.n528 VPWR.n527 9.33404
R10993 VPWR.n2283 VPWR.n2282 9.33404
R10994 VPWR.n2279 VPWR.n2278 9.33404
R10995 VPWR.n2273 VPWR.n2272 9.33404
R10996 VPWR.n2269 VPWR.n2268 9.33404
R10997 VPWR.n2259 VPWR.n2258 9.33404
R10998 VPWR.n2253 VPWR.n2252 9.33404
R10999 VPWR.n2249 VPWR.n2248 9.33404
R11000 VPWR.n2243 VPWR.n2242 9.33404
R11001 VPWR.n2239 VPWR.n2238 9.33404
R11002 VPWR.n2233 VPWR.n2232 9.33404
R11003 VPWR.n2229 VPWR.n2228 9.33404
R11004 VPWR.n2223 VPWR.n2222 9.33404
R11005 VPWR.n2219 VPWR.n2218 9.33404
R11006 VPWR.n2213 VPWR.n2212 9.33404
R11007 VPWR.n2210 VPWR.n2209 9.33404
R11008 VPWR.n2263 VPWR.n2262 9.33404
R11009 VPWR.n581 VPWR.n580 9.33404
R11010 VPWR.n585 VPWR.n584 9.33404
R11011 VPWR.n589 VPWR.n588 9.33404
R11012 VPWR.n593 VPWR.n592 9.33404
R11013 VPWR.n601 VPWR.n600 9.33404
R11014 VPWR.n605 VPWR.n604 9.33404
R11015 VPWR.n609 VPWR.n608 9.33404
R11016 VPWR.n613 VPWR.n612 9.33404
R11017 VPWR.n617 VPWR.n616 9.33404
R11018 VPWR.n621 VPWR.n620 9.33404
R11019 VPWR.n625 VPWR.n624 9.33404
R11020 VPWR.n629 VPWR.n628 9.33404
R11021 VPWR.n633 VPWR.n632 9.33404
R11022 VPWR.n637 VPWR.n636 9.33404
R11023 VPWR.n640 VPWR.n639 9.33404
R11024 VPWR.n597 VPWR.n596 9.33404
R11025 VPWR.n2112 VPWR.n2111 9.33404
R11026 VPWR.n2116 VPWR.n2115 9.33404
R11027 VPWR.n2122 VPWR.n2121 9.33404
R11028 VPWR.n2126 VPWR.n2125 9.33404
R11029 VPWR.n2136 VPWR.n2135 9.33404
R11030 VPWR.n2142 VPWR.n2141 9.33404
R11031 VPWR.n2146 VPWR.n2145 9.33404
R11032 VPWR.n2152 VPWR.n2151 9.33404
R11033 VPWR.n2156 VPWR.n2155 9.33404
R11034 VPWR.n2162 VPWR.n2161 9.33404
R11035 VPWR.n2166 VPWR.n2165 9.33404
R11036 VPWR.n2172 VPWR.n2171 9.33404
R11037 VPWR.n2176 VPWR.n2175 9.33404
R11038 VPWR.n2182 VPWR.n2181 9.33404
R11039 VPWR.n2185 VPWR.n2184 9.33404
R11040 VPWR.n2132 VPWR.n2131 9.33404
R11041 VPWR.n736 VPWR.n735 9.33404
R11042 VPWR.n732 VPWR.n731 9.33404
R11043 VPWR.n728 VPWR.n727 9.33404
R11044 VPWR.n724 VPWR.n723 9.33404
R11045 VPWR.n716 VPWR.n715 9.33404
R11046 VPWR.n712 VPWR.n711 9.33404
R11047 VPWR.n708 VPWR.n707 9.33404
R11048 VPWR.n704 VPWR.n703 9.33404
R11049 VPWR.n700 VPWR.n699 9.33404
R11050 VPWR.n696 VPWR.n695 9.33404
R11051 VPWR.n692 VPWR.n691 9.33404
R11052 VPWR.n688 VPWR.n687 9.33404
R11053 VPWR.n684 VPWR.n683 9.33404
R11054 VPWR.n680 VPWR.n679 9.33404
R11055 VPWR.n677 VPWR.n676 9.33404
R11056 VPWR.n720 VPWR.n719 9.33404
R11057 VPWR.n2087 VPWR.n2086 9.33404
R11058 VPWR.n2083 VPWR.n2082 9.33404
R11059 VPWR.n2077 VPWR.n2076 9.33404
R11060 VPWR.n2073 VPWR.n2072 9.33404
R11061 VPWR.n2063 VPWR.n2062 9.33404
R11062 VPWR.n2057 VPWR.n2056 9.33404
R11063 VPWR.n2053 VPWR.n2052 9.33404
R11064 VPWR.n2047 VPWR.n2046 9.33404
R11065 VPWR.n2043 VPWR.n2042 9.33404
R11066 VPWR.n2037 VPWR.n2036 9.33404
R11067 VPWR.n2033 VPWR.n2032 9.33404
R11068 VPWR.n2027 VPWR.n2026 9.33404
R11069 VPWR.n2023 VPWR.n2022 9.33404
R11070 VPWR.n2017 VPWR.n2016 9.33404
R11071 VPWR.n2014 VPWR.n2013 9.33404
R11072 VPWR.n2067 VPWR.n2066 9.33404
R11073 VPWR.n773 VPWR.n772 9.33404
R11074 VPWR.n777 VPWR.n776 9.33404
R11075 VPWR.n781 VPWR.n780 9.33404
R11076 VPWR.n785 VPWR.n784 9.33404
R11077 VPWR.n793 VPWR.n792 9.33404
R11078 VPWR.n797 VPWR.n796 9.33404
R11079 VPWR.n801 VPWR.n800 9.33404
R11080 VPWR.n805 VPWR.n804 9.33404
R11081 VPWR.n809 VPWR.n808 9.33404
R11082 VPWR.n813 VPWR.n812 9.33404
R11083 VPWR.n817 VPWR.n816 9.33404
R11084 VPWR.n821 VPWR.n820 9.33404
R11085 VPWR.n825 VPWR.n824 9.33404
R11086 VPWR.n829 VPWR.n828 9.33404
R11087 VPWR.n832 VPWR.n831 9.33404
R11088 VPWR.n789 VPWR.n788 9.33404
R11089 VPWR.n1916 VPWR.n1915 9.33404
R11090 VPWR.n1920 VPWR.n1919 9.33404
R11091 VPWR.n1926 VPWR.n1925 9.33404
R11092 VPWR.n1930 VPWR.n1929 9.33404
R11093 VPWR.n1940 VPWR.n1939 9.33404
R11094 VPWR.n1946 VPWR.n1945 9.33404
R11095 VPWR.n1950 VPWR.n1949 9.33404
R11096 VPWR.n1956 VPWR.n1955 9.33404
R11097 VPWR.n1960 VPWR.n1959 9.33404
R11098 VPWR.n1966 VPWR.n1965 9.33404
R11099 VPWR.n1970 VPWR.n1969 9.33404
R11100 VPWR.n1976 VPWR.n1975 9.33404
R11101 VPWR.n1980 VPWR.n1979 9.33404
R11102 VPWR.n1986 VPWR.n1985 9.33404
R11103 VPWR.n1989 VPWR.n1988 9.33404
R11104 VPWR.n1936 VPWR.n1935 9.33404
R11105 VPWR.n928 VPWR.n927 9.33404
R11106 VPWR.n924 VPWR.n923 9.33404
R11107 VPWR.n920 VPWR.n919 9.33404
R11108 VPWR.n916 VPWR.n915 9.33404
R11109 VPWR.n908 VPWR.n907 9.33404
R11110 VPWR.n904 VPWR.n903 9.33404
R11111 VPWR.n900 VPWR.n899 9.33404
R11112 VPWR.n896 VPWR.n895 9.33404
R11113 VPWR.n892 VPWR.n891 9.33404
R11114 VPWR.n888 VPWR.n887 9.33404
R11115 VPWR.n884 VPWR.n883 9.33404
R11116 VPWR.n880 VPWR.n879 9.33404
R11117 VPWR.n876 VPWR.n875 9.33404
R11118 VPWR.n872 VPWR.n871 9.33404
R11119 VPWR.n869 VPWR.n868 9.33404
R11120 VPWR.n912 VPWR.n911 9.33404
R11121 VPWR.n1871 VPWR.n1870 9.33404
R11122 VPWR.n981 VPWR.n980 9.33404
R11123 VPWR.n1495 VPWR.n1494 9.33404
R11124 VPWR.n401 VPWR.n400 9.33404
R11125 VPWR.n2465 VPWR.n2464 9.33404
R11126 VPWR.n340 VPWR.n339 9.33404
R11127 VPWR.n977 VPWR.n976 9.33404
R11128 VPWR.n1491 VPWR.n1490 9.33404
R11129 VPWR.n1867 VPWR.n1866 9.33404
R11130 VPWR.n985 VPWR.n984 9.33404
R11131 VPWR.n1505 VPWR.n1504 9.33404
R11132 VPWR.n409 VPWR.n408 9.33404
R11133 VPWR.n417 VPWR.n416 9.33404
R11134 VPWR.n421 VPWR.n420 9.33404
R11135 VPWR.n425 VPWR.n424 9.33404
R11136 VPWR.n429 VPWR.n428 9.33404
R11137 VPWR.n433 VPWR.n432 9.33404
R11138 VPWR.n437 VPWR.n436 9.33404
R11139 VPWR.n441 VPWR.n440 9.33404
R11140 VPWR.n445 VPWR.n444 9.33404
R11141 VPWR.n448 VPWR.n447 9.33404
R11142 VPWR.n413 VPWR.n412 9.33404
R11143 VPWR.n2449 VPWR.n2448 9.33404
R11144 VPWR.n328 VPWR.n327 9.33404
R11145 VPWR.n989 VPWR.n988 9.33404
R11146 VPWR.n1509 VPWR.n1508 9.33404
R11147 VPWR.n1861 VPWR.n1860 9.33404
R11148 VPWR.n1851 VPWR.n1850 9.33404
R11149 VPWR.n1847 VPWR.n1846 9.33404
R11150 VPWR.n1841 VPWR.n1840 9.33404
R11151 VPWR.n1837 VPWR.n1836 9.33404
R11152 VPWR.n1831 VPWR.n1830 9.33404
R11153 VPWR.n1827 VPWR.n1826 9.33404
R11154 VPWR.n1821 VPWR.n1820 9.33404
R11155 VPWR.n1818 VPWR.n1817 9.33404
R11156 VPWR.n1857 VPWR.n1856 9.33404
R11157 VPWR.n993 VPWR.n992 9.33404
R11158 VPWR.n1519 VPWR.n1518 9.33404
R11159 VPWR.n2469 VPWR.n2468 9.33404
R11160 VPWR.n344 VPWR.n343 9.33404
R11161 VPWR.n1480 VPWR.n1130 9.33404
R11162 VPWR.n997 VPWR.n996 9.33404
R11163 VPWR.n1523 VPWR.n1522 9.33404
R11164 VPWR.n2439 VPWR.n2438 9.33404
R11165 VPWR.n2429 VPWR.n2428 9.33404
R11166 VPWR.n2425 VPWR.n2424 9.33404
R11167 VPWR.n2419 VPWR.n2418 9.33404
R11168 VPWR.n2415 VPWR.n2414 9.33404
R11169 VPWR.n2409 VPWR.n2408 9.33404
R11170 VPWR.n2406 VPWR.n2405 9.33404
R11171 VPWR.n2435 VPWR.n2434 9.33404
R11172 VPWR.n316 VPWR.n315 9.33404
R11173 VPWR.n1538 VPWR.n1537 9.33404
R11174 VPWR.n1001 VPWR.n1000 9.33404
R11175 VPWR.n1005 VPWR.n1004 9.33404
R11176 VPWR.n1009 VPWR.n1008 9.33404
R11177 VPWR.n1013 VPWR.n1012 9.33404
R11178 VPWR.n1017 VPWR.n1016 9.33404
R11179 VPWR.n1021 VPWR.n1020 9.33404
R11180 VPWR.n1024 VPWR.n1023 9.33404
R11181 VPWR.n969 VPWR.n968 9.33404
R11182 VPWR.n1474 VPWR.n1473 9.33404
R11183 VPWR.n312 VPWR.n311 9.33404
R11184 VPWR.n1763 VPWR.n1762 9.33404
R11185 VPWR.n308 VPWR.n307 9.33404
R11186 VPWR.n304 VPWR.n303 9.33404
R11187 VPWR.n296 VPWR.n295 9.33404
R11188 VPWR.n293 VPWR.n292 9.33404
R11189 VPWR.n300 VPWR.n299 9.33404
R11190 VPWR.n1751 VPWR.n1750 9.33404
R11191 VPWR.n1790 VPWR.n1789 9.33404
R11192 VPWR.n1793 VPWR.n1792 9.33404
R11193 VPWR.n1759 VPWR.n1758 9.33404
R11194 VPWR.n2714 VPWR 9.32394
R11195 VPWR.n2677 VPWR 9.32394
R11196 VPWR.n2640 VPWR 9.32394
R11197 VPWR VPWR.n2607 9.32394
R11198 VPWR.n18 VPWR.n17 9.3005
R11199 VPWR.n15 VPWR.n14 9.3005
R11200 VPWR.n13 VPWR.n2 9.3005
R11201 VPWR.n10 VPWR.n9 9.3005
R11202 VPWR.n8 VPWR.n3 9.3005
R11203 VPWR.n12 VPWR.n11 9.3005
R11204 VPWR.n16 VPWR.n0 9.3005
R11205 VPWR.n1254 VPWR.n1253 9.3005
R11206 VPWR.n1251 VPWR.n1250 9.3005
R11207 VPWR.n1249 VPWR.n1236 9.3005
R11208 VPWR.n1246 VPWR.n1244 9.3005
R11209 VPWR.n1243 VPWR.n1237 9.3005
R11210 VPWR.n1248 VPWR.n1247 9.3005
R11211 VPWR.n1252 VPWR.n1233 9.3005
R11212 VPWR.n1278 VPWR.n1277 9.3005
R11213 VPWR.n1272 VPWR.n1259 9.3005
R11214 VPWR.n1269 VPWR.n1267 9.3005
R11215 VPWR.n1266 VPWR.n1260 9.3005
R11216 VPWR.n1271 VPWR.n1270 9.3005
R11217 VPWR.n1274 VPWR.n1273 9.3005
R11218 VPWR.n1276 VPWR.n1256 9.3005
R11219 VPWR.n1301 VPWR.n1300 9.3005
R11220 VPWR.n1296 VPWR.n1283 9.3005
R11221 VPWR.n1293 VPWR.n1291 9.3005
R11222 VPWR.n1290 VPWR.n1284 9.3005
R11223 VPWR.n1295 VPWR.n1294 9.3005
R11224 VPWR.n1298 VPWR.n1297 9.3005
R11225 VPWR.n1299 VPWR.n1280 9.3005
R11226 VPWR.n1332 VPWR.n1303 9.3005
R11227 VPWR.n1331 VPWR.n1330 9.3005
R11228 VPWR.n1311 VPWR.n1310 9.3005
R11229 VPWR.n1313 VPWR.n1312 9.3005
R11230 VPWR.n1315 VPWR.n1309 9.3005
R11231 VPWR.n1317 VPWR.n1316 9.3005
R11232 VPWR.n1318 VPWR.n1308 9.3005
R11233 VPWR.n1320 VPWR.n1319 9.3005
R11234 VPWR.n1324 VPWR.n1305 9.3005
R11235 VPWR.n1326 VPWR.n1325 9.3005
R11236 VPWR.n1328 VPWR.n1327 9.3005
R11237 VPWR.n1334 VPWR.n1333 9.3005
R11238 VPWR.n1336 VPWR.n1335 9.3005
R11239 VPWR.n1375 VPWR.n1374 9.3005
R11240 VPWR.n1370 VPWR.n1338 9.3005
R11241 VPWR.n1369 VPWR.n1368 9.3005
R11242 VPWR.n1347 VPWR.n1346 9.3005
R11243 VPWR.n1349 VPWR.n1348 9.3005
R11244 VPWR.n1352 VPWR.n1342 9.3005
R11245 VPWR.n1354 VPWR.n1353 9.3005
R11246 VPWR.n1355 VPWR.n1341 9.3005
R11247 VPWR.n1357 VPWR.n1356 9.3005
R11248 VPWR.n1361 VPWR.n1340 9.3005
R11249 VPWR.n1363 VPWR.n1362 9.3005
R11250 VPWR.n1365 VPWR.n1364 9.3005
R11251 VPWR.n1372 VPWR.n1371 9.3005
R11252 VPWR.n1408 VPWR.n1407 9.3005
R11253 VPWR.n1386 VPWR.n1385 9.3005
R11254 VPWR.n1388 VPWR.n1387 9.3005
R11255 VPWR.n1391 VPWR.n1381 9.3005
R11256 VPWR.n1393 VPWR.n1392 9.3005
R11257 VPWR.n1394 VPWR.n1380 9.3005
R11258 VPWR.n1396 VPWR.n1395 9.3005
R11259 VPWR.n1400 VPWR.n1379 9.3005
R11260 VPWR.n1402 VPWR.n1401 9.3005
R11261 VPWR.n1404 VPWR.n1403 9.3005
R11262 VPWR.n1409 VPWR.n1377 9.3005
R11263 VPWR.n1411 VPWR.n1410 9.3005
R11264 VPWR.n1445 VPWR.n1444 9.3005
R11265 VPWR.n1423 VPWR.n1422 9.3005
R11266 VPWR.n1425 VPWR.n1424 9.3005
R11267 VPWR.n1428 VPWR.n1418 9.3005
R11268 VPWR.n1430 VPWR.n1429 9.3005
R11269 VPWR.n1431 VPWR.n1417 9.3005
R11270 VPWR.n1433 VPWR.n1432 9.3005
R11271 VPWR.n1437 VPWR.n1416 9.3005
R11272 VPWR.n1439 VPWR.n1438 9.3005
R11273 VPWR.n1441 VPWR.n1440 9.3005
R11274 VPWR.n2807 VPWR.n2806 9.3005
R11275 VPWR.n2808 VPWR.n2800 9.3005
R11276 VPWR.n2809 VPWR.n2799 9.3005
R11277 VPWR.n2810 VPWR.n2798 9.3005
R11278 VPWR.n2812 VPWR.n2811 9.3005
R11279 VPWR.n2796 VPWR.n2795 9.3005
R11280 VPWR.n2790 VPWR.n2789 9.3005
R11281 VPWR.n2791 VPWR.n2781 9.3005
R11282 VPWR.n2793 VPWR.n2792 9.3005
R11283 VPWR.n2794 VPWR.n2779 9.3005
R11284 VPWR.n2777 VPWR.n2776 9.3005
R11285 VPWR.n2775 VPWR.n2759 9.3005
R11286 VPWR.n2770 VPWR.n2769 9.3005
R11287 VPWR.n2771 VPWR.n2761 9.3005
R11288 VPWR.n2773 VPWR.n2772 9.3005
R11289 VPWR.n2757 VPWR.n2756 9.3005
R11290 VPWR.n2751 VPWR.n2750 9.3005
R11291 VPWR.n2752 VPWR.n2742 9.3005
R11292 VPWR.n2754 VPWR.n2753 9.3005
R11293 VPWR.n2755 VPWR.n2740 9.3005
R11294 VPWR.n2738 VPWR.n2737 9.3005
R11295 VPWR.n2718 VPWR.n2717 9.3005
R11296 VPWR.n2719 VPWR.n2713 9.3005
R11297 VPWR.n2721 VPWR.n2720 9.3005
R11298 VPWR.n2723 VPWR.n2711 9.3005
R11299 VPWR.n2725 VPWR.n2724 9.3005
R11300 VPWR.n2727 VPWR.n2726 9.3005
R11301 VPWR.n2728 VPWR.n2707 9.3005
R11302 VPWR.n2732 VPWR.n2731 9.3005
R11303 VPWR.n2733 VPWR.n2706 9.3005
R11304 VPWR.n2735 VPWR.n2734 9.3005
R11305 VPWR.n2736 VPWR.n2704 9.3005
R11306 VPWR.n2702 VPWR.n2701 9.3005
R11307 VPWR.n2682 VPWR.n2681 9.3005
R11308 VPWR.n2683 VPWR.n2676 9.3005
R11309 VPWR.n2685 VPWR.n2684 9.3005
R11310 VPWR.n2687 VPWR.n2673 9.3005
R11311 VPWR.n2689 VPWR.n2688 9.3005
R11312 VPWR.n2691 VPWR.n2690 9.3005
R11313 VPWR.n2692 VPWR.n2669 9.3005
R11314 VPWR.n2695 VPWR.n2694 9.3005
R11315 VPWR.n2696 VPWR.n2668 9.3005
R11316 VPWR.n2698 VPWR.n2697 9.3005
R11317 VPWR.n2699 VPWR.n2666 9.3005
R11318 VPWR.n2645 VPWR.n2644 9.3005
R11319 VPWR.n2646 VPWR.n2639 9.3005
R11320 VPWR.n2648 VPWR.n2647 9.3005
R11321 VPWR.n2650 VPWR.n2636 9.3005
R11322 VPWR.n2652 VPWR.n2651 9.3005
R11323 VPWR.n2654 VPWR.n2653 9.3005
R11324 VPWR.n2655 VPWR.n2632 9.3005
R11325 VPWR.n2658 VPWR.n2657 9.3005
R11326 VPWR.n2659 VPWR.n2631 9.3005
R11327 VPWR.n2661 VPWR.n2660 9.3005
R11328 VPWR.n2662 VPWR.n2629 9.3005
R11329 VPWR.n2627 VPWR.n2626 9.3005
R11330 VPWR.n2609 VPWR.n2608 9.3005
R11331 VPWR.n2611 VPWR.n2604 9.3005
R11332 VPWR.n2616 VPWR.n2615 9.3005
R11333 VPWR.n2617 VPWR.n2603 9.3005
R11334 VPWR.n2619 VPWR.n2618 9.3005
R11335 VPWR.n2621 VPWR.n2600 9.3005
R11336 VPWR.n2623 VPWR.n2622 9.3005
R11337 VPWR.n2625 VPWR.n2624 9.3005
R11338 VPWR.n2505 VPWR.n2504 9.3005
R11339 VPWR.n2569 VPWR.n2568 9.3005
R11340 VPWR.n2509 VPWR.n2508 9.3005
R11341 VPWR.n2553 VPWR.n2552 9.3005
R11342 VPWR.n2545 VPWR.n2544 9.3005
R11343 VPWR.n2533 VPWR.n2532 9.3005
R11344 VPWR.n2529 VPWR.n2528 9.3005
R11345 VPWR.n1222 VPWR.n1221 9.3005
R11346 VPWR.n2521 VPWR.n2520 9.3005
R11347 VPWR.n1184 VPWR.n1102 9.3005
R11348 VPWR.n1218 VPWR.n1094 9.3005
R11349 VPWR.n2541 VPWR.n2540 9.3005
R11350 VPWR.n1215 VPWR.n1092 9.3005
R11351 VPWR.n1212 VPWR.n1211 9.3005
R11352 VPWR.n2517 VPWR.n2516 9.3005
R11353 VPWR.n1181 VPWR.n1104 9.3005
R11354 VPWR.n1204 VPWR.n1084 9.3005
R11355 VPWR.n2557 VPWR.n2556 9.3005
R11356 VPWR.n1201 VPWR.n1082 9.3005
R11357 VPWR.n1592 VPWR.n1591 9.3005
R11358 VPWR.n2565 VPWR.n2564 9.3005
R11359 VPWR.n1198 VPWR.n1197 9.3005
R11360 VPWR.n1190 VPWR.n1074 9.3005
R11361 VPWR.n1742 VPWR.n1741 9.3005
R11362 VPWR.n1187 VPWR.n1071 9.3005
R11363 VPWR.n2577 VPWR.n2576 9.3005
R11364 VPWR.n2581 VPWR.n2580 9.3005
R11365 VPWR.n2592 VPWR.n2591 9.3005
R11366 VPWR.n2589 VPWR.n2588 9.3005
R11367 VPWR.n1738 VPWR.n1737 9.3005
R11368 VPWR.n1063 VPWR.n1062 9.3005
R11369 VPWR.n1596 VPWR.n1595 9.3005
R11370 VPWR.n1275 VPWR.n1274 8.28285
R11371 VPWR.n2774 VPWR.n2773 8.28285
R11372 VPWR.n1607 VPWR.n1109 8.25914
R11373 VPWR.n1728 VPWR.n1727 8.25914
R11374 VPWR.n281 VPWR.n113 8.25914
R11375 VPWR.n136 VPWR.n124 8.25914
R11376 VPWR.n1780 VPWR.n1779 7.91351
R11377 VPWR.n1771 VPWR.n1770 7.9105
R11378 VPWR.n1042 VPWR.n1041 7.9105
R11379 VPWR.n1546 VPWR.n1545 7.9105
R11380 VPWR.n1551 VPWR.n1550 7.9105
R11381 VPWR.n1556 VPWR.n1555 7.9105
R11382 VPWR.n1561 VPWR.n1560 7.9105
R11383 VPWR.n1566 VPWR.n1565 7.9105
R11384 VPWR.n1571 VPWR.n1570 7.9105
R11385 VPWR.n1576 VPWR.n1575 7.9105
R11386 VPWR.n1581 VPWR.n1580 7.9105
R11387 VPWR.n1136 VPWR.n1135 7.9105
R11388 VPWR.n1461 VPWR.n1460 7.9105
R11389 VPWR.n1456 VPWR.n1455 7.9105
R11390 VPWR.n1776 VPWR.n1775 7.9105
R11391 VPWR.n1784 VPWR.n1783 7.9105
R11392 VPWR.n282 VPWR.n281 7.9105
R11393 VPWR.n280 VPWR.n279 7.9105
R11394 VPWR.n268 VPWR.n267 7.9105
R11395 VPWR.n256 VPWR.n255 7.9105
R11396 VPWR.n244 VPWR.n243 7.9105
R11397 VPWR.n232 VPWR.n231 7.9105
R11398 VPWR.n220 VPWR.n219 7.9105
R11399 VPWR.n208 VPWR.n207 7.9105
R11400 VPWR.n196 VPWR.n195 7.9105
R11401 VPWR.n184 VPWR.n183 7.9105
R11402 VPWR.n172 VPWR.n171 7.9105
R11403 VPWR.n160 VPWR.n159 7.9105
R11404 VPWR.n148 VPWR.n147 7.9105
R11405 VPWR.n136 VPWR.n135 7.9105
R11406 VPWR.n1727 VPWR.n1726 7.9105
R11407 VPWR.n1715 VPWR.n1714 7.9105
R11408 VPWR.n1701 VPWR.n1068 7.9105
R11409 VPWR.n1690 VPWR.n1689 7.9105
R11410 VPWR.n1688 VPWR.n1687 7.9105
R11411 VPWR.n1674 VPWR.n1079 7.9105
R11412 VPWR.n1663 VPWR.n1662 7.9105
R11413 VPWR.n1661 VPWR.n1660 7.9105
R11414 VPWR.n1647 VPWR.n1089 7.9105
R11415 VPWR.n1636 VPWR.n1635 7.9105
R11416 VPWR.n1634 VPWR.n1633 7.9105
R11417 VPWR.n1620 VPWR.n1099 7.9105
R11418 VPWR.n1609 VPWR.n1608 7.9105
R11419 VPWR.n1607 VPWR.n1606 7.9105
R11420 VPWR.n26 VPWR.n24 7.8627
R11421 VPWR.n7 VPWR.n6 7.56315
R11422 VPWR.n1242 VPWR.n1241 7.56315
R11423 VPWR.n1265 VPWR.n1264 7.56315
R11424 VPWR.n1289 VPWR.n1288 7.56315
R11425 VPWR.n2805 VPWR.n2803 6.4511
R11426 VPWR.n2788 VPWR.n2785 6.4511
R11427 VPWR.n2768 VPWR.n2765 6.4511
R11428 VPWR.n2749 VPWR.n2746 6.4511
R11429 VPWR.n1362 VPWR.n1339 6.4005
R11430 VPWR.n1401 VPWR.n1378 6.4005
R11431 VPWR.n1438 VPWR.n1415 6.4005
R11432 VPWR.n2723 VPWR.n2722 6.4005
R11433 VPWR.n2693 VPWR.n2692 6.4005
R11434 VPWR.n2656 VPWR.n2655 6.4005
R11435 VPWR.n2622 VPWR.n2599 6.4005
R11436 VPWR.n1595 VPWR.n1122 6.04494
R11437 VPWR.n2505 VPWR.n99 6.04494
R11438 VPWR.n1467 VPWR.n1231 6.04494
R11439 VPWR.n351 VPWR.n290 6.04494
R11440 VPWR.n2568 VPWR.n68 6.04494
R11441 VPWR.n1534 VPWR.n1153 6.04494
R11442 VPWR.n348 VPWR.n346 6.04494
R11443 VPWR.n2508 VPWR.n98 6.04494
R11444 VPWR.n965 VPWR.n963 6.04494
R11445 VPWR.n2478 VPWR.n356 6.04494
R11446 VPWR.n2475 VPWR.n357 6.04494
R11447 VPWR.n320 VPWR.n318 6.04494
R11448 VPWR.n2553 VPWR.n75 6.04494
R11449 VPWR.n973 VPWR.n971 6.04494
R11450 VPWR.n2445 VPWR.n369 6.04494
R11451 VPWR.n324 VPWR.n322 6.04494
R11452 VPWR.n2544 VPWR.n80 6.04494
R11453 VPWR.n1890 VPWR.n932 6.04494
R11454 VPWR.n1887 VPWR.n933 6.04494
R11455 VPWR.n1880 VPWR.n936 6.04494
R11456 VPWR.n389 VPWR.n387 6.04494
R11457 VPWR.n393 VPWR.n391 6.04494
R11458 VPWR.n397 VPWR.n395 6.04494
R11459 VPWR.n2455 VPWR.n365 6.04494
R11460 VPWR.n332 VPWR.n330 6.04494
R11461 VPWR.n2532 VPWR.n86 6.04494
R11462 VPWR.n1877 VPWR.n937 6.04494
R11463 VPWR.n405 VPWR.n403 6.04494
R11464 VPWR.n2458 VPWR.n364 6.04494
R11465 VPWR.n336 VPWR.n334 6.04494
R11466 VPWR.n2529 VPWR.n87 6.04494
R11467 VPWR.n2308 VPWR.n481 6.04494
R11468 VPWR.n2311 VPWR.n480 6.04494
R11469 VPWR.n2318 VPWR.n477 6.04494
R11470 VPWR.n2321 VPWR.n476 6.04494
R11471 VPWR.n2331 VPWR.n472 6.04494
R11472 VPWR.n2338 VPWR.n469 6.04494
R11473 VPWR.n2341 VPWR.n468 6.04494
R11474 VPWR.n2348 VPWR.n465 6.04494
R11475 VPWR.n2351 VPWR.n464 6.04494
R11476 VPWR.n2358 VPWR.n461 6.04494
R11477 VPWR.n2361 VPWR.n460 6.04494
R11478 VPWR.n2368 VPWR.n457 6.04494
R11479 VPWR.n2371 VPWR.n456 6.04494
R11480 VPWR.n2378 VPWR.n453 6.04494
R11481 VPWR.n2380 VPWR.n452 6.04494
R11482 VPWR.n2328 VPWR.n473 6.04494
R11483 VPWR.n543 VPWR.n482 6.04494
R11484 VPWR.n540 VPWR.n538 6.04494
R11485 VPWR.n536 VPWR.n534 6.04494
R11486 VPWR.n532 VPWR.n530 6.04494
R11487 VPWR.n524 VPWR.n522 6.04494
R11488 VPWR.n520 VPWR.n518 6.04494
R11489 VPWR.n516 VPWR.n514 6.04494
R11490 VPWR.n512 VPWR.n510 6.04494
R11491 VPWR.n508 VPWR.n506 6.04494
R11492 VPWR.n504 VPWR.n502 6.04494
R11493 VPWR.n500 VPWR.n498 6.04494
R11494 VPWR.n496 VPWR.n494 6.04494
R11495 VPWR.n492 VPWR.n490 6.04494
R11496 VPWR.n488 VPWR.n486 6.04494
R11497 VPWR.n485 VPWR.n483 6.04494
R11498 VPWR.n528 VPWR.n526 6.04494
R11499 VPWR.n2282 VPWR.n548 6.04494
R11500 VPWR.n2279 VPWR.n549 6.04494
R11501 VPWR.n2272 VPWR.n552 6.04494
R11502 VPWR.n2269 VPWR.n553 6.04494
R11503 VPWR.n2259 VPWR.n557 6.04494
R11504 VPWR.n2252 VPWR.n560 6.04494
R11505 VPWR.n2249 VPWR.n561 6.04494
R11506 VPWR.n2242 VPWR.n564 6.04494
R11507 VPWR.n2239 VPWR.n565 6.04494
R11508 VPWR.n2232 VPWR.n568 6.04494
R11509 VPWR.n2229 VPWR.n569 6.04494
R11510 VPWR.n2222 VPWR.n572 6.04494
R11511 VPWR.n2219 VPWR.n573 6.04494
R11512 VPWR.n2212 VPWR.n576 6.04494
R11513 VPWR.n2210 VPWR.n577 6.04494
R11514 VPWR.n2262 VPWR.n556 6.04494
R11515 VPWR.n581 VPWR.n579 6.04494
R11516 VPWR.n585 VPWR.n583 6.04494
R11517 VPWR.n589 VPWR.n587 6.04494
R11518 VPWR.n593 VPWR.n591 6.04494
R11519 VPWR.n601 VPWR.n599 6.04494
R11520 VPWR.n605 VPWR.n603 6.04494
R11521 VPWR.n609 VPWR.n607 6.04494
R11522 VPWR.n613 VPWR.n611 6.04494
R11523 VPWR.n617 VPWR.n615 6.04494
R11524 VPWR.n621 VPWR.n619 6.04494
R11525 VPWR.n625 VPWR.n623 6.04494
R11526 VPWR.n629 VPWR.n627 6.04494
R11527 VPWR.n633 VPWR.n631 6.04494
R11528 VPWR.n637 VPWR.n635 6.04494
R11529 VPWR.n639 VPWR.n578 6.04494
R11530 VPWR.n597 VPWR.n595 6.04494
R11531 VPWR.n2112 VPWR.n673 6.04494
R11532 VPWR.n2115 VPWR.n672 6.04494
R11533 VPWR.n2122 VPWR.n669 6.04494
R11534 VPWR.n2125 VPWR.n668 6.04494
R11535 VPWR.n2135 VPWR.n664 6.04494
R11536 VPWR.n2142 VPWR.n661 6.04494
R11537 VPWR.n2145 VPWR.n660 6.04494
R11538 VPWR.n2152 VPWR.n657 6.04494
R11539 VPWR.n2155 VPWR.n656 6.04494
R11540 VPWR.n2162 VPWR.n653 6.04494
R11541 VPWR.n2165 VPWR.n652 6.04494
R11542 VPWR.n2172 VPWR.n649 6.04494
R11543 VPWR.n2175 VPWR.n648 6.04494
R11544 VPWR.n2182 VPWR.n645 6.04494
R11545 VPWR.n2184 VPWR.n644 6.04494
R11546 VPWR.n2132 VPWR.n665 6.04494
R11547 VPWR.n735 VPWR.n674 6.04494
R11548 VPWR.n732 VPWR.n730 6.04494
R11549 VPWR.n728 VPWR.n726 6.04494
R11550 VPWR.n724 VPWR.n722 6.04494
R11551 VPWR.n716 VPWR.n714 6.04494
R11552 VPWR.n712 VPWR.n710 6.04494
R11553 VPWR.n708 VPWR.n706 6.04494
R11554 VPWR.n704 VPWR.n702 6.04494
R11555 VPWR.n700 VPWR.n698 6.04494
R11556 VPWR.n696 VPWR.n694 6.04494
R11557 VPWR.n692 VPWR.n690 6.04494
R11558 VPWR.n688 VPWR.n686 6.04494
R11559 VPWR.n684 VPWR.n682 6.04494
R11560 VPWR.n680 VPWR.n678 6.04494
R11561 VPWR.n677 VPWR.n675 6.04494
R11562 VPWR.n720 VPWR.n718 6.04494
R11563 VPWR.n2086 VPWR.n740 6.04494
R11564 VPWR.n2083 VPWR.n741 6.04494
R11565 VPWR.n2076 VPWR.n744 6.04494
R11566 VPWR.n2073 VPWR.n745 6.04494
R11567 VPWR.n2063 VPWR.n749 6.04494
R11568 VPWR.n2056 VPWR.n752 6.04494
R11569 VPWR.n2053 VPWR.n753 6.04494
R11570 VPWR.n2046 VPWR.n756 6.04494
R11571 VPWR.n2043 VPWR.n757 6.04494
R11572 VPWR.n2036 VPWR.n760 6.04494
R11573 VPWR.n2033 VPWR.n761 6.04494
R11574 VPWR.n2026 VPWR.n764 6.04494
R11575 VPWR.n2023 VPWR.n765 6.04494
R11576 VPWR.n2016 VPWR.n768 6.04494
R11577 VPWR.n2014 VPWR.n769 6.04494
R11578 VPWR.n2066 VPWR.n748 6.04494
R11579 VPWR.n773 VPWR.n771 6.04494
R11580 VPWR.n777 VPWR.n775 6.04494
R11581 VPWR.n781 VPWR.n779 6.04494
R11582 VPWR.n785 VPWR.n783 6.04494
R11583 VPWR.n793 VPWR.n791 6.04494
R11584 VPWR.n797 VPWR.n795 6.04494
R11585 VPWR.n801 VPWR.n799 6.04494
R11586 VPWR.n805 VPWR.n803 6.04494
R11587 VPWR.n809 VPWR.n807 6.04494
R11588 VPWR.n813 VPWR.n811 6.04494
R11589 VPWR.n817 VPWR.n815 6.04494
R11590 VPWR.n821 VPWR.n819 6.04494
R11591 VPWR.n825 VPWR.n823 6.04494
R11592 VPWR.n829 VPWR.n827 6.04494
R11593 VPWR.n831 VPWR.n770 6.04494
R11594 VPWR.n789 VPWR.n787 6.04494
R11595 VPWR.n1916 VPWR.n865 6.04494
R11596 VPWR.n1919 VPWR.n864 6.04494
R11597 VPWR.n1926 VPWR.n861 6.04494
R11598 VPWR.n1929 VPWR.n860 6.04494
R11599 VPWR.n1939 VPWR.n856 6.04494
R11600 VPWR.n1946 VPWR.n853 6.04494
R11601 VPWR.n1949 VPWR.n852 6.04494
R11602 VPWR.n1956 VPWR.n849 6.04494
R11603 VPWR.n1959 VPWR.n848 6.04494
R11604 VPWR.n1966 VPWR.n845 6.04494
R11605 VPWR.n1969 VPWR.n844 6.04494
R11606 VPWR.n1976 VPWR.n841 6.04494
R11607 VPWR.n1979 VPWR.n840 6.04494
R11608 VPWR.n1986 VPWR.n837 6.04494
R11609 VPWR.n1988 VPWR.n836 6.04494
R11610 VPWR.n1936 VPWR.n857 6.04494
R11611 VPWR.n927 VPWR.n866 6.04494
R11612 VPWR.n924 VPWR.n922 6.04494
R11613 VPWR.n920 VPWR.n918 6.04494
R11614 VPWR.n916 VPWR.n914 6.04494
R11615 VPWR.n908 VPWR.n906 6.04494
R11616 VPWR.n904 VPWR.n902 6.04494
R11617 VPWR.n900 VPWR.n898 6.04494
R11618 VPWR.n896 VPWR.n894 6.04494
R11619 VPWR.n892 VPWR.n890 6.04494
R11620 VPWR.n888 VPWR.n886 6.04494
R11621 VPWR.n884 VPWR.n882 6.04494
R11622 VPWR.n880 VPWR.n878 6.04494
R11623 VPWR.n876 VPWR.n874 6.04494
R11624 VPWR.n872 VPWR.n870 6.04494
R11625 VPWR.n869 VPWR.n867 6.04494
R11626 VPWR.n912 VPWR.n910 6.04494
R11627 VPWR.n1870 VPWR.n940 6.04494
R11628 VPWR.n981 VPWR.n979 6.04494
R11629 VPWR.n1494 VPWR.n1227 6.04494
R11630 VPWR.n1221 VPWR.n1179 6.04494
R11631 VPWR.n401 VPWR.n399 6.04494
R11632 VPWR.n2465 VPWR.n361 6.04494
R11633 VPWR.n340 VPWR.n338 6.04494
R11634 VPWR.n2520 VPWR.n92 6.04494
R11635 VPWR.n977 VPWR.n975 6.04494
R11636 VPWR.n1491 VPWR.n1485 6.04494
R11637 VPWR.n1184 VPWR.n1183 6.04494
R11638 VPWR.n1867 VPWR.n941 6.04494
R11639 VPWR.n985 VPWR.n983 6.04494
R11640 VPWR.n1505 VPWR.n1173 6.04494
R11641 VPWR.n1218 VPWR.n1217 6.04494
R11642 VPWR.n409 VPWR.n407 6.04494
R11643 VPWR.n417 VPWR.n415 6.04494
R11644 VPWR.n421 VPWR.n419 6.04494
R11645 VPWR.n425 VPWR.n423 6.04494
R11646 VPWR.n429 VPWR.n427 6.04494
R11647 VPWR.n433 VPWR.n431 6.04494
R11648 VPWR.n437 VPWR.n435 6.04494
R11649 VPWR.n441 VPWR.n439 6.04494
R11650 VPWR.n445 VPWR.n443 6.04494
R11651 VPWR.n447 VPWR.n386 6.04494
R11652 VPWR.n413 VPWR.n411 6.04494
R11653 VPWR.n2448 VPWR.n368 6.04494
R11654 VPWR.n328 VPWR.n326 6.04494
R11655 VPWR.n2541 VPWR.n81 6.04494
R11656 VPWR.n989 VPWR.n987 6.04494
R11657 VPWR.n1508 VPWR.n1169 6.04494
R11658 VPWR.n1215 VPWR.n1214 6.04494
R11659 VPWR.n1860 VPWR.n944 6.04494
R11660 VPWR.n1850 VPWR.n948 6.04494
R11661 VPWR.n1847 VPWR.n949 6.04494
R11662 VPWR.n1840 VPWR.n952 6.04494
R11663 VPWR.n1837 VPWR.n953 6.04494
R11664 VPWR.n1830 VPWR.n956 6.04494
R11665 VPWR.n1827 VPWR.n957 6.04494
R11666 VPWR.n1820 VPWR.n960 6.04494
R11667 VPWR.n1818 VPWR.n961 6.04494
R11668 VPWR.n1857 VPWR.n945 6.04494
R11669 VPWR.n993 VPWR.n991 6.04494
R11670 VPWR.n1519 VPWR.n1163 6.04494
R11671 VPWR.n1212 VPWR.n1206 6.04494
R11672 VPWR.n2468 VPWR.n360 6.04494
R11673 VPWR.n344 VPWR.n342 6.04494
R11674 VPWR.n2517 VPWR.n93 6.04494
R11675 VPWR.n1480 VPWR.n1479 6.04494
R11676 VPWR.n1181 VPWR.n1180 6.04494
R11677 VPWR.n997 VPWR.n995 6.04494
R11678 VPWR.n1522 VPWR.n1159 6.04494
R11679 VPWR.n1204 VPWR.n1203 6.04494
R11680 VPWR.n2438 VPWR.n372 6.04494
R11681 VPWR.n2428 VPWR.n376 6.04494
R11682 VPWR.n2425 VPWR.n377 6.04494
R11683 VPWR.n2418 VPWR.n380 6.04494
R11684 VPWR.n2415 VPWR.n381 6.04494
R11685 VPWR.n2408 VPWR.n384 6.04494
R11686 VPWR.n2406 VPWR.n385 6.04494
R11687 VPWR.n2435 VPWR.n373 6.04494
R11688 VPWR.n316 VPWR.n314 6.04494
R11689 VPWR.n2556 VPWR.n74 6.04494
R11690 VPWR.n1537 VPWR.n1149 6.04494
R11691 VPWR.n1201 VPWR.n1200 6.04494
R11692 VPWR.n1001 VPWR.n999 6.04494
R11693 VPWR.n1005 VPWR.n1003 6.04494
R11694 VPWR.n1009 VPWR.n1007 6.04494
R11695 VPWR.n1013 VPWR.n1011 6.04494
R11696 VPWR.n1017 VPWR.n1015 6.04494
R11697 VPWR.n1021 VPWR.n1019 6.04494
R11698 VPWR.n1023 VPWR.n962 6.04494
R11699 VPWR.n969 VPWR.n967 6.04494
R11700 VPWR.n1474 VPWR.n1472 6.04494
R11701 VPWR.n1592 VPWR.n1123 6.04494
R11702 VPWR.n312 VPWR.n310 6.04494
R11703 VPWR.n2565 VPWR.n69 6.04494
R11704 VPWR.n1198 VPWR.n1192 6.04494
R11705 VPWR.n1762 VPWR.n1049 6.04494
R11706 VPWR.n1190 VPWR.n1189 6.04494
R11707 VPWR.n308 VPWR.n306 6.04494
R11708 VPWR.n304 VPWR.n302 6.04494
R11709 VPWR.n296 VPWR.n294 6.04494
R11710 VPWR.n293 VPWR.n291 6.04494
R11711 VPWR.n300 VPWR.n298 6.04494
R11712 VPWR.n1741 VPWR.n1058 6.04494
R11713 VPWR.n1750 VPWR.n1748 6.04494
R11714 VPWR.n1790 VPWR.n1036 6.04494
R11715 VPWR.n1792 VPWR.n1032 6.04494
R11716 VPWR.n1759 VPWR.n1053 6.04494
R11717 VPWR.n1187 VPWR.n1186 6.04494
R11718 VPWR.n2577 VPWR.n63 6.04494
R11719 VPWR.n2580 VPWR.n62 6.04494
R11720 VPWR.n2589 VPWR.n57 6.04494
R11721 VPWR.n2591 VPWR.n56 6.04494
R11722 VPWR.n1738 VPWR.n1059 6.04494
R11723 VPWR.n1062 VPWR.n1061 6.04494
R11724 VPWR.n2785 VPWR.n2784 5.39628
R11725 VPWR.n2765 VPWR.n2764 5.39628
R11726 VPWR.n2746 VPWR.n2745 5.39628
R11727 VPWR.n54 VPWR 4.72593
R11728 VPWR.n52 VPWR 4.72593
R11729 VPWR.n50 VPWR 4.72593
R11730 VPWR.n48 VPWR 4.72593
R11731 VPWR.n46 VPWR 4.72593
R11732 VPWR.n44 VPWR 4.72593
R11733 VPWR.n42 VPWR 4.72593
R11734 VPWR.n40 VPWR 4.72593
R11735 VPWR.n38 VPWR 4.72593
R11736 VPWR.n36 VPWR 4.72593
R11737 VPWR.n34 VPWR 4.72593
R11738 VPWR.n32 VPWR 4.72593
R11739 VPWR.n30 VPWR 4.72593
R11740 VPWR.n28 VPWR 4.72593
R11741 VPWR.n26 VPWR 4.72593
R11742 VPWR.n1446 VPWR.n1445 4.55954
R11743 VPWR.n2571 VPWR.n2570 4.5005
R11744 VPWR.n2511 VPWR.n2510 4.5005
R11745 VPWR.n2551 VPWR.n2550 4.5005
R11746 VPWR.n319 VPWR.n77 4.5005
R11747 VPWR.n2547 VPWR.n2546 4.5005
R11748 VPWR.n323 VPWR.n78 4.5005
R11749 VPWR.n2535 VPWR.n2534 4.5005
R11750 VPWR.n331 VPWR.n84 4.5005
R11751 VPWR.n2454 VPWR.n2453 4.5005
R11752 VPWR.n2527 VPWR.n2526 4.5005
R11753 VPWR.n335 VPWR.n89 4.5005
R11754 VPWR.n2460 VPWR.n2459 4.5005
R11755 VPWR.n1498 VPWR.n1223 4.5005
R11756 VPWR.n1497 VPWR.n1495 4.5005
R11757 VPWR.n980 VPWR.n939 4.5005
R11758 VPWR.n1872 VPWR.n1871 4.5005
R11759 VPWR.n911 VPWR.n858 4.5005
R11760 VPWR.n1935 VPWR.n1934 4.5005
R11761 VPWR.n788 VPWR.n747 4.5005
R11762 VPWR.n2068 VPWR.n2067 4.5005
R11763 VPWR.n719 VPWR.n666 4.5005
R11764 VPWR.n2131 VPWR.n2130 4.5005
R11765 VPWR.n596 VPWR.n555 4.5005
R11766 VPWR.n2264 VPWR.n2263 4.5005
R11767 VPWR.n527 VPWR.n474 4.5005
R11768 VPWR.n2327 VPWR.n2326 4.5005
R11769 VPWR.n404 VPWR.n363 4.5005
R11770 VPWR.n2523 VPWR.n2522 4.5005
R11771 VPWR.n339 VPWR.n90 4.5005
R11772 VPWR.n2464 VPWR.n2463 4.5005
R11773 VPWR.n400 VPWR.n362 4.5005
R11774 VPWR.n2323 VPWR.n2322 4.5005
R11775 VPWR.n531 VPWR.n475 4.5005
R11776 VPWR.n2268 VPWR.n2267 4.5005
R11777 VPWR.n592 VPWR.n554 4.5005
R11778 VPWR.n2127 VPWR.n2126 4.5005
R11779 VPWR.n723 VPWR.n667 4.5005
R11780 VPWR.n2072 VPWR.n2071 4.5005
R11781 VPWR.n784 VPWR.n746 4.5005
R11782 VPWR.n1931 VPWR.n1930 4.5005
R11783 VPWR.n915 VPWR.n859 4.5005
R11784 VPWR.n1488 VPWR.n1486 4.5005
R11785 VPWR.n1490 VPWR.n1489 4.5005
R11786 VPWR.n976 VPWR.n938 4.5005
R11787 VPWR.n1876 VPWR.n1875 4.5005
R11788 VPWR.n1501 VPWR.n1174 4.5005
R11789 VPWR.n1504 VPWR.n1503 4.5005
R11790 VPWR.n984 VPWR.n942 4.5005
R11791 VPWR.n1866 VPWR.n1865 4.5005
R11792 VPWR.n907 VPWR.n855 4.5005
R11793 VPWR.n1941 VPWR.n1940 4.5005
R11794 VPWR.n792 VPWR.n750 4.5005
R11795 VPWR.n2062 VPWR.n2061 4.5005
R11796 VPWR.n715 VPWR.n663 4.5005
R11797 VPWR.n2137 VPWR.n2136 4.5005
R11798 VPWR.n600 VPWR.n558 4.5005
R11799 VPWR.n2258 VPWR.n2257 4.5005
R11800 VPWR.n523 VPWR.n471 4.5005
R11801 VPWR.n2333 VPWR.n2332 4.5005
R11802 VPWR.n408 VPWR.n366 4.5005
R11803 VPWR.n2539 VPWR.n2538 4.5005
R11804 VPWR.n327 VPWR.n83 4.5005
R11805 VPWR.n2450 VPWR.n2449 4.5005
R11806 VPWR.n412 VPWR.n367 4.5005
R11807 VPWR.n2337 VPWR.n2336 4.5005
R11808 VPWR.n519 VPWR.n470 4.5005
R11809 VPWR.n2254 VPWR.n2253 4.5005
R11810 VPWR.n604 VPWR.n559 4.5005
R11811 VPWR.n2141 VPWR.n2140 4.5005
R11812 VPWR.n711 VPWR.n662 4.5005
R11813 VPWR.n2058 VPWR.n2057 4.5005
R11814 VPWR.n796 VPWR.n751 4.5005
R11815 VPWR.n1945 VPWR.n1944 4.5005
R11816 VPWR.n903 VPWR.n854 4.5005
R11817 VPWR.n1512 VPWR.n1165 4.5005
R11818 VPWR.n1511 VPWR.n1509 4.5005
R11819 VPWR.n988 VPWR.n943 4.5005
R11820 VPWR.n1862 VPWR.n1861 4.5005
R11821 VPWR.n1515 VPWR.n1164 4.5005
R11822 VPWR.n1518 VPWR.n1517 4.5005
R11823 VPWR.n992 VPWR.n946 4.5005
R11824 VPWR.n1856 VPWR.n1855 4.5005
R11825 VPWR.n899 VPWR.n851 4.5005
R11826 VPWR.n1951 VPWR.n1950 4.5005
R11827 VPWR.n800 VPWR.n754 4.5005
R11828 VPWR.n2052 VPWR.n2051 4.5005
R11829 VPWR.n707 VPWR.n659 4.5005
R11830 VPWR.n2147 VPWR.n2146 4.5005
R11831 VPWR.n608 VPWR.n562 4.5005
R11832 VPWR.n2248 VPWR.n2247 4.5005
R11833 VPWR.n515 VPWR.n467 4.5005
R11834 VPWR.n2343 VPWR.n2342 4.5005
R11835 VPWR.n416 VPWR.n370 4.5005
R11836 VPWR.n2444 VPWR.n2443 4.5005
R11837 VPWR.n2515 VPWR.n2514 4.5005
R11838 VPWR.n343 VPWR.n95 4.5005
R11839 VPWR.n2470 VPWR.n2469 4.5005
R11840 VPWR.n396 VPWR.n359 4.5005
R11841 VPWR.n2317 VPWR.n2316 4.5005
R11842 VPWR.n535 VPWR.n478 4.5005
R11843 VPWR.n2274 VPWR.n2273 4.5005
R11844 VPWR.n588 VPWR.n551 4.5005
R11845 VPWR.n2121 VPWR.n2120 4.5005
R11846 VPWR.n727 VPWR.n670 4.5005
R11847 VPWR.n2078 VPWR.n2077 4.5005
R11848 VPWR.n780 VPWR.n743 4.5005
R11849 VPWR.n1925 VPWR.n1924 4.5005
R11850 VPWR.n919 VPWR.n862 4.5005
R11851 VPWR.n1882 VPWR.n1881 4.5005
R11852 VPWR.n1586 VPWR.n1129 4.5005
R11853 VPWR.n1585 VPWR.n1130 4.5005
R11854 VPWR.n972 VPWR.n935 4.5005
R11855 VPWR.n1526 VPWR.n1155 4.5005
R11856 VPWR.n1525 VPWR.n1523 4.5005
R11857 VPWR.n996 VPWR.n947 4.5005
R11858 VPWR.n1852 VPWR.n1851 4.5005
R11859 VPWR.n895 VPWR.n850 4.5005
R11860 VPWR.n1955 VPWR.n1954 4.5005
R11861 VPWR.n804 VPWR.n755 4.5005
R11862 VPWR.n2048 VPWR.n2047 4.5005
R11863 VPWR.n703 VPWR.n658 4.5005
R11864 VPWR.n2151 VPWR.n2150 4.5005
R11865 VPWR.n612 VPWR.n563 4.5005
R11866 VPWR.n2244 VPWR.n2243 4.5005
R11867 VPWR.n511 VPWR.n466 4.5005
R11868 VPWR.n2347 VPWR.n2346 4.5005
R11869 VPWR.n420 VPWR.n371 4.5005
R11870 VPWR.n2440 VPWR.n2439 4.5005
R11871 VPWR.n2559 VPWR.n2558 4.5005
R11872 VPWR.n315 VPWR.n72 4.5005
R11873 VPWR.n2434 VPWR.n2433 4.5005
R11874 VPWR.n424 VPWR.n374 4.5005
R11875 VPWR.n2353 VPWR.n2352 4.5005
R11876 VPWR.n507 VPWR.n463 4.5005
R11877 VPWR.n2238 VPWR.n2237 4.5005
R11878 VPWR.n616 VPWR.n566 4.5005
R11879 VPWR.n2157 VPWR.n2156 4.5005
R11880 VPWR.n699 VPWR.n655 4.5005
R11881 VPWR.n2042 VPWR.n2041 4.5005
R11882 VPWR.n808 VPWR.n758 4.5005
R11883 VPWR.n1961 VPWR.n1960 4.5005
R11884 VPWR.n891 VPWR.n847 4.5005
R11885 VPWR.n1846 VPWR.n1845 4.5005
R11886 VPWR.n1145 VPWR.n1144 4.5005
R11887 VPWR.n1539 VPWR.n1538 4.5005
R11888 VPWR.n1000 VPWR.n950 4.5005
R11889 VPWR.n1590 VPWR.n1589 4.5005
R11890 VPWR.n1473 VPWR.n1128 4.5005
R11891 VPWR.n968 VPWR.n934 4.5005
R11892 VPWR.n1886 VPWR.n1885 4.5005
R11893 VPWR.n923 VPWR.n863 4.5005
R11894 VPWR.n1921 VPWR.n1920 4.5005
R11895 VPWR.n776 VPWR.n742 4.5005
R11896 VPWR.n2082 VPWR.n2081 4.5005
R11897 VPWR.n731 VPWR.n671 4.5005
R11898 VPWR.n2117 VPWR.n2116 4.5005
R11899 VPWR.n584 VPWR.n550 4.5005
R11900 VPWR.n2278 VPWR.n2277 4.5005
R11901 VPWR.n539 VPWR.n479 4.5005
R11902 VPWR.n2313 VPWR.n2312 4.5005
R11903 VPWR.n392 VPWR.n358 4.5005
R11904 VPWR.n2474 VPWR.n2473 4.5005
R11905 VPWR.n347 VPWR.n96 4.5005
R11906 VPWR.n2563 VPWR.n2562 4.5005
R11907 VPWR.n311 VPWR.n71 4.5005
R11908 VPWR.n2430 VPWR.n2429 4.5005
R11909 VPWR.n428 VPWR.n375 4.5005
R11910 VPWR.n2357 VPWR.n2356 4.5005
R11911 VPWR.n503 VPWR.n462 4.5005
R11912 VPWR.n2234 VPWR.n2233 4.5005
R11913 VPWR.n620 VPWR.n567 4.5005
R11914 VPWR.n2161 VPWR.n2160 4.5005
R11915 VPWR.n695 VPWR.n654 4.5005
R11916 VPWR.n2038 VPWR.n2037 4.5005
R11917 VPWR.n812 VPWR.n759 4.5005
R11918 VPWR.n1965 VPWR.n1964 4.5005
R11919 VPWR.n887 VPWR.n846 4.5005
R11920 VPWR.n1842 VPWR.n1841 4.5005
R11921 VPWR.n1004 VPWR.n951 4.5005
R11922 VPWR.n1531 VPWR.n1154 4.5005
R11923 VPWR.n1533 VPWR.n1532 4.5005
R11924 VPWR.n1073 VPWR.n1045 4.5005
R11925 VPWR.n1764 VPWR.n1763 4.5005
R11926 VPWR.n1008 VPWR.n954 4.5005
R11927 VPWR.n1836 VPWR.n1835 4.5005
R11928 VPWR.n883 VPWR.n843 4.5005
R11929 VPWR.n1971 VPWR.n1970 4.5005
R11930 VPWR.n816 VPWR.n762 4.5005
R11931 VPWR.n2032 VPWR.n2031 4.5005
R11932 VPWR.n691 VPWR.n651 4.5005
R11933 VPWR.n2167 VPWR.n2166 4.5005
R11934 VPWR.n624 VPWR.n570 4.5005
R11935 VPWR.n2228 VPWR.n2227 4.5005
R11936 VPWR.n499 VPWR.n459 4.5005
R11937 VPWR.n2363 VPWR.n2362 4.5005
R11938 VPWR.n432 VPWR.n378 4.5005
R11939 VPWR.n2424 VPWR.n2423 4.5005
R11940 VPWR.n307 VPWR.n66 4.5005
R11941 VPWR.n299 VPWR.n60 4.5005
R11942 VPWR.n2414 VPWR.n2413 4.5005
R11943 VPWR.n440 VPWR.n382 4.5005
R11944 VPWR.n2373 VPWR.n2372 4.5005
R11945 VPWR.n491 VPWR.n455 4.5005
R11946 VPWR.n2218 VPWR.n2217 4.5005
R11947 VPWR.n632 VPWR.n574 4.5005
R11948 VPWR.n2177 VPWR.n2176 4.5005
R11949 VPWR.n683 VPWR.n647 4.5005
R11950 VPWR.n2022 VPWR.n2021 4.5005
R11951 VPWR.n824 VPWR.n766 4.5005
R11952 VPWR.n1981 VPWR.n1980 4.5005
R11953 VPWR.n875 VPWR.n839 4.5005
R11954 VPWR.n1826 VPWR.n1825 4.5005
R11955 VPWR.n1016 VPWR.n958 4.5005
R11956 VPWR.n1753 VPWR.n1743 4.5005
R11957 VPWR.n1752 VPWR.n1751 4.5005
R11958 VPWR.n1756 VPWR.n1054 4.5005
R11959 VPWR.n1758 VPWR.n1757 4.5005
R11960 VPWR.n1012 VPWR.n955 4.5005
R11961 VPWR.n1832 VPWR.n1831 4.5005
R11962 VPWR.n879 VPWR.n842 4.5005
R11963 VPWR.n1975 VPWR.n1974 4.5005
R11964 VPWR.n820 VPWR.n763 4.5005
R11965 VPWR.n2028 VPWR.n2027 4.5005
R11966 VPWR.n687 VPWR.n650 4.5005
R11967 VPWR.n2171 VPWR.n2170 4.5005
R11968 VPWR.n628 VPWR.n571 4.5005
R11969 VPWR.n2224 VPWR.n2223 4.5005
R11970 VPWR.n495 VPWR.n458 4.5005
R11971 VPWR.n2367 VPWR.n2366 4.5005
R11972 VPWR.n436 VPWR.n379 4.5005
R11973 VPWR.n2420 VPWR.n2419 4.5005
R11974 VPWR.n303 VPWR.n65 4.5005
R11975 VPWR.n2575 VPWR.n2574 4.5005
R11976 VPWR.n2583 VPWR.n2582 4.5005
R11977 VPWR.n2587 VPWR.n2586 4.5005
R11978 VPWR.n295 VPWR.n59 4.5005
R11979 VPWR.n2410 VPWR.n2409 4.5005
R11980 VPWR.n444 VPWR.n383 4.5005
R11981 VPWR.n2377 VPWR.n2376 4.5005
R11982 VPWR.n487 VPWR.n454 4.5005
R11983 VPWR.n2214 VPWR.n2213 4.5005
R11984 VPWR.n636 VPWR.n575 4.5005
R11985 VPWR.n2181 VPWR.n2180 4.5005
R11986 VPWR.n679 VPWR.n646 4.5005
R11987 VPWR.n2018 VPWR.n2017 4.5005
R11988 VPWR.n828 VPWR.n767 4.5005
R11989 VPWR.n1985 VPWR.n1984 4.5005
R11990 VPWR.n871 VPWR.n838 4.5005
R11991 VPWR.n1822 VPWR.n1821 4.5005
R11992 VPWR.n1020 VPWR.n959 4.5005
R11993 VPWR.n1789 VPWR.n1788 4.5005
R11994 VPWR.n1736 VPWR.n1037 4.5005
R11995 VPWR.n1232 VPWR.n1121 4.5005
R11996 VPWR.n1466 VPWR.n1465 4.5005
R11997 VPWR.n964 VPWR.n931 4.5005
R11998 VPWR.n1892 VPWR.n1891 4.5005
R11999 VPWR.n929 VPWR.n928 4.5005
R12000 VPWR.n1915 VPWR.n1914 4.5005
R12001 VPWR.n772 VPWR.n739 4.5005
R12002 VPWR.n2088 VPWR.n2087 4.5005
R12003 VPWR.n737 VPWR.n736 4.5005
R12004 VPWR.n2111 VPWR.n2110 4.5005
R12005 VPWR.n580 VPWR.n547 4.5005
R12006 VPWR.n2284 VPWR.n2283 4.5005
R12007 VPWR.n545 VPWR.n544 4.5005
R12008 VPWR.n2307 VPWR.n2306 4.5005
R12009 VPWR.n388 VPWR.n355 4.5005
R12010 VPWR.n2480 VPWR.n2479 4.5005
R12011 VPWR.n353 VPWR.n352 4.5005
R12012 VPWR.n2503 VPWR.n2502 4.5005
R12013 VPWR.n2594 VPWR.n2593 4.5005
R12014 VPWR.n292 VPWR.n22 4.5005
R12015 VPWR.n2405 VPWR.n2404 4.5005
R12016 VPWR.n449 VPWR.n448 4.5005
R12017 VPWR.n2382 VPWR.n2381 4.5005
R12018 VPWR.n484 VPWR.n451 4.5005
R12019 VPWR.n2209 VPWR.n2208 4.5005
R12020 VPWR.n641 VPWR.n640 4.5005
R12021 VPWR.n2186 VPWR.n2185 4.5005
R12022 VPWR.n676 VPWR.n643 4.5005
R12023 VPWR.n2013 VPWR.n2012 4.5005
R12024 VPWR.n833 VPWR.n832 4.5005
R12025 VPWR.n1990 VPWR.n1989 4.5005
R12026 VPWR.n868 VPWR.n835 4.5005
R12027 VPWR.n1817 VPWR.n1816 4.5005
R12028 VPWR.n1025 VPWR.n1024 4.5005
R12029 VPWR.n1794 VPWR.n1793 4.5005
R12030 VPWR.n1060 VPWR.n1028 4.5005
R12031 VPWR.n2628 VPWR 4.49965
R12032 VPWR.n19 VPWR.n18 4.20017
R12033 VPWR.n1255 VPWR.n1254 4.20017
R12034 VPWR.n1279 VPWR.n1278 4.20017
R12035 VPWR.n1302 VPWR.n1301 4.20017
R12036 VPWR.n1337 VPWR.n1336 4.20017
R12037 VPWR.n1376 VPWR.n1375 4.20017
R12038 VPWR.n1414 VPWR.n1413 4.20017
R12039 VPWR.n2813 VPWR 4.14027
R12040 VPWR.n2797 VPWR 4.14027
R12041 VPWR.n2778 VPWR 4.14027
R12042 VPWR.n2758 VPWR 4.14027
R12043 VPWR.n2739 VPWR 4.14027
R12044 VPWR.n2703 VPWR 4.14027
R12045 VPWR.n2665 VPWR 4.14027
R12046 VPWR.n55 VPWR.n54 4.0005
R12047 VPWR.n2716 VPWR.n2713 3.76521
R12048 VPWR.n2680 VPWR.n2676 3.76521
R12049 VPWR.n2643 VPWR.n2639 3.76521
R12050 VPWR.n2611 VPWR.n2610 3.76521
R12051 VPWR.n1906 VPWR.n858 3.4105
R12052 VPWR.n1934 VPWR.n1933 3.4105
R12053 VPWR.n1997 VPWR.n747 3.4105
R12054 VPWR.n2069 VPWR.n2068 3.4105
R12055 VPWR.n2102 VPWR.n666 3.4105
R12056 VPWR.n2130 VPWR.n2129 3.4105
R12057 VPWR.n2193 VPWR.n555 3.4105
R12058 VPWR.n2265 VPWR.n2264 3.4105
R12059 VPWR.n2298 VPWR.n474 3.4105
R12060 VPWR.n2326 VPWR.n2325 3.4105
R12061 VPWR.n2389 VPWR.n363 3.4105
R12062 VPWR.n2388 VPWR.n362 3.4105
R12063 VPWR.n2324 VPWR.n2323 3.4105
R12064 VPWR.n2299 VPWR.n475 3.4105
R12065 VPWR.n2267 VPWR.n2266 3.4105
R12066 VPWR.n2192 VPWR.n554 3.4105
R12067 VPWR.n2128 VPWR.n2127 3.4105
R12068 VPWR.n2103 VPWR.n667 3.4105
R12069 VPWR.n2071 VPWR.n2070 3.4105
R12070 VPWR.n1996 VPWR.n746 3.4105
R12071 VPWR.n1932 VPWR.n1931 3.4105
R12072 VPWR.n1907 VPWR.n859 3.4105
R12073 VPWR.n1875 VPWR.n1874 3.4105
R12074 VPWR.n1873 VPWR.n1872 3.4105
R12075 VPWR.n1865 VPWR.n1864 3.4105
R12076 VPWR.n1905 VPWR.n855 3.4105
R12077 VPWR.n1942 VPWR.n1941 3.4105
R12078 VPWR.n1998 VPWR.n750 3.4105
R12079 VPWR.n2061 VPWR.n2060 3.4105
R12080 VPWR.n2101 VPWR.n663 3.4105
R12081 VPWR.n2138 VPWR.n2137 3.4105
R12082 VPWR.n2194 VPWR.n558 3.4105
R12083 VPWR.n2257 VPWR.n2256 3.4105
R12084 VPWR.n2297 VPWR.n471 3.4105
R12085 VPWR.n2334 VPWR.n2333 3.4105
R12086 VPWR.n2390 VPWR.n366 3.4105
R12087 VPWR.n2391 VPWR.n367 3.4105
R12088 VPWR.n2336 VPWR.n2335 3.4105
R12089 VPWR.n2296 VPWR.n470 3.4105
R12090 VPWR.n2255 VPWR.n2254 3.4105
R12091 VPWR.n2195 VPWR.n559 3.4105
R12092 VPWR.n2140 VPWR.n2139 3.4105
R12093 VPWR.n2100 VPWR.n662 3.4105
R12094 VPWR.n2059 VPWR.n2058 3.4105
R12095 VPWR.n1999 VPWR.n751 3.4105
R12096 VPWR.n1944 VPWR.n1943 3.4105
R12097 VPWR.n1904 VPWR.n854 3.4105
R12098 VPWR.n1863 VPWR.n1862 3.4105
R12099 VPWR.n1855 VPWR.n1854 3.4105
R12100 VPWR.n1903 VPWR.n851 3.4105
R12101 VPWR.n1952 VPWR.n1951 3.4105
R12102 VPWR.n2000 VPWR.n754 3.4105
R12103 VPWR.n2051 VPWR.n2050 3.4105
R12104 VPWR.n2099 VPWR.n659 3.4105
R12105 VPWR.n2148 VPWR.n2147 3.4105
R12106 VPWR.n2196 VPWR.n562 3.4105
R12107 VPWR.n2247 VPWR.n2246 3.4105
R12108 VPWR.n2295 VPWR.n467 3.4105
R12109 VPWR.n2344 VPWR.n2343 3.4105
R12110 VPWR.n2392 VPWR.n370 3.4105
R12111 VPWR.n2443 VPWR.n2442 3.4105
R12112 VPWR.n2451 VPWR.n2450 3.4105
R12113 VPWR.n2453 VPWR.n2452 3.4105
R12114 VPWR.n2461 VPWR.n2460 3.4105
R12115 VPWR.n2463 VPWR.n2462 3.4105
R12116 VPWR.n2471 VPWR.n2470 3.4105
R12117 VPWR.n2387 VPWR.n359 3.4105
R12118 VPWR.n2316 VPWR.n2315 3.4105
R12119 VPWR.n2300 VPWR.n478 3.4105
R12120 VPWR.n2275 VPWR.n2274 3.4105
R12121 VPWR.n2191 VPWR.n551 3.4105
R12122 VPWR.n2120 VPWR.n2119 3.4105
R12123 VPWR.n2104 VPWR.n670 3.4105
R12124 VPWR.n2079 VPWR.n2078 3.4105
R12125 VPWR.n1995 VPWR.n743 3.4105
R12126 VPWR.n1924 VPWR.n1923 3.4105
R12127 VPWR.n1908 VPWR.n862 3.4105
R12128 VPWR.n1883 VPWR.n1882 3.4105
R12129 VPWR.n1799 VPWR.n935 3.4105
R12130 VPWR.n1800 VPWR.n938 3.4105
R12131 VPWR.n1801 VPWR.n939 3.4105
R12132 VPWR.n1802 VPWR.n942 3.4105
R12133 VPWR.n1803 VPWR.n943 3.4105
R12134 VPWR.n1804 VPWR.n946 3.4105
R12135 VPWR.n1805 VPWR.n947 3.4105
R12136 VPWR.n1853 VPWR.n1852 3.4105
R12137 VPWR.n1902 VPWR.n850 3.4105
R12138 VPWR.n1954 VPWR.n1953 3.4105
R12139 VPWR.n2001 VPWR.n755 3.4105
R12140 VPWR.n2049 VPWR.n2048 3.4105
R12141 VPWR.n2098 VPWR.n658 3.4105
R12142 VPWR.n2150 VPWR.n2149 3.4105
R12143 VPWR.n2197 VPWR.n563 3.4105
R12144 VPWR.n2245 VPWR.n2244 3.4105
R12145 VPWR.n2294 VPWR.n466 3.4105
R12146 VPWR.n2346 VPWR.n2345 3.4105
R12147 VPWR.n2393 VPWR.n371 3.4105
R12148 VPWR.n2441 VPWR.n2440 3.4105
R12149 VPWR.n2433 VPWR.n2432 3.4105
R12150 VPWR.n2394 VPWR.n374 3.4105
R12151 VPWR.n2354 VPWR.n2353 3.4105
R12152 VPWR.n2293 VPWR.n463 3.4105
R12153 VPWR.n2237 VPWR.n2236 3.4105
R12154 VPWR.n2198 VPWR.n566 3.4105
R12155 VPWR.n2158 VPWR.n2157 3.4105
R12156 VPWR.n2097 VPWR.n655 3.4105
R12157 VPWR.n2041 VPWR.n2040 3.4105
R12158 VPWR.n2002 VPWR.n758 3.4105
R12159 VPWR.n1962 VPWR.n1961 3.4105
R12160 VPWR.n1901 VPWR.n847 3.4105
R12161 VPWR.n1845 VPWR.n1844 3.4105
R12162 VPWR.n1806 VPWR.n950 3.4105
R12163 VPWR.n1798 VPWR.n934 3.4105
R12164 VPWR.n1885 VPWR.n1884 3.4105
R12165 VPWR.n1909 VPWR.n863 3.4105
R12166 VPWR.n1922 VPWR.n1921 3.4105
R12167 VPWR.n1994 VPWR.n742 3.4105
R12168 VPWR.n2081 VPWR.n2080 3.4105
R12169 VPWR.n2105 VPWR.n671 3.4105
R12170 VPWR.n2118 VPWR.n2117 3.4105
R12171 VPWR.n2190 VPWR.n550 3.4105
R12172 VPWR.n2277 VPWR.n2276 3.4105
R12173 VPWR.n2301 VPWR.n479 3.4105
R12174 VPWR.n2314 VPWR.n2313 3.4105
R12175 VPWR.n2386 VPWR.n358 3.4105
R12176 VPWR.n2473 VPWR.n2472 3.4105
R12177 VPWR.n2497 VPWR.n96 3.4105
R12178 VPWR.n2496 VPWR.n95 3.4105
R12179 VPWR.n2495 VPWR.n90 3.4105
R12180 VPWR.n2494 VPWR.n89 3.4105
R12181 VPWR.n2493 VPWR.n84 3.4105
R12182 VPWR.n2492 VPWR.n83 3.4105
R12183 VPWR.n2491 VPWR.n78 3.4105
R12184 VPWR.n2490 VPWR.n77 3.4105
R12185 VPWR.n2489 VPWR.n72 3.4105
R12186 VPWR.n2488 VPWR.n71 3.4105
R12187 VPWR.n2431 VPWR.n2430 3.4105
R12188 VPWR.n2395 VPWR.n375 3.4105
R12189 VPWR.n2356 VPWR.n2355 3.4105
R12190 VPWR.n2292 VPWR.n462 3.4105
R12191 VPWR.n2235 VPWR.n2234 3.4105
R12192 VPWR.n2199 VPWR.n567 3.4105
R12193 VPWR.n2160 VPWR.n2159 3.4105
R12194 VPWR.n2096 VPWR.n654 3.4105
R12195 VPWR.n2039 VPWR.n2038 3.4105
R12196 VPWR.n2003 VPWR.n759 3.4105
R12197 VPWR.n1964 VPWR.n1963 3.4105
R12198 VPWR.n1900 VPWR.n846 3.4105
R12199 VPWR.n1843 VPWR.n1842 3.4105
R12200 VPWR.n1807 VPWR.n951 3.4105
R12201 VPWR.n1532 VPWR.n1143 3.4105
R12202 VPWR.n1540 VPWR.n1539 3.4105
R12203 VPWR.n1525 VPWR.n1524 3.4105
R12204 VPWR.n1517 VPWR.n1516 3.4105
R12205 VPWR.n1511 VPWR.n1510 3.4105
R12206 VPWR.n1503 VPWR.n1502 3.4105
R12207 VPWR.n1497 VPWR.n1496 3.4105
R12208 VPWR.n1489 VPWR.n1132 3.4105
R12209 VPWR.n1585 VPWR.n1584 3.4105
R12210 VPWR.n1452 VPWR.n1128 3.4105
R12211 VPWR.n1765 VPWR.n1764 3.4105
R12212 VPWR.n1808 VPWR.n954 3.4105
R12213 VPWR.n1835 VPWR.n1834 3.4105
R12214 VPWR.n1899 VPWR.n843 3.4105
R12215 VPWR.n1972 VPWR.n1971 3.4105
R12216 VPWR.n2004 VPWR.n762 3.4105
R12217 VPWR.n2031 VPWR.n2030 3.4105
R12218 VPWR.n2095 VPWR.n651 3.4105
R12219 VPWR.n2168 VPWR.n2167 3.4105
R12220 VPWR.n2200 VPWR.n570 3.4105
R12221 VPWR.n2227 VPWR.n2226 3.4105
R12222 VPWR.n2291 VPWR.n459 3.4105
R12223 VPWR.n2364 VPWR.n2363 3.4105
R12224 VPWR.n2396 VPWR.n378 3.4105
R12225 VPWR.n2423 VPWR.n2422 3.4105
R12226 VPWR.n2487 VPWR.n66 3.4105
R12227 VPWR.n2485 VPWR.n60 3.4105
R12228 VPWR.n2413 VPWR.n2412 3.4105
R12229 VPWR.n2398 VPWR.n382 3.4105
R12230 VPWR.n2374 VPWR.n2373 3.4105
R12231 VPWR.n2289 VPWR.n455 3.4105
R12232 VPWR.n2217 VPWR.n2216 3.4105
R12233 VPWR.n2202 VPWR.n574 3.4105
R12234 VPWR.n2178 VPWR.n2177 3.4105
R12235 VPWR.n2093 VPWR.n647 3.4105
R12236 VPWR.n2021 VPWR.n2020 3.4105
R12237 VPWR.n2006 VPWR.n766 3.4105
R12238 VPWR.n1982 VPWR.n1981 3.4105
R12239 VPWR.n1897 VPWR.n839 3.4105
R12240 VPWR.n1825 VPWR.n1824 3.4105
R12241 VPWR.n1810 VPWR.n958 3.4105
R12242 VPWR.n1752 VPWR.n1744 3.4105
R12243 VPWR.n1757 VPWR.n1043 3.4105
R12244 VPWR.n1809 VPWR.n955 3.4105
R12245 VPWR.n1833 VPWR.n1832 3.4105
R12246 VPWR.n1898 VPWR.n842 3.4105
R12247 VPWR.n1974 VPWR.n1973 3.4105
R12248 VPWR.n2005 VPWR.n763 3.4105
R12249 VPWR.n2029 VPWR.n2028 3.4105
R12250 VPWR.n2094 VPWR.n650 3.4105
R12251 VPWR.n2170 VPWR.n2169 3.4105
R12252 VPWR.n2201 VPWR.n571 3.4105
R12253 VPWR.n2225 VPWR.n2224 3.4105
R12254 VPWR.n2290 VPWR.n458 3.4105
R12255 VPWR.n2366 VPWR.n2365 3.4105
R12256 VPWR.n2397 VPWR.n379 3.4105
R12257 VPWR.n2421 VPWR.n2420 3.4105
R12258 VPWR.n2486 VPWR.n65 3.4105
R12259 VPWR.n2484 VPWR.n59 3.4105
R12260 VPWR.n2411 VPWR.n2410 3.4105
R12261 VPWR.n2399 VPWR.n383 3.4105
R12262 VPWR.n2376 VPWR.n2375 3.4105
R12263 VPWR.n2288 VPWR.n454 3.4105
R12264 VPWR.n2215 VPWR.n2214 3.4105
R12265 VPWR.n2203 VPWR.n575 3.4105
R12266 VPWR.n2180 VPWR.n2179 3.4105
R12267 VPWR.n2092 VPWR.n646 3.4105
R12268 VPWR.n2019 VPWR.n2018 3.4105
R12269 VPWR.n2007 VPWR.n767 3.4105
R12270 VPWR.n1984 VPWR.n1983 3.4105
R12271 VPWR.n1896 VPWR.n838 3.4105
R12272 VPWR.n1823 VPWR.n1822 3.4105
R12273 VPWR.n1811 VPWR.n959 3.4105
R12274 VPWR.n1788 VPWR.n1787 3.4105
R12275 VPWR.n1465 VPWR.n1464 3.4105
R12276 VPWR.n1797 VPWR.n931 3.4105
R12277 VPWR.n1893 VPWR.n1892 3.4105
R12278 VPWR.n1910 VPWR.n929 3.4105
R12279 VPWR.n1914 VPWR.n1913 3.4105
R12280 VPWR.n1993 VPWR.n739 3.4105
R12281 VPWR.n2089 VPWR.n2088 3.4105
R12282 VPWR.n2106 VPWR.n737 3.4105
R12283 VPWR.n2110 VPWR.n2109 3.4105
R12284 VPWR.n2189 VPWR.n547 3.4105
R12285 VPWR.n2285 VPWR.n2284 3.4105
R12286 VPWR.n2302 VPWR.n545 3.4105
R12287 VPWR.n2306 VPWR.n2305 3.4105
R12288 VPWR.n2385 VPWR.n355 3.4105
R12289 VPWR.n2481 VPWR.n2480 3.4105
R12290 VPWR.n2498 VPWR.n353 3.4105
R12291 VPWR.n2502 VPWR.n2501 3.4105
R12292 VPWR.n2512 VPWR.n2511 3.4105
R12293 VPWR.n2514 VPWR.n2513 3.4105
R12294 VPWR.n2524 VPWR.n2523 3.4105
R12295 VPWR.n2526 VPWR.n2525 3.4105
R12296 VPWR.n2536 VPWR.n2535 3.4105
R12297 VPWR.n2538 VPWR.n2537 3.4105
R12298 VPWR.n2548 VPWR.n2547 3.4105
R12299 VPWR.n2550 VPWR.n2549 3.4105
R12300 VPWR.n2560 VPWR.n2559 3.4105
R12301 VPWR.n2562 VPWR.n2561 3.4105
R12302 VPWR.n2572 VPWR.n2571 3.4105
R12303 VPWR.n2574 VPWR.n2573 3.4105
R12304 VPWR.n2584 VPWR.n2583 3.4105
R12305 VPWR.n2586 VPWR.n2585 3.4105
R12306 VPWR.n2595 VPWR.n2594 3.4105
R12307 VPWR.n2483 VPWR.n22 3.4105
R12308 VPWR.n2404 VPWR.n2403 3.4105
R12309 VPWR.n2400 VPWR.n449 3.4105
R12310 VPWR.n2383 VPWR.n2382 3.4105
R12311 VPWR.n2287 VPWR.n451 3.4105
R12312 VPWR.n2208 VPWR.n2207 3.4105
R12313 VPWR.n2204 VPWR.n641 3.4105
R12314 VPWR.n2187 VPWR.n2186 3.4105
R12315 VPWR.n2091 VPWR.n643 3.4105
R12316 VPWR.n2012 VPWR.n2011 3.4105
R12317 VPWR.n2008 VPWR.n833 3.4105
R12318 VPWR.n1991 VPWR.n1990 3.4105
R12319 VPWR.n1895 VPWR.n835 3.4105
R12320 VPWR.n1816 VPWR.n1815 3.4105
R12321 VPWR.n1812 VPWR.n1025 3.4105
R12322 VPWR.n1795 VPWR.n1794 3.4105
R12323 VPWR.n1055 VPWR.n1028 3.4105
R12324 VPWR.n1056 VPWR.n1037 3.4105
R12325 VPWR.n1754 VPWR.n1753 3.4105
R12326 VPWR.n1756 VPWR.n1755 3.4105
R12327 VPWR.n1529 VPWR.n1045 3.4105
R12328 VPWR.n1531 VPWR.n1530 3.4105
R12329 VPWR.n1528 VPWR.n1145 3.4105
R12330 VPWR.n1527 VPWR.n1526 3.4105
R12331 VPWR.n1515 VPWR.n1514 3.4105
R12332 VPWR.n1513 VPWR.n1512 3.4105
R12333 VPWR.n1501 VPWR.n1500 3.4105
R12334 VPWR.n1499 VPWR.n1498 3.4105
R12335 VPWR.n1488 VPWR.n1487 3.4105
R12336 VPWR.n1587 VPWR.n1586 3.4105
R12337 VPWR.n1589 VPWR.n1588 3.4105
R12338 VPWR.n1448 VPWR.n1232 3.4105
R12339 VPWR.n1345 VPWR.n1341 3.38874
R12340 VPWR.n1384 VPWR.n1380 3.38874
R12341 VPWR.n1421 VPWR.n1417 3.38874
R12342 VPWR.n28 VPWR.n26 3.36211
R12343 VPWR.n30 VPWR.n28 3.36211
R12344 VPWR.n32 VPWR.n30 3.36211
R12345 VPWR.n34 VPWR.n32 3.36211
R12346 VPWR.n36 VPWR.n34 3.36211
R12347 VPWR.n38 VPWR.n36 3.36211
R12348 VPWR.n40 VPWR.n38 3.36211
R12349 VPWR.n42 VPWR.n40 3.36211
R12350 VPWR.n44 VPWR.n42 3.36211
R12351 VPWR.n46 VPWR.n44 3.36211
R12352 VPWR.n48 VPWR.n46 3.36211
R12353 VPWR.n50 VPWR.n48 3.36211
R12354 VPWR.n52 VPWR.n50 3.36211
R12355 VPWR.n54 VPWR.n52 3.36211
R12356 VPWR.t1250 VPWR.t998 3.35739
R12357 VPWR.t994 VPWR.t228 3.35739
R12358 VPWR.n2571 VPWR.n66 3.28012
R12359 VPWR.n2511 VPWR.n96 3.28012
R12360 VPWR.n2550 VPWR.n77 3.28012
R12361 VPWR.n2440 VPWR.n77 3.28012
R12362 VPWR.n2547 VPWR.n78 3.28012
R12363 VPWR.n2443 VPWR.n78 3.28012
R12364 VPWR.n2535 VPWR.n84 3.28012
R12365 VPWR.n2453 VPWR.n84 3.28012
R12366 VPWR.n2453 VPWR.n366 3.28012
R12367 VPWR.n2526 VPWR.n89 3.28012
R12368 VPWR.n2460 VPWR.n89 3.28012
R12369 VPWR.n2460 VPWR.n363 3.28012
R12370 VPWR.n1498 VPWR.n1497 3.28012
R12371 VPWR.n1497 VPWR.n939 3.28012
R12372 VPWR.n1872 VPWR.n939 3.28012
R12373 VPWR.n1872 VPWR.n858 3.28012
R12374 VPWR.n1934 VPWR.n858 3.28012
R12375 VPWR.n1934 VPWR.n747 3.28012
R12376 VPWR.n2068 VPWR.n747 3.28012
R12377 VPWR.n2068 VPWR.n666 3.28012
R12378 VPWR.n2130 VPWR.n666 3.28012
R12379 VPWR.n2130 VPWR.n555 3.28012
R12380 VPWR.n2264 VPWR.n555 3.28012
R12381 VPWR.n2264 VPWR.n474 3.28012
R12382 VPWR.n2326 VPWR.n474 3.28012
R12383 VPWR.n2326 VPWR.n363 3.28012
R12384 VPWR.n2523 VPWR.n90 3.28012
R12385 VPWR.n2463 VPWR.n90 3.28012
R12386 VPWR.n2463 VPWR.n362 3.28012
R12387 VPWR.n2323 VPWR.n362 3.28012
R12388 VPWR.n2323 VPWR.n475 3.28012
R12389 VPWR.n2267 VPWR.n475 3.28012
R12390 VPWR.n2267 VPWR.n554 3.28012
R12391 VPWR.n2127 VPWR.n554 3.28012
R12392 VPWR.n2127 VPWR.n667 3.28012
R12393 VPWR.n2071 VPWR.n667 3.28012
R12394 VPWR.n2071 VPWR.n746 3.28012
R12395 VPWR.n1931 VPWR.n746 3.28012
R12396 VPWR.n1931 VPWR.n859 3.28012
R12397 VPWR.n1875 VPWR.n859 3.28012
R12398 VPWR.n1489 VPWR.n1488 3.28012
R12399 VPWR.n1489 VPWR.n938 3.28012
R12400 VPWR.n1875 VPWR.n938 3.28012
R12401 VPWR.n1503 VPWR.n1501 3.28012
R12402 VPWR.n1503 VPWR.n942 3.28012
R12403 VPWR.n1865 VPWR.n942 3.28012
R12404 VPWR.n1865 VPWR.n855 3.28012
R12405 VPWR.n1941 VPWR.n855 3.28012
R12406 VPWR.n1941 VPWR.n750 3.28012
R12407 VPWR.n2061 VPWR.n750 3.28012
R12408 VPWR.n2061 VPWR.n663 3.28012
R12409 VPWR.n2137 VPWR.n663 3.28012
R12410 VPWR.n2137 VPWR.n558 3.28012
R12411 VPWR.n2257 VPWR.n558 3.28012
R12412 VPWR.n2257 VPWR.n471 3.28012
R12413 VPWR.n2333 VPWR.n471 3.28012
R12414 VPWR.n2333 VPWR.n366 3.28012
R12415 VPWR.n2538 VPWR.n83 3.28012
R12416 VPWR.n2450 VPWR.n83 3.28012
R12417 VPWR.n2450 VPWR.n367 3.28012
R12418 VPWR.n2336 VPWR.n367 3.28012
R12419 VPWR.n2336 VPWR.n470 3.28012
R12420 VPWR.n2254 VPWR.n470 3.28012
R12421 VPWR.n2254 VPWR.n559 3.28012
R12422 VPWR.n2140 VPWR.n559 3.28012
R12423 VPWR.n2140 VPWR.n662 3.28012
R12424 VPWR.n2058 VPWR.n662 3.28012
R12425 VPWR.n2058 VPWR.n751 3.28012
R12426 VPWR.n1944 VPWR.n751 3.28012
R12427 VPWR.n1944 VPWR.n854 3.28012
R12428 VPWR.n1862 VPWR.n854 3.28012
R12429 VPWR.n1512 VPWR.n1511 3.28012
R12430 VPWR.n1511 VPWR.n943 3.28012
R12431 VPWR.n1862 VPWR.n943 3.28012
R12432 VPWR.n1517 VPWR.n1515 3.28012
R12433 VPWR.n1517 VPWR.n946 3.28012
R12434 VPWR.n1855 VPWR.n946 3.28012
R12435 VPWR.n1855 VPWR.n851 3.28012
R12436 VPWR.n1951 VPWR.n851 3.28012
R12437 VPWR.n1951 VPWR.n754 3.28012
R12438 VPWR.n2051 VPWR.n754 3.28012
R12439 VPWR.n2051 VPWR.n659 3.28012
R12440 VPWR.n2147 VPWR.n659 3.28012
R12441 VPWR.n2147 VPWR.n562 3.28012
R12442 VPWR.n2247 VPWR.n562 3.28012
R12443 VPWR.n2247 VPWR.n467 3.28012
R12444 VPWR.n2343 VPWR.n467 3.28012
R12445 VPWR.n2343 VPWR.n370 3.28012
R12446 VPWR.n2443 VPWR.n370 3.28012
R12447 VPWR.n2514 VPWR.n95 3.28012
R12448 VPWR.n2470 VPWR.n95 3.28012
R12449 VPWR.n2470 VPWR.n359 3.28012
R12450 VPWR.n2316 VPWR.n359 3.28012
R12451 VPWR.n2316 VPWR.n478 3.28012
R12452 VPWR.n2274 VPWR.n478 3.28012
R12453 VPWR.n2274 VPWR.n551 3.28012
R12454 VPWR.n2120 VPWR.n551 3.28012
R12455 VPWR.n2120 VPWR.n670 3.28012
R12456 VPWR.n2078 VPWR.n670 3.28012
R12457 VPWR.n2078 VPWR.n743 3.28012
R12458 VPWR.n1924 VPWR.n743 3.28012
R12459 VPWR.n1924 VPWR.n862 3.28012
R12460 VPWR.n1882 VPWR.n862 3.28012
R12461 VPWR.n1882 VPWR.n935 3.28012
R12462 VPWR.n1586 VPWR.n1585 3.28012
R12463 VPWR.n1585 VPWR.n935 3.28012
R12464 VPWR.n1526 VPWR.n1525 3.28012
R12465 VPWR.n1525 VPWR.n947 3.28012
R12466 VPWR.n1852 VPWR.n947 3.28012
R12467 VPWR.n1852 VPWR.n850 3.28012
R12468 VPWR.n1954 VPWR.n850 3.28012
R12469 VPWR.n1954 VPWR.n755 3.28012
R12470 VPWR.n2048 VPWR.n755 3.28012
R12471 VPWR.n2048 VPWR.n658 3.28012
R12472 VPWR.n2150 VPWR.n658 3.28012
R12473 VPWR.n2150 VPWR.n563 3.28012
R12474 VPWR.n2244 VPWR.n563 3.28012
R12475 VPWR.n2244 VPWR.n466 3.28012
R12476 VPWR.n2346 VPWR.n466 3.28012
R12477 VPWR.n2346 VPWR.n371 3.28012
R12478 VPWR.n2440 VPWR.n371 3.28012
R12479 VPWR.n2559 VPWR.n72 3.28012
R12480 VPWR.n2433 VPWR.n72 3.28012
R12481 VPWR.n2433 VPWR.n374 3.28012
R12482 VPWR.n2353 VPWR.n374 3.28012
R12483 VPWR.n2353 VPWR.n463 3.28012
R12484 VPWR.n2237 VPWR.n463 3.28012
R12485 VPWR.n2237 VPWR.n566 3.28012
R12486 VPWR.n2157 VPWR.n566 3.28012
R12487 VPWR.n2157 VPWR.n655 3.28012
R12488 VPWR.n2041 VPWR.n655 3.28012
R12489 VPWR.n2041 VPWR.n758 3.28012
R12490 VPWR.n1961 VPWR.n758 3.28012
R12491 VPWR.n1961 VPWR.n847 3.28012
R12492 VPWR.n1845 VPWR.n847 3.28012
R12493 VPWR.n1845 VPWR.n950 3.28012
R12494 VPWR.n1539 VPWR.n1145 3.28012
R12495 VPWR.n1539 VPWR.n950 3.28012
R12496 VPWR.n1589 VPWR.n1128 3.28012
R12497 VPWR.n1128 VPWR.n934 3.28012
R12498 VPWR.n1885 VPWR.n934 3.28012
R12499 VPWR.n1885 VPWR.n863 3.28012
R12500 VPWR.n1921 VPWR.n863 3.28012
R12501 VPWR.n1921 VPWR.n742 3.28012
R12502 VPWR.n2081 VPWR.n742 3.28012
R12503 VPWR.n2081 VPWR.n671 3.28012
R12504 VPWR.n2117 VPWR.n671 3.28012
R12505 VPWR.n2117 VPWR.n550 3.28012
R12506 VPWR.n2277 VPWR.n550 3.28012
R12507 VPWR.n2277 VPWR.n479 3.28012
R12508 VPWR.n2313 VPWR.n479 3.28012
R12509 VPWR.n2313 VPWR.n358 3.28012
R12510 VPWR.n2473 VPWR.n358 3.28012
R12511 VPWR.n2473 VPWR.n96 3.28012
R12512 VPWR.n2562 VPWR.n71 3.28012
R12513 VPWR.n2430 VPWR.n71 3.28012
R12514 VPWR.n2430 VPWR.n375 3.28012
R12515 VPWR.n2356 VPWR.n375 3.28012
R12516 VPWR.n2356 VPWR.n462 3.28012
R12517 VPWR.n2234 VPWR.n462 3.28012
R12518 VPWR.n2234 VPWR.n567 3.28012
R12519 VPWR.n2160 VPWR.n567 3.28012
R12520 VPWR.n2160 VPWR.n654 3.28012
R12521 VPWR.n2038 VPWR.n654 3.28012
R12522 VPWR.n2038 VPWR.n759 3.28012
R12523 VPWR.n1964 VPWR.n759 3.28012
R12524 VPWR.n1964 VPWR.n846 3.28012
R12525 VPWR.n1842 VPWR.n846 3.28012
R12526 VPWR.n1842 VPWR.n951 3.28012
R12527 VPWR.n1532 VPWR.n951 3.28012
R12528 VPWR.n1532 VPWR.n1531 3.28012
R12529 VPWR.n1764 VPWR.n1045 3.28012
R12530 VPWR.n1764 VPWR.n954 3.28012
R12531 VPWR.n1835 VPWR.n954 3.28012
R12532 VPWR.n1835 VPWR.n843 3.28012
R12533 VPWR.n1971 VPWR.n843 3.28012
R12534 VPWR.n1971 VPWR.n762 3.28012
R12535 VPWR.n2031 VPWR.n762 3.28012
R12536 VPWR.n2031 VPWR.n651 3.28012
R12537 VPWR.n2167 VPWR.n651 3.28012
R12538 VPWR.n2167 VPWR.n570 3.28012
R12539 VPWR.n2227 VPWR.n570 3.28012
R12540 VPWR.n2227 VPWR.n459 3.28012
R12541 VPWR.n2363 VPWR.n459 3.28012
R12542 VPWR.n2363 VPWR.n378 3.28012
R12543 VPWR.n2423 VPWR.n378 3.28012
R12544 VPWR.n2423 VPWR.n66 3.28012
R12545 VPWR.n2583 VPWR.n60 3.28012
R12546 VPWR.n2413 VPWR.n60 3.28012
R12547 VPWR.n2413 VPWR.n382 3.28012
R12548 VPWR.n2373 VPWR.n382 3.28012
R12549 VPWR.n2373 VPWR.n455 3.28012
R12550 VPWR.n2217 VPWR.n455 3.28012
R12551 VPWR.n2217 VPWR.n574 3.28012
R12552 VPWR.n2177 VPWR.n574 3.28012
R12553 VPWR.n2177 VPWR.n647 3.28012
R12554 VPWR.n2021 VPWR.n647 3.28012
R12555 VPWR.n2021 VPWR.n766 3.28012
R12556 VPWR.n1981 VPWR.n766 3.28012
R12557 VPWR.n1981 VPWR.n839 3.28012
R12558 VPWR.n1825 VPWR.n839 3.28012
R12559 VPWR.n1825 VPWR.n958 3.28012
R12560 VPWR.n1752 VPWR.n958 3.28012
R12561 VPWR.n1753 VPWR.n1752 3.28012
R12562 VPWR.n1757 VPWR.n1756 3.28012
R12563 VPWR.n1757 VPWR.n955 3.28012
R12564 VPWR.n1832 VPWR.n955 3.28012
R12565 VPWR.n1832 VPWR.n842 3.28012
R12566 VPWR.n1974 VPWR.n842 3.28012
R12567 VPWR.n1974 VPWR.n763 3.28012
R12568 VPWR.n2028 VPWR.n763 3.28012
R12569 VPWR.n2028 VPWR.n650 3.28012
R12570 VPWR.n2170 VPWR.n650 3.28012
R12571 VPWR.n2170 VPWR.n571 3.28012
R12572 VPWR.n2224 VPWR.n571 3.28012
R12573 VPWR.n2224 VPWR.n458 3.28012
R12574 VPWR.n2366 VPWR.n458 3.28012
R12575 VPWR.n2366 VPWR.n379 3.28012
R12576 VPWR.n2420 VPWR.n379 3.28012
R12577 VPWR.n2420 VPWR.n65 3.28012
R12578 VPWR.n2574 VPWR.n65 3.28012
R12579 VPWR.n2586 VPWR.n59 3.28012
R12580 VPWR.n2410 VPWR.n59 3.28012
R12581 VPWR.n2410 VPWR.n383 3.28012
R12582 VPWR.n2376 VPWR.n383 3.28012
R12583 VPWR.n2376 VPWR.n454 3.28012
R12584 VPWR.n2214 VPWR.n454 3.28012
R12585 VPWR.n2214 VPWR.n575 3.28012
R12586 VPWR.n2180 VPWR.n575 3.28012
R12587 VPWR.n2180 VPWR.n646 3.28012
R12588 VPWR.n2018 VPWR.n646 3.28012
R12589 VPWR.n2018 VPWR.n767 3.28012
R12590 VPWR.n1984 VPWR.n767 3.28012
R12591 VPWR.n1984 VPWR.n838 3.28012
R12592 VPWR.n1822 VPWR.n838 3.28012
R12593 VPWR.n1822 VPWR.n959 3.28012
R12594 VPWR.n1788 VPWR.n959 3.28012
R12595 VPWR.n1788 VPWR.n1037 3.28012
R12596 VPWR.n1465 VPWR.n1232 3.28012
R12597 VPWR.n1465 VPWR.n931 3.28012
R12598 VPWR.n1892 VPWR.n931 3.28012
R12599 VPWR.n1892 VPWR.n929 3.28012
R12600 VPWR.n1914 VPWR.n929 3.28012
R12601 VPWR.n1914 VPWR.n739 3.28012
R12602 VPWR.n2088 VPWR.n739 3.28012
R12603 VPWR.n2088 VPWR.n737 3.28012
R12604 VPWR.n2110 VPWR.n737 3.28012
R12605 VPWR.n2110 VPWR.n547 3.28012
R12606 VPWR.n2284 VPWR.n547 3.28012
R12607 VPWR.n2284 VPWR.n545 3.28012
R12608 VPWR.n2306 VPWR.n545 3.28012
R12609 VPWR.n2306 VPWR.n355 3.28012
R12610 VPWR.n2480 VPWR.n355 3.28012
R12611 VPWR.n2480 VPWR.n353 3.28012
R12612 VPWR.n2502 VPWR.n353 3.28012
R12613 VPWR.n2404 VPWR.n22 3.28012
R12614 VPWR.n2404 VPWR.n449 3.28012
R12615 VPWR.n2382 VPWR.n449 3.28012
R12616 VPWR.n2382 VPWR.n451 3.28012
R12617 VPWR.n2208 VPWR.n451 3.28012
R12618 VPWR.n2208 VPWR.n641 3.28012
R12619 VPWR.n2186 VPWR.n641 3.28012
R12620 VPWR.n2186 VPWR.n643 3.28012
R12621 VPWR.n2012 VPWR.n643 3.28012
R12622 VPWR.n2012 VPWR.n833 3.28012
R12623 VPWR.n1990 VPWR.n833 3.28012
R12624 VPWR.n1990 VPWR.n835 3.28012
R12625 VPWR.n1816 VPWR.n835 3.28012
R12626 VPWR.n1816 VPWR.n1025 3.28012
R12627 VPWR.n1794 VPWR.n1025 3.28012
R12628 VPWR.n1794 VPWR.n1028 3.28012
R12629 VPWR.n2594 VPWR.n22 3.26393
R12630 VPWR.n2832 VPWR.n2831 3.1005
R12631 VPWR.n2826 VPWR.n2825 3.1005
R12632 VPWR.n2846 VPWR.n2815 3.1005
R12633 VPWR.n1324 VPWR.n1322 3.01226
R12634 VPWR.n2863 VPWR 2.83761
R12635 VPWR.n1328 VPWR.n1304 2.63579
R12636 VPWR.n2731 VPWR.n2730 2.25932
R12637 VPWR.n1447 VPWR.n1446 2.01514
R12638 VPWR.n1447 VPWR.n1026 1.65255
R12639 VPWR.n2384 VPWR.n2383 1.32852
R12640 VPWR.n2287 VPWR.n450 1.32852
R12641 VPWR.n2207 VPWR.n2206 1.32852
R12642 VPWR.n2205 VPWR.n2204 1.32852
R12643 VPWR.n2188 VPWR.n2187 1.32852
R12644 VPWR.n2091 VPWR.n642 1.32852
R12645 VPWR.n2011 VPWR.n2010 1.32852
R12646 VPWR.n2009 VPWR.n2008 1.32852
R12647 VPWR.n1992 VPWR.n1991 1.32852
R12648 VPWR.n1895 VPWR.n834 1.32852
R12649 VPWR.n2401 VPWR.n2400 1.32852
R12650 VPWR.n1815 VPWR.n1814 1.32852
R12651 VPWR.n2403 VPWR.n2402 1.32852
R12652 VPWR.n1813 VPWR.n1812 1.32852
R12653 VPWR.n2483 VPWR.n21 1.32852
R12654 VPWR.n1796 VPWR.n1795 1.32852
R12655 VPWR.n2596 VPWR.n2595 1.32852
R12656 VPWR.n1055 VPWR.n1026 1.32852
R12657 VPWR.n2482 VPWR 1.25994
R12658 VPWR VPWR.n354 1.25994
R12659 VPWR VPWR.n2304 1.25994
R12660 VPWR.n2303 VPWR 1.25994
R12661 VPWR.n2286 VPWR 1.25994
R12662 VPWR VPWR.n546 1.25994
R12663 VPWR VPWR.n2108 1.25994
R12664 VPWR.n2107 VPWR 1.25994
R12665 VPWR.n2090 VPWR 1.25994
R12666 VPWR VPWR.n738 1.25994
R12667 VPWR VPWR.n1912 1.25994
R12668 VPWR.n1911 VPWR 1.25994
R12669 VPWR.n1894 VPWR 1.25994
R12670 VPWR VPWR.n930 1.25994
R12671 VPWR.n2499 VPWR 1.25994
R12672 VPWR VPWR.n1450 1.25994
R12673 VPWR VPWR.n2500 1.25994
R12674 VPWR.n1449 VPWR 1.25994
R12675 VPWR.n2597 VPWR.n2596 1.144
R12676 VPWR.n2861 VPWR.n2860 0.936724
R12677 VPWR.n2592 VPWR 0.925943
R12678 VPWR VPWR.n1063 0.925943
R12679 VPWR.n2860 VPWR.n2816 0.925245
R12680 VPWR.n2569 VPWR.n67 0.904391
R12681 VPWR.n2509 VPWR.n97 0.904391
R12682 VPWR.n2552 VPWR.n76 0.904391
R12683 VPWR.n2545 VPWR.n79 0.904391
R12684 VPWR.n2533 VPWR.n85 0.904391
R12685 VPWR.n2528 VPWR.n88 0.904391
R12686 VPWR.n1222 VPWR.n1178 0.904391
R12687 VPWR.n2521 VPWR.n91 0.904391
R12688 VPWR.n1624 VPWR.n1102 0.904391
R12689 VPWR.n1640 VPWR.n1094 0.904391
R12690 VPWR.n2540 VPWR.n82 0.904391
R12691 VPWR.n1651 VPWR.n1092 0.904391
R12692 VPWR.n1211 VPWR.n1210 0.904391
R12693 VPWR.n2516 VPWR.n94 0.904391
R12694 VPWR.n1613 VPWR.n1104 0.904391
R12695 VPWR.n1667 VPWR.n1084 0.904391
R12696 VPWR.n2557 VPWR.n73 0.904391
R12697 VPWR.n1678 VPWR.n1082 0.904391
R12698 VPWR.n1591 VPWR.n1127 0.904391
R12699 VPWR.n2564 VPWR.n70 0.904391
R12700 VPWR.n1197 VPWR.n1196 0.904391
R12701 VPWR.n1694 VPWR.n1074 0.904391
R12702 VPWR.n1742 VPWR.n1057 0.904391
R12703 VPWR.n1705 VPWR.n1071 0.904391
R12704 VPWR.n2581 VPWR.n61 0.904391
R12705 VPWR.n2588 VPWR.n58 0.904391
R12706 VPWR.n1737 VPWR.n1735 0.904391
R12707 VPWR.n1597 VPWR.n1596 0.904391
R12708 VPWR.n2504 VPWR.n289 0.904391
R12709 VPWR.n2576 VPWR.n64 0.904391
R12710 VPWR VPWR.n2863 0.812229
R12711 VPWR.n140 VPWR.n64 0.675548
R12712 VPWR.n152 VPWR.n67 0.675548
R12713 VPWR.n164 VPWR.n70 0.675548
R12714 VPWR.n176 VPWR.n73 0.675548
R12715 VPWR.n188 VPWR.n76 0.675548
R12716 VPWR.n200 VPWR.n79 0.675548
R12717 VPWR.n212 VPWR.n82 0.675548
R12718 VPWR.n224 VPWR.n85 0.675548
R12719 VPWR.n236 VPWR.n88 0.675548
R12720 VPWR.n248 VPWR.n91 0.675548
R12721 VPWR.n260 VPWR.n94 0.675548
R12722 VPWR.n272 VPWR.n97 0.675548
R12723 VPWR.n289 VPWR.n288 0.675548
R12724 VPWR.n128 VPWR.n61 0.675548
R12725 VPWR.n117 VPWR.n58 0.675548
R12726 VPWR.n1735 VPWR.n1734 0.675548
R12727 VPWR.n1719 VPWR.n1057 0.675548
R12728 VPWR.n1707 VPWR.n1705 0.675548
R12729 VPWR.n1696 VPWR.n1694 0.675548
R12730 VPWR.n1196 VPWR.n1195 0.675548
R12731 VPWR.n1680 VPWR.n1678 0.675548
R12732 VPWR.n1669 VPWR.n1667 0.675548
R12733 VPWR.n1210 VPWR.n1209 0.675548
R12734 VPWR.n1653 VPWR.n1651 0.675548
R12735 VPWR.n1642 VPWR.n1640 0.675548
R12736 VPWR.n1178 VPWR.n1177 0.675548
R12737 VPWR.n1626 VPWR.n1624 0.675548
R12738 VPWR.n1615 VPWR.n1613 0.675548
R12739 VPWR.n1127 VPWR.n1126 0.675548
R12740 VPWR.n1599 VPWR.n1597 0.675548
R12741 VPWR.n2806 VPWR.n2805 0.672385
R12742 VPWR.n2790 VPWR.n2785 0.672385
R12743 VPWR.n2770 VPWR.n2765 0.672385
R12744 VPWR.n2751 VPWR.n2746 0.672385
R12745 VPWR.n7 VPWR 0.63497
R12746 VPWR.n1242 VPWR 0.63497
R12747 VPWR.n1265 VPWR 0.63497
R12748 VPWR.n1289 VPWR 0.63497
R12749 VPWR.n24 VPWR 0.499542
R12750 VPWR.n2814 VPWR.n2813 0.442692
R12751 VPWR.n1120 VPWR.n1118 0.404056
R12752 VPWR.n144 VPWR.n138 0.404056
R12753 VPWR.n156 VPWR.n150 0.404056
R12754 VPWR.n168 VPWR.n162 0.404056
R12755 VPWR.n180 VPWR.n174 0.404056
R12756 VPWR.n192 VPWR.n186 0.404056
R12757 VPWR.n204 VPWR.n198 0.404056
R12758 VPWR.n216 VPWR.n210 0.404056
R12759 VPWR.n228 VPWR.n222 0.404056
R12760 VPWR.n240 VPWR.n234 0.404056
R12761 VPWR.n252 VPWR.n246 0.404056
R12762 VPWR.n264 VPWR.n258 0.404056
R12763 VPWR.n276 VPWR.n270 0.404056
R12764 VPWR.n283 VPWR.n101 0.404056
R12765 VPWR.n110 VPWR.n105 0.404056
R12766 VPWR.n132 VPWR.n126 0.404056
R12767 VPWR.n121 VPWR.n115 0.404056
R12768 VPWR.n1729 VPWR.n1065 0.404056
R12769 VPWR.n1723 VPWR.n1717 0.404056
R12770 VPWR.n1711 VPWR.n1070 0.404056
R12771 VPWR.n1704 VPWR.n1702 0.404056
R12772 VPWR.n1693 VPWR.n1691 0.404056
R12773 VPWR.n1684 VPWR.n1081 0.404056
R12774 VPWR.n1677 VPWR.n1675 0.404056
R12775 VPWR.n1666 VPWR.n1664 0.404056
R12776 VPWR.n1657 VPWR.n1091 0.404056
R12777 VPWR.n1650 VPWR.n1648 0.404056
R12778 VPWR.n1639 VPWR.n1637 0.404056
R12779 VPWR.n1630 VPWR.n1101 0.404056
R12780 VPWR.n1623 VPWR.n1621 0.404056
R12781 VPWR.n1612 VPWR.n1610 0.404056
R12782 VPWR.n1603 VPWR.n1111 0.404056
R12783 VPWR.n2860 VPWR.n2859 0.388
R12784 VPWR.n1608 VPWR.n1607 0.349144
R12785 VPWR.n1608 VPWR.n1099 0.349144
R12786 VPWR.n1634 VPWR.n1099 0.349144
R12787 VPWR.n1635 VPWR.n1634 0.349144
R12788 VPWR.n1635 VPWR.n1089 0.349144
R12789 VPWR.n1661 VPWR.n1089 0.349144
R12790 VPWR.n1662 VPWR.n1661 0.349144
R12791 VPWR.n1662 VPWR.n1079 0.349144
R12792 VPWR.n1688 VPWR.n1079 0.349144
R12793 VPWR.n1689 VPWR.n1688 0.349144
R12794 VPWR.n1689 VPWR.n1068 0.349144
R12795 VPWR.n1715 VPWR.n1068 0.349144
R12796 VPWR.n1727 VPWR.n1715 0.349144
R12797 VPWR.n281 VPWR.n280 0.349144
R12798 VPWR.n280 VPWR.n268 0.349144
R12799 VPWR.n268 VPWR.n256 0.349144
R12800 VPWR.n256 VPWR.n244 0.349144
R12801 VPWR.n244 VPWR.n232 0.349144
R12802 VPWR.n232 VPWR.n220 0.349144
R12803 VPWR.n220 VPWR.n208 0.349144
R12804 VPWR.n208 VPWR.n196 0.349144
R12805 VPWR.n196 VPWR.n184 0.349144
R12806 VPWR.n184 VPWR.n172 0.349144
R12807 VPWR.n172 VPWR.n160 0.349144
R12808 VPWR.n160 VPWR.n148 0.349144
R12809 VPWR.n148 VPWR.n136 0.349144
R12810 VPWR.n1462 VPWR.n1456 0.346131
R12811 VPWR.n1461 VPWR.n1457 0.346131
R12812 VPWR.n1582 VPWR.n1136 0.346131
R12813 VPWR.n1581 VPWR.n1577 0.346131
R12814 VPWR.n1576 VPWR.n1572 0.346131
R12815 VPWR.n1571 VPWR.n1567 0.346131
R12816 VPWR.n1566 VPWR.n1562 0.346131
R12817 VPWR.n1561 VPWR.n1557 0.346131
R12818 VPWR.n1556 VPWR.n1552 0.346131
R12819 VPWR.n1551 VPWR.n1547 0.346131
R12820 VPWR.n1546 VPWR.n1542 0.346131
R12821 VPWR.n1767 VPWR.n1042 0.346131
R12822 VPWR.n1784 VPWR.n1780 0.346131
R12823 VPWR.n1785 VPWR.n1776 0.346131
R12824 VPWR.n1772 VPWR.n1771 0.346131
R12825 VPWR.n2862 VPWR.n2861 0.304571
R12826 VPWR.n2594 VPWR.n55 0.300179
R12827 VPWR.n1118 VPWR.n1113 0.286958
R12828 VPWR.n145 VPWR.n144 0.286958
R12829 VPWR.n157 VPWR.n156 0.286958
R12830 VPWR.n169 VPWR.n168 0.286958
R12831 VPWR.n181 VPWR.n180 0.286958
R12832 VPWR.n193 VPWR.n192 0.286958
R12833 VPWR.n205 VPWR.n204 0.286958
R12834 VPWR.n217 VPWR.n216 0.286958
R12835 VPWR.n229 VPWR.n228 0.286958
R12836 VPWR.n241 VPWR.n240 0.286958
R12837 VPWR.n253 VPWR.n252 0.286958
R12838 VPWR.n265 VPWR.n264 0.286958
R12839 VPWR.n277 VPWR.n276 0.286958
R12840 VPWR.n283 VPWR.n102 0.286958
R12841 VPWR.n111 VPWR.n110 0.286958
R12842 VPWR.n133 VPWR.n132 0.286958
R12843 VPWR.n122 VPWR.n121 0.286958
R12844 VPWR.n1729 VPWR.n1066 0.286958
R12845 VPWR.n1724 VPWR.n1723 0.286958
R12846 VPWR.n1712 VPWR.n1711 0.286958
R12847 VPWR.n1702 VPWR.n1072 0.286958
R12848 VPWR.n1691 VPWR.n1075 0.286958
R12849 VPWR.n1685 VPWR.n1684 0.286958
R12850 VPWR.n1675 VPWR.n1083 0.286958
R12851 VPWR.n1664 VPWR.n1085 0.286958
R12852 VPWR.n1658 VPWR.n1657 0.286958
R12853 VPWR.n1648 VPWR.n1093 0.286958
R12854 VPWR.n1637 VPWR.n1095 0.286958
R12855 VPWR.n1631 VPWR.n1630 0.286958
R12856 VPWR.n1621 VPWR.n1103 0.286958
R12857 VPWR.n1610 VPWR.n1105 0.286958
R12858 VPWR.n1604 VPWR.n1603 0.286958
R12859 VPWR.n55 VPWR 0.2505
R12860 VPWR VPWR.n2481 0.249238
R12861 VPWR.n2472 VPWR 0.249238
R12862 VPWR VPWR.n2471 0.249238
R12863 VPWR.n2385 VPWR 0.249238
R12864 VPWR.n2386 VPWR 0.249238
R12865 VPWR.n2387 VPWR 0.249238
R12866 VPWR.n2388 VPWR 0.249238
R12867 VPWR.n2305 VPWR 0.249238
R12868 VPWR.n2314 VPWR 0.249238
R12869 VPWR.n2315 VPWR 0.249238
R12870 VPWR.n2324 VPWR 0.249238
R12871 VPWR.n2325 VPWR 0.249238
R12872 VPWR.n2383 VPWR 0.249238
R12873 VPWR.n2375 VPWR 0.249238
R12874 VPWR.n2374 VPWR 0.249238
R12875 VPWR.n2365 VPWR 0.249238
R12876 VPWR.n2364 VPWR 0.249238
R12877 VPWR.n2355 VPWR 0.249238
R12878 VPWR.n2354 VPWR 0.249238
R12879 VPWR.n2345 VPWR 0.249238
R12880 VPWR.n2344 VPWR 0.249238
R12881 VPWR.n2335 VPWR 0.249238
R12882 VPWR.n2334 VPWR 0.249238
R12883 VPWR VPWR.n2302 0.249238
R12884 VPWR VPWR.n2301 0.249238
R12885 VPWR VPWR.n2300 0.249238
R12886 VPWR VPWR.n2299 0.249238
R12887 VPWR VPWR.n2298 0.249238
R12888 VPWR VPWR.n2287 0.249238
R12889 VPWR VPWR.n2288 0.249238
R12890 VPWR VPWR.n2289 0.249238
R12891 VPWR VPWR.n2290 0.249238
R12892 VPWR VPWR.n2291 0.249238
R12893 VPWR VPWR.n2292 0.249238
R12894 VPWR VPWR.n2293 0.249238
R12895 VPWR VPWR.n2294 0.249238
R12896 VPWR VPWR.n2295 0.249238
R12897 VPWR VPWR.n2296 0.249238
R12898 VPWR VPWR.n2297 0.249238
R12899 VPWR VPWR.n2285 0.249238
R12900 VPWR.n2276 VPWR 0.249238
R12901 VPWR VPWR.n2275 0.249238
R12902 VPWR.n2266 VPWR 0.249238
R12903 VPWR VPWR.n2265 0.249238
R12904 VPWR.n2207 VPWR 0.249238
R12905 VPWR VPWR.n2215 0.249238
R12906 VPWR.n2216 VPWR 0.249238
R12907 VPWR VPWR.n2225 0.249238
R12908 VPWR.n2226 VPWR 0.249238
R12909 VPWR VPWR.n2235 0.249238
R12910 VPWR.n2236 VPWR 0.249238
R12911 VPWR VPWR.n2245 0.249238
R12912 VPWR.n2246 VPWR 0.249238
R12913 VPWR VPWR.n2255 0.249238
R12914 VPWR.n2256 VPWR 0.249238
R12915 VPWR.n2189 VPWR 0.249238
R12916 VPWR.n2190 VPWR 0.249238
R12917 VPWR.n2191 VPWR 0.249238
R12918 VPWR.n2192 VPWR 0.249238
R12919 VPWR.n2193 VPWR 0.249238
R12920 VPWR.n2204 VPWR 0.249238
R12921 VPWR.n2203 VPWR 0.249238
R12922 VPWR.n2202 VPWR 0.249238
R12923 VPWR.n2201 VPWR 0.249238
R12924 VPWR.n2200 VPWR 0.249238
R12925 VPWR.n2199 VPWR 0.249238
R12926 VPWR.n2198 VPWR 0.249238
R12927 VPWR.n2197 VPWR 0.249238
R12928 VPWR.n2196 VPWR 0.249238
R12929 VPWR.n2195 VPWR 0.249238
R12930 VPWR.n2194 VPWR 0.249238
R12931 VPWR.n2109 VPWR 0.249238
R12932 VPWR.n2118 VPWR 0.249238
R12933 VPWR.n2119 VPWR 0.249238
R12934 VPWR.n2128 VPWR 0.249238
R12935 VPWR.n2129 VPWR 0.249238
R12936 VPWR.n2187 VPWR 0.249238
R12937 VPWR.n2179 VPWR 0.249238
R12938 VPWR.n2178 VPWR 0.249238
R12939 VPWR.n2169 VPWR 0.249238
R12940 VPWR.n2168 VPWR 0.249238
R12941 VPWR.n2159 VPWR 0.249238
R12942 VPWR.n2158 VPWR 0.249238
R12943 VPWR.n2149 VPWR 0.249238
R12944 VPWR.n2148 VPWR 0.249238
R12945 VPWR.n2139 VPWR 0.249238
R12946 VPWR.n2138 VPWR 0.249238
R12947 VPWR VPWR.n2106 0.249238
R12948 VPWR VPWR.n2105 0.249238
R12949 VPWR VPWR.n2104 0.249238
R12950 VPWR VPWR.n2103 0.249238
R12951 VPWR VPWR.n2102 0.249238
R12952 VPWR VPWR.n2091 0.249238
R12953 VPWR VPWR.n2092 0.249238
R12954 VPWR VPWR.n2093 0.249238
R12955 VPWR VPWR.n2094 0.249238
R12956 VPWR VPWR.n2095 0.249238
R12957 VPWR VPWR.n2096 0.249238
R12958 VPWR VPWR.n2097 0.249238
R12959 VPWR VPWR.n2098 0.249238
R12960 VPWR VPWR.n2099 0.249238
R12961 VPWR VPWR.n2100 0.249238
R12962 VPWR VPWR.n2101 0.249238
R12963 VPWR VPWR.n2089 0.249238
R12964 VPWR.n2080 VPWR 0.249238
R12965 VPWR VPWR.n2079 0.249238
R12966 VPWR.n2070 VPWR 0.249238
R12967 VPWR VPWR.n2069 0.249238
R12968 VPWR.n2011 VPWR 0.249238
R12969 VPWR VPWR.n2019 0.249238
R12970 VPWR.n2020 VPWR 0.249238
R12971 VPWR VPWR.n2029 0.249238
R12972 VPWR.n2030 VPWR 0.249238
R12973 VPWR VPWR.n2039 0.249238
R12974 VPWR.n2040 VPWR 0.249238
R12975 VPWR VPWR.n2049 0.249238
R12976 VPWR.n2050 VPWR 0.249238
R12977 VPWR VPWR.n2059 0.249238
R12978 VPWR.n2060 VPWR 0.249238
R12979 VPWR.n1993 VPWR 0.249238
R12980 VPWR.n1994 VPWR 0.249238
R12981 VPWR.n1995 VPWR 0.249238
R12982 VPWR.n1996 VPWR 0.249238
R12983 VPWR.n1997 VPWR 0.249238
R12984 VPWR.n2008 VPWR 0.249238
R12985 VPWR.n2007 VPWR 0.249238
R12986 VPWR.n2006 VPWR 0.249238
R12987 VPWR.n2005 VPWR 0.249238
R12988 VPWR.n2004 VPWR 0.249238
R12989 VPWR.n2003 VPWR 0.249238
R12990 VPWR.n2002 VPWR 0.249238
R12991 VPWR.n2001 VPWR 0.249238
R12992 VPWR.n2000 VPWR 0.249238
R12993 VPWR.n1999 VPWR 0.249238
R12994 VPWR.n1998 VPWR 0.249238
R12995 VPWR.n1913 VPWR 0.249238
R12996 VPWR.n1922 VPWR 0.249238
R12997 VPWR.n1923 VPWR 0.249238
R12998 VPWR.n1932 VPWR 0.249238
R12999 VPWR.n1933 VPWR 0.249238
R13000 VPWR.n1991 VPWR 0.249238
R13001 VPWR.n1983 VPWR 0.249238
R13002 VPWR.n1982 VPWR 0.249238
R13003 VPWR.n1973 VPWR 0.249238
R13004 VPWR.n1972 VPWR 0.249238
R13005 VPWR.n1963 VPWR 0.249238
R13006 VPWR.n1962 VPWR 0.249238
R13007 VPWR.n1953 VPWR 0.249238
R13008 VPWR.n1952 VPWR 0.249238
R13009 VPWR.n1943 VPWR 0.249238
R13010 VPWR.n1942 VPWR 0.249238
R13011 VPWR VPWR.n1910 0.249238
R13012 VPWR VPWR.n1909 0.249238
R13013 VPWR VPWR.n1908 0.249238
R13014 VPWR VPWR.n1907 0.249238
R13015 VPWR VPWR.n1906 0.249238
R13016 VPWR VPWR.n1895 0.249238
R13017 VPWR VPWR.n1896 0.249238
R13018 VPWR VPWR.n1897 0.249238
R13019 VPWR VPWR.n1898 0.249238
R13020 VPWR VPWR.n1899 0.249238
R13021 VPWR VPWR.n1900 0.249238
R13022 VPWR VPWR.n1901 0.249238
R13023 VPWR VPWR.n1902 0.249238
R13024 VPWR VPWR.n1903 0.249238
R13025 VPWR VPWR.n1904 0.249238
R13026 VPWR VPWR.n1905 0.249238
R13027 VPWR.n2400 VPWR 0.249238
R13028 VPWR.n2399 VPWR 0.249238
R13029 VPWR.n2398 VPWR 0.249238
R13030 VPWR.n2397 VPWR 0.249238
R13031 VPWR.n2396 VPWR 0.249238
R13032 VPWR.n2395 VPWR 0.249238
R13033 VPWR.n2394 VPWR 0.249238
R13034 VPWR.n2393 VPWR 0.249238
R13035 VPWR.n2392 VPWR 0.249238
R13036 VPWR.n2391 VPWR 0.249238
R13037 VPWR.n2390 VPWR 0.249238
R13038 VPWR.n2389 VPWR 0.249238
R13039 VPWR VPWR.n1893 0.249238
R13040 VPWR.n1884 VPWR 0.249238
R13041 VPWR VPWR.n1883 0.249238
R13042 VPWR.n1874 VPWR 0.249238
R13043 VPWR VPWR.n1873 0.249238
R13044 VPWR.n1864 VPWR 0.249238
R13045 VPWR.n1815 VPWR 0.249238
R13046 VPWR VPWR.n1823 0.249238
R13047 VPWR.n1824 VPWR 0.249238
R13048 VPWR VPWR.n1833 0.249238
R13049 VPWR.n1834 VPWR 0.249238
R13050 VPWR VPWR.n1843 0.249238
R13051 VPWR.n1844 VPWR 0.249238
R13052 VPWR VPWR.n1853 0.249238
R13053 VPWR.n1854 VPWR 0.249238
R13054 VPWR VPWR.n1863 0.249238
R13055 VPWR.n2403 VPWR 0.249238
R13056 VPWR VPWR.n2411 0.249238
R13057 VPWR.n2412 VPWR 0.249238
R13058 VPWR VPWR.n2421 0.249238
R13059 VPWR.n2422 VPWR 0.249238
R13060 VPWR VPWR.n2431 0.249238
R13061 VPWR.n2432 VPWR 0.249238
R13062 VPWR VPWR.n2441 0.249238
R13063 VPWR.n2442 VPWR 0.249238
R13064 VPWR VPWR.n2451 0.249238
R13065 VPWR.n2452 VPWR 0.249238
R13066 VPWR VPWR.n2461 0.249238
R13067 VPWR.n2462 VPWR 0.249238
R13068 VPWR.n1797 VPWR 0.249238
R13069 VPWR.n1798 VPWR 0.249238
R13070 VPWR.n1799 VPWR 0.249238
R13071 VPWR.n1800 VPWR 0.249238
R13072 VPWR.n1801 VPWR 0.249238
R13073 VPWR.n1802 VPWR 0.249238
R13074 VPWR.n1803 VPWR 0.249238
R13075 VPWR.n1804 VPWR 0.249238
R13076 VPWR.n1805 VPWR 0.249238
R13077 VPWR.n1812 VPWR 0.249238
R13078 VPWR.n1811 VPWR 0.249238
R13079 VPWR.n1810 VPWR 0.249238
R13080 VPWR.n1809 VPWR 0.249238
R13081 VPWR.n1808 VPWR 0.249238
R13082 VPWR.n1807 VPWR 0.249238
R13083 VPWR.n1806 VPWR 0.249238
R13084 VPWR VPWR.n2498 0.249238
R13085 VPWR VPWR.n2497 0.249238
R13086 VPWR VPWR.n2496 0.249238
R13087 VPWR VPWR.n2495 0.249238
R13088 VPWR VPWR.n2494 0.249238
R13089 VPWR VPWR.n2493 0.249238
R13090 VPWR VPWR.n2492 0.249238
R13091 VPWR VPWR.n2491 0.249238
R13092 VPWR VPWR.n2490 0.249238
R13093 VPWR VPWR.n2489 0.249238
R13094 VPWR VPWR.n2488 0.249238
R13095 VPWR VPWR.n2483 0.249238
R13096 VPWR VPWR.n2484 0.249238
R13097 VPWR VPWR.n2485 0.249238
R13098 VPWR VPWR.n2486 0.249238
R13099 VPWR VPWR.n2487 0.249238
R13100 VPWR.n2501 VPWR 0.249238
R13101 VPWR.n2512 VPWR 0.249238
R13102 VPWR.n2513 VPWR 0.249238
R13103 VPWR.n2524 VPWR 0.249238
R13104 VPWR.n2525 VPWR 0.249238
R13105 VPWR.n2536 VPWR 0.249238
R13106 VPWR.n2537 VPWR 0.249238
R13107 VPWR.n2548 VPWR 0.249238
R13108 VPWR.n2549 VPWR 0.249238
R13109 VPWR.n2560 VPWR 0.249238
R13110 VPWR.n2561 VPWR 0.249238
R13111 VPWR.n2572 VPWR 0.249238
R13112 VPWR.n2573 VPWR 0.249238
R13113 VPWR.n2584 VPWR 0.249238
R13114 VPWR.n2585 VPWR 0.249238
R13115 VPWR.n2595 VPWR 0.249238
R13116 VPWR VPWR.n1055 0.249238
R13117 VPWR VPWR.n1056 0.249238
R13118 VPWR VPWR.n1754 0.249238
R13119 VPWR.n1755 VPWR 0.249238
R13120 VPWR VPWR.n1529 0.249238
R13121 VPWR.n1530 VPWR 0.249238
R13122 VPWR.n1528 VPWR 0.249238
R13123 VPWR.n1527 VPWR 0.249238
R13124 VPWR.n1514 VPWR 0.249238
R13125 VPWR.n1513 VPWR 0.249238
R13126 VPWR.n1500 VPWR 0.249238
R13127 VPWR.n1499 VPWR 0.249238
R13128 VPWR.n1487 VPWR 0.249238
R13129 VPWR VPWR.n1587 0.249238
R13130 VPWR.n1588 VPWR 0.249238
R13131 VPWR VPWR.n1448 0.249238
R13132 VPWR.n2861 VPWR.n2815 0.245065
R13133 VPWR.n2813 VPWR.n2797 0.213567
R13134 VPWR.n2797 VPWR.n2778 0.213567
R13135 VPWR.n2778 VPWR.n2758 0.213567
R13136 VPWR.n2758 VPWR.n2739 0.213567
R13137 VPWR.n2739 VPWR.n2703 0.213567
R13138 VPWR.n2703 VPWR.n2665 0.213567
R13139 VPWR.n2665 VPWR.n2628 0.213567
R13140 VPWR.n1446 VPWR.n1414 0.213567
R13141 VPWR.n1414 VPWR.n1376 0.213567
R13142 VPWR.n1376 VPWR.n1337 0.213567
R13143 VPWR.n1337 VPWR.n1302 0.213567
R13144 VPWR.n1302 VPWR.n1279 0.213567
R13145 VPWR.n1279 VPWR.n1255 0.213567
R13146 VPWR.n1255 VPWR.n19 0.213567
R13147 VPWR VPWR.n2862 0.204304
R13148 VPWR.n1449 VPWR.n1447 0.182233
R13149 VPWR.n1450 VPWR.n1449 0.154425
R13150 VPWR.n1450 VPWR.n930 0.154425
R13151 VPWR.n1894 VPWR.n930 0.154425
R13152 VPWR.n1911 VPWR.n1894 0.154425
R13153 VPWR.n1912 VPWR.n1911 0.154425
R13154 VPWR.n1912 VPWR.n738 0.154425
R13155 VPWR.n2090 VPWR.n738 0.154425
R13156 VPWR.n2107 VPWR.n2090 0.154425
R13157 VPWR.n2108 VPWR.n2107 0.154425
R13158 VPWR.n2108 VPWR.n546 0.154425
R13159 VPWR.n2286 VPWR.n546 0.154425
R13160 VPWR.n2303 VPWR.n2286 0.154425
R13161 VPWR.n2304 VPWR.n2303 0.154425
R13162 VPWR.n2304 VPWR.n354 0.154425
R13163 VPWR.n2482 VPWR.n354 0.154425
R13164 VPWR.n2499 VPWR.n2482 0.154425
R13165 VPWR.n2500 VPWR.n2499 0.154425
R13166 VPWR.n1796 VPWR.n1026 0.154425
R13167 VPWR.n1813 VPWR.n1796 0.154425
R13168 VPWR.n1814 VPWR.n1813 0.154425
R13169 VPWR.n1814 VPWR.n834 0.154425
R13170 VPWR.n1992 VPWR.n834 0.154425
R13171 VPWR.n2009 VPWR.n1992 0.154425
R13172 VPWR.n2010 VPWR.n2009 0.154425
R13173 VPWR.n2010 VPWR.n642 0.154425
R13174 VPWR.n2188 VPWR.n642 0.154425
R13175 VPWR.n2205 VPWR.n2188 0.154425
R13176 VPWR.n2206 VPWR.n2205 0.154425
R13177 VPWR.n2206 VPWR.n450 0.154425
R13178 VPWR.n2384 VPWR.n450 0.154425
R13179 VPWR.n2401 VPWR.n2384 0.154425
R13180 VPWR.n2402 VPWR.n2401 0.154425
R13181 VPWR.n2402 VPWR.n21 0.154425
R13182 VPWR.n2596 VPWR.n21 0.154425
R13183 VPWR.n8 VPWR.n7 0.147771
R13184 VPWR.n1243 VPWR.n1242 0.147771
R13185 VPWR.n1266 VPWR.n1265 0.147771
R13186 VPWR.n1290 VPWR.n1289 0.147771
R13187 VPWR.n1113 VPWR 0.135917
R13188 VPWR.n145 VPWR 0.135917
R13189 VPWR.n157 VPWR 0.135917
R13190 VPWR.n169 VPWR 0.135917
R13191 VPWR.n181 VPWR 0.135917
R13192 VPWR.n193 VPWR 0.135917
R13193 VPWR.n205 VPWR 0.135917
R13194 VPWR.n217 VPWR 0.135917
R13195 VPWR.n229 VPWR 0.135917
R13196 VPWR.n241 VPWR 0.135917
R13197 VPWR.n253 VPWR 0.135917
R13198 VPWR.n265 VPWR 0.135917
R13199 VPWR.n277 VPWR 0.135917
R13200 VPWR.n102 VPWR 0.135917
R13201 VPWR.n111 VPWR 0.135917
R13202 VPWR.n133 VPWR 0.135917
R13203 VPWR.n122 VPWR 0.135917
R13204 VPWR.n1066 VPWR 0.135917
R13205 VPWR.n1724 VPWR 0.135917
R13206 VPWR.n1712 VPWR 0.135917
R13207 VPWR.n1072 VPWR 0.135917
R13208 VPWR.n1075 VPWR 0.135917
R13209 VPWR.n1685 VPWR 0.135917
R13210 VPWR.n1083 VPWR 0.135917
R13211 VPWR.n1085 VPWR 0.135917
R13212 VPWR.n1658 VPWR 0.135917
R13213 VPWR.n1093 VPWR 0.135917
R13214 VPWR.n1095 VPWR 0.135917
R13215 VPWR.n1631 VPWR 0.135917
R13216 VPWR.n1103 VPWR 0.135917
R13217 VPWR.n1105 VPWR 0.135917
R13218 VPWR.n1604 VPWR 0.135917
R13219 VPWR.n2863 VPWR.n2814 0.127988
R13220 VPWR.n2825 VPWR.n2816 0.1255
R13221 VPWR.n2831 VPWR.n2816 0.1255
R13222 VPWR.n18 VPWR.n0 0.120292
R13223 VPWR.n14 VPWR.n0 0.120292
R13224 VPWR.n9 VPWR.n8 0.120292
R13225 VPWR.n1254 VPWR.n1233 0.120292
R13226 VPWR.n1250 VPWR.n1233 0.120292
R13227 VPWR.n1244 VPWR.n1243 0.120292
R13228 VPWR.n1278 VPWR.n1256 0.120292
R13229 VPWR.n1273 VPWR.n1256 0.120292
R13230 VPWR.n1267 VPWR.n1266 0.120292
R13231 VPWR.n1301 VPWR.n1280 0.120292
R13232 VPWR.n1297 VPWR.n1280 0.120292
R13233 VPWR.n1291 VPWR.n1290 0.120292
R13234 VPWR.n1333 VPWR.n1332 0.120292
R13235 VPWR.n1326 VPWR.n1305 0.120292
R13236 VPWR.n1319 VPWR.n1305 0.120292
R13237 VPWR.n1319 VPWR.n1318 0.120292
R13238 VPWR.n1317 VPWR.n1309 0.120292
R13239 VPWR.n1312 VPWR.n1309 0.120292
R13240 VPWR.n1312 VPWR.n1311 0.120292
R13241 VPWR.n1371 VPWR.n1370 0.120292
R13242 VPWR.n1364 VPWR.n1363 0.120292
R13243 VPWR.n1363 VPWR.n1340 0.120292
R13244 VPWR.n1356 VPWR.n1340 0.120292
R13245 VPWR.n1356 VPWR.n1355 0.120292
R13246 VPWR.n1355 VPWR.n1354 0.120292
R13247 VPWR.n1354 VPWR.n1342 0.120292
R13248 VPWR.n1348 VPWR.n1342 0.120292
R13249 VPWR.n1348 VPWR.n1347 0.120292
R13250 VPWR.n1410 VPWR.n1409 0.120292
R13251 VPWR.n1403 VPWR.n1402 0.120292
R13252 VPWR.n1402 VPWR.n1379 0.120292
R13253 VPWR.n1395 VPWR.n1379 0.120292
R13254 VPWR.n1395 VPWR.n1394 0.120292
R13255 VPWR.n1394 VPWR.n1393 0.120292
R13256 VPWR.n1393 VPWR.n1381 0.120292
R13257 VPWR.n1387 VPWR.n1381 0.120292
R13258 VPWR.n1387 VPWR.n1386 0.120292
R13259 VPWR.n1440 VPWR.n1439 0.120292
R13260 VPWR.n1439 VPWR.n1416 0.120292
R13261 VPWR.n1432 VPWR.n1416 0.120292
R13262 VPWR.n1432 VPWR.n1431 0.120292
R13263 VPWR.n1431 VPWR.n1430 0.120292
R13264 VPWR.n1430 VPWR.n1418 0.120292
R13265 VPWR.n1424 VPWR.n1418 0.120292
R13266 VPWR.n1424 VPWR.n1423 0.120292
R13267 VPWR.n2812 VPWR.n2798 0.120292
R13268 VPWR.n2796 VPWR.n2779 0.120292
R13269 VPWR.n2777 VPWR.n2759 0.120292
R13270 VPWR.n2757 VPWR.n2740 0.120292
R13271 VPWR.n2719 VPWR.n2718 0.120292
R13272 VPWR.n2720 VPWR.n2719 0.120292
R13273 VPWR.n2720 VPWR.n2711 0.120292
R13274 VPWR.n2725 VPWR.n2711 0.120292
R13275 VPWR.n2726 VPWR.n2725 0.120292
R13276 VPWR.n2726 VPWR.n2707 0.120292
R13277 VPWR.n2732 VPWR.n2707 0.120292
R13278 VPWR.n2734 VPWR.n2704 0.120292
R13279 VPWR.n2738 VPWR.n2704 0.120292
R13280 VPWR.n2683 VPWR.n2682 0.120292
R13281 VPWR.n2684 VPWR.n2683 0.120292
R13282 VPWR.n2684 VPWR.n2673 0.120292
R13283 VPWR.n2689 VPWR.n2673 0.120292
R13284 VPWR.n2690 VPWR.n2689 0.120292
R13285 VPWR.n2690 VPWR.n2669 0.120292
R13286 VPWR.n2695 VPWR.n2669 0.120292
R13287 VPWR.n2697 VPWR.n2666 0.120292
R13288 VPWR.n2702 VPWR.n2666 0.120292
R13289 VPWR.n2646 VPWR.n2645 0.120292
R13290 VPWR.n2647 VPWR.n2646 0.120292
R13291 VPWR.n2647 VPWR.n2636 0.120292
R13292 VPWR.n2652 VPWR.n2636 0.120292
R13293 VPWR.n2653 VPWR.n2652 0.120292
R13294 VPWR.n2653 VPWR.n2632 0.120292
R13295 VPWR.n2658 VPWR.n2632 0.120292
R13296 VPWR.n2660 VPWR.n2629 0.120292
R13297 VPWR.n2664 VPWR.n2629 0.120292
R13298 VPWR.n2608 VPWR.n2604 0.120292
R13299 VPWR.n2616 VPWR.n2604 0.120292
R13300 VPWR.n2617 VPWR.n2616 0.120292
R13301 VPWR.n2618 VPWR.n2617 0.120292
R13302 VPWR.n2618 VPWR.n2600 0.120292
R13303 VPWR.n2623 VPWR.n2600 0.120292
R13304 VPWR.n2624 VPWR.n2623 0.120292
R13305 VPWR.n1605 VPWR 0.118556
R13306 VPWR.n1108 VPWR 0.118556
R13307 VPWR.n1619 VPWR 0.118556
R13308 VPWR.n1632 VPWR 0.118556
R13309 VPWR.n1098 VPWR 0.118556
R13310 VPWR.n1646 VPWR 0.118556
R13311 VPWR.n1659 VPWR 0.118556
R13312 VPWR.n1088 VPWR 0.118556
R13313 VPWR.n1673 VPWR 0.118556
R13314 VPWR.n1686 VPWR 0.118556
R13315 VPWR.n1078 VPWR 0.118556
R13316 VPWR.n1700 VPWR 0.118556
R13317 VPWR.n1713 VPWR 0.118556
R13318 VPWR.n1725 VPWR 0.118556
R13319 VPWR VPWR.n1112 0.118556
R13320 VPWR.n1067 VPWR 0.118556
R13321 VPWR.n123 VPWR 0.118556
R13322 VPWR.n112 VPWR 0.118556
R13323 VPWR.n103 VPWR 0.118556
R13324 VPWR.n278 VPWR 0.118556
R13325 VPWR.n266 VPWR 0.118556
R13326 VPWR.n254 VPWR 0.118556
R13327 VPWR.n242 VPWR 0.118556
R13328 VPWR.n230 VPWR 0.118556
R13329 VPWR.n218 VPWR 0.118556
R13330 VPWR.n206 VPWR 0.118556
R13331 VPWR.n194 VPWR 0.118556
R13332 VPWR.n182 VPWR 0.118556
R13333 VPWR.n170 VPWR 0.118556
R13334 VPWR.n158 VPWR 0.118556
R13335 VPWR.n146 VPWR 0.118556
R13336 VPWR.n134 VPWR 0.118556
R13337 VPWR.n1765 VPWR.n1044 0.108238
R13338 VPWR.n1541 VPWR.n1143 0.108238
R13339 VPWR.n1540 VPWR.n1142 0.108238
R13340 VPWR.n1524 VPWR.n1141 0.108238
R13341 VPWR.n1516 VPWR.n1140 0.108238
R13342 VPWR.n1510 VPWR.n1139 0.108238
R13343 VPWR.n1502 VPWR.n1138 0.108238
R13344 VPWR.n1496 VPWR.n1137 0.108238
R13345 VPWR.n1583 VPWR.n1132 0.108238
R13346 VPWR.n1584 VPWR.n1131 0.108238
R13347 VPWR.n1463 VPWR.n1452 0.108238
R13348 VPWR.n1464 VPWR.n1451 0.108238
R13349 VPWR.n1795 VPWR.n1027 0.108238
R13350 VPWR.n1766 VPWR.n1043 0.108238
R13351 VPWR.n1744 VPWR.n1038 0.108238
R13352 VPWR.n1787 VPWR.n1786 0.108238
R13353 VPWR.n2481 VPWR 0.100405
R13354 VPWR.n2472 VPWR 0.100405
R13355 VPWR VPWR.n2385 0.100405
R13356 VPWR VPWR.n2386 0.100405
R13357 VPWR VPWR.n2387 0.100405
R13358 VPWR.n2305 VPWR 0.100405
R13359 VPWR VPWR.n2314 0.100405
R13360 VPWR.n2315 VPWR 0.100405
R13361 VPWR VPWR.n2324 0.100405
R13362 VPWR.n2375 VPWR 0.100405
R13363 VPWR VPWR.n2374 0.100405
R13364 VPWR.n2365 VPWR 0.100405
R13365 VPWR VPWR.n2364 0.100405
R13366 VPWR.n2355 VPWR 0.100405
R13367 VPWR VPWR.n2354 0.100405
R13368 VPWR.n2345 VPWR 0.100405
R13369 VPWR VPWR.n2344 0.100405
R13370 VPWR.n2335 VPWR 0.100405
R13371 VPWR VPWR.n2334 0.100405
R13372 VPWR.n2325 VPWR 0.100405
R13373 VPWR.n2302 VPWR 0.100405
R13374 VPWR.n2301 VPWR 0.100405
R13375 VPWR.n2300 VPWR 0.100405
R13376 VPWR.n2299 VPWR 0.100405
R13377 VPWR.n2288 VPWR 0.100405
R13378 VPWR.n2289 VPWR 0.100405
R13379 VPWR.n2290 VPWR 0.100405
R13380 VPWR.n2291 VPWR 0.100405
R13381 VPWR.n2292 VPWR 0.100405
R13382 VPWR.n2293 VPWR 0.100405
R13383 VPWR.n2294 VPWR 0.100405
R13384 VPWR.n2295 VPWR 0.100405
R13385 VPWR.n2296 VPWR 0.100405
R13386 VPWR.n2297 VPWR 0.100405
R13387 VPWR.n2298 VPWR 0.100405
R13388 VPWR.n2285 VPWR 0.100405
R13389 VPWR.n2276 VPWR 0.100405
R13390 VPWR.n2275 VPWR 0.100405
R13391 VPWR.n2266 VPWR 0.100405
R13392 VPWR.n2215 VPWR 0.100405
R13393 VPWR.n2216 VPWR 0.100405
R13394 VPWR.n2225 VPWR 0.100405
R13395 VPWR.n2226 VPWR 0.100405
R13396 VPWR.n2235 VPWR 0.100405
R13397 VPWR.n2236 VPWR 0.100405
R13398 VPWR.n2245 VPWR 0.100405
R13399 VPWR.n2246 VPWR 0.100405
R13400 VPWR.n2255 VPWR 0.100405
R13401 VPWR.n2256 VPWR 0.100405
R13402 VPWR.n2265 VPWR 0.100405
R13403 VPWR VPWR.n2189 0.100405
R13404 VPWR VPWR.n2190 0.100405
R13405 VPWR VPWR.n2191 0.100405
R13406 VPWR VPWR.n2192 0.100405
R13407 VPWR VPWR.n2203 0.100405
R13408 VPWR VPWR.n2202 0.100405
R13409 VPWR VPWR.n2201 0.100405
R13410 VPWR VPWR.n2200 0.100405
R13411 VPWR VPWR.n2199 0.100405
R13412 VPWR VPWR.n2198 0.100405
R13413 VPWR VPWR.n2197 0.100405
R13414 VPWR VPWR.n2196 0.100405
R13415 VPWR VPWR.n2195 0.100405
R13416 VPWR VPWR.n2194 0.100405
R13417 VPWR VPWR.n2193 0.100405
R13418 VPWR.n2109 VPWR 0.100405
R13419 VPWR VPWR.n2118 0.100405
R13420 VPWR.n2119 VPWR 0.100405
R13421 VPWR VPWR.n2128 0.100405
R13422 VPWR.n2179 VPWR 0.100405
R13423 VPWR VPWR.n2178 0.100405
R13424 VPWR.n2169 VPWR 0.100405
R13425 VPWR VPWR.n2168 0.100405
R13426 VPWR.n2159 VPWR 0.100405
R13427 VPWR VPWR.n2158 0.100405
R13428 VPWR.n2149 VPWR 0.100405
R13429 VPWR VPWR.n2148 0.100405
R13430 VPWR.n2139 VPWR 0.100405
R13431 VPWR VPWR.n2138 0.100405
R13432 VPWR.n2129 VPWR 0.100405
R13433 VPWR.n2106 VPWR 0.100405
R13434 VPWR.n2105 VPWR 0.100405
R13435 VPWR.n2104 VPWR 0.100405
R13436 VPWR.n2103 VPWR 0.100405
R13437 VPWR.n2092 VPWR 0.100405
R13438 VPWR.n2093 VPWR 0.100405
R13439 VPWR.n2094 VPWR 0.100405
R13440 VPWR.n2095 VPWR 0.100405
R13441 VPWR.n2096 VPWR 0.100405
R13442 VPWR.n2097 VPWR 0.100405
R13443 VPWR.n2098 VPWR 0.100405
R13444 VPWR.n2099 VPWR 0.100405
R13445 VPWR.n2100 VPWR 0.100405
R13446 VPWR.n2101 VPWR 0.100405
R13447 VPWR.n2102 VPWR 0.100405
R13448 VPWR.n2089 VPWR 0.100405
R13449 VPWR.n2080 VPWR 0.100405
R13450 VPWR.n2079 VPWR 0.100405
R13451 VPWR.n2070 VPWR 0.100405
R13452 VPWR.n2019 VPWR 0.100405
R13453 VPWR.n2020 VPWR 0.100405
R13454 VPWR.n2029 VPWR 0.100405
R13455 VPWR.n2030 VPWR 0.100405
R13456 VPWR.n2039 VPWR 0.100405
R13457 VPWR.n2040 VPWR 0.100405
R13458 VPWR.n2049 VPWR 0.100405
R13459 VPWR.n2050 VPWR 0.100405
R13460 VPWR.n2059 VPWR 0.100405
R13461 VPWR.n2060 VPWR 0.100405
R13462 VPWR.n2069 VPWR 0.100405
R13463 VPWR VPWR.n1993 0.100405
R13464 VPWR VPWR.n1994 0.100405
R13465 VPWR VPWR.n1995 0.100405
R13466 VPWR VPWR.n1996 0.100405
R13467 VPWR VPWR.n2007 0.100405
R13468 VPWR VPWR.n2006 0.100405
R13469 VPWR VPWR.n2005 0.100405
R13470 VPWR VPWR.n2004 0.100405
R13471 VPWR VPWR.n2003 0.100405
R13472 VPWR VPWR.n2002 0.100405
R13473 VPWR VPWR.n2001 0.100405
R13474 VPWR VPWR.n2000 0.100405
R13475 VPWR VPWR.n1999 0.100405
R13476 VPWR VPWR.n1998 0.100405
R13477 VPWR VPWR.n1997 0.100405
R13478 VPWR.n1913 VPWR 0.100405
R13479 VPWR VPWR.n1922 0.100405
R13480 VPWR.n1923 VPWR 0.100405
R13481 VPWR VPWR.n1932 0.100405
R13482 VPWR.n1983 VPWR 0.100405
R13483 VPWR VPWR.n1982 0.100405
R13484 VPWR.n1973 VPWR 0.100405
R13485 VPWR VPWR.n1972 0.100405
R13486 VPWR.n1963 VPWR 0.100405
R13487 VPWR VPWR.n1962 0.100405
R13488 VPWR.n1953 VPWR 0.100405
R13489 VPWR VPWR.n1952 0.100405
R13490 VPWR.n1943 VPWR 0.100405
R13491 VPWR VPWR.n1942 0.100405
R13492 VPWR.n1933 VPWR 0.100405
R13493 VPWR.n1910 VPWR 0.100405
R13494 VPWR.n1909 VPWR 0.100405
R13495 VPWR.n1908 VPWR 0.100405
R13496 VPWR.n1907 VPWR 0.100405
R13497 VPWR.n1896 VPWR 0.100405
R13498 VPWR.n1897 VPWR 0.100405
R13499 VPWR.n1898 VPWR 0.100405
R13500 VPWR.n1899 VPWR 0.100405
R13501 VPWR.n1900 VPWR 0.100405
R13502 VPWR.n1901 VPWR 0.100405
R13503 VPWR.n1902 VPWR 0.100405
R13504 VPWR.n1903 VPWR 0.100405
R13505 VPWR.n1904 VPWR 0.100405
R13506 VPWR.n1905 VPWR 0.100405
R13507 VPWR.n1906 VPWR 0.100405
R13508 VPWR VPWR.n2399 0.100405
R13509 VPWR VPWR.n2398 0.100405
R13510 VPWR VPWR.n2397 0.100405
R13511 VPWR VPWR.n2396 0.100405
R13512 VPWR VPWR.n2395 0.100405
R13513 VPWR VPWR.n2394 0.100405
R13514 VPWR VPWR.n2393 0.100405
R13515 VPWR VPWR.n2392 0.100405
R13516 VPWR VPWR.n2391 0.100405
R13517 VPWR VPWR.n2390 0.100405
R13518 VPWR VPWR.n2389 0.100405
R13519 VPWR VPWR.n2388 0.100405
R13520 VPWR.n1893 VPWR 0.100405
R13521 VPWR.n1884 VPWR 0.100405
R13522 VPWR.n1883 VPWR 0.100405
R13523 VPWR.n1874 VPWR 0.100405
R13524 VPWR.n1873 VPWR 0.100405
R13525 VPWR.n1823 VPWR 0.100405
R13526 VPWR.n1824 VPWR 0.100405
R13527 VPWR.n1833 VPWR 0.100405
R13528 VPWR.n1834 VPWR 0.100405
R13529 VPWR.n1843 VPWR 0.100405
R13530 VPWR.n1844 VPWR 0.100405
R13531 VPWR.n1853 VPWR 0.100405
R13532 VPWR.n1854 VPWR 0.100405
R13533 VPWR.n1863 VPWR 0.100405
R13534 VPWR.n1864 VPWR 0.100405
R13535 VPWR.n2411 VPWR 0.100405
R13536 VPWR.n2412 VPWR 0.100405
R13537 VPWR.n2421 VPWR 0.100405
R13538 VPWR.n2422 VPWR 0.100405
R13539 VPWR.n2431 VPWR 0.100405
R13540 VPWR.n2432 VPWR 0.100405
R13541 VPWR.n2441 VPWR 0.100405
R13542 VPWR.n2442 VPWR 0.100405
R13543 VPWR.n2451 VPWR 0.100405
R13544 VPWR.n2452 VPWR 0.100405
R13545 VPWR.n2461 VPWR 0.100405
R13546 VPWR.n2462 VPWR 0.100405
R13547 VPWR.n2471 VPWR 0.100405
R13548 VPWR VPWR.n1797 0.100405
R13549 VPWR VPWR.n1798 0.100405
R13550 VPWR VPWR.n1799 0.100405
R13551 VPWR VPWR.n1800 0.100405
R13552 VPWR VPWR.n1801 0.100405
R13553 VPWR VPWR.n1802 0.100405
R13554 VPWR VPWR.n1803 0.100405
R13555 VPWR VPWR.n1804 0.100405
R13556 VPWR VPWR.n1811 0.100405
R13557 VPWR VPWR.n1810 0.100405
R13558 VPWR VPWR.n1809 0.100405
R13559 VPWR VPWR.n1808 0.100405
R13560 VPWR VPWR.n1807 0.100405
R13561 VPWR VPWR.n1806 0.100405
R13562 VPWR VPWR.n1805 0.100405
R13563 VPWR.n2498 VPWR 0.100405
R13564 VPWR.n2497 VPWR 0.100405
R13565 VPWR.n2496 VPWR 0.100405
R13566 VPWR.n2495 VPWR 0.100405
R13567 VPWR.n2494 VPWR 0.100405
R13568 VPWR.n2493 VPWR 0.100405
R13569 VPWR.n2492 VPWR 0.100405
R13570 VPWR.n2491 VPWR 0.100405
R13571 VPWR.n2490 VPWR 0.100405
R13572 VPWR.n2489 VPWR 0.100405
R13573 VPWR.n2484 VPWR 0.100405
R13574 VPWR.n2485 VPWR 0.100405
R13575 VPWR.n2486 VPWR 0.100405
R13576 VPWR.n2487 VPWR 0.100405
R13577 VPWR.n2488 VPWR 0.100405
R13578 VPWR.n1143 VPWR 0.100405
R13579 VPWR VPWR.n1540 0.100405
R13580 VPWR.n1524 VPWR 0.100405
R13581 VPWR.n1516 VPWR 0.100405
R13582 VPWR.n1510 VPWR 0.100405
R13583 VPWR.n1502 VPWR 0.100405
R13584 VPWR.n1496 VPWR 0.100405
R13585 VPWR VPWR.n1132 0.100405
R13586 VPWR.n1584 VPWR 0.100405
R13587 VPWR.n1452 VPWR 0.100405
R13588 VPWR.n1464 VPWR 0.100405
R13589 VPWR.n1043 VPWR 0.100405
R13590 VPWR.n1744 VPWR 0.100405
R13591 VPWR.n1787 VPWR 0.100405
R13592 VPWR VPWR.n1765 0.100405
R13593 VPWR.n2501 VPWR 0.100405
R13594 VPWR VPWR.n2512 0.100405
R13595 VPWR.n2513 VPWR 0.100405
R13596 VPWR VPWR.n2524 0.100405
R13597 VPWR.n2525 VPWR 0.100405
R13598 VPWR VPWR.n2536 0.100405
R13599 VPWR.n2537 VPWR 0.100405
R13600 VPWR VPWR.n2548 0.100405
R13601 VPWR.n2549 VPWR 0.100405
R13602 VPWR VPWR.n2560 0.100405
R13603 VPWR.n2561 VPWR 0.100405
R13604 VPWR VPWR.n2572 0.100405
R13605 VPWR.n2573 VPWR 0.100405
R13606 VPWR VPWR.n2584 0.100405
R13607 VPWR.n2585 VPWR 0.100405
R13608 VPWR.n1056 VPWR 0.100405
R13609 VPWR.n1754 VPWR 0.100405
R13610 VPWR.n1755 VPWR 0.100405
R13611 VPWR.n1529 VPWR 0.100405
R13612 VPWR.n1530 VPWR 0.100405
R13613 VPWR VPWR.n1528 0.100405
R13614 VPWR VPWR.n1527 0.100405
R13615 VPWR.n1514 VPWR 0.100405
R13616 VPWR VPWR.n1513 0.100405
R13617 VPWR.n1500 VPWR 0.100405
R13618 VPWR VPWR.n1499 0.100405
R13619 VPWR.n1487 VPWR 0.100405
R13620 VPWR.n1587 VPWR 0.100405
R13621 VPWR.n1588 VPWR 0.100405
R13622 VPWR.n1448 VPWR 0.100405
R13623 VPWR VPWR.n2798 0.0994583
R13624 VPWR VPWR.n2779 0.0994583
R13625 VPWR VPWR.n1326 0.0981562
R13626 VPWR.n1371 VPWR 0.0981562
R13627 VPWR.n1410 VPWR 0.0981562
R13628 VPWR.n9 VPWR 0.0968542
R13629 VPWR.n1244 VPWR 0.0968542
R13630 VPWR.n1267 VPWR 0.0968542
R13631 VPWR.n1291 VPWR 0.0968542
R13632 VPWR.n1333 VPWR 0.0968542
R13633 VPWR VPWR.n2759 0.0968542
R13634 VPWR VPWR.n2740 0.0968542
R13635 VPWR.n2718 VPWR 0.0968542
R13636 VPWR.n2682 VPWR 0.0968542
R13637 VPWR.n2645 VPWR 0.0968542
R13638 VPWR.n2608 VPWR 0.0968542
R13639 VPWR VPWR.n1044 0.0945
R13640 VPWR.n1541 VPWR 0.0945
R13641 VPWR VPWR.n1142 0.0945
R13642 VPWR VPWR.n1141 0.0945
R13643 VPWR VPWR.n1140 0.0945
R13644 VPWR VPWR.n1139 0.0945
R13645 VPWR VPWR.n1138 0.0945
R13646 VPWR.n1137 VPWR 0.0945
R13647 VPWR VPWR.n1583 0.0945
R13648 VPWR VPWR.n1131 0.0945
R13649 VPWR VPWR.n1463 0.0945
R13650 VPWR.n1451 VPWR 0.0945
R13651 VPWR VPWR.n1038 0.0945
R13652 VPWR.n1786 VPWR 0.0945
R13653 VPWR VPWR.n1027 0.0945
R13654 VPWR.n1766 VPWR 0.0945
R13655 VPWR.n1117 VPWR 0.093504
R13656 VPWR.n109 VPWR 0.093504
R13657 VPWR.n143 VPWR 0.093504
R13658 VPWR.n155 VPWR 0.093504
R13659 VPWR.n167 VPWR 0.093504
R13660 VPWR.n179 VPWR 0.093504
R13661 VPWR.n191 VPWR 0.093504
R13662 VPWR.n203 VPWR 0.093504
R13663 VPWR.n215 VPWR 0.093504
R13664 VPWR.n227 VPWR 0.093504
R13665 VPWR.n239 VPWR 0.093504
R13666 VPWR.n251 VPWR 0.093504
R13667 VPWR.n263 VPWR 0.093504
R13668 VPWR.n275 VPWR 0.093504
R13669 VPWR VPWR.n285 0.093504
R13670 VPWR.n131 VPWR 0.093504
R13671 VPWR.n120 VPWR 0.093504
R13672 VPWR VPWR.n1731 0.093504
R13673 VPWR.n1722 VPWR 0.093504
R13674 VPWR.n1710 VPWR 0.093504
R13675 VPWR.n1699 VPWR 0.093504
R13676 VPWR VPWR.n1077 0.093504
R13677 VPWR.n1683 VPWR 0.093504
R13678 VPWR.n1672 VPWR 0.093504
R13679 VPWR VPWR.n1087 0.093504
R13680 VPWR.n1656 VPWR 0.093504
R13681 VPWR.n1645 VPWR 0.093504
R13682 VPWR VPWR.n1097 0.093504
R13683 VPWR.n1629 VPWR 0.093504
R13684 VPWR.n1618 VPWR 0.093504
R13685 VPWR VPWR.n1107 0.093504
R13686 VPWR.n1602 VPWR 0.093504
R13687 VPWR.n2598 VPWR 0.0849042
R13688 VPWR.n1112 VPWR.n1109 0.0845517
R13689 VPWR.n147 VPWR.n146 0.0845517
R13690 VPWR.n159 VPWR.n158 0.0845517
R13691 VPWR.n171 VPWR.n170 0.0845517
R13692 VPWR.n183 VPWR.n182 0.0845517
R13693 VPWR.n195 VPWR.n194 0.0845517
R13694 VPWR.n207 VPWR.n206 0.0845517
R13695 VPWR.n219 VPWR.n218 0.0845517
R13696 VPWR.n231 VPWR.n230 0.0845517
R13697 VPWR.n243 VPWR.n242 0.0845517
R13698 VPWR.n255 VPWR.n254 0.0845517
R13699 VPWR.n267 VPWR.n266 0.0845517
R13700 VPWR.n279 VPWR.n278 0.0845517
R13701 VPWR.n282 VPWR.n103 0.0845517
R13702 VPWR.n113 VPWR.n112 0.0845517
R13703 VPWR.n135 VPWR.n134 0.0845517
R13704 VPWR.n124 VPWR.n123 0.0845517
R13705 VPWR.n1728 VPWR.n1067 0.0845517
R13706 VPWR.n1726 VPWR.n1725 0.0845517
R13707 VPWR.n1714 VPWR.n1713 0.0845517
R13708 VPWR.n1701 VPWR.n1700 0.0845517
R13709 VPWR.n1690 VPWR.n1078 0.0845517
R13710 VPWR.n1687 VPWR.n1686 0.0845517
R13711 VPWR.n1674 VPWR.n1673 0.0845517
R13712 VPWR.n1663 VPWR.n1088 0.0845517
R13713 VPWR.n1660 VPWR.n1659 0.0845517
R13714 VPWR.n1647 VPWR.n1646 0.0845517
R13715 VPWR.n1636 VPWR.n1098 0.0845517
R13716 VPWR.n1633 VPWR.n1632 0.0845517
R13717 VPWR.n1620 VPWR.n1619 0.0845517
R13718 VPWR.n1609 VPWR.n1108 0.0845517
R13719 VPWR.n1606 VPWR.n1605 0.0845517
R13720 VPWR.n1456 VPWR.n1451 0.0740128
R13721 VPWR.n1542 VPWR.n1044 0.071
R13722 VPWR.n1547 VPWR.n1541 0.071
R13723 VPWR.n1552 VPWR.n1142 0.071
R13724 VPWR.n1557 VPWR.n1141 0.071
R13725 VPWR.n1562 VPWR.n1140 0.071
R13726 VPWR.n1567 VPWR.n1139 0.071
R13727 VPWR.n1572 VPWR.n1138 0.071
R13728 VPWR.n1577 VPWR.n1137 0.071
R13729 VPWR.n1583 VPWR.n1582 0.071
R13730 VPWR.n1457 VPWR.n1131 0.071
R13731 VPWR.n1463 VPWR.n1462 0.071
R13732 VPWR.n1772 VPWR.n1038 0.071
R13733 VPWR.n1786 VPWR.n1785 0.071
R13734 VPWR.n1780 VPWR.n1027 0.071
R13735 VPWR.n1767 VPWR.n1766 0.071
R13736 VPWR VPWR.n1115 0.0678077
R13737 VPWR VPWR.n107 0.0678077
R13738 VPWR VPWR.n141 0.0678077
R13739 VPWR VPWR.n153 0.0678077
R13740 VPWR VPWR.n165 0.0678077
R13741 VPWR VPWR.n177 0.0678077
R13742 VPWR VPWR.n189 0.0678077
R13743 VPWR VPWR.n201 0.0678077
R13744 VPWR VPWR.n213 0.0678077
R13745 VPWR VPWR.n225 0.0678077
R13746 VPWR VPWR.n237 0.0678077
R13747 VPWR VPWR.n249 0.0678077
R13748 VPWR VPWR.n261 0.0678077
R13749 VPWR VPWR.n273 0.0678077
R13750 VPWR.n286 VPWR 0.0678077
R13751 VPWR VPWR.n129 0.0678077
R13752 VPWR VPWR.n118 0.0678077
R13753 VPWR.n1732 VPWR 0.0678077
R13754 VPWR VPWR.n1720 0.0678077
R13755 VPWR VPWR.n1708 0.0678077
R13756 VPWR VPWR.n1697 0.0678077
R13757 VPWR.n1193 VPWR 0.0678077
R13758 VPWR VPWR.n1681 0.0678077
R13759 VPWR VPWR.n1670 0.0678077
R13760 VPWR.n1207 VPWR 0.0678077
R13761 VPWR VPWR.n1654 0.0678077
R13762 VPWR VPWR.n1643 0.0678077
R13763 VPWR.n1175 VPWR 0.0678077
R13764 VPWR VPWR.n1627 0.0678077
R13765 VPWR VPWR.n1616 0.0678077
R13766 VPWR.n1124 VPWR 0.0678077
R13767 VPWR VPWR.n1600 0.0678077
R13768 VPWR.n150 VPWR 0.063
R13769 VPWR.n162 VPWR 0.063
R13770 VPWR.n174 VPWR 0.063
R13771 VPWR.n186 VPWR 0.063
R13772 VPWR.n198 VPWR 0.063
R13773 VPWR.n210 VPWR 0.063
R13774 VPWR.n222 VPWR 0.063
R13775 VPWR.n234 VPWR 0.063
R13776 VPWR.n246 VPWR 0.063
R13777 VPWR.n258 VPWR 0.063
R13778 VPWR.n270 VPWR 0.063
R13779 VPWR.n101 VPWR 0.063
R13780 VPWR.n105 VPWR 0.063
R13781 VPWR.n138 VPWR 0.063
R13782 VPWR.n115 VPWR 0.063
R13783 VPWR.n126 VPWR 0.063
R13784 VPWR.n1065 VPWR 0.063
R13785 VPWR.n1717 VPWR 0.063
R13786 VPWR.n1070 VPWR 0.063
R13787 VPWR VPWR.n1704 0.063
R13788 VPWR VPWR.n1693 0.063
R13789 VPWR VPWR.n1081 0.063
R13790 VPWR VPWR.n1677 0.063
R13791 VPWR VPWR.n1666 0.063
R13792 VPWR VPWR.n1091 0.063
R13793 VPWR VPWR.n1650 0.063
R13794 VPWR VPWR.n1639 0.063
R13795 VPWR VPWR.n1101 0.063
R13796 VPWR VPWR.n1623 0.063
R13797 VPWR VPWR.n1612 0.063
R13798 VPWR VPWR.n1111 0.063
R13799 VPWR VPWR.n1120 0.063
R13800 VPWR.n1115 VPWR 0.0608448
R13801 VPWR.n107 VPWR 0.0608448
R13802 VPWR.n141 VPWR 0.0608448
R13803 VPWR.n153 VPWR 0.0608448
R13804 VPWR.n165 VPWR 0.0608448
R13805 VPWR.n177 VPWR 0.0608448
R13806 VPWR.n189 VPWR 0.0608448
R13807 VPWR.n201 VPWR 0.0608448
R13808 VPWR.n213 VPWR 0.0608448
R13809 VPWR.n225 VPWR 0.0608448
R13810 VPWR.n237 VPWR 0.0608448
R13811 VPWR.n249 VPWR 0.0608448
R13812 VPWR.n261 VPWR 0.0608448
R13813 VPWR.n273 VPWR 0.0608448
R13814 VPWR.n286 VPWR 0.0608448
R13815 VPWR.n129 VPWR 0.0608448
R13816 VPWR.n118 VPWR 0.0608448
R13817 VPWR.n1732 VPWR 0.0608448
R13818 VPWR.n1720 VPWR 0.0608448
R13819 VPWR.n1708 VPWR 0.0608448
R13820 VPWR.n1697 VPWR 0.0608448
R13821 VPWR.n1193 VPWR 0.0608448
R13822 VPWR.n1681 VPWR 0.0608448
R13823 VPWR.n1670 VPWR 0.0608448
R13824 VPWR.n1207 VPWR 0.0608448
R13825 VPWR.n1654 VPWR 0.0608448
R13826 VPWR.n1643 VPWR 0.0608448
R13827 VPWR.n1175 VPWR 0.0608448
R13828 VPWR.n1627 VPWR 0.0608448
R13829 VPWR.n1616 VPWR 0.0608448
R13830 VPWR.n1124 VPWR 0.0608448
R13831 VPWR.n1600 VPWR 0.0608448
R13832 VPWR VPWR.n13 0.0603958
R13833 VPWR VPWR.n12 0.0603958
R13834 VPWR VPWR.n1249 0.0603958
R13835 VPWR VPWR.n1248 0.0603958
R13836 VPWR VPWR.n1272 0.0603958
R13837 VPWR VPWR.n1271 0.0603958
R13838 VPWR VPWR.n1296 0.0603958
R13839 VPWR VPWR.n1295 0.0603958
R13840 VPWR.n1332 VPWR 0.0603958
R13841 VPWR VPWR.n1331 0.0603958
R13842 VPWR.n1327 VPWR 0.0603958
R13843 VPWR.n1318 VPWR 0.0603958
R13844 VPWR VPWR.n1317 0.0603958
R13845 VPWR.n1370 VPWR 0.0603958
R13846 VPWR VPWR.n1369 0.0603958
R13847 VPWR.n1364 VPWR 0.0603958
R13848 VPWR.n1409 VPWR 0.0603958
R13849 VPWR VPWR.n1408 0.0603958
R13850 VPWR.n1403 VPWR 0.0603958
R13851 VPWR.n1440 VPWR 0.0603958
R13852 VPWR VPWR.n2800 0.0603958
R13853 VPWR VPWR.n2799 0.0603958
R13854 VPWR VPWR.n2812 0.0603958
R13855 VPWR.n2791 VPWR 0.0603958
R13856 VPWR.n2792 VPWR 0.0603958
R13857 VPWR VPWR.n2796 0.0603958
R13858 VPWR.n2771 VPWR 0.0603958
R13859 VPWR.n2772 VPWR 0.0603958
R13860 VPWR VPWR.n2777 0.0603958
R13861 VPWR.n2752 VPWR 0.0603958
R13862 VPWR.n2753 VPWR 0.0603958
R13863 VPWR VPWR.n2757 0.0603958
R13864 VPWR.n2733 VPWR 0.0603958
R13865 VPWR.n2734 VPWR 0.0603958
R13866 VPWR VPWR.n2695 0.0603958
R13867 VPWR.n2696 VPWR 0.0603958
R13868 VPWR.n2697 VPWR 0.0603958
R13869 VPWR VPWR.n2658 0.0603958
R13870 VPWR.n2659 VPWR 0.0603958
R13871 VPWR.n2660 VPWR 0.0603958
R13872 VPWR.n2624 VPWR 0.0603958
R13873 VPWR.n2627 VPWR 0.0603958
R13874 VPWR.n1770 VPWR.n1769 0.0599512
R13875 VPWR.n1041 VPWR.n1040 0.0599512
R13876 VPWR.n1545 VPWR.n1544 0.0599512
R13877 VPWR.n1550 VPWR.n1549 0.0599512
R13878 VPWR.n1555 VPWR.n1554 0.0599512
R13879 VPWR.n1560 VPWR.n1559 0.0599512
R13880 VPWR.n1565 VPWR.n1564 0.0599512
R13881 VPWR.n1570 VPWR.n1569 0.0599512
R13882 VPWR.n1575 VPWR.n1574 0.0599512
R13883 VPWR.n1580 VPWR.n1579 0.0599512
R13884 VPWR.n1135 VPWR.n1134 0.0599512
R13885 VPWR.n1460 VPWR.n1459 0.0599512
R13886 VPWR.n1455 VPWR.n1454 0.0599512
R13887 VPWR.n1775 VPWR.n1774 0.0599512
R13888 VPWR.n1783 VPWR.n1782 0.0599512
R13889 VPWR.n1779 VPWR.n1778 0.0599512
R13890 VPWR.n1118 VPWR.n1117 0.0565345
R13891 VPWR.n1112 VPWR 0.0565345
R13892 VPWR.n144 VPWR.n143 0.0565345
R13893 VPWR.n146 VPWR 0.0565345
R13894 VPWR.n156 VPWR.n155 0.0565345
R13895 VPWR.n158 VPWR 0.0565345
R13896 VPWR.n168 VPWR.n167 0.0565345
R13897 VPWR.n170 VPWR 0.0565345
R13898 VPWR.n180 VPWR.n179 0.0565345
R13899 VPWR.n182 VPWR 0.0565345
R13900 VPWR.n192 VPWR.n191 0.0565345
R13901 VPWR.n194 VPWR 0.0565345
R13902 VPWR.n204 VPWR.n203 0.0565345
R13903 VPWR.n206 VPWR 0.0565345
R13904 VPWR.n216 VPWR.n215 0.0565345
R13905 VPWR.n218 VPWR 0.0565345
R13906 VPWR.n228 VPWR.n227 0.0565345
R13907 VPWR.n230 VPWR 0.0565345
R13908 VPWR.n240 VPWR.n239 0.0565345
R13909 VPWR.n242 VPWR 0.0565345
R13910 VPWR.n252 VPWR.n251 0.0565345
R13911 VPWR.n254 VPWR 0.0565345
R13912 VPWR.n264 VPWR.n263 0.0565345
R13913 VPWR.n266 VPWR 0.0565345
R13914 VPWR.n276 VPWR.n275 0.0565345
R13915 VPWR.n278 VPWR 0.0565345
R13916 VPWR.n285 VPWR.n283 0.0565345
R13917 VPWR.n103 VPWR 0.0565345
R13918 VPWR.n110 VPWR.n109 0.0565345
R13919 VPWR.n112 VPWR 0.0565345
R13920 VPWR.n132 VPWR.n131 0.0565345
R13921 VPWR.n134 VPWR 0.0565345
R13922 VPWR.n121 VPWR.n120 0.0565345
R13923 VPWR.n123 VPWR 0.0565345
R13924 VPWR.n1731 VPWR.n1729 0.0565345
R13925 VPWR.n1067 VPWR 0.0565345
R13926 VPWR.n1723 VPWR.n1722 0.0565345
R13927 VPWR.n1725 VPWR 0.0565345
R13928 VPWR.n1711 VPWR.n1710 0.0565345
R13929 VPWR.n1713 VPWR 0.0565345
R13930 VPWR.n1702 VPWR.n1699 0.0565345
R13931 VPWR.n1700 VPWR 0.0565345
R13932 VPWR.n1691 VPWR.n1077 0.0565345
R13933 VPWR.n1078 VPWR 0.0565345
R13934 VPWR.n1684 VPWR.n1683 0.0565345
R13935 VPWR.n1686 VPWR 0.0565345
R13936 VPWR.n1675 VPWR.n1672 0.0565345
R13937 VPWR.n1673 VPWR 0.0565345
R13938 VPWR.n1664 VPWR.n1087 0.0565345
R13939 VPWR.n1088 VPWR 0.0565345
R13940 VPWR.n1657 VPWR.n1656 0.0565345
R13941 VPWR.n1659 VPWR 0.0565345
R13942 VPWR.n1648 VPWR.n1645 0.0565345
R13943 VPWR.n1646 VPWR 0.0565345
R13944 VPWR.n1637 VPWR.n1097 0.0565345
R13945 VPWR.n1098 VPWR 0.0565345
R13946 VPWR.n1630 VPWR.n1629 0.0565345
R13947 VPWR.n1632 VPWR 0.0565345
R13948 VPWR.n1621 VPWR.n1618 0.0565345
R13949 VPWR.n1619 VPWR 0.0565345
R13950 VPWR.n1610 VPWR.n1107 0.0565345
R13951 VPWR.n1108 VPWR 0.0565345
R13952 VPWR.n1603 VPWR.n1602 0.0565345
R13953 VPWR.n1605 VPWR 0.0565345
R13954 VPWR.n1769 VPWR 0.0469286
R13955 VPWR.n1040 VPWR 0.0469286
R13956 VPWR.n1544 VPWR 0.0469286
R13957 VPWR.n1549 VPWR 0.0469286
R13958 VPWR.n1554 VPWR 0.0469286
R13959 VPWR.n1559 VPWR 0.0469286
R13960 VPWR.n1564 VPWR 0.0469286
R13961 VPWR.n1569 VPWR 0.0469286
R13962 VPWR.n1574 VPWR 0.0469286
R13963 VPWR.n1579 VPWR 0.0469286
R13964 VPWR.n1134 VPWR 0.0469286
R13965 VPWR.n1459 VPWR 0.0469286
R13966 VPWR.n1454 VPWR 0.0469286
R13967 VPWR.n1774 VPWR 0.0469286
R13968 VPWR.n1782 VPWR 0.0469286
R13969 VPWR.n1778 VPWR 0.0469286
R13970 VPWR.n1769 VPWR 0.0401341
R13971 VPWR.n1040 VPWR 0.0401341
R13972 VPWR.n1544 VPWR 0.0401341
R13973 VPWR.n1549 VPWR 0.0401341
R13974 VPWR.n1554 VPWR 0.0401341
R13975 VPWR.n1559 VPWR 0.0401341
R13976 VPWR.n1564 VPWR 0.0401341
R13977 VPWR.n1569 VPWR 0.0401341
R13978 VPWR.n1574 VPWR 0.0401341
R13979 VPWR.n1579 VPWR 0.0401341
R13980 VPWR.n1134 VPWR 0.0401341
R13981 VPWR.n1459 VPWR 0.0401341
R13982 VPWR.n1454 VPWR 0.0401341
R13983 VPWR.n1774 VPWR 0.0401341
R13984 VPWR.n1782 VPWR 0.0401341
R13985 VPWR.n1778 VPWR 0.0401341
R13986 VPWR.n13 VPWR 0.0382604
R13987 VPWR.n1249 VPWR 0.0382604
R13988 VPWR.n1272 VPWR 0.0382604
R13989 VPWR.n1296 VPWR 0.0382604
R13990 VPWR.n1331 VPWR 0.0382604
R13991 VPWR.n1369 VPWR 0.0382604
R13992 VPWR.n1408 VPWR 0.0382604
R13993 VPWR.n1445 VPWR 0.0382604
R13994 VPWR.n20 VPWR 0.0375125
R13995 VPWR.n20 VPWR 0.0373589
R13996 VPWR.n1118 VPWR.n1109 0.0349828
R13997 VPWR.n147 VPWR.n144 0.0349828
R13998 VPWR.n159 VPWR.n156 0.0349828
R13999 VPWR.n171 VPWR.n168 0.0349828
R14000 VPWR.n183 VPWR.n180 0.0349828
R14001 VPWR.n195 VPWR.n192 0.0349828
R14002 VPWR.n207 VPWR.n204 0.0349828
R14003 VPWR.n219 VPWR.n216 0.0349828
R14004 VPWR.n231 VPWR.n228 0.0349828
R14005 VPWR.n243 VPWR.n240 0.0349828
R14006 VPWR.n255 VPWR.n252 0.0349828
R14007 VPWR.n267 VPWR.n264 0.0349828
R14008 VPWR.n279 VPWR.n276 0.0349828
R14009 VPWR.n283 VPWR.n282 0.0349828
R14010 VPWR.n113 VPWR.n110 0.0349828
R14011 VPWR.n135 VPWR.n132 0.0349828
R14012 VPWR.n124 VPWR.n121 0.0349828
R14013 VPWR.n1729 VPWR.n1728 0.0349828
R14014 VPWR.n1726 VPWR.n1723 0.0349828
R14015 VPWR.n1714 VPWR.n1711 0.0349828
R14016 VPWR.n1702 VPWR.n1701 0.0349828
R14017 VPWR.n1691 VPWR.n1690 0.0349828
R14018 VPWR.n1687 VPWR.n1684 0.0349828
R14019 VPWR.n1675 VPWR.n1674 0.0349828
R14020 VPWR.n1664 VPWR.n1663 0.0349828
R14021 VPWR.n1660 VPWR.n1657 0.0349828
R14022 VPWR.n1648 VPWR.n1647 0.0349828
R14023 VPWR.n1637 VPWR.n1636 0.0349828
R14024 VPWR.n1633 VPWR.n1630 0.0349828
R14025 VPWR.n1621 VPWR.n1620 0.0349828
R14026 VPWR.n1610 VPWR.n1609 0.0349828
R14027 VPWR.n1606 VPWR.n1603 0.0349828
R14028 VPWR.n2504 VPWR.n2503 0.0340366
R14029 VPWR.n2570 VPWR.n2569 0.0340366
R14030 VPWR.n2510 VPWR.n2509 0.0340366
R14031 VPWR.n2552 VPWR.n2551 0.0340366
R14032 VPWR.n2546 VPWR.n2545 0.0340366
R14033 VPWR.n2534 VPWR.n2533 0.0340366
R14034 VPWR.n2528 VPWR.n2527 0.0340366
R14035 VPWR.n1223 VPWR.n1222 0.0340366
R14036 VPWR.n2522 VPWR.n2521 0.0340366
R14037 VPWR.n1486 VPWR.n1102 0.0340366
R14038 VPWR.n1174 VPWR.n1094 0.0340366
R14039 VPWR.n2540 VPWR.n2539 0.0340366
R14040 VPWR.n1165 VPWR.n1092 0.0340366
R14041 VPWR.n1211 VPWR.n1164 0.0340366
R14042 VPWR.n2516 VPWR.n2515 0.0340366
R14043 VPWR.n1129 VPWR.n1104 0.0340366
R14044 VPWR.n1155 VPWR.n1084 0.0340366
R14045 VPWR.n2558 VPWR.n2557 0.0340366
R14046 VPWR.n1144 VPWR.n1082 0.0340366
R14047 VPWR.n1591 VPWR.n1590 0.0340366
R14048 VPWR.n2564 VPWR.n2563 0.0340366
R14049 VPWR.n1197 VPWR.n1154 0.0340366
R14050 VPWR.n1074 VPWR.n1073 0.0340366
R14051 VPWR.n1743 VPWR.n1742 0.0340366
R14052 VPWR.n1071 VPWR.n1054 0.0340366
R14053 VPWR.n2576 VPWR.n2575 0.0340366
R14054 VPWR.n2582 VPWR.n2581 0.0340366
R14055 VPWR.n2593 VPWR.n2592 0.0340366
R14056 VPWR.n2588 VPWR.n2587 0.0340366
R14057 VPWR.n1737 VPWR.n1736 0.0340366
R14058 VPWR.n1063 VPWR.n1060 0.0340366
R14059 VPWR.n1596 VPWR.n1121 0.0340366
R14060 VPWR.n2628 VPWR.n2598 0.0320292
R14061 VPWR.n2800 VPWR 0.03175
R14062 VPWR VPWR.n2791 0.03175
R14063 VPWR VPWR.n2771 0.03175
R14064 VPWR VPWR.n2752 0.03175
R14065 VPWR VPWR.n2733 0.03175
R14066 VPWR VPWR.n2696 0.03175
R14067 VPWR VPWR.n2659 0.03175
R14068 VPWR VPWR.n2627 0.03175
R14069 VPWR.n2598 VPWR.n2597 0.0240975
R14070 VPWR.n2597 VPWR.n20 0.0240975
R14071 VPWR.n2814 VPWR 0.024
R14072 VPWR.n14 VPWR 0.0239375
R14073 VPWR.n12 VPWR 0.0239375
R14074 VPWR.n1250 VPWR 0.0239375
R14075 VPWR.n1248 VPWR 0.0239375
R14076 VPWR.n1271 VPWR 0.0239375
R14077 VPWR.n1295 VPWR 0.0239375
R14078 VPWR.n2753 VPWR 0.0239375
R14079 VPWR.n2503 VPWR 0.0233659
R14080 VPWR.n1466 VPWR 0.0233659
R14081 VPWR.n352 VPWR 0.0233659
R14082 VPWR.n2570 VPWR 0.0233659
R14083 VPWR.n1533 VPWR 0.0233659
R14084 VPWR.n347 VPWR 0.0233659
R14085 VPWR.n2510 VPWR 0.0233659
R14086 VPWR.n964 VPWR 0.0233659
R14087 VPWR.n2479 VPWR 0.0233659
R14088 VPWR.n2474 VPWR 0.0233659
R14089 VPWR.n319 VPWR 0.0233659
R14090 VPWR.n2551 VPWR 0.0233659
R14091 VPWR.n972 VPWR 0.0233659
R14092 VPWR.n2444 VPWR 0.0233659
R14093 VPWR.n323 VPWR 0.0233659
R14094 VPWR.n2546 VPWR 0.0233659
R14095 VPWR.n1891 VPWR 0.0233659
R14096 VPWR.n1886 VPWR 0.0233659
R14097 VPWR.n1881 VPWR 0.0233659
R14098 VPWR.n388 VPWR 0.0233659
R14099 VPWR.n392 VPWR 0.0233659
R14100 VPWR.n396 VPWR 0.0233659
R14101 VPWR.n2454 VPWR 0.0233659
R14102 VPWR.n331 VPWR 0.0233659
R14103 VPWR.n2534 VPWR 0.0233659
R14104 VPWR.n1876 VPWR 0.0233659
R14105 VPWR.n404 VPWR 0.0233659
R14106 VPWR.n2459 VPWR 0.0233659
R14107 VPWR.n335 VPWR 0.0233659
R14108 VPWR.n2527 VPWR 0.0233659
R14109 VPWR.n2307 VPWR 0.0233659
R14110 VPWR.n2312 VPWR 0.0233659
R14111 VPWR.n2317 VPWR 0.0233659
R14112 VPWR.n2322 VPWR 0.0233659
R14113 VPWR.n2332 VPWR 0.0233659
R14114 VPWR.n2337 VPWR 0.0233659
R14115 VPWR.n2342 VPWR 0.0233659
R14116 VPWR.n2347 VPWR 0.0233659
R14117 VPWR.n2352 VPWR 0.0233659
R14118 VPWR.n2357 VPWR 0.0233659
R14119 VPWR.n2362 VPWR 0.0233659
R14120 VPWR.n2367 VPWR 0.0233659
R14121 VPWR.n2372 VPWR 0.0233659
R14122 VPWR.n2377 VPWR 0.0233659
R14123 VPWR.n2381 VPWR 0.0233659
R14124 VPWR.n2327 VPWR 0.0233659
R14125 VPWR.n544 VPWR 0.0233659
R14126 VPWR.n539 VPWR 0.0233659
R14127 VPWR.n535 VPWR 0.0233659
R14128 VPWR.n531 VPWR 0.0233659
R14129 VPWR.n523 VPWR 0.0233659
R14130 VPWR.n519 VPWR 0.0233659
R14131 VPWR.n515 VPWR 0.0233659
R14132 VPWR.n511 VPWR 0.0233659
R14133 VPWR.n507 VPWR 0.0233659
R14134 VPWR.n503 VPWR 0.0233659
R14135 VPWR.n499 VPWR 0.0233659
R14136 VPWR.n495 VPWR 0.0233659
R14137 VPWR.n491 VPWR 0.0233659
R14138 VPWR.n487 VPWR 0.0233659
R14139 VPWR.n484 VPWR 0.0233659
R14140 VPWR.n527 VPWR 0.0233659
R14141 VPWR.n2283 VPWR 0.0233659
R14142 VPWR.n2278 VPWR 0.0233659
R14143 VPWR.n2273 VPWR 0.0233659
R14144 VPWR.n2268 VPWR 0.0233659
R14145 VPWR.n2258 VPWR 0.0233659
R14146 VPWR.n2253 VPWR 0.0233659
R14147 VPWR.n2248 VPWR 0.0233659
R14148 VPWR.n2243 VPWR 0.0233659
R14149 VPWR.n2238 VPWR 0.0233659
R14150 VPWR.n2233 VPWR 0.0233659
R14151 VPWR.n2228 VPWR 0.0233659
R14152 VPWR.n2223 VPWR 0.0233659
R14153 VPWR.n2218 VPWR 0.0233659
R14154 VPWR.n2213 VPWR 0.0233659
R14155 VPWR.n2209 VPWR 0.0233659
R14156 VPWR.n2263 VPWR 0.0233659
R14157 VPWR.n580 VPWR 0.0233659
R14158 VPWR.n584 VPWR 0.0233659
R14159 VPWR.n588 VPWR 0.0233659
R14160 VPWR.n592 VPWR 0.0233659
R14161 VPWR.n600 VPWR 0.0233659
R14162 VPWR.n604 VPWR 0.0233659
R14163 VPWR.n608 VPWR 0.0233659
R14164 VPWR.n612 VPWR 0.0233659
R14165 VPWR.n616 VPWR 0.0233659
R14166 VPWR.n620 VPWR 0.0233659
R14167 VPWR.n624 VPWR 0.0233659
R14168 VPWR.n628 VPWR 0.0233659
R14169 VPWR.n632 VPWR 0.0233659
R14170 VPWR.n636 VPWR 0.0233659
R14171 VPWR.n640 VPWR 0.0233659
R14172 VPWR.n596 VPWR 0.0233659
R14173 VPWR.n2111 VPWR 0.0233659
R14174 VPWR.n2116 VPWR 0.0233659
R14175 VPWR.n2121 VPWR 0.0233659
R14176 VPWR.n2126 VPWR 0.0233659
R14177 VPWR.n2136 VPWR 0.0233659
R14178 VPWR.n2141 VPWR 0.0233659
R14179 VPWR.n2146 VPWR 0.0233659
R14180 VPWR.n2151 VPWR 0.0233659
R14181 VPWR.n2156 VPWR 0.0233659
R14182 VPWR.n2161 VPWR 0.0233659
R14183 VPWR.n2166 VPWR 0.0233659
R14184 VPWR.n2171 VPWR 0.0233659
R14185 VPWR.n2176 VPWR 0.0233659
R14186 VPWR.n2181 VPWR 0.0233659
R14187 VPWR.n2185 VPWR 0.0233659
R14188 VPWR.n2131 VPWR 0.0233659
R14189 VPWR.n736 VPWR 0.0233659
R14190 VPWR.n731 VPWR 0.0233659
R14191 VPWR.n727 VPWR 0.0233659
R14192 VPWR.n723 VPWR 0.0233659
R14193 VPWR.n715 VPWR 0.0233659
R14194 VPWR.n711 VPWR 0.0233659
R14195 VPWR.n707 VPWR 0.0233659
R14196 VPWR.n703 VPWR 0.0233659
R14197 VPWR.n699 VPWR 0.0233659
R14198 VPWR.n695 VPWR 0.0233659
R14199 VPWR.n691 VPWR 0.0233659
R14200 VPWR.n687 VPWR 0.0233659
R14201 VPWR.n683 VPWR 0.0233659
R14202 VPWR.n679 VPWR 0.0233659
R14203 VPWR.n676 VPWR 0.0233659
R14204 VPWR.n719 VPWR 0.0233659
R14205 VPWR.n2087 VPWR 0.0233659
R14206 VPWR.n2082 VPWR 0.0233659
R14207 VPWR.n2077 VPWR 0.0233659
R14208 VPWR.n2072 VPWR 0.0233659
R14209 VPWR.n2062 VPWR 0.0233659
R14210 VPWR.n2057 VPWR 0.0233659
R14211 VPWR.n2052 VPWR 0.0233659
R14212 VPWR.n2047 VPWR 0.0233659
R14213 VPWR.n2042 VPWR 0.0233659
R14214 VPWR.n2037 VPWR 0.0233659
R14215 VPWR.n2032 VPWR 0.0233659
R14216 VPWR.n2027 VPWR 0.0233659
R14217 VPWR.n2022 VPWR 0.0233659
R14218 VPWR.n2017 VPWR 0.0233659
R14219 VPWR.n2013 VPWR 0.0233659
R14220 VPWR.n2067 VPWR 0.0233659
R14221 VPWR.n772 VPWR 0.0233659
R14222 VPWR.n776 VPWR 0.0233659
R14223 VPWR.n780 VPWR 0.0233659
R14224 VPWR.n784 VPWR 0.0233659
R14225 VPWR.n792 VPWR 0.0233659
R14226 VPWR.n796 VPWR 0.0233659
R14227 VPWR.n800 VPWR 0.0233659
R14228 VPWR.n804 VPWR 0.0233659
R14229 VPWR.n808 VPWR 0.0233659
R14230 VPWR.n812 VPWR 0.0233659
R14231 VPWR.n816 VPWR 0.0233659
R14232 VPWR.n820 VPWR 0.0233659
R14233 VPWR.n824 VPWR 0.0233659
R14234 VPWR.n828 VPWR 0.0233659
R14235 VPWR.n832 VPWR 0.0233659
R14236 VPWR.n788 VPWR 0.0233659
R14237 VPWR.n1915 VPWR 0.0233659
R14238 VPWR.n1920 VPWR 0.0233659
R14239 VPWR.n1925 VPWR 0.0233659
R14240 VPWR.n1930 VPWR 0.0233659
R14241 VPWR.n1940 VPWR 0.0233659
R14242 VPWR.n1945 VPWR 0.0233659
R14243 VPWR.n1950 VPWR 0.0233659
R14244 VPWR.n1955 VPWR 0.0233659
R14245 VPWR.n1960 VPWR 0.0233659
R14246 VPWR.n1965 VPWR 0.0233659
R14247 VPWR.n1970 VPWR 0.0233659
R14248 VPWR.n1975 VPWR 0.0233659
R14249 VPWR.n1980 VPWR 0.0233659
R14250 VPWR.n1985 VPWR 0.0233659
R14251 VPWR.n1989 VPWR 0.0233659
R14252 VPWR.n1935 VPWR 0.0233659
R14253 VPWR.n928 VPWR 0.0233659
R14254 VPWR.n923 VPWR 0.0233659
R14255 VPWR.n919 VPWR 0.0233659
R14256 VPWR.n915 VPWR 0.0233659
R14257 VPWR.n907 VPWR 0.0233659
R14258 VPWR.n903 VPWR 0.0233659
R14259 VPWR.n899 VPWR 0.0233659
R14260 VPWR.n895 VPWR 0.0233659
R14261 VPWR.n891 VPWR 0.0233659
R14262 VPWR.n887 VPWR 0.0233659
R14263 VPWR.n883 VPWR 0.0233659
R14264 VPWR.n879 VPWR 0.0233659
R14265 VPWR.n875 VPWR 0.0233659
R14266 VPWR.n871 VPWR 0.0233659
R14267 VPWR.n868 VPWR 0.0233659
R14268 VPWR.n911 VPWR 0.0233659
R14269 VPWR.n1871 VPWR 0.0233659
R14270 VPWR.n980 VPWR 0.0233659
R14271 VPWR.n1495 VPWR 0.0233659
R14272 VPWR.n1223 VPWR 0.0233659
R14273 VPWR.n400 VPWR 0.0233659
R14274 VPWR.n2464 VPWR 0.0233659
R14275 VPWR.n339 VPWR 0.0233659
R14276 VPWR.n2522 VPWR 0.0233659
R14277 VPWR.n976 VPWR 0.0233659
R14278 VPWR.n1490 VPWR 0.0233659
R14279 VPWR.n1486 VPWR 0.0233659
R14280 VPWR.n1866 VPWR 0.0233659
R14281 VPWR.n984 VPWR 0.0233659
R14282 VPWR.n1504 VPWR 0.0233659
R14283 VPWR.n1174 VPWR 0.0233659
R14284 VPWR.n408 VPWR 0.0233659
R14285 VPWR.n416 VPWR 0.0233659
R14286 VPWR.n420 VPWR 0.0233659
R14287 VPWR.n424 VPWR 0.0233659
R14288 VPWR.n428 VPWR 0.0233659
R14289 VPWR.n432 VPWR 0.0233659
R14290 VPWR.n436 VPWR 0.0233659
R14291 VPWR.n440 VPWR 0.0233659
R14292 VPWR.n444 VPWR 0.0233659
R14293 VPWR.n448 VPWR 0.0233659
R14294 VPWR.n412 VPWR 0.0233659
R14295 VPWR.n2449 VPWR 0.0233659
R14296 VPWR.n327 VPWR 0.0233659
R14297 VPWR.n2539 VPWR 0.0233659
R14298 VPWR.n988 VPWR 0.0233659
R14299 VPWR.n1509 VPWR 0.0233659
R14300 VPWR.n1165 VPWR 0.0233659
R14301 VPWR.n1861 VPWR 0.0233659
R14302 VPWR.n1851 VPWR 0.0233659
R14303 VPWR.n1846 VPWR 0.0233659
R14304 VPWR.n1841 VPWR 0.0233659
R14305 VPWR.n1836 VPWR 0.0233659
R14306 VPWR.n1831 VPWR 0.0233659
R14307 VPWR.n1826 VPWR 0.0233659
R14308 VPWR.n1821 VPWR 0.0233659
R14309 VPWR.n1817 VPWR 0.0233659
R14310 VPWR.n1856 VPWR 0.0233659
R14311 VPWR.n992 VPWR 0.0233659
R14312 VPWR.n1518 VPWR 0.0233659
R14313 VPWR.n1164 VPWR 0.0233659
R14314 VPWR.n2469 VPWR 0.0233659
R14315 VPWR.n343 VPWR 0.0233659
R14316 VPWR.n2515 VPWR 0.0233659
R14317 VPWR.n1130 VPWR 0.0233659
R14318 VPWR.n1129 VPWR 0.0233659
R14319 VPWR.n996 VPWR 0.0233659
R14320 VPWR.n1523 VPWR 0.0233659
R14321 VPWR.n1155 VPWR 0.0233659
R14322 VPWR.n2439 VPWR 0.0233659
R14323 VPWR.n2429 VPWR 0.0233659
R14324 VPWR.n2424 VPWR 0.0233659
R14325 VPWR.n2419 VPWR 0.0233659
R14326 VPWR.n2414 VPWR 0.0233659
R14327 VPWR.n2409 VPWR 0.0233659
R14328 VPWR.n2405 VPWR 0.0233659
R14329 VPWR.n2434 VPWR 0.0233659
R14330 VPWR.n315 VPWR 0.0233659
R14331 VPWR.n2558 VPWR 0.0233659
R14332 VPWR.n1538 VPWR 0.0233659
R14333 VPWR.n1144 VPWR 0.0233659
R14334 VPWR.n1000 VPWR 0.0233659
R14335 VPWR.n1004 VPWR 0.0233659
R14336 VPWR.n1008 VPWR 0.0233659
R14337 VPWR.n1012 VPWR 0.0233659
R14338 VPWR.n1016 VPWR 0.0233659
R14339 VPWR.n1020 VPWR 0.0233659
R14340 VPWR.n1024 VPWR 0.0233659
R14341 VPWR.n968 VPWR 0.0233659
R14342 VPWR.n1473 VPWR 0.0233659
R14343 VPWR.n1590 VPWR 0.0233659
R14344 VPWR.n311 VPWR 0.0233659
R14345 VPWR.n2563 VPWR 0.0233659
R14346 VPWR.n1154 VPWR 0.0233659
R14347 VPWR.n1763 VPWR 0.0233659
R14348 VPWR.n1073 VPWR 0.0233659
R14349 VPWR.n307 VPWR 0.0233659
R14350 VPWR.n303 VPWR 0.0233659
R14351 VPWR.n295 VPWR 0.0233659
R14352 VPWR.n292 VPWR 0.0233659
R14353 VPWR.n299 VPWR 0.0233659
R14354 VPWR.n1743 VPWR 0.0233659
R14355 VPWR.n1751 VPWR 0.0233659
R14356 VPWR.n1789 VPWR 0.0233659
R14357 VPWR.n1793 VPWR 0.0233659
R14358 VPWR.n1758 VPWR 0.0233659
R14359 VPWR.n1054 VPWR 0.0233659
R14360 VPWR.n2575 VPWR 0.0233659
R14361 VPWR.n2582 VPWR 0.0233659
R14362 VPWR.n2593 VPWR 0.0233659
R14363 VPWR.n2587 VPWR 0.0233659
R14364 VPWR.n1736 VPWR 0.0233659
R14365 VPWR.n1060 VPWR 0.0233659
R14366 VPWR.n1121 VPWR 0.0233659
R14367 VPWR.n1336 VPWR 0.0226354
R14368 VPWR.n1327 VPWR 0.0226354
R14369 VPWR.n1413 VPWR 0.0226354
R14370 VPWR.n2772 VPWR 0.0226354
R14371 VPWR VPWR.n2732 0.0226354
R14372 VPWR VPWR.n2702 0.0226354
R14373 VPWR VPWR.n2664 0.0226354
R14374 VPWR VPWR.n64 0.0220517
R14375 VPWR VPWR.n67 0.0220517
R14376 VPWR VPWR.n70 0.0220517
R14377 VPWR VPWR.n73 0.0220517
R14378 VPWR VPWR.n76 0.0220517
R14379 VPWR VPWR.n79 0.0220517
R14380 VPWR VPWR.n82 0.0220517
R14381 VPWR VPWR.n85 0.0220517
R14382 VPWR VPWR.n88 0.0220517
R14383 VPWR VPWR.n91 0.0220517
R14384 VPWR VPWR.n94 0.0220517
R14385 VPWR VPWR.n97 0.0220517
R14386 VPWR.n289 VPWR 0.0220517
R14387 VPWR VPWR.n61 0.0220517
R14388 VPWR VPWR.n58 0.0220517
R14389 VPWR.n1735 VPWR 0.0220517
R14390 VPWR VPWR.n1057 0.0220517
R14391 VPWR.n1705 VPWR 0.0220517
R14392 VPWR.n1694 VPWR 0.0220517
R14393 VPWR.n1196 VPWR 0.0220517
R14394 VPWR.n1678 VPWR 0.0220517
R14395 VPWR.n1667 VPWR 0.0220517
R14396 VPWR.n1210 VPWR 0.0220517
R14397 VPWR.n1651 VPWR 0.0220517
R14398 VPWR.n1640 VPWR 0.0220517
R14399 VPWR.n1178 VPWR 0.0220517
R14400 VPWR.n1624 VPWR 0.0220517
R14401 VPWR.n1613 VPWR 0.0220517
R14402 VPWR.n1127 VPWR 0.0220517
R14403 VPWR.n1597 VPWR 0.0220517
R14404 VPWR.n1273 VPWR 0.0213333
R14405 VPWR.n1297 VPWR 0.0213333
R14406 VPWR.n1311 VPWR 0.0213333
R14407 VPWR.n1375 VPWR 0.0213333
R14408 VPWR.n1347 VPWR 0.0213333
R14409 VPWR.n1386 VPWR 0.0213333
R14410 VPWR.n1423 VPWR 0.0213333
R14411 VPWR.n2806 VPWR 0.0213333
R14412 VPWR.n2799 VPWR 0.0213333
R14413 VPWR VPWR.n2790 0.0213333
R14414 VPWR.n2792 VPWR 0.0213333
R14415 VPWR VPWR.n2770 0.0213333
R14416 VPWR VPWR.n2751 0.0213333
R14417 VPWR VPWR.n2738 0.0213333
R14418 VPWR.n2500 VPWR 0.0196917
R14419 VPWR.n24 VPWR 0.0143889
R14420 VPWR VPWR.n19 0.0099
R14421 VPWR VPWR.n1604 0.00397222
R14422 VPWR VPWR.n1105 0.00397222
R14423 VPWR VPWR.n1103 0.00397222
R14424 VPWR VPWR.n1631 0.00397222
R14425 VPWR VPWR.n1095 0.00397222
R14426 VPWR VPWR.n1093 0.00397222
R14427 VPWR VPWR.n1658 0.00397222
R14428 VPWR VPWR.n1085 0.00397222
R14429 VPWR VPWR.n1083 0.00397222
R14430 VPWR VPWR.n1685 0.00397222
R14431 VPWR VPWR.n1075 0.00397222
R14432 VPWR VPWR.n1072 0.00397222
R14433 VPWR VPWR.n1712 0.00397222
R14434 VPWR VPWR.n1724 0.00397222
R14435 VPWR.n1113 VPWR 0.00397222
R14436 VPWR VPWR.n1066 0.00397222
R14437 VPWR VPWR.n122 0.00397222
R14438 VPWR VPWR.n111 0.00397222
R14439 VPWR VPWR.n102 0.00397222
R14440 VPWR VPWR.n277 0.00397222
R14441 VPWR VPWR.n265 0.00397222
R14442 VPWR VPWR.n253 0.00397222
R14443 VPWR VPWR.n241 0.00397222
R14444 VPWR VPWR.n229 0.00397222
R14445 VPWR VPWR.n217 0.00397222
R14446 VPWR VPWR.n205 0.00397222
R14447 VPWR VPWR.n193 0.00397222
R14448 VPWR VPWR.n181 0.00397222
R14449 VPWR VPWR.n169 0.00397222
R14450 VPWR VPWR.n157 0.00397222
R14451 VPWR VPWR.n145 0.00397222
R14452 VPWR VPWR.n133 0.00397222
R14453 VPWR.n1462 VPWR.n1461 0.00351282
R14454 VPWR.n1457 VPWR.n1136 0.00351282
R14455 VPWR.n1582 VPWR.n1581 0.00351282
R14456 VPWR.n1577 VPWR.n1576 0.00351282
R14457 VPWR.n1572 VPWR.n1571 0.00351282
R14458 VPWR.n1567 VPWR.n1566 0.00351282
R14459 VPWR.n1562 VPWR.n1561 0.00351282
R14460 VPWR.n1557 VPWR.n1556 0.00351282
R14461 VPWR.n1552 VPWR.n1551 0.00351282
R14462 VPWR.n1547 VPWR.n1546 0.00351282
R14463 VPWR.n1542 VPWR.n1042 0.00351282
R14464 VPWR.n1785 VPWR.n1784 0.00351282
R14465 VPWR.n1776 VPWR.n1772 0.00351282
R14466 VPWR.n1771 VPWR.n1767 0.00351282
R14467 VPWR.n141 VPWR.n140 0.00265517
R14468 VPWR.n153 VPWR.n152 0.00265517
R14469 VPWR.n165 VPWR.n164 0.00265517
R14470 VPWR.n177 VPWR.n176 0.00265517
R14471 VPWR.n189 VPWR.n188 0.00265517
R14472 VPWR.n201 VPWR.n200 0.00265517
R14473 VPWR.n213 VPWR.n212 0.00265517
R14474 VPWR.n225 VPWR.n224 0.00265517
R14475 VPWR.n237 VPWR.n236 0.00265517
R14476 VPWR.n249 VPWR.n248 0.00265517
R14477 VPWR.n261 VPWR.n260 0.00265517
R14478 VPWR.n273 VPWR.n272 0.00265517
R14479 VPWR.n288 VPWR.n286 0.00265517
R14480 VPWR.n129 VPWR.n128 0.00265517
R14481 VPWR.n118 VPWR.n117 0.00265517
R14482 VPWR.n1734 VPWR.n1732 0.00265517
R14483 VPWR.n1720 VPWR.n1719 0.00265517
R14484 VPWR.n1708 VPWR.n1707 0.00265517
R14485 VPWR.n1697 VPWR.n1696 0.00265517
R14486 VPWR.n1195 VPWR.n1193 0.00265517
R14487 VPWR.n1681 VPWR.n1680 0.00265517
R14488 VPWR.n1670 VPWR.n1669 0.00265517
R14489 VPWR.n1209 VPWR.n1207 0.00265517
R14490 VPWR.n1654 VPWR.n1653 0.00265517
R14491 VPWR.n1643 VPWR.n1642 0.00265517
R14492 VPWR.n1177 VPWR.n1175 0.00265517
R14493 VPWR.n1627 VPWR.n1626 0.00265517
R14494 VPWR.n1616 VPWR.n1615 0.00265517
R14495 VPWR.n1126 VPWR.n1124 0.00265517
R14496 VPWR.n1600 VPWR.n1599 0.00265517
R14497 Iout.n1020 Iout.t144 239.927
R14498 Iout.n509 Iout.t98 239.927
R14499 Iout.n513 Iout.t130 239.927
R14500 Iout.n507 Iout.t171 239.927
R14501 Iout.n504 Iout.t115 239.927
R14502 Iout.n500 Iout.t23 239.927
R14503 Iout.n192 Iout.t233 239.927
R14504 Iout.n195 Iout.t167 239.927
R14505 Iout.n199 Iout.t57 239.927
R14506 Iout.n202 Iout.t19 239.927
R14507 Iout.n206 Iout.t226 239.927
R14508 Iout.n210 Iout.t131 239.927
R14509 Iout.n214 Iout.t91 239.927
R14510 Iout.n218 Iout.t146 239.927
R14511 Iout.n222 Iout.t32 239.927
R14512 Iout.n226 Iout.t117 239.927
R14513 Iout.n232 Iout.t172 239.927
R14514 Iout.n235 Iout.t178 239.927
R14515 Iout.n238 Iout.t3 239.927
R14516 Iout.n241 Iout.t119 239.927
R14517 Iout.n244 Iout.t50 239.927
R14518 Iout.n247 Iout.t13 239.927
R14519 Iout.n250 Iout.t5 239.927
R14520 Iout.n255 Iout.t157 239.927
R14521 Iout.n252 Iout.t99 239.927
R14522 Iout.n489 Iout.t8 239.927
R14523 Iout.n494 Iout.t197 239.927
R14524 Iout.n491 Iout.t145 239.927
R14525 Iout.n519 Iout.t212 239.927
R14526 Iout.n149 Iout.t16 239.927
R14527 Iout.n146 Iout.t79 239.927
R14528 Iout.n1010 Iout.t189 239.927
R14529 Iout.n1007 Iout.t15 239.927
R14530 Iout.n140 Iout.t118 239.927
R14531 Iout.n143 Iout.t64 239.927
R14532 Iout.n525 Iout.t22 239.927
R14533 Iout.n480 Iout.t186 239.927
R14534 Iout.n483 Iout.t169 239.927
R14535 Iout.n478 Iout.t17 239.927
R14536 Iout.n259 Iout.t147 239.927
R14537 Iout.n186 Iout.t33 239.927
R14538 Iout.n271 Iout.t107 239.927
R14539 Iout.n180 Iout.t235 239.927
R14540 Iout.n283 Iout.t225 239.927
R14541 Iout.n174 Iout.t137 239.927
R14542 Iout.n168 Iout.t239 239.927
R14543 Iout.n301 Iout.t74 239.927
R14544 Iout.n289 Iout.t222 239.927
R14545 Iout.n177 Iout.t1 239.927
R14546 Iout.n277 Iout.t53 239.927
R14547 Iout.n183 Iout.t88 239.927
R14548 Iout.n265 Iout.t238 239.927
R14549 Iout.n189 Iout.t182 239.927
R14550 Iout.n472 Iout.t149 239.927
R14551 Iout.n469 Iout.t77 239.927
R14552 Iout.n156 Iout.t72 239.927
R14553 Iout.n531 Iout.t35 239.927
R14554 Iout.n534 Iout.t111 239.927
R14555 Iout.n536 Iout.t92 239.927
R14556 Iout.n133 Iout.t21 239.927
R14557 Iout.n136 Iout.t100 239.927
R14558 Iout.n542 Iout.t123 239.927
R14559 Iout.n460 Iout.t188 239.927
R14560 Iout.n463 Iout.t20 239.927
R14561 Iout.n458 Iout.t241 239.927
R14562 Iout.n305 Iout.t102 239.927
R14563 Iout.n308 Iout.t87 239.927
R14564 Iout.n311 Iout.t175 239.927
R14565 Iout.n314 Iout.t204 239.927
R14566 Iout.n317 Iout.t28 239.927
R14567 Iout.n320 Iout.t94 239.927
R14568 Iout.n392 Iout.t247 239.927
R14569 Iout.n378 Iout.t38 239.927
R14570 Iout.n376 Iout.t231 239.927
R14571 Iout.n394 Iout.t7 239.927
R14572 Iout.n408 Iout.t10 239.927
R14573 Iout.n410 Iout.t135 239.927
R14574 Iout.n424 Iout.t105 239.927
R14575 Iout.n426 Iout.t45 239.927
R14576 Iout.n447 Iout.t67 239.927
R14577 Iout.n452 Iout.t248 239.927
R14578 Iout.n449 Iout.t127 239.927
R14579 Iout.n548 Iout.t54 239.927
R14580 Iout.n130 Iout.t103 239.927
R14581 Iout.n559 Iout.t63 239.927
R14582 Iout.n557 Iout.t114 239.927
R14583 Iout.n554 Iout.t195 239.927
R14584 Iout.n434 Iout.t140 239.927
R14585 Iout.n438 Iout.t192 239.927
R14586 Iout.n441 Iout.t213 239.927
R14587 Iout.n432 Iout.t240 239.927
R14588 Iout.n418 Iout.t143 239.927
R14589 Iout.n416 Iout.t132 239.927
R14590 Iout.n402 Iout.t196 239.927
R14591 Iout.n357 Iout.t252 239.927
R14592 Iout.n360 Iout.t158 239.927
R14593 Iout.n363 Iout.t148 239.927
R14594 Iout.n366 Iout.t89 239.927
R14595 Iout.n354 Iout.t136 239.927
R14596 Iout.n351 Iout.t108 239.927
R14597 Iout.n348 Iout.t26 239.927
R14598 Iout.n345 Iout.t207 239.927
R14599 Iout.n342 Iout.t124 239.927
R14600 Iout.n339 Iout.t223 239.927
R14601 Iout.n336 Iout.t253 239.927
R14602 Iout.n333 Iout.t191 239.927
R14603 Iout.n117 Iout.t206 239.927
R14604 Iout.n582 Iout.t184 239.927
R14605 Iout.n111 Iout.t255 239.927
R14606 Iout.n594 Iout.t71 239.927
R14607 Iout.n105 Iout.t237 239.927
R14608 Iout.n606 Iout.t101 239.927
R14609 Iout.n99 Iout.t249 239.927
R14610 Iout.n618 Iout.t160 239.927
R14611 Iout.n624 Iout.t168 239.927
R14612 Iout.n90 Iout.t113 239.927
R14613 Iout.n636 Iout.t155 239.927
R14614 Iout.n81 Iout.t62 239.927
R14615 Iout.n648 Iout.t120 239.927
R14616 Iout.n96 Iout.t112 239.927
R14617 Iout.n612 Iout.t61 239.927
R14618 Iout.n102 Iout.t156 239.927
R14619 Iout.n600 Iout.t78 239.927
R14620 Iout.n108 Iout.t229 239.927
R14621 Iout.n588 Iout.t30 239.927
R14622 Iout.n687 Iout.t211 239.927
R14623 Iout.n684 Iout.t161 239.927
R14624 Iout.n681 Iout.t106 239.927
R14625 Iout.n678 Iout.t202 239.927
R14626 Iout.n675 Iout.t34 239.927
R14627 Iout.n672 Iout.t173 239.927
R14628 Iout.n747 Iout.t4 239.927
R14629 Iout.n50 Iout.t209 239.927
R14630 Iout.n759 Iout.t25 239.927
R14631 Iout.n44 Iout.t215 239.927
R14632 Iout.n771 Iout.t84 239.927
R14633 Iout.n42 Iout.t125 239.927
R14634 Iout.n56 Iout.t109 239.927
R14635 Iout.n735 Iout.t218 239.927
R14636 Iout.n62 Iout.t27 239.927
R14637 Iout.n723 Iout.t210 239.927
R14638 Iout.n717 Iout.t44 239.927
R14639 Iout.n65 Iout.t224 239.927
R14640 Iout.n729 Iout.t90 239.927
R14641 Iout.n59 Iout.t185 239.927
R14642 Iout.n805 Iout.t42 239.927
R14643 Iout.n808 Iout.t242 239.927
R14644 Iout.n811 Iout.t31 239.927
R14645 Iout.n814 Iout.t153 239.927
R14646 Iout.n817 Iout.t52 239.927
R14647 Iout.n820 Iout.t40 239.927
R14648 Iout.n823 Iout.t232 239.927
R14649 Iout.n802 Iout.t246 239.927
R14650 Iout.n799 Iout.t174 239.927
R14651 Iout.n890 Iout.t110 239.927
R14652 Iout.n888 Iout.t29 239.927
R14653 Iout.n881 Iout.t183 239.927
R14654 Iout.n869 Iout.t214 239.927
R14655 Iout.n867 Iout.t43 239.927
R14656 Iout.n855 Iout.t181 239.927
R14657 Iout.n853 Iout.t141 239.927
R14658 Iout.n841 Iout.t65 239.927
R14659 Iout.n839 Iout.t0 239.927
R14660 Iout.n827 Iout.t251 239.927
R14661 Iout.n883 Iout.t126 239.927
R14662 Iout.n895 Iout.t236 239.927
R14663 Iout.n897 Iout.t14 239.927
R14664 Iout.n909 Iout.t49 239.927
R14665 Iout.n911 Iout.t39 239.927
R14666 Iout.n923 Iout.t250 239.927
R14667 Iout.n926 Iout.t219 239.927
R14668 Iout.n22 Iout.t150 239.927
R14669 Iout.n876 Iout.t69 239.927
R14670 Iout.n874 Iout.t95 239.927
R14671 Iout.n862 Iout.t70 239.927
R14672 Iout.n860 Iout.t76 239.927
R14673 Iout.n848 Iout.t180 239.927
R14674 Iout.n846 Iout.t151 239.927
R14675 Iout.n834 Iout.t199 239.927
R14676 Iout.n832 Iout.t243 239.927
R14677 Iout.n902 Iout.t85 239.927
R14678 Iout.n904 Iout.t228 239.927
R14679 Iout.n916 Iout.t176 239.927
R14680 Iout.n918 Iout.t12 239.927
R14681 Iout.n931 Iout.t82 239.927
R14682 Iout.n934 Iout.t234 239.927
R14683 Iout.n796 Iout.t51 239.927
R14684 Iout.n793 Iout.t166 239.927
R14685 Iout.n790 Iout.t133 239.927
R14686 Iout.n787 Iout.t6 239.927
R14687 Iout.n784 Iout.t121 239.927
R14688 Iout.n781 Iout.t221 239.927
R14689 Iout.n938 Iout.t60 239.927
R14690 Iout.n741 Iout.t122 239.927
R14691 Iout.n53 Iout.t205 239.927
R14692 Iout.n753 Iout.t104 239.927
R14693 Iout.n47 Iout.t227 239.927
R14694 Iout.n765 Iout.t97 239.927
R14695 Iout.n38 Iout.t59 239.927
R14696 Iout.n777 Iout.t152 239.927
R14697 Iout.n71 Iout.t83 239.927
R14698 Iout.n705 Iout.t208 239.927
R14699 Iout.n77 Iout.t194 239.927
R14700 Iout.n944 Iout.t75 239.927
R14701 Iout.n19 Iout.t142 239.927
R14702 Iout.n68 Iout.t179 239.927
R14703 Iout.n711 Iout.t193 239.927
R14704 Iout.n74 Iout.t24 239.927
R14705 Iout.n699 Iout.t47 239.927
R14706 Iout.n950 Iout.t230 239.927
R14707 Iout.n953 Iout.t68 239.927
R14708 Iout.n669 Iout.t138 239.927
R14709 Iout.n666 Iout.t56 239.927
R14710 Iout.n663 Iout.t93 239.927
R14711 Iout.n660 Iout.t73 239.927
R14712 Iout.n657 Iout.t11 239.927
R14713 Iout.n654 Iout.t2 239.927
R14714 Iout.n690 Iout.t245 239.927
R14715 Iout.n695 Iout.t200 239.927
R14716 Iout.n692 Iout.t177 239.927
R14717 Iout.n957 Iout.t159 239.927
R14718 Iout.n114 Iout.t216 239.927
R14719 Iout.n576 Iout.t198 239.927
R14720 Iout.n573 Iout.t187 239.927
R14721 Iout.n963 Iout.t203 239.927
R14722 Iout.n14 Iout.t162 239.927
R14723 Iout.n93 Iout.t36 239.927
R14724 Iout.n630 Iout.t163 239.927
R14725 Iout.n87 Iout.t18 239.927
R14726 Iout.n642 Iout.t116 239.927
R14727 Iout.n85 Iout.t41 239.927
R14728 Iout.n563 Iout.t96 239.927
R14729 Iout.n969 Iout.t129 239.927
R14730 Iout.n972 Iout.t165 239.927
R14731 Iout.n569 Iout.t86 239.927
R14732 Iout.n123 Iout.t220 239.927
R14733 Iout.n120 Iout.t164 239.927
R14734 Iout.n976 Iout.t190 239.927
R14735 Iout.n400 Iout.t128 239.927
R14736 Iout.n386 Iout.t66 239.927
R14737 Iout.n384 Iout.t170 239.927
R14738 Iout.n370 Iout.t217 239.927
R14739 Iout.n982 Iout.t9 239.927
R14740 Iout.n9 Iout.t244 239.927
R14741 Iout.n127 Iout.t139 239.927
R14742 Iout.n988 Iout.t80 239.927
R14743 Iout.n991 Iout.t37 239.927
R14744 Iout.n323 Iout.t134 239.927
R14745 Iout.n326 Iout.t55 239.927
R14746 Iout.n329 Iout.t254 239.927
R14747 Iout.n995 Iout.t201 239.927
R14748 Iout.n1001 Iout.t46 239.927
R14749 Iout.n4 Iout.t58 239.927
R14750 Iout.n295 Iout.t81 239.927
R14751 Iout.n172 Iout.t154 239.927
R14752 Iout.n1014 Iout.t48 239.927
R14753 Iout.n1021 Iout.n1020 7.9105
R14754 Iout.n510 Iout.n509 7.9105
R14755 Iout.n514 Iout.n513 7.9105
R14756 Iout.n508 Iout.n507 7.9105
R14757 Iout.n505 Iout.n504 7.9105
R14758 Iout.n501 Iout.n500 7.9105
R14759 Iout.n193 Iout.n192 7.9105
R14760 Iout.n196 Iout.n195 7.9105
R14761 Iout.n200 Iout.n199 7.9105
R14762 Iout.n203 Iout.n202 7.9105
R14763 Iout.n207 Iout.n206 7.9105
R14764 Iout.n211 Iout.n210 7.9105
R14765 Iout.n215 Iout.n214 7.9105
R14766 Iout.n219 Iout.n218 7.9105
R14767 Iout.n223 Iout.n222 7.9105
R14768 Iout.n227 Iout.n226 7.9105
R14769 Iout.n233 Iout.n232 7.9105
R14770 Iout.n236 Iout.n235 7.9105
R14771 Iout.n239 Iout.n238 7.9105
R14772 Iout.n242 Iout.n241 7.9105
R14773 Iout.n245 Iout.n244 7.9105
R14774 Iout.n248 Iout.n247 7.9105
R14775 Iout.n251 Iout.n250 7.9105
R14776 Iout.n256 Iout.n255 7.9105
R14777 Iout.n253 Iout.n252 7.9105
R14778 Iout.n490 Iout.n489 7.9105
R14779 Iout.n495 Iout.n494 7.9105
R14780 Iout.n492 Iout.n491 7.9105
R14781 Iout.n520 Iout.n519 7.9105
R14782 Iout.n150 Iout.n149 7.9105
R14783 Iout.n147 Iout.n146 7.9105
R14784 Iout.n1011 Iout.n1010 7.9105
R14785 Iout.n1008 Iout.n1007 7.9105
R14786 Iout.n141 Iout.n140 7.9105
R14787 Iout.n144 Iout.n143 7.9105
R14788 Iout.n526 Iout.n525 7.9105
R14789 Iout.n481 Iout.n480 7.9105
R14790 Iout.n484 Iout.n483 7.9105
R14791 Iout.n479 Iout.n478 7.9105
R14792 Iout.n260 Iout.n259 7.9105
R14793 Iout.n187 Iout.n186 7.9105
R14794 Iout.n272 Iout.n271 7.9105
R14795 Iout.n181 Iout.n180 7.9105
R14796 Iout.n284 Iout.n283 7.9105
R14797 Iout.n175 Iout.n174 7.9105
R14798 Iout.n169 Iout.n168 7.9105
R14799 Iout.n302 Iout.n301 7.9105
R14800 Iout.n290 Iout.n289 7.9105
R14801 Iout.n178 Iout.n177 7.9105
R14802 Iout.n278 Iout.n277 7.9105
R14803 Iout.n184 Iout.n183 7.9105
R14804 Iout.n266 Iout.n265 7.9105
R14805 Iout.n190 Iout.n189 7.9105
R14806 Iout.n473 Iout.n472 7.9105
R14807 Iout.n470 Iout.n469 7.9105
R14808 Iout.n157 Iout.n156 7.9105
R14809 Iout.n532 Iout.n531 7.9105
R14810 Iout.n535 Iout.n534 7.9105
R14811 Iout.n537 Iout.n536 7.9105
R14812 Iout.n134 Iout.n133 7.9105
R14813 Iout.n137 Iout.n136 7.9105
R14814 Iout.n543 Iout.n542 7.9105
R14815 Iout.n461 Iout.n460 7.9105
R14816 Iout.n464 Iout.n463 7.9105
R14817 Iout.n459 Iout.n458 7.9105
R14818 Iout.n306 Iout.n305 7.9105
R14819 Iout.n309 Iout.n308 7.9105
R14820 Iout.n312 Iout.n311 7.9105
R14821 Iout.n315 Iout.n314 7.9105
R14822 Iout.n318 Iout.n317 7.9105
R14823 Iout.n321 Iout.n320 7.9105
R14824 Iout.n393 Iout.n392 7.9105
R14825 Iout.n379 Iout.n378 7.9105
R14826 Iout.n377 Iout.n376 7.9105
R14827 Iout.n395 Iout.n394 7.9105
R14828 Iout.n409 Iout.n408 7.9105
R14829 Iout.n411 Iout.n410 7.9105
R14830 Iout.n425 Iout.n424 7.9105
R14831 Iout.n427 Iout.n426 7.9105
R14832 Iout.n448 Iout.n447 7.9105
R14833 Iout.n453 Iout.n452 7.9105
R14834 Iout.n450 Iout.n449 7.9105
R14835 Iout.n549 Iout.n548 7.9105
R14836 Iout.n131 Iout.n130 7.9105
R14837 Iout.n560 Iout.n559 7.9105
R14838 Iout.n558 Iout.n557 7.9105
R14839 Iout.n555 Iout.n554 7.9105
R14840 Iout.n435 Iout.n434 7.9105
R14841 Iout.n439 Iout.n438 7.9105
R14842 Iout.n442 Iout.n441 7.9105
R14843 Iout.n433 Iout.n432 7.9105
R14844 Iout.n419 Iout.n418 7.9105
R14845 Iout.n417 Iout.n416 7.9105
R14846 Iout.n403 Iout.n402 7.9105
R14847 Iout.n358 Iout.n357 7.9105
R14848 Iout.n361 Iout.n360 7.9105
R14849 Iout.n364 Iout.n363 7.9105
R14850 Iout.n367 Iout.n366 7.9105
R14851 Iout.n355 Iout.n354 7.9105
R14852 Iout.n352 Iout.n351 7.9105
R14853 Iout.n349 Iout.n348 7.9105
R14854 Iout.n346 Iout.n345 7.9105
R14855 Iout.n343 Iout.n342 7.9105
R14856 Iout.n340 Iout.n339 7.9105
R14857 Iout.n337 Iout.n336 7.9105
R14858 Iout.n334 Iout.n333 7.9105
R14859 Iout.n118 Iout.n117 7.9105
R14860 Iout.n583 Iout.n582 7.9105
R14861 Iout.n112 Iout.n111 7.9105
R14862 Iout.n595 Iout.n594 7.9105
R14863 Iout.n106 Iout.n105 7.9105
R14864 Iout.n607 Iout.n606 7.9105
R14865 Iout.n100 Iout.n99 7.9105
R14866 Iout.n619 Iout.n618 7.9105
R14867 Iout.n625 Iout.n624 7.9105
R14868 Iout.n91 Iout.n90 7.9105
R14869 Iout.n637 Iout.n636 7.9105
R14870 Iout.n82 Iout.n81 7.9105
R14871 Iout.n649 Iout.n648 7.9105
R14872 Iout.n97 Iout.n96 7.9105
R14873 Iout.n613 Iout.n612 7.9105
R14874 Iout.n103 Iout.n102 7.9105
R14875 Iout.n601 Iout.n600 7.9105
R14876 Iout.n109 Iout.n108 7.9105
R14877 Iout.n589 Iout.n588 7.9105
R14878 Iout.n688 Iout.n687 7.9105
R14879 Iout.n685 Iout.n684 7.9105
R14880 Iout.n682 Iout.n681 7.9105
R14881 Iout.n679 Iout.n678 7.9105
R14882 Iout.n676 Iout.n675 7.9105
R14883 Iout.n673 Iout.n672 7.9105
R14884 Iout.n748 Iout.n747 7.9105
R14885 Iout.n51 Iout.n50 7.9105
R14886 Iout.n760 Iout.n759 7.9105
R14887 Iout.n45 Iout.n44 7.9105
R14888 Iout.n772 Iout.n771 7.9105
R14889 Iout.n43 Iout.n42 7.9105
R14890 Iout.n57 Iout.n56 7.9105
R14891 Iout.n736 Iout.n735 7.9105
R14892 Iout.n63 Iout.n62 7.9105
R14893 Iout.n724 Iout.n723 7.9105
R14894 Iout.n718 Iout.n717 7.9105
R14895 Iout.n66 Iout.n65 7.9105
R14896 Iout.n730 Iout.n729 7.9105
R14897 Iout.n60 Iout.n59 7.9105
R14898 Iout.n806 Iout.n805 7.9105
R14899 Iout.n809 Iout.n808 7.9105
R14900 Iout.n812 Iout.n811 7.9105
R14901 Iout.n815 Iout.n814 7.9105
R14902 Iout.n818 Iout.n817 7.9105
R14903 Iout.n821 Iout.n820 7.9105
R14904 Iout.n824 Iout.n823 7.9105
R14905 Iout.n803 Iout.n802 7.9105
R14906 Iout.n800 Iout.n799 7.9105
R14907 Iout.n891 Iout.n890 7.9105
R14908 Iout.n889 Iout.n888 7.9105
R14909 Iout.n882 Iout.n881 7.9105
R14910 Iout.n870 Iout.n869 7.9105
R14911 Iout.n868 Iout.n867 7.9105
R14912 Iout.n856 Iout.n855 7.9105
R14913 Iout.n854 Iout.n853 7.9105
R14914 Iout.n842 Iout.n841 7.9105
R14915 Iout.n840 Iout.n839 7.9105
R14916 Iout.n828 Iout.n827 7.9105
R14917 Iout.n884 Iout.n883 7.9105
R14918 Iout.n896 Iout.n895 7.9105
R14919 Iout.n898 Iout.n897 7.9105
R14920 Iout.n910 Iout.n909 7.9105
R14921 Iout.n912 Iout.n911 7.9105
R14922 Iout.n924 Iout.n923 7.9105
R14923 Iout.n927 Iout.n926 7.9105
R14924 Iout.n23 Iout.n22 7.9105
R14925 Iout.n877 Iout.n876 7.9105
R14926 Iout.n875 Iout.n874 7.9105
R14927 Iout.n863 Iout.n862 7.9105
R14928 Iout.n861 Iout.n860 7.9105
R14929 Iout.n849 Iout.n848 7.9105
R14930 Iout.n847 Iout.n846 7.9105
R14931 Iout.n835 Iout.n834 7.9105
R14932 Iout.n833 Iout.n832 7.9105
R14933 Iout.n903 Iout.n902 7.9105
R14934 Iout.n905 Iout.n904 7.9105
R14935 Iout.n917 Iout.n916 7.9105
R14936 Iout.n919 Iout.n918 7.9105
R14937 Iout.n932 Iout.n931 7.9105
R14938 Iout.n935 Iout.n934 7.9105
R14939 Iout.n797 Iout.n796 7.9105
R14940 Iout.n794 Iout.n793 7.9105
R14941 Iout.n791 Iout.n790 7.9105
R14942 Iout.n788 Iout.n787 7.9105
R14943 Iout.n785 Iout.n784 7.9105
R14944 Iout.n782 Iout.n781 7.9105
R14945 Iout.n939 Iout.n938 7.9105
R14946 Iout.n742 Iout.n741 7.9105
R14947 Iout.n54 Iout.n53 7.9105
R14948 Iout.n754 Iout.n753 7.9105
R14949 Iout.n48 Iout.n47 7.9105
R14950 Iout.n766 Iout.n765 7.9105
R14951 Iout.n39 Iout.n38 7.9105
R14952 Iout.n778 Iout.n777 7.9105
R14953 Iout.n72 Iout.n71 7.9105
R14954 Iout.n706 Iout.n705 7.9105
R14955 Iout.n78 Iout.n77 7.9105
R14956 Iout.n945 Iout.n944 7.9105
R14957 Iout.n20 Iout.n19 7.9105
R14958 Iout.n69 Iout.n68 7.9105
R14959 Iout.n712 Iout.n711 7.9105
R14960 Iout.n75 Iout.n74 7.9105
R14961 Iout.n700 Iout.n699 7.9105
R14962 Iout.n951 Iout.n950 7.9105
R14963 Iout.n954 Iout.n953 7.9105
R14964 Iout.n670 Iout.n669 7.9105
R14965 Iout.n667 Iout.n666 7.9105
R14966 Iout.n664 Iout.n663 7.9105
R14967 Iout.n661 Iout.n660 7.9105
R14968 Iout.n658 Iout.n657 7.9105
R14969 Iout.n655 Iout.n654 7.9105
R14970 Iout.n691 Iout.n690 7.9105
R14971 Iout.n696 Iout.n695 7.9105
R14972 Iout.n693 Iout.n692 7.9105
R14973 Iout.n958 Iout.n957 7.9105
R14974 Iout.n115 Iout.n114 7.9105
R14975 Iout.n577 Iout.n576 7.9105
R14976 Iout.n574 Iout.n573 7.9105
R14977 Iout.n964 Iout.n963 7.9105
R14978 Iout.n15 Iout.n14 7.9105
R14979 Iout.n94 Iout.n93 7.9105
R14980 Iout.n631 Iout.n630 7.9105
R14981 Iout.n88 Iout.n87 7.9105
R14982 Iout.n643 Iout.n642 7.9105
R14983 Iout.n86 Iout.n85 7.9105
R14984 Iout.n564 Iout.n563 7.9105
R14985 Iout.n970 Iout.n969 7.9105
R14986 Iout.n973 Iout.n972 7.9105
R14987 Iout.n570 Iout.n569 7.9105
R14988 Iout.n124 Iout.n123 7.9105
R14989 Iout.n121 Iout.n120 7.9105
R14990 Iout.n977 Iout.n976 7.9105
R14991 Iout.n401 Iout.n400 7.9105
R14992 Iout.n387 Iout.n386 7.9105
R14993 Iout.n385 Iout.n384 7.9105
R14994 Iout.n371 Iout.n370 7.9105
R14995 Iout.n983 Iout.n982 7.9105
R14996 Iout.n10 Iout.n9 7.9105
R14997 Iout.n128 Iout.n127 7.9105
R14998 Iout.n989 Iout.n988 7.9105
R14999 Iout.n992 Iout.n991 7.9105
R15000 Iout.n324 Iout.n323 7.9105
R15001 Iout.n327 Iout.n326 7.9105
R15002 Iout.n330 Iout.n329 7.9105
R15003 Iout.n996 Iout.n995 7.9105
R15004 Iout.n1002 Iout.n1001 7.9105
R15005 Iout.n5 Iout.n4 7.9105
R15006 Iout.n296 Iout.n295 7.9105
R15007 Iout.n173 Iout.n172 7.9105
R15008 Iout.n1015 Iout.n1014 7.9105
R15009 Iout.n886 Iout.n885 3.86101
R15010 Iout.n880 Iout.n879 3.86101
R15011 Iout.n894 Iout.n893 3.86101
R15012 Iout.n872 Iout.n871 3.86101
R15013 Iout.n900 Iout.n899 3.86101
R15014 Iout.n866 Iout.n865 3.86101
R15015 Iout.n908 Iout.n907 3.86101
R15016 Iout.n858 Iout.n857 3.86101
R15017 Iout.n914 Iout.n913 3.86101
R15018 Iout.n852 Iout.n851 3.86101
R15019 Iout.n922 Iout.n921 3.86101
R15020 Iout.n844 Iout.n843 3.86101
R15021 Iout.n929 Iout.n928 3.86101
R15022 Iout.n838 Iout.n837 3.86101
R15023 Iout.n925 Iout.n21 3.86101
R15024 Iout.n830 Iout.n829 3.86101
R15025 Iout.n879 Iout.n878 3.4105
R15026 Iout.n887 Iout.n886 3.4105
R15027 Iout.n893 Iout.n892 3.4105
R15028 Iout.n798 Iout.n28 3.4105
R15029 Iout.n801 Iout.n29 3.4105
R15030 Iout.n804 Iout.n30 3.4105
R15031 Iout.n807 Iout.n31 3.4105
R15032 Iout.n873 Iout.n872 3.4105
R15033 Iout.n744 Iout.n743 3.4105
R15034 Iout.n740 Iout.n739 3.4105
R15035 Iout.n732 Iout.n731 3.4105
R15036 Iout.n728 Iout.n727 3.4105
R15037 Iout.n720 Iout.n719 3.4105
R15038 Iout.n795 Iout.n27 3.4105
R15039 Iout.n901 Iout.n900 3.4105
R15040 Iout.n722 Iout.n721 3.4105
R15041 Iout.n726 Iout.n725 3.4105
R15042 Iout.n734 Iout.n733 3.4105
R15043 Iout.n738 Iout.n737 3.4105
R15044 Iout.n746 Iout.n745 3.4105
R15045 Iout.n750 Iout.n749 3.4105
R15046 Iout.n752 Iout.n751 3.4105
R15047 Iout.n810 Iout.n32 3.4105
R15048 Iout.n865 Iout.n864 3.4105
R15049 Iout.n668 Iout.n55 3.4105
R15050 Iout.n671 Iout.n58 3.4105
R15051 Iout.n674 Iout.n61 3.4105
R15052 Iout.n677 Iout.n64 3.4105
R15053 Iout.n680 Iout.n67 3.4105
R15054 Iout.n683 Iout.n70 3.4105
R15055 Iout.n686 Iout.n73 3.4105
R15056 Iout.n714 Iout.n713 3.4105
R15057 Iout.n716 Iout.n715 3.4105
R15058 Iout.n792 Iout.n26 3.4105
R15059 Iout.n907 Iout.n906 3.4105
R15060 Iout.n587 Iout.n586 3.4105
R15061 Iout.n591 Iout.n590 3.4105
R15062 Iout.n599 Iout.n598 3.4105
R15063 Iout.n603 Iout.n602 3.4105
R15064 Iout.n611 Iout.n610 3.4105
R15065 Iout.n615 Iout.n614 3.4105
R15066 Iout.n623 Iout.n622 3.4105
R15067 Iout.n627 Iout.n626 3.4105
R15068 Iout.n665 Iout.n52 3.4105
R15069 Iout.n758 Iout.n757 3.4105
R15070 Iout.n756 Iout.n755 3.4105
R15071 Iout.n813 Iout.n33 3.4105
R15072 Iout.n859 Iout.n858 3.4105
R15073 Iout.n629 Iout.n628 3.4105
R15074 Iout.n621 Iout.n620 3.4105
R15075 Iout.n617 Iout.n616 3.4105
R15076 Iout.n609 Iout.n608 3.4105
R15077 Iout.n605 Iout.n604 3.4105
R15078 Iout.n597 Iout.n596 3.4105
R15079 Iout.n593 Iout.n592 3.4105
R15080 Iout.n585 Iout.n584 3.4105
R15081 Iout.n581 Iout.n580 3.4105
R15082 Iout.n579 Iout.n578 3.4105
R15083 Iout.n689 Iout.n76 3.4105
R15084 Iout.n710 Iout.n709 3.4105
R15085 Iout.n708 Iout.n707 3.4105
R15086 Iout.n789 Iout.n25 3.4105
R15087 Iout.n915 Iout.n914 3.4105
R15088 Iout.n572 Iout.n571 3.4105
R15089 Iout.n335 Iout.n116 3.4105
R15090 Iout.n338 Iout.n113 3.4105
R15091 Iout.n341 Iout.n110 3.4105
R15092 Iout.n344 Iout.n107 3.4105
R15093 Iout.n347 Iout.n104 3.4105
R15094 Iout.n350 Iout.n101 3.4105
R15095 Iout.n353 Iout.n98 3.4105
R15096 Iout.n356 Iout.n95 3.4105
R15097 Iout.n359 Iout.n92 3.4105
R15098 Iout.n633 Iout.n632 3.4105
R15099 Iout.n635 Iout.n634 3.4105
R15100 Iout.n662 Iout.n49 3.4105
R15101 Iout.n762 Iout.n761 3.4105
R15102 Iout.n764 Iout.n763 3.4105
R15103 Iout.n816 Iout.n34 3.4105
R15104 Iout.n851 Iout.n850 3.4105
R15105 Iout.n399 Iout.n398 3.4105
R15106 Iout.n405 Iout.n404 3.4105
R15107 Iout.n415 Iout.n414 3.4105
R15108 Iout.n421 Iout.n420 3.4105
R15109 Iout.n431 Iout.n430 3.4105
R15110 Iout.n444 Iout.n443 3.4105
R15111 Iout.n440 Iout.n159 3.4105
R15112 Iout.n437 Iout.n436 3.4105
R15113 Iout.n553 Iout.n552 3.4105
R15114 Iout.n556 Iout.n119 3.4105
R15115 Iout.n562 Iout.n561 3.4105
R15116 Iout.n568 Iout.n567 3.4105
R15117 Iout.n566 Iout.n565 3.4105
R15118 Iout.n575 Iout.n79 3.4105
R15119 Iout.n698 Iout.n697 3.4105
R15120 Iout.n702 Iout.n701 3.4105
R15121 Iout.n704 Iout.n703 3.4105
R15122 Iout.n786 Iout.n24 3.4105
R15123 Iout.n921 Iout.n920 3.4105
R15124 Iout.n129 Iout.n125 3.4105
R15125 Iout.n547 Iout.n546 3.4105
R15126 Iout.n551 Iout.n550 3.4105
R15127 Iout.n451 Iout.n158 3.4105
R15128 Iout.n455 Iout.n454 3.4105
R15129 Iout.n446 Iout.n445 3.4105
R15130 Iout.n429 Iout.n428 3.4105
R15131 Iout.n423 Iout.n422 3.4105
R15132 Iout.n413 Iout.n412 3.4105
R15133 Iout.n407 Iout.n406 3.4105
R15134 Iout.n397 Iout.n396 3.4105
R15135 Iout.n391 Iout.n390 3.4105
R15136 Iout.n389 Iout.n388 3.4105
R15137 Iout.n362 Iout.n89 3.4105
R15138 Iout.n641 Iout.n640 3.4105
R15139 Iout.n639 Iout.n638 3.4105
R15140 Iout.n659 Iout.n46 3.4105
R15141 Iout.n770 Iout.n769 3.4105
R15142 Iout.n768 Iout.n767 3.4105
R15143 Iout.n819 Iout.n35 3.4105
R15144 Iout.n845 Iout.n844 3.4105
R15145 Iout.n325 Iout.n165 3.4105
R15146 Iout.n322 Iout.n164 3.4105
R15147 Iout.n319 Iout.n163 3.4105
R15148 Iout.n316 Iout.n162 3.4105
R15149 Iout.n313 Iout.n161 3.4105
R15150 Iout.n310 Iout.n160 3.4105
R15151 Iout.n307 Iout.n155 3.4105
R15152 Iout.n457 Iout.n456 3.4105
R15153 Iout.n466 Iout.n465 3.4105
R15154 Iout.n462 Iout.n126 3.4105
R15155 Iout.n545 Iout.n544 3.4105
R15156 Iout.n541 Iout.n540 3.4105
R15157 Iout.n135 Iout.n3 3.4105
R15158 Iout.n987 Iout.n986 3.4105
R15159 Iout.n985 Iout.n984 3.4105
R15160 Iout.n122 Iout.n8 3.4105
R15161 Iout.n968 Iout.n967 3.4105
R15162 Iout.n966 Iout.n965 3.4105
R15163 Iout.n694 Iout.n13 3.4105
R15164 Iout.n949 Iout.n948 3.4105
R15165 Iout.n947 Iout.n946 3.4105
R15166 Iout.n783 Iout.n18 3.4105
R15167 Iout.n930 Iout.n929 3.4105
R15168 Iout.n1004 Iout.n1003 3.4105
R15169 Iout.n539 Iout.n538 3.4105
R15170 Iout.n533 Iout.n132 3.4105
R15171 Iout.n530 Iout.n529 3.4105
R15172 Iout.n468 Iout.n467 3.4105
R15173 Iout.n471 Iout.n153 3.4105
R15174 Iout.n475 Iout.n474 3.4105
R15175 Iout.n264 Iout.n263 3.4105
R15176 Iout.n268 Iout.n267 3.4105
R15177 Iout.n276 Iout.n275 3.4105
R15178 Iout.n280 Iout.n279 3.4105
R15179 Iout.n288 Iout.n287 3.4105
R15180 Iout.n292 Iout.n291 3.4105
R15181 Iout.n300 Iout.n299 3.4105
R15182 Iout.n328 Iout.n166 3.4105
R15183 Iout.n381 Iout.n380 3.4105
R15184 Iout.n383 Iout.n382 3.4105
R15185 Iout.n365 Iout.n83 3.4105
R15186 Iout.n645 Iout.n644 3.4105
R15187 Iout.n647 Iout.n646 3.4105
R15188 Iout.n656 Iout.n40 3.4105
R15189 Iout.n774 Iout.n773 3.4105
R15190 Iout.n776 Iout.n775 3.4105
R15191 Iout.n822 Iout.n36 3.4105
R15192 Iout.n837 Iout.n836 3.4105
R15193 Iout.n298 Iout.n297 3.4105
R15194 Iout.n294 Iout.n293 3.4105
R15195 Iout.n286 Iout.n285 3.4105
R15196 Iout.n282 Iout.n281 3.4105
R15197 Iout.n274 Iout.n273 3.4105
R15198 Iout.n270 Iout.n269 3.4105
R15199 Iout.n262 Iout.n261 3.4105
R15200 Iout.n477 Iout.n476 3.4105
R15201 Iout.n486 Iout.n485 3.4105
R15202 Iout.n482 Iout.n151 3.4105
R15203 Iout.n528 Iout.n527 3.4105
R15204 Iout.n524 Iout.n523 3.4105
R15205 Iout.n142 Iout.n138 3.4105
R15206 Iout.n1006 Iout.n1005 3.4105
R15207 Iout.n1009 Iout.n0 3.4105
R15208 Iout.n1000 Iout.n999 3.4105
R15209 Iout.n998 Iout.n997 3.4105
R15210 Iout.n990 Iout.n6 3.4105
R15211 Iout.n981 Iout.n980 3.4105
R15212 Iout.n979 Iout.n978 3.4105
R15213 Iout.n971 Iout.n11 3.4105
R15214 Iout.n962 Iout.n961 3.4105
R15215 Iout.n960 Iout.n959 3.4105
R15216 Iout.n952 Iout.n16 3.4105
R15217 Iout.n943 Iout.n942 3.4105
R15218 Iout.n941 Iout.n940 3.4105
R15219 Iout.n933 Iout.n21 3.4105
R15220 Iout.n1017 Iout.n1016 3.4105
R15221 Iout.n148 Iout.n2 3.4105
R15222 Iout.n518 Iout.n517 3.4105
R15223 Iout.n522 Iout.n521 3.4105
R15224 Iout.n493 Iout.n139 3.4105
R15225 Iout.n497 Iout.n496 3.4105
R15226 Iout.n488 Iout.n487 3.4105
R15227 Iout.n254 Iout.n154 3.4105
R15228 Iout.n258 Iout.n257 3.4105
R15229 Iout.n249 Iout.n188 3.4105
R15230 Iout.n246 Iout.n185 3.4105
R15231 Iout.n243 Iout.n182 3.4105
R15232 Iout.n240 Iout.n179 3.4105
R15233 Iout.n237 Iout.n176 3.4105
R15234 Iout.n234 Iout.n170 3.4105
R15235 Iout.n231 Iout.n230 3.4105
R15236 Iout.n171 Iout.n167 3.4105
R15237 Iout.n304 Iout.n303 3.4105
R15238 Iout.n332 Iout.n331 3.4105
R15239 Iout.n375 Iout.n374 3.4105
R15240 Iout.n373 Iout.n372 3.4105
R15241 Iout.n369 Iout.n368 3.4105
R15242 Iout.n84 Iout.n80 3.4105
R15243 Iout.n651 Iout.n650 3.4105
R15244 Iout.n653 Iout.n652 3.4105
R15245 Iout.n41 Iout.n37 3.4105
R15246 Iout.n780 Iout.n779 3.4105
R15247 Iout.n826 Iout.n825 3.4105
R15248 Iout.n831 Iout.n830 3.4105
R15249 Iout.n229 Iout.n228 3.4105
R15250 Iout.n225 Iout.n224 3.4105
R15251 Iout.n221 Iout.n220 3.4105
R15252 Iout.n217 Iout.n216 3.4105
R15253 Iout.n213 Iout.n212 3.4105
R15254 Iout.n209 Iout.n208 3.4105
R15255 Iout.n205 Iout.n204 3.4105
R15256 Iout.n201 Iout.n191 3.4105
R15257 Iout.n198 Iout.n197 3.4105
R15258 Iout.n194 Iout.n152 3.4105
R15259 Iout.n499 Iout.n498 3.4105
R15260 Iout.n503 Iout.n502 3.4105
R15261 Iout.n506 Iout.n145 3.4105
R15262 Iout.n516 Iout.n515 3.4105
R15263 Iout.n512 Iout.n511 3.4105
R15264 Iout.n1019 Iout.n1018 3.4105
R15265 Iout.n936 Iout.n23 1.43848
R15266 Iout.n936 Iout.n935 1.34612
R15267 Iout.n939 Iout.n937 1.34612
R15268 Iout.n20 Iout.n17 1.34612
R15269 Iout.n955 Iout.n954 1.34612
R15270 Iout.n958 Iout.n956 1.34612
R15271 Iout.n15 Iout.n12 1.34612
R15272 Iout.n974 Iout.n973 1.34612
R15273 Iout.n977 Iout.n975 1.34612
R15274 Iout.n10 Iout.n7 1.34612
R15275 Iout.n993 Iout.n992 1.34612
R15276 Iout.n996 Iout.n994 1.34612
R15277 Iout.n5 Iout.n1 1.34612
R15278 Iout.n1012 Iout.n1011 1.34612
R15279 Iout.n1015 Iout.n1013 1.34612
R15280 Iout.n1022 Iout.n1021 1.34612
R15281 Iout.n197 Iout.n154 0.451012
R15282 Iout.n476 Iout.n154 0.451012
R15283 Iout.n476 Iout.n475 0.451012
R15284 Iout.n475 Iout.n155 0.451012
R15285 Iout.n445 Iout.n155 0.451012
R15286 Iout.n445 Iout.n444 0.451012
R15287 Iout.n444 Iout.n107 0.451012
R15288 Iout.n604 Iout.n107 0.451012
R15289 Iout.n604 Iout.n603 0.451012
R15290 Iout.n603 Iout.n64 0.451012
R15291 Iout.n733 Iout.n64 0.451012
R15292 Iout.n733 Iout.n732 0.451012
R15293 Iout.n732 Iout.n29 0.451012
R15294 Iout.n886 Iout.n29 0.451012
R15295 Iout.n258 Iout.n191 0.451012
R15296 Iout.n262 Iout.n258 0.451012
R15297 Iout.n263 Iout.n262 0.451012
R15298 Iout.n263 Iout.n160 0.451012
R15299 Iout.n429 Iout.n160 0.451012
R15300 Iout.n430 Iout.n429 0.451012
R15301 Iout.n430 Iout.n104 0.451012
R15302 Iout.n609 Iout.n104 0.451012
R15303 Iout.n610 Iout.n609 0.451012
R15304 Iout.n610 Iout.n61 0.451012
R15305 Iout.n738 Iout.n61 0.451012
R15306 Iout.n739 Iout.n738 0.451012
R15307 Iout.n739 Iout.n30 0.451012
R15308 Iout.n879 Iout.n30 0.451012
R15309 Iout.n487 Iout.n152 0.451012
R15310 Iout.n487 Iout.n486 0.451012
R15311 Iout.n486 Iout.n153 0.451012
R15312 Iout.n456 Iout.n153 0.451012
R15313 Iout.n456 Iout.n455 0.451012
R15314 Iout.n455 Iout.n159 0.451012
R15315 Iout.n159 Iout.n110 0.451012
R15316 Iout.n597 Iout.n110 0.451012
R15317 Iout.n598 Iout.n597 0.451012
R15318 Iout.n598 Iout.n67 0.451012
R15319 Iout.n726 Iout.n67 0.451012
R15320 Iout.n727 Iout.n726 0.451012
R15321 Iout.n727 Iout.n28 0.451012
R15322 Iout.n893 Iout.n28 0.451012
R15323 Iout.n204 Iout.n188 0.451012
R15324 Iout.n269 Iout.n188 0.451012
R15325 Iout.n269 Iout.n268 0.451012
R15326 Iout.n268 Iout.n161 0.451012
R15327 Iout.n422 Iout.n161 0.451012
R15328 Iout.n422 Iout.n421 0.451012
R15329 Iout.n421 Iout.n101 0.451012
R15330 Iout.n616 Iout.n101 0.451012
R15331 Iout.n616 Iout.n615 0.451012
R15332 Iout.n615 Iout.n58 0.451012
R15333 Iout.n745 Iout.n58 0.451012
R15334 Iout.n745 Iout.n744 0.451012
R15335 Iout.n744 Iout.n31 0.451012
R15336 Iout.n872 Iout.n31 0.451012
R15337 Iout.n498 Iout.n497 0.451012
R15338 Iout.n497 Iout.n151 0.451012
R15339 Iout.n467 Iout.n151 0.451012
R15340 Iout.n467 Iout.n466 0.451012
R15341 Iout.n466 Iout.n158 0.451012
R15342 Iout.n436 Iout.n158 0.451012
R15343 Iout.n436 Iout.n113 0.451012
R15344 Iout.n592 Iout.n113 0.451012
R15345 Iout.n592 Iout.n591 0.451012
R15346 Iout.n591 Iout.n70 0.451012
R15347 Iout.n721 Iout.n70 0.451012
R15348 Iout.n721 Iout.n720 0.451012
R15349 Iout.n720 Iout.n27 0.451012
R15350 Iout.n900 Iout.n27 0.451012
R15351 Iout.n208 Iout.n185 0.451012
R15352 Iout.n274 Iout.n185 0.451012
R15353 Iout.n275 Iout.n274 0.451012
R15354 Iout.n275 Iout.n162 0.451012
R15355 Iout.n413 Iout.n162 0.451012
R15356 Iout.n414 Iout.n413 0.451012
R15357 Iout.n414 Iout.n98 0.451012
R15358 Iout.n621 Iout.n98 0.451012
R15359 Iout.n622 Iout.n621 0.451012
R15360 Iout.n622 Iout.n55 0.451012
R15361 Iout.n750 Iout.n55 0.451012
R15362 Iout.n751 Iout.n750 0.451012
R15363 Iout.n751 Iout.n32 0.451012
R15364 Iout.n865 Iout.n32 0.451012
R15365 Iout.n502 Iout.n139 0.451012
R15366 Iout.n528 Iout.n139 0.451012
R15367 Iout.n529 Iout.n528 0.451012
R15368 Iout.n529 Iout.n126 0.451012
R15369 Iout.n551 Iout.n126 0.451012
R15370 Iout.n552 Iout.n551 0.451012
R15371 Iout.n552 Iout.n116 0.451012
R15372 Iout.n585 Iout.n116 0.451012
R15373 Iout.n586 Iout.n585 0.451012
R15374 Iout.n586 Iout.n73 0.451012
R15375 Iout.n714 Iout.n73 0.451012
R15376 Iout.n715 Iout.n714 0.451012
R15377 Iout.n715 Iout.n26 0.451012
R15378 Iout.n907 Iout.n26 0.451012
R15379 Iout.n212 Iout.n182 0.451012
R15380 Iout.n281 Iout.n182 0.451012
R15381 Iout.n281 Iout.n280 0.451012
R15382 Iout.n280 Iout.n163 0.451012
R15383 Iout.n406 Iout.n163 0.451012
R15384 Iout.n406 Iout.n405 0.451012
R15385 Iout.n405 Iout.n95 0.451012
R15386 Iout.n628 Iout.n95 0.451012
R15387 Iout.n628 Iout.n627 0.451012
R15388 Iout.n627 Iout.n52 0.451012
R15389 Iout.n757 Iout.n52 0.451012
R15390 Iout.n757 Iout.n756 0.451012
R15391 Iout.n756 Iout.n33 0.451012
R15392 Iout.n858 Iout.n33 0.451012
R15393 Iout.n522 Iout.n145 0.451012
R15394 Iout.n523 Iout.n522 0.451012
R15395 Iout.n523 Iout.n132 0.451012
R15396 Iout.n545 Iout.n132 0.451012
R15397 Iout.n546 Iout.n545 0.451012
R15398 Iout.n546 Iout.n119 0.451012
R15399 Iout.n572 Iout.n119 0.451012
R15400 Iout.n580 Iout.n572 0.451012
R15401 Iout.n580 Iout.n579 0.451012
R15402 Iout.n579 Iout.n76 0.451012
R15403 Iout.n709 Iout.n76 0.451012
R15404 Iout.n709 Iout.n708 0.451012
R15405 Iout.n708 Iout.n25 0.451012
R15406 Iout.n914 Iout.n25 0.451012
R15407 Iout.n216 Iout.n179 0.451012
R15408 Iout.n286 Iout.n179 0.451012
R15409 Iout.n287 Iout.n286 0.451012
R15410 Iout.n287 Iout.n164 0.451012
R15411 Iout.n397 Iout.n164 0.451012
R15412 Iout.n398 Iout.n397 0.451012
R15413 Iout.n398 Iout.n92 0.451012
R15414 Iout.n633 Iout.n92 0.451012
R15415 Iout.n634 Iout.n633 0.451012
R15416 Iout.n634 Iout.n49 0.451012
R15417 Iout.n762 Iout.n49 0.451012
R15418 Iout.n763 Iout.n762 0.451012
R15419 Iout.n763 Iout.n34 0.451012
R15420 Iout.n851 Iout.n34 0.451012
R15421 Iout.n517 Iout.n516 0.451012
R15422 Iout.n517 Iout.n138 0.451012
R15423 Iout.n539 Iout.n138 0.451012
R15424 Iout.n540 Iout.n539 0.451012
R15425 Iout.n540 Iout.n125 0.451012
R15426 Iout.n562 Iout.n125 0.451012
R15427 Iout.n567 Iout.n562 0.451012
R15428 Iout.n567 Iout.n566 0.451012
R15429 Iout.n566 Iout.n79 0.451012
R15430 Iout.n698 Iout.n79 0.451012
R15431 Iout.n702 Iout.n698 0.451012
R15432 Iout.n703 Iout.n702 0.451012
R15433 Iout.n703 Iout.n24 0.451012
R15434 Iout.n921 Iout.n24 0.451012
R15435 Iout.n220 Iout.n176 0.451012
R15436 Iout.n293 Iout.n176 0.451012
R15437 Iout.n293 Iout.n292 0.451012
R15438 Iout.n292 Iout.n165 0.451012
R15439 Iout.n390 Iout.n165 0.451012
R15440 Iout.n390 Iout.n389 0.451012
R15441 Iout.n389 Iout.n89 0.451012
R15442 Iout.n640 Iout.n89 0.451012
R15443 Iout.n640 Iout.n639 0.451012
R15444 Iout.n639 Iout.n46 0.451012
R15445 Iout.n769 Iout.n46 0.451012
R15446 Iout.n769 Iout.n768 0.451012
R15447 Iout.n768 Iout.n35 0.451012
R15448 Iout.n844 Iout.n35 0.451012
R15449 Iout.n511 Iout.n2 0.451012
R15450 Iout.n1005 Iout.n2 0.451012
R15451 Iout.n1005 Iout.n1004 0.451012
R15452 Iout.n1004 Iout.n3 0.451012
R15453 Iout.n986 Iout.n3 0.451012
R15454 Iout.n986 Iout.n985 0.451012
R15455 Iout.n985 Iout.n8 0.451012
R15456 Iout.n967 Iout.n8 0.451012
R15457 Iout.n967 Iout.n966 0.451012
R15458 Iout.n966 Iout.n13 0.451012
R15459 Iout.n948 Iout.n13 0.451012
R15460 Iout.n948 Iout.n947 0.451012
R15461 Iout.n947 Iout.n18 0.451012
R15462 Iout.n929 Iout.n18 0.451012
R15463 Iout.n224 Iout.n170 0.451012
R15464 Iout.n298 Iout.n170 0.451012
R15465 Iout.n299 Iout.n298 0.451012
R15466 Iout.n299 Iout.n166 0.451012
R15467 Iout.n381 Iout.n166 0.451012
R15468 Iout.n382 Iout.n381 0.451012
R15469 Iout.n382 Iout.n83 0.451012
R15470 Iout.n645 Iout.n83 0.451012
R15471 Iout.n646 Iout.n645 0.451012
R15472 Iout.n646 Iout.n40 0.451012
R15473 Iout.n774 Iout.n40 0.451012
R15474 Iout.n775 Iout.n774 0.451012
R15475 Iout.n775 Iout.n36 0.451012
R15476 Iout.n837 Iout.n36 0.451012
R15477 Iout.n1018 Iout.n1017 0.451012
R15478 Iout.n1017 Iout.n0 0.451012
R15479 Iout.n999 Iout.n0 0.451012
R15480 Iout.n999 Iout.n998 0.451012
R15481 Iout.n998 Iout.n6 0.451012
R15482 Iout.n980 Iout.n6 0.451012
R15483 Iout.n980 Iout.n979 0.451012
R15484 Iout.n979 Iout.n11 0.451012
R15485 Iout.n961 Iout.n11 0.451012
R15486 Iout.n961 Iout.n960 0.451012
R15487 Iout.n960 Iout.n16 0.451012
R15488 Iout.n942 Iout.n16 0.451012
R15489 Iout.n942 Iout.n941 0.451012
R15490 Iout.n941 Iout.n21 0.451012
R15491 Iout.n230 Iout.n229 0.451012
R15492 Iout.n230 Iout.n167 0.451012
R15493 Iout.n304 Iout.n167 0.451012
R15494 Iout.n332 Iout.n304 0.451012
R15495 Iout.n374 Iout.n332 0.451012
R15496 Iout.n374 Iout.n373 0.451012
R15497 Iout.n373 Iout.n369 0.451012
R15498 Iout.n369 Iout.n80 0.451012
R15499 Iout.n651 Iout.n80 0.451012
R15500 Iout.n652 Iout.n651 0.451012
R15501 Iout.n652 Iout.n37 0.451012
R15502 Iout.n780 Iout.n37 0.451012
R15503 Iout.n826 Iout.n780 0.451012
R15504 Iout.n830 Iout.n826 0.451012
R15505 Iout.n231 Iout 0.2919
R15506 Iout.n303 Iout 0.2919
R15507 Iout Iout.n300 0.2919
R15508 Iout.n375 Iout 0.2919
R15509 Iout.n380 Iout 0.2919
R15510 Iout.n391 Iout 0.2919
R15511 Iout.n368 Iout 0.2919
R15512 Iout Iout.n365 0.2919
R15513 Iout Iout.n362 0.2919
R15514 Iout Iout.n359 0.2919
R15515 Iout.n650 Iout 0.2919
R15516 Iout Iout.n647 0.2919
R15517 Iout.n638 Iout 0.2919
R15518 Iout Iout.n635 0.2919
R15519 Iout.n626 Iout 0.2919
R15520 Iout.n41 Iout 0.2919
R15521 Iout.n773 Iout 0.2919
R15522 Iout Iout.n770 0.2919
R15523 Iout.n761 Iout 0.2919
R15524 Iout Iout.n758 0.2919
R15525 Iout.n749 Iout 0.2919
R15526 Iout.n825 Iout 0.2919
R15527 Iout Iout.n822 0.2919
R15528 Iout Iout.n819 0.2919
R15529 Iout Iout.n816 0.2919
R15530 Iout Iout.n813 0.2919
R15531 Iout Iout.n810 0.2919
R15532 Iout Iout.n807 0.2919
R15533 Iout.n829 Iout 0.2919
R15534 Iout.n838 Iout 0.2919
R15535 Iout.n843 Iout 0.2919
R15536 Iout.n852 Iout 0.2919
R15537 Iout.n857 Iout 0.2919
R15538 Iout.n866 Iout 0.2919
R15539 Iout.n871 Iout 0.2919
R15540 Iout.n880 Iout 0.2919
R15541 Iout Iout.n925 0.2919
R15542 Iout.n928 Iout 0.2919
R15543 Iout.n922 Iout 0.2919
R15544 Iout.n913 Iout 0.2919
R15545 Iout.n908 Iout 0.2919
R15546 Iout.n899 Iout 0.2919
R15547 Iout.n894 Iout 0.2919
R15548 Iout.n885 Iout 0.2919
R15549 Iout.n831 Iout 0.2919
R15550 Iout.n836 Iout 0.2919
R15551 Iout.n845 Iout 0.2919
R15552 Iout.n850 Iout 0.2919
R15553 Iout.n859 Iout 0.2919
R15554 Iout.n864 Iout 0.2919
R15555 Iout.n873 Iout 0.2919
R15556 Iout.n878 Iout 0.2919
R15557 Iout.n887 Iout 0.2919
R15558 Iout.n892 Iout 0.2919
R15559 Iout.n933 Iout 0.2919
R15560 Iout.n930 Iout 0.2919
R15561 Iout.n920 Iout 0.2919
R15562 Iout.n915 Iout 0.2919
R15563 Iout.n906 Iout 0.2919
R15564 Iout.n901 Iout 0.2919
R15565 Iout.n940 Iout 0.2919
R15566 Iout Iout.n783 0.2919
R15567 Iout Iout.n786 0.2919
R15568 Iout Iout.n789 0.2919
R15569 Iout Iout.n792 0.2919
R15570 Iout Iout.n795 0.2919
R15571 Iout Iout.n798 0.2919
R15572 Iout Iout.n801 0.2919
R15573 Iout Iout.n804 0.2919
R15574 Iout.n779 Iout 0.2919
R15575 Iout Iout.n776 0.2919
R15576 Iout.n767 Iout 0.2919
R15577 Iout Iout.n764 0.2919
R15578 Iout.n755 Iout 0.2919
R15579 Iout Iout.n752 0.2919
R15580 Iout.n743 Iout 0.2919
R15581 Iout Iout.n740 0.2919
R15582 Iout.n731 Iout 0.2919
R15583 Iout Iout.n728 0.2919
R15584 Iout.n719 Iout 0.2919
R15585 Iout Iout.n943 0.2919
R15586 Iout.n946 Iout 0.2919
R15587 Iout Iout.n704 0.2919
R15588 Iout.n707 Iout 0.2919
R15589 Iout Iout.n716 0.2919
R15590 Iout.n952 Iout 0.2919
R15591 Iout.n949 Iout 0.2919
R15592 Iout.n701 Iout 0.2919
R15593 Iout Iout.n710 0.2919
R15594 Iout.n713 Iout 0.2919
R15595 Iout Iout.n722 0.2919
R15596 Iout.n725 Iout 0.2919
R15597 Iout Iout.n734 0.2919
R15598 Iout.n737 Iout 0.2919
R15599 Iout Iout.n746 0.2919
R15600 Iout.n653 Iout 0.2919
R15601 Iout.n656 Iout 0.2919
R15602 Iout.n659 Iout 0.2919
R15603 Iout.n662 Iout 0.2919
R15604 Iout.n665 Iout 0.2919
R15605 Iout.n668 Iout 0.2919
R15606 Iout.n671 Iout 0.2919
R15607 Iout.n674 Iout 0.2919
R15608 Iout.n677 Iout 0.2919
R15609 Iout.n680 Iout 0.2919
R15610 Iout.n683 Iout 0.2919
R15611 Iout.n686 Iout 0.2919
R15612 Iout.n959 Iout 0.2919
R15613 Iout Iout.n694 0.2919
R15614 Iout.n697 Iout 0.2919
R15615 Iout.n689 Iout 0.2919
R15616 Iout Iout.n962 0.2919
R15617 Iout.n965 Iout 0.2919
R15618 Iout Iout.n575 0.2919
R15619 Iout.n578 Iout 0.2919
R15620 Iout Iout.n587 0.2919
R15621 Iout.n590 Iout 0.2919
R15622 Iout Iout.n599 0.2919
R15623 Iout.n602 Iout 0.2919
R15624 Iout Iout.n611 0.2919
R15625 Iout.n614 Iout 0.2919
R15626 Iout Iout.n623 0.2919
R15627 Iout.n84 Iout 0.2919
R15628 Iout.n644 Iout 0.2919
R15629 Iout Iout.n641 0.2919
R15630 Iout.n632 Iout 0.2919
R15631 Iout Iout.n629 0.2919
R15632 Iout.n620 Iout 0.2919
R15633 Iout Iout.n617 0.2919
R15634 Iout.n608 Iout 0.2919
R15635 Iout Iout.n605 0.2919
R15636 Iout.n596 Iout 0.2919
R15637 Iout Iout.n593 0.2919
R15638 Iout.n584 Iout 0.2919
R15639 Iout Iout.n581 0.2919
R15640 Iout.n971 Iout 0.2919
R15641 Iout.n968 Iout 0.2919
R15642 Iout.n565 Iout 0.2919
R15643 Iout.n978 Iout 0.2919
R15644 Iout Iout.n122 0.2919
R15645 Iout Iout.n568 0.2919
R15646 Iout.n571 Iout 0.2919
R15647 Iout Iout.n335 0.2919
R15648 Iout Iout.n338 0.2919
R15649 Iout Iout.n341 0.2919
R15650 Iout Iout.n344 0.2919
R15651 Iout Iout.n347 0.2919
R15652 Iout Iout.n350 0.2919
R15653 Iout Iout.n353 0.2919
R15654 Iout Iout.n356 0.2919
R15655 Iout.n372 Iout 0.2919
R15656 Iout.n383 Iout 0.2919
R15657 Iout.n388 Iout 0.2919
R15658 Iout.n399 Iout 0.2919
R15659 Iout.n404 Iout 0.2919
R15660 Iout.n415 Iout 0.2919
R15661 Iout.n420 Iout 0.2919
R15662 Iout.n431 Iout 0.2919
R15663 Iout.n443 Iout 0.2919
R15664 Iout Iout.n440 0.2919
R15665 Iout Iout.n437 0.2919
R15666 Iout.n553 Iout 0.2919
R15667 Iout.n556 Iout 0.2919
R15668 Iout.n561 Iout 0.2919
R15669 Iout Iout.n981 0.2919
R15670 Iout.n984 Iout 0.2919
R15671 Iout.n990 Iout 0.2919
R15672 Iout.n987 Iout 0.2919
R15673 Iout Iout.n129 0.2919
R15674 Iout Iout.n547 0.2919
R15675 Iout.n550 Iout 0.2919
R15676 Iout Iout.n451 0.2919
R15677 Iout.n454 Iout 0.2919
R15678 Iout.n446 Iout 0.2919
R15679 Iout.n428 Iout 0.2919
R15680 Iout.n423 Iout 0.2919
R15681 Iout.n412 Iout 0.2919
R15682 Iout.n407 Iout 0.2919
R15683 Iout.n396 Iout 0.2919
R15684 Iout.n331 Iout 0.2919
R15685 Iout Iout.n328 0.2919
R15686 Iout Iout.n325 0.2919
R15687 Iout Iout.n322 0.2919
R15688 Iout Iout.n319 0.2919
R15689 Iout Iout.n316 0.2919
R15690 Iout Iout.n313 0.2919
R15691 Iout Iout.n310 0.2919
R15692 Iout Iout.n307 0.2919
R15693 Iout.n457 Iout 0.2919
R15694 Iout.n465 Iout 0.2919
R15695 Iout Iout.n462 0.2919
R15696 Iout.n544 Iout 0.2919
R15697 Iout Iout.n541 0.2919
R15698 Iout Iout.n135 0.2919
R15699 Iout.n997 Iout 0.2919
R15700 Iout Iout.n1000 0.2919
R15701 Iout.n1003 Iout 0.2919
R15702 Iout.n538 Iout 0.2919
R15703 Iout.n533 Iout 0.2919
R15704 Iout.n530 Iout 0.2919
R15705 Iout Iout.n468 0.2919
R15706 Iout Iout.n471 0.2919
R15707 Iout.n474 Iout 0.2919
R15708 Iout Iout.n264 0.2919
R15709 Iout.n267 Iout 0.2919
R15710 Iout Iout.n276 0.2919
R15711 Iout.n279 Iout 0.2919
R15712 Iout Iout.n288 0.2919
R15713 Iout.n291 Iout 0.2919
R15714 Iout.n171 Iout 0.2919
R15715 Iout.n297 Iout 0.2919
R15716 Iout Iout.n294 0.2919
R15717 Iout.n285 Iout 0.2919
R15718 Iout Iout.n282 0.2919
R15719 Iout.n273 Iout 0.2919
R15720 Iout Iout.n270 0.2919
R15721 Iout.n261 Iout 0.2919
R15722 Iout.n477 Iout 0.2919
R15723 Iout.n485 Iout 0.2919
R15724 Iout Iout.n482 0.2919
R15725 Iout.n527 Iout 0.2919
R15726 Iout Iout.n524 0.2919
R15727 Iout Iout.n142 0.2919
R15728 Iout.n1006 Iout 0.2919
R15729 Iout.n1009 Iout 0.2919
R15730 Iout.n1016 Iout 0.2919
R15731 Iout Iout.n148 0.2919
R15732 Iout Iout.n518 0.2919
R15733 Iout.n521 Iout 0.2919
R15734 Iout Iout.n493 0.2919
R15735 Iout.n496 Iout 0.2919
R15736 Iout.n488 Iout 0.2919
R15737 Iout Iout.n254 0.2919
R15738 Iout.n257 Iout 0.2919
R15739 Iout.n249 Iout 0.2919
R15740 Iout.n246 Iout 0.2919
R15741 Iout.n243 Iout 0.2919
R15742 Iout.n240 Iout 0.2919
R15743 Iout.n237 Iout 0.2919
R15744 Iout.n234 Iout 0.2919
R15745 Iout.n228 Iout 0.2919
R15746 Iout Iout.n225 0.2919
R15747 Iout Iout.n221 0.2919
R15748 Iout Iout.n217 0.2919
R15749 Iout Iout.n213 0.2919
R15750 Iout Iout.n209 0.2919
R15751 Iout Iout.n205 0.2919
R15752 Iout Iout.n201 0.2919
R15753 Iout Iout.n198 0.2919
R15754 Iout Iout.n194 0.2919
R15755 Iout.n499 Iout 0.2919
R15756 Iout.n503 Iout 0.2919
R15757 Iout.n506 Iout 0.2919
R15758 Iout.n515 Iout 0.2919
R15759 Iout Iout.n512 0.2919
R15760 Iout.n1019 Iout 0.2919
R15761 Iout.n1013 Iout.n1012 0.092855
R15762 Iout.n1012 Iout.n1 0.092855
R15763 Iout.n994 Iout.n1 0.092855
R15764 Iout.n994 Iout.n993 0.092855
R15765 Iout.n993 Iout.n7 0.092855
R15766 Iout.n975 Iout.n7 0.092855
R15767 Iout.n975 Iout.n974 0.092855
R15768 Iout.n974 Iout.n12 0.092855
R15769 Iout.n956 Iout.n12 0.092855
R15770 Iout.n956 Iout.n955 0.092855
R15771 Iout.n955 Iout.n17 0.092855
R15772 Iout.n937 Iout.n17 0.092855
R15773 Iout.n937 Iout.n936 0.092855
R15774 Iout.n197 Iout 0.0818902
R15775 Iout.n191 Iout 0.0818902
R15776 Iout.n152 Iout 0.0818902
R15777 Iout.n204 Iout 0.0818902
R15778 Iout.n498 Iout 0.0818902
R15779 Iout.n208 Iout 0.0818902
R15780 Iout.n502 Iout 0.0818902
R15781 Iout.n212 Iout 0.0818902
R15782 Iout.n145 Iout 0.0818902
R15783 Iout.n216 Iout 0.0818902
R15784 Iout.n516 Iout 0.0818902
R15785 Iout.n220 Iout 0.0818902
R15786 Iout.n511 Iout 0.0818902
R15787 Iout.n224 Iout 0.0818902
R15788 Iout.n1018 Iout 0.0818902
R15789 Iout.n229 Iout 0.0818902
R15790 Iout.n1013 Iout 0.072645
R15791 Iout.n302 Iout 0.0532071
R15792 Iout Iout.n377 0.0532071
R15793 Iout.n379 Iout 0.0532071
R15794 Iout.n367 Iout 0.0532071
R15795 Iout.n364 Iout 0.0532071
R15796 Iout.n361 Iout 0.0532071
R15797 Iout.n649 Iout 0.0532071
R15798 Iout Iout.n82 0.0532071
R15799 Iout.n637 Iout 0.0532071
R15800 Iout Iout.n91 0.0532071
R15801 Iout Iout.n43 0.0532071
R15802 Iout.n772 Iout 0.0532071
R15803 Iout Iout.n45 0.0532071
R15804 Iout.n760 Iout 0.0532071
R15805 Iout Iout.n51 0.0532071
R15806 Iout.n824 Iout 0.0532071
R15807 Iout.n821 Iout 0.0532071
R15808 Iout.n818 Iout 0.0532071
R15809 Iout.n815 Iout 0.0532071
R15810 Iout.n812 Iout 0.0532071
R15811 Iout.n809 Iout 0.0532071
R15812 Iout.n828 Iout 0.0532071
R15813 Iout Iout.n840 0.0532071
R15814 Iout.n842 Iout 0.0532071
R15815 Iout Iout.n854 0.0532071
R15816 Iout.n856 Iout 0.0532071
R15817 Iout Iout.n868 0.0532071
R15818 Iout.n870 Iout 0.0532071
R15819 Iout.n927 Iout 0.0532071
R15820 Iout Iout.n924 0.0532071
R15821 Iout.n912 Iout 0.0532071
R15822 Iout Iout.n910 0.0532071
R15823 Iout.n898 Iout 0.0532071
R15824 Iout Iout.n896 0.0532071
R15825 Iout.n884 Iout 0.0532071
R15826 Iout Iout.n882 0.0532071
R15827 Iout Iout.n833 0.0532071
R15828 Iout.n835 Iout 0.0532071
R15829 Iout Iout.n847 0.0532071
R15830 Iout.n849 Iout 0.0532071
R15831 Iout Iout.n861 0.0532071
R15832 Iout.n863 Iout 0.0532071
R15833 Iout Iout.n875 0.0532071
R15834 Iout.n877 Iout 0.0532071
R15835 Iout Iout.n889 0.0532071
R15836 Iout Iout.n932 0.0532071
R15837 Iout.n919 Iout 0.0532071
R15838 Iout Iout.n917 0.0532071
R15839 Iout.n905 Iout 0.0532071
R15840 Iout Iout.n903 0.0532071
R15841 Iout.n891 Iout 0.0532071
R15842 Iout.n782 Iout 0.0532071
R15843 Iout.n785 Iout 0.0532071
R15844 Iout.n788 Iout 0.0532071
R15845 Iout.n791 Iout 0.0532071
R15846 Iout.n794 Iout 0.0532071
R15847 Iout.n797 Iout 0.0532071
R15848 Iout.n800 Iout 0.0532071
R15849 Iout.n803 Iout 0.0532071
R15850 Iout.n806 Iout 0.0532071
R15851 Iout.n778 Iout 0.0532071
R15852 Iout Iout.n39 0.0532071
R15853 Iout.n766 Iout 0.0532071
R15854 Iout Iout.n48 0.0532071
R15855 Iout.n754 Iout 0.0532071
R15856 Iout Iout.n54 0.0532071
R15857 Iout.n742 Iout 0.0532071
R15858 Iout Iout.n60 0.0532071
R15859 Iout.n730 Iout 0.0532071
R15860 Iout Iout.n66 0.0532071
R15861 Iout.n945 Iout 0.0532071
R15862 Iout.n78 Iout 0.0532071
R15863 Iout.n706 Iout 0.0532071
R15864 Iout Iout.n72 0.0532071
R15865 Iout.n718 Iout 0.0532071
R15866 Iout Iout.n951 0.0532071
R15867 Iout.n700 Iout 0.0532071
R15868 Iout Iout.n75 0.0532071
R15869 Iout.n712 Iout 0.0532071
R15870 Iout Iout.n69 0.0532071
R15871 Iout.n724 Iout 0.0532071
R15872 Iout Iout.n63 0.0532071
R15873 Iout.n736 Iout 0.0532071
R15874 Iout Iout.n57 0.0532071
R15875 Iout.n748 Iout 0.0532071
R15876 Iout Iout.n655 0.0532071
R15877 Iout Iout.n658 0.0532071
R15878 Iout Iout.n661 0.0532071
R15879 Iout Iout.n664 0.0532071
R15880 Iout Iout.n667 0.0532071
R15881 Iout Iout.n670 0.0532071
R15882 Iout Iout.n673 0.0532071
R15883 Iout Iout.n676 0.0532071
R15884 Iout Iout.n679 0.0532071
R15885 Iout Iout.n682 0.0532071
R15886 Iout Iout.n685 0.0532071
R15887 Iout.n693 Iout 0.0532071
R15888 Iout.n696 Iout 0.0532071
R15889 Iout Iout.n691 0.0532071
R15890 Iout Iout.n688 0.0532071
R15891 Iout.n964 Iout 0.0532071
R15892 Iout.n574 Iout 0.0532071
R15893 Iout.n577 Iout 0.0532071
R15894 Iout Iout.n115 0.0532071
R15895 Iout.n589 Iout 0.0532071
R15896 Iout Iout.n109 0.0532071
R15897 Iout.n601 Iout 0.0532071
R15898 Iout Iout.n103 0.0532071
R15899 Iout.n613 Iout 0.0532071
R15900 Iout Iout.n97 0.0532071
R15901 Iout.n625 Iout 0.0532071
R15902 Iout Iout.n86 0.0532071
R15903 Iout.n643 Iout 0.0532071
R15904 Iout Iout.n88 0.0532071
R15905 Iout.n631 Iout 0.0532071
R15906 Iout Iout.n94 0.0532071
R15907 Iout.n619 Iout 0.0532071
R15908 Iout Iout.n100 0.0532071
R15909 Iout.n607 Iout 0.0532071
R15910 Iout Iout.n106 0.0532071
R15911 Iout.n595 Iout 0.0532071
R15912 Iout Iout.n112 0.0532071
R15913 Iout.n583 Iout 0.0532071
R15914 Iout Iout.n970 0.0532071
R15915 Iout.n564 Iout 0.0532071
R15916 Iout Iout.n118 0.0532071
R15917 Iout.n121 Iout 0.0532071
R15918 Iout.n124 Iout 0.0532071
R15919 Iout.n570 Iout 0.0532071
R15920 Iout.n334 Iout 0.0532071
R15921 Iout.n337 Iout 0.0532071
R15922 Iout.n340 Iout 0.0532071
R15923 Iout.n343 Iout 0.0532071
R15924 Iout.n346 Iout 0.0532071
R15925 Iout.n349 Iout 0.0532071
R15926 Iout.n352 Iout 0.0532071
R15927 Iout.n355 Iout 0.0532071
R15928 Iout.n358 Iout 0.0532071
R15929 Iout.n371 Iout 0.0532071
R15930 Iout Iout.n385 0.0532071
R15931 Iout.n387 Iout 0.0532071
R15932 Iout Iout.n401 0.0532071
R15933 Iout.n403 Iout 0.0532071
R15934 Iout Iout.n417 0.0532071
R15935 Iout.n419 Iout 0.0532071
R15936 Iout Iout.n433 0.0532071
R15937 Iout.n442 Iout 0.0532071
R15938 Iout.n439 Iout 0.0532071
R15939 Iout.n435 Iout 0.0532071
R15940 Iout Iout.n555 0.0532071
R15941 Iout Iout.n558 0.0532071
R15942 Iout.n983 Iout 0.0532071
R15943 Iout.n560 Iout 0.0532071
R15944 Iout Iout.n989 0.0532071
R15945 Iout.n128 Iout 0.0532071
R15946 Iout.n131 Iout 0.0532071
R15947 Iout.n549 Iout 0.0532071
R15948 Iout.n450 Iout 0.0532071
R15949 Iout.n453 Iout 0.0532071
R15950 Iout Iout.n448 0.0532071
R15951 Iout.n427 Iout 0.0532071
R15952 Iout Iout.n425 0.0532071
R15953 Iout.n411 Iout 0.0532071
R15954 Iout Iout.n409 0.0532071
R15955 Iout.n395 Iout 0.0532071
R15956 Iout Iout.n393 0.0532071
R15957 Iout.n330 Iout 0.0532071
R15958 Iout.n327 Iout 0.0532071
R15959 Iout.n324 Iout 0.0532071
R15960 Iout.n321 Iout 0.0532071
R15961 Iout.n318 Iout 0.0532071
R15962 Iout.n315 Iout 0.0532071
R15963 Iout.n312 Iout 0.0532071
R15964 Iout.n309 Iout 0.0532071
R15965 Iout.n306 Iout 0.0532071
R15966 Iout Iout.n459 0.0532071
R15967 Iout.n464 Iout 0.0532071
R15968 Iout.n461 Iout 0.0532071
R15969 Iout.n543 Iout 0.0532071
R15970 Iout.n137 Iout 0.0532071
R15971 Iout.n134 Iout 0.0532071
R15972 Iout.n1002 Iout 0.0532071
R15973 Iout.n537 Iout 0.0532071
R15974 Iout Iout.n535 0.0532071
R15975 Iout Iout.n532 0.0532071
R15976 Iout.n157 Iout 0.0532071
R15977 Iout.n470 Iout 0.0532071
R15978 Iout.n473 Iout 0.0532071
R15979 Iout.n190 Iout 0.0532071
R15980 Iout.n266 Iout 0.0532071
R15981 Iout Iout.n184 0.0532071
R15982 Iout.n278 Iout 0.0532071
R15983 Iout Iout.n178 0.0532071
R15984 Iout.n290 Iout 0.0532071
R15985 Iout Iout.n169 0.0532071
R15986 Iout Iout.n173 0.0532071
R15987 Iout.n296 Iout 0.0532071
R15988 Iout Iout.n175 0.0532071
R15989 Iout.n284 Iout 0.0532071
R15990 Iout Iout.n181 0.0532071
R15991 Iout.n272 Iout 0.0532071
R15992 Iout Iout.n187 0.0532071
R15993 Iout.n260 Iout 0.0532071
R15994 Iout Iout.n479 0.0532071
R15995 Iout.n484 Iout 0.0532071
R15996 Iout.n481 Iout 0.0532071
R15997 Iout.n526 Iout 0.0532071
R15998 Iout.n144 Iout 0.0532071
R15999 Iout.n141 Iout 0.0532071
R16000 Iout Iout.n1008 0.0532071
R16001 Iout.n147 Iout 0.0532071
R16002 Iout.n150 Iout 0.0532071
R16003 Iout.n520 Iout 0.0532071
R16004 Iout.n492 Iout 0.0532071
R16005 Iout.n495 Iout 0.0532071
R16006 Iout Iout.n490 0.0532071
R16007 Iout.n253 Iout 0.0532071
R16008 Iout.n256 Iout 0.0532071
R16009 Iout Iout.n251 0.0532071
R16010 Iout Iout.n248 0.0532071
R16011 Iout Iout.n245 0.0532071
R16012 Iout Iout.n242 0.0532071
R16013 Iout Iout.n239 0.0532071
R16014 Iout Iout.n236 0.0532071
R16015 Iout Iout.n233 0.0532071
R16016 Iout.n227 Iout 0.0532071
R16017 Iout.n223 Iout 0.0532071
R16018 Iout.n219 Iout 0.0532071
R16019 Iout.n215 Iout 0.0532071
R16020 Iout.n211 Iout 0.0532071
R16021 Iout.n207 Iout 0.0532071
R16022 Iout.n203 Iout 0.0532071
R16023 Iout.n200 Iout 0.0532071
R16024 Iout.n196 Iout 0.0532071
R16025 Iout.n193 Iout 0.0532071
R16026 Iout Iout.n501 0.0532071
R16027 Iout Iout.n505 0.0532071
R16028 Iout Iout.n508 0.0532071
R16029 Iout.n514 Iout 0.0532071
R16030 Iout.n510 Iout 0.0532071
R16031 Iout.n1020 Iout 0.03925
R16032 Iout.n509 Iout 0.03925
R16033 Iout.n513 Iout 0.03925
R16034 Iout.n507 Iout 0.03925
R16035 Iout.n504 Iout 0.03925
R16036 Iout.n500 Iout 0.03925
R16037 Iout.n192 Iout 0.03925
R16038 Iout.n195 Iout 0.03925
R16039 Iout.n199 Iout 0.03925
R16040 Iout.n202 Iout 0.03925
R16041 Iout.n206 Iout 0.03925
R16042 Iout.n210 Iout 0.03925
R16043 Iout.n214 Iout 0.03925
R16044 Iout.n218 Iout 0.03925
R16045 Iout.n222 Iout 0.03925
R16046 Iout.n226 Iout 0.03925
R16047 Iout.n232 Iout 0.03925
R16048 Iout.n235 Iout 0.03925
R16049 Iout.n238 Iout 0.03925
R16050 Iout.n241 Iout 0.03925
R16051 Iout.n244 Iout 0.03925
R16052 Iout.n247 Iout 0.03925
R16053 Iout.n250 Iout 0.03925
R16054 Iout.n255 Iout 0.03925
R16055 Iout.n252 Iout 0.03925
R16056 Iout.n489 Iout 0.03925
R16057 Iout.n494 Iout 0.03925
R16058 Iout.n491 Iout 0.03925
R16059 Iout.n519 Iout 0.03925
R16060 Iout.n149 Iout 0.03925
R16061 Iout.n146 Iout 0.03925
R16062 Iout.n1010 Iout 0.03925
R16063 Iout.n1007 Iout 0.03925
R16064 Iout.n140 Iout 0.03925
R16065 Iout.n143 Iout 0.03925
R16066 Iout.n525 Iout 0.03925
R16067 Iout.n480 Iout 0.03925
R16068 Iout.n483 Iout 0.03925
R16069 Iout.n478 Iout 0.03925
R16070 Iout.n259 Iout 0.03925
R16071 Iout.n186 Iout 0.03925
R16072 Iout.n271 Iout 0.03925
R16073 Iout.n180 Iout 0.03925
R16074 Iout.n283 Iout 0.03925
R16075 Iout.n174 Iout 0.03925
R16076 Iout.n168 Iout 0.03925
R16077 Iout.n301 Iout 0.03925
R16078 Iout.n289 Iout 0.03925
R16079 Iout.n177 Iout 0.03925
R16080 Iout.n277 Iout 0.03925
R16081 Iout.n183 Iout 0.03925
R16082 Iout.n265 Iout 0.03925
R16083 Iout.n189 Iout 0.03925
R16084 Iout.n472 Iout 0.03925
R16085 Iout.n469 Iout 0.03925
R16086 Iout.n156 Iout 0.03925
R16087 Iout.n531 Iout 0.03925
R16088 Iout.n534 Iout 0.03925
R16089 Iout.n536 Iout 0.03925
R16090 Iout.n133 Iout 0.03925
R16091 Iout.n136 Iout 0.03925
R16092 Iout.n542 Iout 0.03925
R16093 Iout.n460 Iout 0.03925
R16094 Iout.n463 Iout 0.03925
R16095 Iout.n458 Iout 0.03925
R16096 Iout.n305 Iout 0.03925
R16097 Iout.n308 Iout 0.03925
R16098 Iout.n311 Iout 0.03925
R16099 Iout.n314 Iout 0.03925
R16100 Iout.n317 Iout 0.03925
R16101 Iout.n320 Iout 0.03925
R16102 Iout.n392 Iout 0.03925
R16103 Iout.n378 Iout 0.03925
R16104 Iout.n376 Iout 0.03925
R16105 Iout.n394 Iout 0.03925
R16106 Iout.n408 Iout 0.03925
R16107 Iout.n410 Iout 0.03925
R16108 Iout.n424 Iout 0.03925
R16109 Iout.n426 Iout 0.03925
R16110 Iout.n447 Iout 0.03925
R16111 Iout.n452 Iout 0.03925
R16112 Iout.n449 Iout 0.03925
R16113 Iout.n548 Iout 0.03925
R16114 Iout.n130 Iout 0.03925
R16115 Iout.n559 Iout 0.03925
R16116 Iout.n557 Iout 0.03925
R16117 Iout.n554 Iout 0.03925
R16118 Iout.n434 Iout 0.03925
R16119 Iout.n438 Iout 0.03925
R16120 Iout.n441 Iout 0.03925
R16121 Iout.n432 Iout 0.03925
R16122 Iout.n418 Iout 0.03925
R16123 Iout.n416 Iout 0.03925
R16124 Iout.n402 Iout 0.03925
R16125 Iout.n357 Iout 0.03925
R16126 Iout.n360 Iout 0.03925
R16127 Iout.n363 Iout 0.03925
R16128 Iout.n366 Iout 0.03925
R16129 Iout.n354 Iout 0.03925
R16130 Iout.n351 Iout 0.03925
R16131 Iout.n348 Iout 0.03925
R16132 Iout.n345 Iout 0.03925
R16133 Iout.n342 Iout 0.03925
R16134 Iout.n339 Iout 0.03925
R16135 Iout.n336 Iout 0.03925
R16136 Iout.n333 Iout 0.03925
R16137 Iout.n117 Iout 0.03925
R16138 Iout.n582 Iout 0.03925
R16139 Iout.n111 Iout 0.03925
R16140 Iout.n594 Iout 0.03925
R16141 Iout.n105 Iout 0.03925
R16142 Iout.n606 Iout 0.03925
R16143 Iout.n99 Iout 0.03925
R16144 Iout.n618 Iout 0.03925
R16145 Iout.n624 Iout 0.03925
R16146 Iout.n90 Iout 0.03925
R16147 Iout.n636 Iout 0.03925
R16148 Iout.n81 Iout 0.03925
R16149 Iout.n648 Iout 0.03925
R16150 Iout.n96 Iout 0.03925
R16151 Iout.n612 Iout 0.03925
R16152 Iout.n102 Iout 0.03925
R16153 Iout.n600 Iout 0.03925
R16154 Iout.n108 Iout 0.03925
R16155 Iout.n588 Iout 0.03925
R16156 Iout.n687 Iout 0.03925
R16157 Iout.n684 Iout 0.03925
R16158 Iout.n681 Iout 0.03925
R16159 Iout.n678 Iout 0.03925
R16160 Iout.n675 Iout 0.03925
R16161 Iout.n672 Iout 0.03925
R16162 Iout.n747 Iout 0.03925
R16163 Iout.n50 Iout 0.03925
R16164 Iout.n759 Iout 0.03925
R16165 Iout.n44 Iout 0.03925
R16166 Iout.n771 Iout 0.03925
R16167 Iout.n42 Iout 0.03925
R16168 Iout.n56 Iout 0.03925
R16169 Iout.n735 Iout 0.03925
R16170 Iout.n62 Iout 0.03925
R16171 Iout.n723 Iout 0.03925
R16172 Iout.n717 Iout 0.03925
R16173 Iout.n65 Iout 0.03925
R16174 Iout.n729 Iout 0.03925
R16175 Iout.n59 Iout 0.03925
R16176 Iout.n805 Iout 0.03925
R16177 Iout.n808 Iout 0.03925
R16178 Iout.n811 Iout 0.03925
R16179 Iout.n814 Iout 0.03925
R16180 Iout.n817 Iout 0.03925
R16181 Iout.n820 Iout 0.03925
R16182 Iout.n823 Iout 0.03925
R16183 Iout.n802 Iout 0.03925
R16184 Iout.n799 Iout 0.03925
R16185 Iout.n890 Iout 0.03925
R16186 Iout.n888 Iout 0.03925
R16187 Iout.n881 Iout 0.03925
R16188 Iout.n869 Iout 0.03925
R16189 Iout.n867 Iout 0.03925
R16190 Iout.n855 Iout 0.03925
R16191 Iout.n853 Iout 0.03925
R16192 Iout.n841 Iout 0.03925
R16193 Iout.n839 Iout 0.03925
R16194 Iout.n827 Iout 0.03925
R16195 Iout.n883 Iout 0.03925
R16196 Iout.n895 Iout 0.03925
R16197 Iout.n897 Iout 0.03925
R16198 Iout.n909 Iout 0.03925
R16199 Iout.n911 Iout 0.03925
R16200 Iout.n923 Iout 0.03925
R16201 Iout.n926 Iout 0.03925
R16202 Iout.n22 Iout 0.03925
R16203 Iout.n876 Iout 0.03925
R16204 Iout.n874 Iout 0.03925
R16205 Iout.n862 Iout 0.03925
R16206 Iout.n860 Iout 0.03925
R16207 Iout.n848 Iout 0.03925
R16208 Iout.n846 Iout 0.03925
R16209 Iout.n834 Iout 0.03925
R16210 Iout.n832 Iout 0.03925
R16211 Iout.n902 Iout 0.03925
R16212 Iout.n904 Iout 0.03925
R16213 Iout.n916 Iout 0.03925
R16214 Iout.n918 Iout 0.03925
R16215 Iout.n931 Iout 0.03925
R16216 Iout.n934 Iout 0.03925
R16217 Iout.n796 Iout 0.03925
R16218 Iout.n793 Iout 0.03925
R16219 Iout.n790 Iout 0.03925
R16220 Iout.n787 Iout 0.03925
R16221 Iout.n784 Iout 0.03925
R16222 Iout.n781 Iout 0.03925
R16223 Iout.n938 Iout 0.03925
R16224 Iout.n741 Iout 0.03925
R16225 Iout.n53 Iout 0.03925
R16226 Iout.n753 Iout 0.03925
R16227 Iout.n47 Iout 0.03925
R16228 Iout.n765 Iout 0.03925
R16229 Iout.n38 Iout 0.03925
R16230 Iout.n777 Iout 0.03925
R16231 Iout.n71 Iout 0.03925
R16232 Iout.n705 Iout 0.03925
R16233 Iout.n77 Iout 0.03925
R16234 Iout.n944 Iout 0.03925
R16235 Iout.n19 Iout 0.03925
R16236 Iout.n68 Iout 0.03925
R16237 Iout.n711 Iout 0.03925
R16238 Iout.n74 Iout 0.03925
R16239 Iout.n699 Iout 0.03925
R16240 Iout.n950 Iout 0.03925
R16241 Iout.n953 Iout 0.03925
R16242 Iout.n669 Iout 0.03925
R16243 Iout.n666 Iout 0.03925
R16244 Iout.n663 Iout 0.03925
R16245 Iout.n660 Iout 0.03925
R16246 Iout.n657 Iout 0.03925
R16247 Iout.n654 Iout 0.03925
R16248 Iout.n690 Iout 0.03925
R16249 Iout.n695 Iout 0.03925
R16250 Iout.n692 Iout 0.03925
R16251 Iout.n957 Iout 0.03925
R16252 Iout.n114 Iout 0.03925
R16253 Iout.n576 Iout 0.03925
R16254 Iout.n573 Iout 0.03925
R16255 Iout.n963 Iout 0.03925
R16256 Iout.n14 Iout 0.03925
R16257 Iout.n93 Iout 0.03925
R16258 Iout.n630 Iout 0.03925
R16259 Iout.n87 Iout 0.03925
R16260 Iout.n642 Iout 0.03925
R16261 Iout.n85 Iout 0.03925
R16262 Iout.n563 Iout 0.03925
R16263 Iout.n969 Iout 0.03925
R16264 Iout.n972 Iout 0.03925
R16265 Iout.n569 Iout 0.03925
R16266 Iout.n123 Iout 0.03925
R16267 Iout.n120 Iout 0.03925
R16268 Iout.n976 Iout 0.03925
R16269 Iout.n400 Iout 0.03925
R16270 Iout.n386 Iout 0.03925
R16271 Iout.n384 Iout 0.03925
R16272 Iout.n370 Iout 0.03925
R16273 Iout.n982 Iout 0.03925
R16274 Iout.n9 Iout 0.03925
R16275 Iout.n127 Iout 0.03925
R16276 Iout.n988 Iout 0.03925
R16277 Iout.n991 Iout 0.03925
R16278 Iout.n323 Iout 0.03925
R16279 Iout.n326 Iout 0.03925
R16280 Iout.n329 Iout 0.03925
R16281 Iout.n995 Iout 0.03925
R16282 Iout.n1001 Iout 0.03925
R16283 Iout.n4 Iout 0.03925
R16284 Iout.n295 Iout 0.03925
R16285 Iout.n172 Iout 0.03925
R16286 Iout.n1014 Iout 0.03925
R16287 Iout.n1022 Iout 0.02071
R16288 Iout Iout.n1022 0.00379
R16289 Iout.n303 Iout.n302 0.00105952
R16290 Iout.n377 Iout.n375 0.00105952
R16291 Iout.n380 Iout.n379 0.00105952
R16292 Iout.n368 Iout.n367 0.00105952
R16293 Iout.n365 Iout.n364 0.00105952
R16294 Iout.n362 Iout.n361 0.00105952
R16295 Iout.n650 Iout.n649 0.00105952
R16296 Iout.n647 Iout.n82 0.00105952
R16297 Iout.n638 Iout.n637 0.00105952
R16298 Iout.n635 Iout.n91 0.00105952
R16299 Iout.n43 Iout.n41 0.00105952
R16300 Iout.n773 Iout.n772 0.00105952
R16301 Iout.n770 Iout.n45 0.00105952
R16302 Iout.n761 Iout.n760 0.00105952
R16303 Iout.n758 Iout.n51 0.00105952
R16304 Iout.n825 Iout.n824 0.00105952
R16305 Iout.n822 Iout.n821 0.00105952
R16306 Iout.n819 Iout.n818 0.00105952
R16307 Iout.n816 Iout.n815 0.00105952
R16308 Iout.n813 Iout.n812 0.00105952
R16309 Iout.n810 Iout.n809 0.00105952
R16310 Iout.n829 Iout.n828 0.00105952
R16311 Iout.n840 Iout.n838 0.00105952
R16312 Iout.n843 Iout.n842 0.00105952
R16313 Iout.n854 Iout.n852 0.00105952
R16314 Iout.n857 Iout.n856 0.00105952
R16315 Iout.n868 Iout.n866 0.00105952
R16316 Iout.n871 Iout.n870 0.00105952
R16317 Iout.n925 Iout.n23 0.00105952
R16318 Iout.n928 Iout.n927 0.00105952
R16319 Iout.n924 Iout.n922 0.00105952
R16320 Iout.n913 Iout.n912 0.00105952
R16321 Iout.n910 Iout.n908 0.00105952
R16322 Iout.n899 Iout.n898 0.00105952
R16323 Iout.n896 Iout.n894 0.00105952
R16324 Iout.n885 Iout.n884 0.00105952
R16325 Iout.n882 Iout.n880 0.00105952
R16326 Iout.n833 Iout.n831 0.00105952
R16327 Iout.n836 Iout.n835 0.00105952
R16328 Iout.n847 Iout.n845 0.00105952
R16329 Iout.n850 Iout.n849 0.00105952
R16330 Iout.n861 Iout.n859 0.00105952
R16331 Iout.n864 Iout.n863 0.00105952
R16332 Iout.n875 Iout.n873 0.00105952
R16333 Iout.n878 Iout.n877 0.00105952
R16334 Iout.n889 Iout.n887 0.00105952
R16335 Iout.n935 Iout.n933 0.00105952
R16336 Iout.n932 Iout.n930 0.00105952
R16337 Iout.n920 Iout.n919 0.00105952
R16338 Iout.n917 Iout.n915 0.00105952
R16339 Iout.n906 Iout.n905 0.00105952
R16340 Iout.n903 Iout.n901 0.00105952
R16341 Iout.n892 Iout.n891 0.00105952
R16342 Iout.n940 Iout.n939 0.00105952
R16343 Iout.n783 Iout.n782 0.00105952
R16344 Iout.n786 Iout.n785 0.00105952
R16345 Iout.n789 Iout.n788 0.00105952
R16346 Iout.n792 Iout.n791 0.00105952
R16347 Iout.n795 Iout.n794 0.00105952
R16348 Iout.n798 Iout.n797 0.00105952
R16349 Iout.n801 Iout.n800 0.00105952
R16350 Iout.n804 Iout.n803 0.00105952
R16351 Iout.n807 Iout.n806 0.00105952
R16352 Iout.n779 Iout.n778 0.00105952
R16353 Iout.n776 Iout.n39 0.00105952
R16354 Iout.n767 Iout.n766 0.00105952
R16355 Iout.n764 Iout.n48 0.00105952
R16356 Iout.n755 Iout.n754 0.00105952
R16357 Iout.n752 Iout.n54 0.00105952
R16358 Iout.n743 Iout.n742 0.00105952
R16359 Iout.n740 Iout.n60 0.00105952
R16360 Iout.n731 Iout.n730 0.00105952
R16361 Iout.n728 Iout.n66 0.00105952
R16362 Iout.n943 Iout.n20 0.00105952
R16363 Iout.n946 Iout.n945 0.00105952
R16364 Iout.n704 Iout.n78 0.00105952
R16365 Iout.n707 Iout.n706 0.00105952
R16366 Iout.n716 Iout.n72 0.00105952
R16367 Iout.n719 Iout.n718 0.00105952
R16368 Iout.n954 Iout.n952 0.00105952
R16369 Iout.n951 Iout.n949 0.00105952
R16370 Iout.n701 Iout.n700 0.00105952
R16371 Iout.n710 Iout.n75 0.00105952
R16372 Iout.n713 Iout.n712 0.00105952
R16373 Iout.n722 Iout.n69 0.00105952
R16374 Iout.n725 Iout.n724 0.00105952
R16375 Iout.n734 Iout.n63 0.00105952
R16376 Iout.n737 Iout.n736 0.00105952
R16377 Iout.n746 Iout.n57 0.00105952
R16378 Iout.n749 Iout.n748 0.00105952
R16379 Iout.n655 Iout.n653 0.00105952
R16380 Iout.n658 Iout.n656 0.00105952
R16381 Iout.n661 Iout.n659 0.00105952
R16382 Iout.n664 Iout.n662 0.00105952
R16383 Iout.n667 Iout.n665 0.00105952
R16384 Iout.n670 Iout.n668 0.00105952
R16385 Iout.n673 Iout.n671 0.00105952
R16386 Iout.n676 Iout.n674 0.00105952
R16387 Iout.n679 Iout.n677 0.00105952
R16388 Iout.n682 Iout.n680 0.00105952
R16389 Iout.n685 Iout.n683 0.00105952
R16390 Iout.n959 Iout.n958 0.00105952
R16391 Iout.n694 Iout.n693 0.00105952
R16392 Iout.n697 Iout.n696 0.00105952
R16393 Iout.n691 Iout.n689 0.00105952
R16394 Iout.n688 Iout.n686 0.00105952
R16395 Iout.n962 Iout.n15 0.00105952
R16396 Iout.n965 Iout.n964 0.00105952
R16397 Iout.n575 Iout.n574 0.00105952
R16398 Iout.n578 Iout.n577 0.00105952
R16399 Iout.n587 Iout.n115 0.00105952
R16400 Iout.n590 Iout.n589 0.00105952
R16401 Iout.n599 Iout.n109 0.00105952
R16402 Iout.n602 Iout.n601 0.00105952
R16403 Iout.n611 Iout.n103 0.00105952
R16404 Iout.n614 Iout.n613 0.00105952
R16405 Iout.n623 Iout.n97 0.00105952
R16406 Iout.n626 Iout.n625 0.00105952
R16407 Iout.n86 Iout.n84 0.00105952
R16408 Iout.n644 Iout.n643 0.00105952
R16409 Iout.n641 Iout.n88 0.00105952
R16410 Iout.n632 Iout.n631 0.00105952
R16411 Iout.n629 Iout.n94 0.00105952
R16412 Iout.n620 Iout.n619 0.00105952
R16413 Iout.n617 Iout.n100 0.00105952
R16414 Iout.n608 Iout.n607 0.00105952
R16415 Iout.n605 Iout.n106 0.00105952
R16416 Iout.n596 Iout.n595 0.00105952
R16417 Iout.n593 Iout.n112 0.00105952
R16418 Iout.n584 Iout.n583 0.00105952
R16419 Iout.n973 Iout.n971 0.00105952
R16420 Iout.n970 Iout.n968 0.00105952
R16421 Iout.n565 Iout.n564 0.00105952
R16422 Iout.n581 Iout.n118 0.00105952
R16423 Iout.n978 Iout.n977 0.00105952
R16424 Iout.n122 Iout.n121 0.00105952
R16425 Iout.n568 Iout.n124 0.00105952
R16426 Iout.n571 Iout.n570 0.00105952
R16427 Iout.n335 Iout.n334 0.00105952
R16428 Iout.n338 Iout.n337 0.00105952
R16429 Iout.n341 Iout.n340 0.00105952
R16430 Iout.n344 Iout.n343 0.00105952
R16431 Iout.n347 Iout.n346 0.00105952
R16432 Iout.n350 Iout.n349 0.00105952
R16433 Iout.n353 Iout.n352 0.00105952
R16434 Iout.n356 Iout.n355 0.00105952
R16435 Iout.n359 Iout.n358 0.00105952
R16436 Iout.n372 Iout.n371 0.00105952
R16437 Iout.n385 Iout.n383 0.00105952
R16438 Iout.n388 Iout.n387 0.00105952
R16439 Iout.n401 Iout.n399 0.00105952
R16440 Iout.n404 Iout.n403 0.00105952
R16441 Iout.n417 Iout.n415 0.00105952
R16442 Iout.n420 Iout.n419 0.00105952
R16443 Iout.n433 Iout.n431 0.00105952
R16444 Iout.n443 Iout.n442 0.00105952
R16445 Iout.n440 Iout.n439 0.00105952
R16446 Iout.n437 Iout.n435 0.00105952
R16447 Iout.n555 Iout.n553 0.00105952
R16448 Iout.n558 Iout.n556 0.00105952
R16449 Iout.n981 Iout.n10 0.00105952
R16450 Iout.n984 Iout.n983 0.00105952
R16451 Iout.n561 Iout.n560 0.00105952
R16452 Iout.n992 Iout.n990 0.00105952
R16453 Iout.n989 Iout.n987 0.00105952
R16454 Iout.n129 Iout.n128 0.00105952
R16455 Iout.n547 Iout.n131 0.00105952
R16456 Iout.n550 Iout.n549 0.00105952
R16457 Iout.n451 Iout.n450 0.00105952
R16458 Iout.n454 Iout.n453 0.00105952
R16459 Iout.n448 Iout.n446 0.00105952
R16460 Iout.n428 Iout.n427 0.00105952
R16461 Iout.n425 Iout.n423 0.00105952
R16462 Iout.n412 Iout.n411 0.00105952
R16463 Iout.n409 Iout.n407 0.00105952
R16464 Iout.n396 Iout.n395 0.00105952
R16465 Iout.n393 Iout.n391 0.00105952
R16466 Iout.n331 Iout.n330 0.00105952
R16467 Iout.n328 Iout.n327 0.00105952
R16468 Iout.n325 Iout.n324 0.00105952
R16469 Iout.n322 Iout.n321 0.00105952
R16470 Iout.n319 Iout.n318 0.00105952
R16471 Iout.n316 Iout.n315 0.00105952
R16472 Iout.n313 Iout.n312 0.00105952
R16473 Iout.n310 Iout.n309 0.00105952
R16474 Iout.n307 Iout.n306 0.00105952
R16475 Iout.n459 Iout.n457 0.00105952
R16476 Iout.n465 Iout.n464 0.00105952
R16477 Iout.n462 Iout.n461 0.00105952
R16478 Iout.n544 Iout.n543 0.00105952
R16479 Iout.n541 Iout.n137 0.00105952
R16480 Iout.n997 Iout.n996 0.00105952
R16481 Iout.n135 Iout.n134 0.00105952
R16482 Iout.n1000 Iout.n5 0.00105952
R16483 Iout.n1003 Iout.n1002 0.00105952
R16484 Iout.n538 Iout.n537 0.00105952
R16485 Iout.n535 Iout.n533 0.00105952
R16486 Iout.n532 Iout.n530 0.00105952
R16487 Iout.n468 Iout.n157 0.00105952
R16488 Iout.n471 Iout.n470 0.00105952
R16489 Iout.n474 Iout.n473 0.00105952
R16490 Iout.n264 Iout.n190 0.00105952
R16491 Iout.n267 Iout.n266 0.00105952
R16492 Iout.n276 Iout.n184 0.00105952
R16493 Iout.n279 Iout.n278 0.00105952
R16494 Iout.n288 Iout.n178 0.00105952
R16495 Iout.n291 Iout.n290 0.00105952
R16496 Iout.n300 Iout.n169 0.00105952
R16497 Iout.n173 Iout.n171 0.00105952
R16498 Iout.n297 Iout.n296 0.00105952
R16499 Iout.n294 Iout.n175 0.00105952
R16500 Iout.n285 Iout.n284 0.00105952
R16501 Iout.n282 Iout.n181 0.00105952
R16502 Iout.n273 Iout.n272 0.00105952
R16503 Iout.n270 Iout.n187 0.00105952
R16504 Iout.n261 Iout.n260 0.00105952
R16505 Iout.n479 Iout.n477 0.00105952
R16506 Iout.n485 Iout.n484 0.00105952
R16507 Iout.n482 Iout.n481 0.00105952
R16508 Iout.n527 Iout.n526 0.00105952
R16509 Iout.n524 Iout.n144 0.00105952
R16510 Iout.n142 Iout.n141 0.00105952
R16511 Iout.n1008 Iout.n1006 0.00105952
R16512 Iout.n1011 Iout.n1009 0.00105952
R16513 Iout.n1016 Iout.n1015 0.00105952
R16514 Iout.n148 Iout.n147 0.00105952
R16515 Iout.n518 Iout.n150 0.00105952
R16516 Iout.n521 Iout.n520 0.00105952
R16517 Iout.n493 Iout.n492 0.00105952
R16518 Iout.n496 Iout.n495 0.00105952
R16519 Iout.n490 Iout.n488 0.00105952
R16520 Iout.n254 Iout.n253 0.00105952
R16521 Iout.n257 Iout.n256 0.00105952
R16522 Iout.n251 Iout.n249 0.00105952
R16523 Iout.n248 Iout.n246 0.00105952
R16524 Iout.n245 Iout.n243 0.00105952
R16525 Iout.n242 Iout.n240 0.00105952
R16526 Iout.n239 Iout.n237 0.00105952
R16527 Iout.n236 Iout.n234 0.00105952
R16528 Iout.n233 Iout.n231 0.00105952
R16529 Iout.n228 Iout.n227 0.00105952
R16530 Iout.n225 Iout.n223 0.00105952
R16531 Iout.n221 Iout.n219 0.00105952
R16532 Iout.n217 Iout.n215 0.00105952
R16533 Iout.n213 Iout.n211 0.00105952
R16534 Iout.n209 Iout.n207 0.00105952
R16535 Iout.n205 Iout.n203 0.00105952
R16536 Iout.n201 Iout.n200 0.00105952
R16537 Iout.n198 Iout.n196 0.00105952
R16538 Iout.n194 Iout.n193 0.00105952
R16539 Iout.n501 Iout.n499 0.00105952
R16540 Iout.n505 Iout.n503 0.00105952
R16541 Iout.n508 Iout.n506 0.00105952
R16542 Iout.n515 Iout.n514 0.00105952
R16543 Iout.n512 Iout.n510 0.00105952
R16544 Iout.n1021 Iout.n1019 0.00105952
R16545 XThC.Tn[10].n71 XThC.Tn[10].n70 256.104
R16546 XThC.Tn[10].n75 XThC.Tn[10].n73 243.68
R16547 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16548 XThC.Tn[10].n75 XThC.Tn[10].n74 205.28
R16549 XThC.Tn[10].n71 XThC.Tn[10].n69 202.095
R16550 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16551 XThC.Tn[10].n65 XThC.Tn[10].n63 161.365
R16552 XThC.Tn[10].n61 XThC.Tn[10].n59 161.365
R16553 XThC.Tn[10].n57 XThC.Tn[10].n55 161.365
R16554 XThC.Tn[10].n53 XThC.Tn[10].n51 161.365
R16555 XThC.Tn[10].n49 XThC.Tn[10].n47 161.365
R16556 XThC.Tn[10].n45 XThC.Tn[10].n43 161.365
R16557 XThC.Tn[10].n41 XThC.Tn[10].n39 161.365
R16558 XThC.Tn[10].n37 XThC.Tn[10].n35 161.365
R16559 XThC.Tn[10].n33 XThC.Tn[10].n31 161.365
R16560 XThC.Tn[10].n29 XThC.Tn[10].n27 161.365
R16561 XThC.Tn[10].n25 XThC.Tn[10].n23 161.365
R16562 XThC.Tn[10].n21 XThC.Tn[10].n19 161.365
R16563 XThC.Tn[10].n17 XThC.Tn[10].n15 161.365
R16564 XThC.Tn[10].n13 XThC.Tn[10].n11 161.365
R16565 XThC.Tn[10].n9 XThC.Tn[10].n7 161.365
R16566 XThC.Tn[10].n6 XThC.Tn[10].n4 161.365
R16567 XThC.Tn[10].n63 XThC.Tn[10].t42 161.202
R16568 XThC.Tn[10].n59 XThC.Tn[10].t32 161.202
R16569 XThC.Tn[10].n55 XThC.Tn[10].t19 161.202
R16570 XThC.Tn[10].n51 XThC.Tn[10].t16 161.202
R16571 XThC.Tn[10].n47 XThC.Tn[10].t40 161.202
R16572 XThC.Tn[10].n43 XThC.Tn[10].t27 161.202
R16573 XThC.Tn[10].n39 XThC.Tn[10].t26 161.202
R16574 XThC.Tn[10].n35 XThC.Tn[10].t39 161.202
R16575 XThC.Tn[10].n31 XThC.Tn[10].t37 161.202
R16576 XThC.Tn[10].n27 XThC.Tn[10].t28 161.202
R16577 XThC.Tn[10].n23 XThC.Tn[10].t15 161.202
R16578 XThC.Tn[10].n19 XThC.Tn[10].t14 161.202
R16579 XThC.Tn[10].n15 XThC.Tn[10].t25 161.202
R16580 XThC.Tn[10].n11 XThC.Tn[10].t23 161.202
R16581 XThC.Tn[10].n7 XThC.Tn[10].t21 161.202
R16582 XThC.Tn[10].n4 XThC.Tn[10].t36 161.202
R16583 XThC.Tn[10].n63 XThC.Tn[10].t13 145.137
R16584 XThC.Tn[10].n59 XThC.Tn[10].t35 145.137
R16585 XThC.Tn[10].n55 XThC.Tn[10].t22 145.137
R16586 XThC.Tn[10].n51 XThC.Tn[10].t20 145.137
R16587 XThC.Tn[10].n47 XThC.Tn[10].t12 145.137
R16588 XThC.Tn[10].n43 XThC.Tn[10].t33 145.137
R16589 XThC.Tn[10].n39 XThC.Tn[10].t31 145.137
R16590 XThC.Tn[10].n35 XThC.Tn[10].t43 145.137
R16591 XThC.Tn[10].n31 XThC.Tn[10].t41 145.137
R16592 XThC.Tn[10].n27 XThC.Tn[10].t34 145.137
R16593 XThC.Tn[10].n23 XThC.Tn[10].t18 145.137
R16594 XThC.Tn[10].n19 XThC.Tn[10].t17 145.137
R16595 XThC.Tn[10].n15 XThC.Tn[10].t30 145.137
R16596 XThC.Tn[10].n11 XThC.Tn[10].t29 145.137
R16597 XThC.Tn[10].n7 XThC.Tn[10].t24 145.137
R16598 XThC.Tn[10].n4 XThC.Tn[10].t38 145.137
R16599 XThC.Tn[10].n73 XThC.Tn[10].t9 26.5955
R16600 XThC.Tn[10].n73 XThC.Tn[10].t10 26.5955
R16601 XThC.Tn[10].n69 XThC.Tn[10].t3 26.5955
R16602 XThC.Tn[10].n69 XThC.Tn[10].t8 26.5955
R16603 XThC.Tn[10].n70 XThC.Tn[10].t5 26.5955
R16604 XThC.Tn[10].n70 XThC.Tn[10].t11 26.5955
R16605 XThC.Tn[10].n74 XThC.Tn[10].t0 26.5955
R16606 XThC.Tn[10].n74 XThC.Tn[10].t1 26.5955
R16607 XThC.Tn[10].n1 XThC.Tn[10].t2 24.9236
R16608 XThC.Tn[10].n1 XThC.Tn[10].t7 24.9236
R16609 XThC.Tn[10].n0 XThC.Tn[10].t6 24.9236
R16610 XThC.Tn[10].n0 XThC.Tn[10].t4 24.9236
R16611 XThC.Tn[10] XThC.Tn[10].n75 22.9652
R16612 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16613 XThC.Tn[10].n72 XThC.Tn[10].n71 13.9299
R16614 XThC.Tn[10] XThC.Tn[10].n72 13.9299
R16615 XThC.Tn[10] XThC.Tn[10].n6 8.0245
R16616 XThC.Tn[10].n66 XThC.Tn[10].n65 7.9105
R16617 XThC.Tn[10].n62 XThC.Tn[10].n61 7.9105
R16618 XThC.Tn[10].n58 XThC.Tn[10].n57 7.9105
R16619 XThC.Tn[10].n54 XThC.Tn[10].n53 7.9105
R16620 XThC.Tn[10].n50 XThC.Tn[10].n49 7.9105
R16621 XThC.Tn[10].n46 XThC.Tn[10].n45 7.9105
R16622 XThC.Tn[10].n42 XThC.Tn[10].n41 7.9105
R16623 XThC.Tn[10].n38 XThC.Tn[10].n37 7.9105
R16624 XThC.Tn[10].n34 XThC.Tn[10].n33 7.9105
R16625 XThC.Tn[10].n30 XThC.Tn[10].n29 7.9105
R16626 XThC.Tn[10].n26 XThC.Tn[10].n25 7.9105
R16627 XThC.Tn[10].n22 XThC.Tn[10].n21 7.9105
R16628 XThC.Tn[10].n18 XThC.Tn[10].n17 7.9105
R16629 XThC.Tn[10].n14 XThC.Tn[10].n13 7.9105
R16630 XThC.Tn[10].n10 XThC.Tn[10].n9 7.9105
R16631 XThC.Tn[10].n68 XThC.Tn[10].n67 7.40985
R16632 XThC.Tn[10].n67 XThC.Tn[10] 4.38575
R16633 XThC.Tn[10].n72 XThC.Tn[10].n68 2.99115
R16634 XThC.Tn[10].n72 XThC.Tn[10] 2.87153
R16635 XThC.Tn[10].n3 XThC.Tn[10] 2.688
R16636 XThC.Tn[10].n68 XThC.Tn[10] 2.2734
R16637 XThC.Tn[10].n67 XThC.Tn[10].n3 0.244922
R16638 XThC.Tn[10].n10 XThC.Tn[10] 0.235138
R16639 XThC.Tn[10].n14 XThC.Tn[10] 0.235138
R16640 XThC.Tn[10].n18 XThC.Tn[10] 0.235138
R16641 XThC.Tn[10].n22 XThC.Tn[10] 0.235138
R16642 XThC.Tn[10].n26 XThC.Tn[10] 0.235138
R16643 XThC.Tn[10].n30 XThC.Tn[10] 0.235138
R16644 XThC.Tn[10].n34 XThC.Tn[10] 0.235138
R16645 XThC.Tn[10].n38 XThC.Tn[10] 0.235138
R16646 XThC.Tn[10].n42 XThC.Tn[10] 0.235138
R16647 XThC.Tn[10].n46 XThC.Tn[10] 0.235138
R16648 XThC.Tn[10].n50 XThC.Tn[10] 0.235138
R16649 XThC.Tn[10].n54 XThC.Tn[10] 0.235138
R16650 XThC.Tn[10].n58 XThC.Tn[10] 0.235138
R16651 XThC.Tn[10].n62 XThC.Tn[10] 0.235138
R16652 XThC.Tn[10].n66 XThC.Tn[10] 0.235138
R16653 XThC.Tn[10].n3 XThC.Tn[10] 0.141947
R16654 XThC.Tn[10] XThC.Tn[10].n10 0.114505
R16655 XThC.Tn[10] XThC.Tn[10].n14 0.114505
R16656 XThC.Tn[10] XThC.Tn[10].n18 0.114505
R16657 XThC.Tn[10] XThC.Tn[10].n22 0.114505
R16658 XThC.Tn[10] XThC.Tn[10].n26 0.114505
R16659 XThC.Tn[10] XThC.Tn[10].n30 0.114505
R16660 XThC.Tn[10] XThC.Tn[10].n34 0.114505
R16661 XThC.Tn[10] XThC.Tn[10].n38 0.114505
R16662 XThC.Tn[10] XThC.Tn[10].n42 0.114505
R16663 XThC.Tn[10] XThC.Tn[10].n46 0.114505
R16664 XThC.Tn[10] XThC.Tn[10].n50 0.114505
R16665 XThC.Tn[10] XThC.Tn[10].n54 0.114505
R16666 XThC.Tn[10] XThC.Tn[10].n58 0.114505
R16667 XThC.Tn[10] XThC.Tn[10].n62 0.114505
R16668 XThC.Tn[10] XThC.Tn[10].n66 0.114505
R16669 XThC.Tn[10].n65 XThC.Tn[10].n64 0.0599512
R16670 XThC.Tn[10].n61 XThC.Tn[10].n60 0.0599512
R16671 XThC.Tn[10].n57 XThC.Tn[10].n56 0.0599512
R16672 XThC.Tn[10].n53 XThC.Tn[10].n52 0.0599512
R16673 XThC.Tn[10].n49 XThC.Tn[10].n48 0.0599512
R16674 XThC.Tn[10].n45 XThC.Tn[10].n44 0.0599512
R16675 XThC.Tn[10].n41 XThC.Tn[10].n40 0.0599512
R16676 XThC.Tn[10].n37 XThC.Tn[10].n36 0.0599512
R16677 XThC.Tn[10].n33 XThC.Tn[10].n32 0.0599512
R16678 XThC.Tn[10].n29 XThC.Tn[10].n28 0.0599512
R16679 XThC.Tn[10].n25 XThC.Tn[10].n24 0.0599512
R16680 XThC.Tn[10].n21 XThC.Tn[10].n20 0.0599512
R16681 XThC.Tn[10].n17 XThC.Tn[10].n16 0.0599512
R16682 XThC.Tn[10].n13 XThC.Tn[10].n12 0.0599512
R16683 XThC.Tn[10].n9 XThC.Tn[10].n8 0.0599512
R16684 XThC.Tn[10].n6 XThC.Tn[10].n5 0.0599512
R16685 XThC.Tn[10].n64 XThC.Tn[10] 0.0469286
R16686 XThC.Tn[10].n60 XThC.Tn[10] 0.0469286
R16687 XThC.Tn[10].n56 XThC.Tn[10] 0.0469286
R16688 XThC.Tn[10].n52 XThC.Tn[10] 0.0469286
R16689 XThC.Tn[10].n48 XThC.Tn[10] 0.0469286
R16690 XThC.Tn[10].n44 XThC.Tn[10] 0.0469286
R16691 XThC.Tn[10].n40 XThC.Tn[10] 0.0469286
R16692 XThC.Tn[10].n36 XThC.Tn[10] 0.0469286
R16693 XThC.Tn[10].n32 XThC.Tn[10] 0.0469286
R16694 XThC.Tn[10].n28 XThC.Tn[10] 0.0469286
R16695 XThC.Tn[10].n24 XThC.Tn[10] 0.0469286
R16696 XThC.Tn[10].n20 XThC.Tn[10] 0.0469286
R16697 XThC.Tn[10].n16 XThC.Tn[10] 0.0469286
R16698 XThC.Tn[10].n12 XThC.Tn[10] 0.0469286
R16699 XThC.Tn[10].n8 XThC.Tn[10] 0.0469286
R16700 XThC.Tn[10].n5 XThC.Tn[10] 0.0469286
R16701 XThC.Tn[10].n64 XThC.Tn[10] 0.0401341
R16702 XThC.Tn[10].n60 XThC.Tn[10] 0.0401341
R16703 XThC.Tn[10].n56 XThC.Tn[10] 0.0401341
R16704 XThC.Tn[10].n52 XThC.Tn[10] 0.0401341
R16705 XThC.Tn[10].n48 XThC.Tn[10] 0.0401341
R16706 XThC.Tn[10].n44 XThC.Tn[10] 0.0401341
R16707 XThC.Tn[10].n40 XThC.Tn[10] 0.0401341
R16708 XThC.Tn[10].n36 XThC.Tn[10] 0.0401341
R16709 XThC.Tn[10].n32 XThC.Tn[10] 0.0401341
R16710 XThC.Tn[10].n28 XThC.Tn[10] 0.0401341
R16711 XThC.Tn[10].n24 XThC.Tn[10] 0.0401341
R16712 XThC.Tn[10].n20 XThC.Tn[10] 0.0401341
R16713 XThC.Tn[10].n16 XThC.Tn[10] 0.0401341
R16714 XThC.Tn[10].n12 XThC.Tn[10] 0.0401341
R16715 XThC.Tn[10].n8 XThC.Tn[10] 0.0401341
R16716 XThC.Tn[10].n5 XThC.Tn[10] 0.0401341
R16717 XThR.TBN.n1 XThR.TBN.t60 212.081
R16718 XThR.TBN.n8 XThR.TBN.t12 212.081
R16719 XThR.TBN.n2 XThR.TBN.t81 212.081
R16720 XThR.TBN.n3 XThR.TBN.t121 212.081
R16721 XThR.TBN.n12 XThR.TBN.t115 212.081
R16722 XThR.TBN.n19 XThR.TBN.t65 212.081
R16723 XThR.TBN.n13 XThR.TBN.t21 212.081
R16724 XThR.TBN.n14 XThR.TBN.t57 212.081
R16725 XThR.TBN.n24 XThR.TBN.t27 212.081
R16726 XThR.TBN.n31 XThR.TBN.t96 212.081
R16727 XThR.TBN.n25 XThR.TBN.t46 212.081
R16728 XThR.TBN.n26 XThR.TBN.t89 212.081
R16729 XThR.TBN.n36 XThR.TBN.t80 212.081
R16730 XThR.TBN.n43 XThR.TBN.t31 212.081
R16731 XThR.TBN.n37 XThR.TBN.t102 212.081
R16732 XThR.TBN.n38 XThR.TBN.t25 212.081
R16733 XThR.TBN.n48 XThR.TBN.t85 212.081
R16734 XThR.TBN.n55 XThR.TBN.t33 212.081
R16735 XThR.TBN.n49 XThR.TBN.t105 212.081
R16736 XThR.TBN.n50 XThR.TBN.t26 212.081
R16737 XThR.TBN.n60 XThR.TBN.t54 212.081
R16738 XThR.TBN.n67 XThR.TBN.t5 212.081
R16739 XThR.TBN.n61 XThR.TBN.t73 212.081
R16740 XThR.TBN.n62 XThR.TBN.t114 212.081
R16741 XThR.TBN.n72 XThR.TBN.t49 212.081
R16742 XThR.TBN.n79 XThR.TBN.t119 212.081
R16743 XThR.TBN.n73 XThR.TBN.t69 212.081
R16744 XThR.TBN.n74 XThR.TBN.t108 212.081
R16745 XThR.TBN.n163 XThR.TBN.t41 212.081
R16746 XThR.TBN.n154 XThR.TBN.t113 212.081
R16747 XThR.TBN.n158 XThR.TBN.t34 212.081
R16748 XThR.TBN.n155 XThR.TBN.t72 212.081
R16749 XThR.TBN.n151 XThR.TBN.t19 212.081
R16750 XThR.TBN.n142 XThR.TBN.t86 212.081
R16751 XThR.TBN.n146 XThR.TBN.t6 212.081
R16752 XThR.TBN.n143 XThR.TBN.t43 212.081
R16753 XThR.TBN.n139 XThR.TBN.t45 212.081
R16754 XThR.TBN.n130 XThR.TBN.t117 212.081
R16755 XThR.TBN.n134 XThR.TBN.t36 212.081
R16756 XThR.TBN.n131 XThR.TBN.t75 212.081
R16757 XThR.TBN.n127 XThR.TBN.t100 212.081
R16758 XThR.TBN.n118 XThR.TBN.t50 212.081
R16759 XThR.TBN.n122 XThR.TBN.t92 212.081
R16760 XThR.TBN.n119 XThR.TBN.t13 212.081
R16761 XThR.TBN.n115 XThR.TBN.t15 212.081
R16762 XThR.TBN.n106 XThR.TBN.t83 212.081
R16763 XThR.TBN.n110 XThR.TBN.t123 212.081
R16764 XThR.TBN.n107 XThR.TBN.t39 212.081
R16765 XThR.TBN.n103 XThR.TBN.t66 212.081
R16766 XThR.TBN.n94 XThR.TBN.t23 212.081
R16767 XThR.TBN.n98 XThR.TBN.t59 212.081
R16768 XThR.TBN.n95 XThR.TBN.t97 212.081
R16769 XThR.TBN.n92 XThR.TBN.t99 212.081
R16770 XThR.TBN.n83 XThR.TBN.t87 212.081
R16771 XThR.TBN.n87 XThR.TBN.t77 212.081
R16772 XThR.TBN.n84 XThR.TBN.t68 212.081
R16773 XThR.TBN.n167 XThR.TBN.t63 212.081
R16774 XThR.TBN.n169 XThR.TBN.t106 212.081
R16775 XThR.TBN.n174 XThR.TBN.t56 212.081
R16776 XThR.TBN.n170 XThR.TBN.t7 212.081
R16777 XThR.TBN XThR.TBN.n180 203.923
R16778 XThR.TBN.n171 XThR.TBN.n170 188.516
R16779 XThR.TBN.n164 XThR.TBN.n163 180.482
R16780 XThR.TBN.n152 XThR.TBN.n151 180.482
R16781 XThR.TBN.n140 XThR.TBN.n139 180.482
R16782 XThR.TBN.n128 XThR.TBN.n127 180.482
R16783 XThR.TBN.n116 XThR.TBN.n115 180.482
R16784 XThR.TBN.n104 XThR.TBN.n103 180.482
R16785 XThR.TBN.n93 XThR.TBN.n92 180.482
R16786 XThR.TBN.n5 XThR.TBN.n4 173.761
R16787 XThR.TBN.n16 XThR.TBN.n15 173.761
R16788 XThR.TBN.n28 XThR.TBN.n27 173.761
R16789 XThR.TBN.n40 XThR.TBN.n39 173.761
R16790 XThR.TBN.n52 XThR.TBN.n51 173.761
R16791 XThR.TBN.n64 XThR.TBN.n63 173.761
R16792 XThR.TBN.n76 XThR.TBN.n75 173.761
R16793 XThR.TBN.n168 XThR.TBN 154.304
R16794 XThR.TBN.n10 XThR.TBN.n9 152
R16795 XThR.TBN.n7 XThR.TBN.n0 152
R16796 XThR.TBN.n6 XThR.TBN.n5 152
R16797 XThR.TBN.n17 XThR.TBN.n16 152
R16798 XThR.TBN.n18 XThR.TBN.n11 152
R16799 XThR.TBN.n21 XThR.TBN.n20 152
R16800 XThR.TBN.n29 XThR.TBN.n28 152
R16801 XThR.TBN.n30 XThR.TBN.n23 152
R16802 XThR.TBN.n33 XThR.TBN.n32 152
R16803 XThR.TBN.n41 XThR.TBN.n40 152
R16804 XThR.TBN.n42 XThR.TBN.n35 152
R16805 XThR.TBN.n45 XThR.TBN.n44 152
R16806 XThR.TBN.n53 XThR.TBN.n52 152
R16807 XThR.TBN.n54 XThR.TBN.n47 152
R16808 XThR.TBN.n57 XThR.TBN.n56 152
R16809 XThR.TBN.n65 XThR.TBN.n64 152
R16810 XThR.TBN.n66 XThR.TBN.n59 152
R16811 XThR.TBN.n69 XThR.TBN.n68 152
R16812 XThR.TBN.n77 XThR.TBN.n76 152
R16813 XThR.TBN.n78 XThR.TBN.n71 152
R16814 XThR.TBN.n81 XThR.TBN.n80 152
R16815 XThR.TBN.n157 XThR.TBN.n156 152
R16816 XThR.TBN.n160 XThR.TBN.n159 152
R16817 XThR.TBN.n162 XThR.TBN.n161 152
R16818 XThR.TBN.n145 XThR.TBN.n144 152
R16819 XThR.TBN.n148 XThR.TBN.n147 152
R16820 XThR.TBN.n150 XThR.TBN.n149 152
R16821 XThR.TBN.n133 XThR.TBN.n132 152
R16822 XThR.TBN.n136 XThR.TBN.n135 152
R16823 XThR.TBN.n138 XThR.TBN.n137 152
R16824 XThR.TBN.n121 XThR.TBN.n120 152
R16825 XThR.TBN.n124 XThR.TBN.n123 152
R16826 XThR.TBN.n126 XThR.TBN.n125 152
R16827 XThR.TBN.n109 XThR.TBN.n108 152
R16828 XThR.TBN.n112 XThR.TBN.n111 152
R16829 XThR.TBN.n114 XThR.TBN.n113 152
R16830 XThR.TBN.n97 XThR.TBN.n96 152
R16831 XThR.TBN.n100 XThR.TBN.n99 152
R16832 XThR.TBN.n102 XThR.TBN.n101 152
R16833 XThR.TBN.n86 XThR.TBN.n85 152
R16834 XThR.TBN.n89 XThR.TBN.n88 152
R16835 XThR.TBN.n91 XThR.TBN.n90 152
R16836 XThR.TBN.n173 XThR.TBN.n172 152
R16837 XThR.TBN.n176 XThR.TBN.n175 152
R16838 XThR.TBN.n1 XThR.TBN.t95 139.78
R16839 XThR.TBN.n8 XThR.TBN.t44 139.78
R16840 XThR.TBN.n2 XThR.TBN.t116 139.78
R16841 XThR.TBN.n3 XThR.TBN.t35 139.78
R16842 XThR.TBN.n12 XThR.TBN.t42 139.78
R16843 XThR.TBN.n19 XThR.TBN.t112 139.78
R16844 XThR.TBN.n13 XThR.TBN.t64 139.78
R16845 XThR.TBN.n14 XThR.TBN.t107 139.78
R16846 XThR.TBN.n24 XThR.TBN.t61 139.78
R16847 XThR.TBN.n31 XThR.TBN.t14 139.78
R16848 XThR.TBN.n25 XThR.TBN.t82 139.78
R16849 XThR.TBN.n26 XThR.TBN.t122 139.78
R16850 XThR.TBN.n36 XThR.TBN.t11 139.78
R16851 XThR.TBN.n43 XThR.TBN.t79 139.78
R16852 XThR.TBN.n37 XThR.TBN.t32 139.78
R16853 XThR.TBN.n38 XThR.TBN.t71 139.78
R16854 XThR.TBN.n48 XThR.TBN.t29 139.78
R16855 XThR.TBN.n55 XThR.TBN.t98 139.78
R16856 XThR.TBN.n49 XThR.TBN.t47 139.78
R16857 XThR.TBN.n50 XThR.TBN.t90 139.78
R16858 XThR.TBN.n60 XThR.TBN.t8 139.78
R16859 XThR.TBN.n67 XThR.TBN.t74 139.78
R16860 XThR.TBN.n61 XThR.TBN.t28 139.78
R16861 XThR.TBN.n62 XThR.TBN.t67 139.78
R16862 XThR.TBN.n72 XThR.TBN.t111 139.78
R16863 XThR.TBN.n79 XThR.TBN.t62 139.78
R16864 XThR.TBN.n73 XThR.TBN.t18 139.78
R16865 XThR.TBN.n74 XThR.TBN.t53 139.78
R16866 XThR.TBN.n163 XThR.TBN.t101 139.78
R16867 XThR.TBN.n154 XThR.TBN.t52 139.78
R16868 XThR.TBN.n158 XThR.TBN.t93 139.78
R16869 XThR.TBN.n155 XThR.TBN.t16 139.78
R16870 XThR.TBN.n151 XThR.TBN.t88 139.78
R16871 XThR.TBN.n142 XThR.TBN.t37 139.78
R16872 XThR.TBN.n146 XThR.TBN.t76 139.78
R16873 XThR.TBN.n143 XThR.TBN.t118 139.78
R16874 XThR.TBN.n139 XThR.TBN.t104 139.78
R16875 XThR.TBN.n130 XThR.TBN.t55 139.78
R16876 XThR.TBN.n134 XThR.TBN.t94 139.78
R16877 XThR.TBN.n131 XThR.TBN.t17 139.78
R16878 XThR.TBN.n127 XThR.TBN.t51 139.78
R16879 XThR.TBN.n118 XThR.TBN.t4 139.78
R16880 XThR.TBN.n122 XThR.TBN.t40 139.78
R16881 XThR.TBN.n119 XThR.TBN.t84 139.78
R16882 XThR.TBN.n115 XThR.TBN.t38 139.78
R16883 XThR.TBN.n106 XThR.TBN.t109 139.78
R16884 XThR.TBN.n110 XThR.TBN.t30 139.78
R16885 XThR.TBN.n107 XThR.TBN.t70 139.78
R16886 XThR.TBN.n103 XThR.TBN.t24 139.78
R16887 XThR.TBN.n94 XThR.TBN.t91 139.78
R16888 XThR.TBN.n98 XThR.TBN.t10 139.78
R16889 XThR.TBN.n95 XThR.TBN.t48 139.78
R16890 XThR.TBN.n92 XThR.TBN.t20 139.78
R16891 XThR.TBN.n83 XThR.TBN.t120 139.78
R16892 XThR.TBN.n87 XThR.TBN.t110 139.78
R16893 XThR.TBN.n84 XThR.TBN.t103 139.78
R16894 XThR.TBN.n167 XThR.TBN.t22 139.78
R16895 XThR.TBN.n169 XThR.TBN.t58 139.78
R16896 XThR.TBN.n174 XThR.TBN.t9 139.78
R16897 XThR.TBN.n170 XThR.TBN.t78 139.78
R16898 XThR.TBN.n184 XThR.TBN.n183 101.489
R16899 XThR.TBN.n179 XThR.TBN 58.2909
R16900 XThR.TBN.n7 XThR.TBN.n6 49.6611
R16901 XThR.TBN.n18 XThR.TBN.n17 49.6611
R16902 XThR.TBN.n30 XThR.TBN.n29 49.6611
R16903 XThR.TBN.n42 XThR.TBN.n41 49.6611
R16904 XThR.TBN.n54 XThR.TBN.n53 49.6611
R16905 XThR.TBN.n66 XThR.TBN.n65 49.6611
R16906 XThR.TBN.n78 XThR.TBN.n77 49.6611
R16907 XThR.TBN.n9 XThR.TBN.n8 44.549
R16908 XThR.TBN.n20 XThR.TBN.n19 44.549
R16909 XThR.TBN.n32 XThR.TBN.n31 44.549
R16910 XThR.TBN.n44 XThR.TBN.n43 44.549
R16911 XThR.TBN.n56 XThR.TBN.n55 44.549
R16912 XThR.TBN.n68 XThR.TBN.n67 44.549
R16913 XThR.TBN.n80 XThR.TBN.n79 44.549
R16914 XThR.TBN.n4 XThR.TBN.n2 43.0884
R16915 XThR.TBN.n15 XThR.TBN.n13 43.0884
R16916 XThR.TBN.n27 XThR.TBN.n25 43.0884
R16917 XThR.TBN.n39 XThR.TBN.n37 43.0884
R16918 XThR.TBN.n51 XThR.TBN.n49 43.0884
R16919 XThR.TBN.n63 XThR.TBN.n61 43.0884
R16920 XThR.TBN.n75 XThR.TBN.n73 43.0884
R16921 XThR.TBN.n163 XThR.TBN.n162 30.6732
R16922 XThR.TBN.n162 XThR.TBN.n154 30.6732
R16923 XThR.TBN.n159 XThR.TBN.n154 30.6732
R16924 XThR.TBN.n159 XThR.TBN.n158 30.6732
R16925 XThR.TBN.n158 XThR.TBN.n157 30.6732
R16926 XThR.TBN.n157 XThR.TBN.n155 30.6732
R16927 XThR.TBN.n151 XThR.TBN.n150 30.6732
R16928 XThR.TBN.n150 XThR.TBN.n142 30.6732
R16929 XThR.TBN.n147 XThR.TBN.n142 30.6732
R16930 XThR.TBN.n147 XThR.TBN.n146 30.6732
R16931 XThR.TBN.n146 XThR.TBN.n145 30.6732
R16932 XThR.TBN.n145 XThR.TBN.n143 30.6732
R16933 XThR.TBN.n139 XThR.TBN.n138 30.6732
R16934 XThR.TBN.n138 XThR.TBN.n130 30.6732
R16935 XThR.TBN.n135 XThR.TBN.n130 30.6732
R16936 XThR.TBN.n135 XThR.TBN.n134 30.6732
R16937 XThR.TBN.n134 XThR.TBN.n133 30.6732
R16938 XThR.TBN.n133 XThR.TBN.n131 30.6732
R16939 XThR.TBN.n127 XThR.TBN.n126 30.6732
R16940 XThR.TBN.n126 XThR.TBN.n118 30.6732
R16941 XThR.TBN.n123 XThR.TBN.n118 30.6732
R16942 XThR.TBN.n123 XThR.TBN.n122 30.6732
R16943 XThR.TBN.n122 XThR.TBN.n121 30.6732
R16944 XThR.TBN.n121 XThR.TBN.n119 30.6732
R16945 XThR.TBN.n115 XThR.TBN.n114 30.6732
R16946 XThR.TBN.n114 XThR.TBN.n106 30.6732
R16947 XThR.TBN.n111 XThR.TBN.n106 30.6732
R16948 XThR.TBN.n111 XThR.TBN.n110 30.6732
R16949 XThR.TBN.n110 XThR.TBN.n109 30.6732
R16950 XThR.TBN.n109 XThR.TBN.n107 30.6732
R16951 XThR.TBN.n103 XThR.TBN.n102 30.6732
R16952 XThR.TBN.n102 XThR.TBN.n94 30.6732
R16953 XThR.TBN.n99 XThR.TBN.n94 30.6732
R16954 XThR.TBN.n99 XThR.TBN.n98 30.6732
R16955 XThR.TBN.n98 XThR.TBN.n97 30.6732
R16956 XThR.TBN.n97 XThR.TBN.n95 30.6732
R16957 XThR.TBN.n92 XThR.TBN.n91 30.6732
R16958 XThR.TBN.n91 XThR.TBN.n83 30.6732
R16959 XThR.TBN.n88 XThR.TBN.n83 30.6732
R16960 XThR.TBN.n88 XThR.TBN.n87 30.6732
R16961 XThR.TBN.n87 XThR.TBN.n86 30.6732
R16962 XThR.TBN.n86 XThR.TBN.n84 30.6732
R16963 XThR.TBN.n168 XThR.TBN.n167 30.6732
R16964 XThR.TBN.n169 XThR.TBN.n168 30.6732
R16965 XThR.TBN.n175 XThR.TBN.n169 30.6732
R16966 XThR.TBN.n175 XThR.TBN.n174 30.6732
R16967 XThR.TBN.n174 XThR.TBN.n173 30.6732
R16968 XThR.TBN.n173 XThR.TBN.n170 30.6732
R16969 XThR.TBN.n180 XThR.TBN.t3 26.5955
R16970 XThR.TBN.n180 XThR.TBN.t2 26.5955
R16971 XThR.TBN.n183 XThR.TBN.t0 24.9236
R16972 XThR.TBN.n183 XThR.TBN.t1 24.9236
R16973 XThR.TBN.n10 XThR.TBN.n0 21.7605
R16974 XThR.TBN.n21 XThR.TBN.n11 21.7605
R16975 XThR.TBN.n33 XThR.TBN.n23 21.7605
R16976 XThR.TBN.n45 XThR.TBN.n35 21.7605
R16977 XThR.TBN.n57 XThR.TBN.n47 21.7605
R16978 XThR.TBN.n69 XThR.TBN.n59 21.7605
R16979 XThR.TBN.n81 XThR.TBN.n71 21.7605
R16980 XThR.TBN.n161 XThR.TBN 18.4325
R16981 XThR.TBN.n149 XThR.TBN 18.4325
R16982 XThR.TBN.n137 XThR.TBN 18.4325
R16983 XThR.TBN.n125 XThR.TBN 18.4325
R16984 XThR.TBN.n113 XThR.TBN 18.4325
R16985 XThR.TBN.n101 XThR.TBN 18.4325
R16986 XThR.TBN.n90 XThR.TBN 18.4325
R16987 XThR.TBN.n4 XThR.TBN.n3 18.2581
R16988 XThR.TBN.n15 XThR.TBN.n14 18.2581
R16989 XThR.TBN.n27 XThR.TBN.n26 18.2581
R16990 XThR.TBN.n39 XThR.TBN.n38 18.2581
R16991 XThR.TBN.n51 XThR.TBN.n50 18.2581
R16992 XThR.TBN.n63 XThR.TBN.n62 18.2581
R16993 XThR.TBN.n75 XThR.TBN.n74 18.2581
R16994 XThR.TBN.n5 XThR.TBN 17.6005
R16995 XThR.TBN.n16 XThR.TBN 17.6005
R16996 XThR.TBN.n28 XThR.TBN 17.6005
R16997 XThR.TBN.n40 XThR.TBN 17.6005
R16998 XThR.TBN.n52 XThR.TBN 17.6005
R16999 XThR.TBN.n64 XThR.TBN 17.6005
R17000 XThR.TBN.n76 XThR.TBN 17.6005
R17001 XThR.TBN.n22 XThR.TBN.n10 17.1655
R17002 XThR.TBN.n172 XThR.TBN 17.1525
R17003 XThR.TBN XThR.TBN.n171 17.1525
R17004 XThR.TBN.n105 XThR.TBN.n93 17.054
R17005 XThR.TBN.n9 XThR.TBN.n1 16.7975
R17006 XThR.TBN.n20 XThR.TBN.n12 16.7975
R17007 XThR.TBN.n32 XThR.TBN.n24 16.7975
R17008 XThR.TBN.n44 XThR.TBN.n36 16.7975
R17009 XThR.TBN.n56 XThR.TBN.n48 16.7975
R17010 XThR.TBN.n68 XThR.TBN.n60 16.7975
R17011 XThR.TBN.n80 XThR.TBN.n72 16.7975
R17012 XThR.TBN XThR.TBN.n160 16.3845
R17013 XThR.TBN XThR.TBN.n148 16.3845
R17014 XThR.TBN XThR.TBN.n136 16.3845
R17015 XThR.TBN XThR.TBN.n124 16.3845
R17016 XThR.TBN XThR.TBN.n112 16.3845
R17017 XThR.TBN XThR.TBN.n100 16.3845
R17018 XThR.TBN XThR.TBN.n89 16.3845
R17019 XThR.TBN.n22 XThR.TBN.n21 16.0405
R17020 XThR.TBN.n34 XThR.TBN.n33 16.0405
R17021 XThR.TBN.n46 XThR.TBN.n45 16.0405
R17022 XThR.TBN.n58 XThR.TBN.n57 16.0405
R17023 XThR.TBN.n70 XThR.TBN.n69 16.0405
R17024 XThR.TBN.n82 XThR.TBN.n81 16.0405
R17025 XThR.TBN.n165 XThR.TBN.n164 15.5925
R17026 XThR.TBN.n153 XThR.TBN.n152 15.5925
R17027 XThR.TBN.n141 XThR.TBN.n140 15.5925
R17028 XThR.TBN.n129 XThR.TBN.n128 15.5925
R17029 XThR.TBN.n117 XThR.TBN.n116 15.5925
R17030 XThR.TBN.n105 XThR.TBN.n104 15.5925
R17031 XThR.TBN.n156 XThR.TBN 14.3365
R17032 XThR.TBN.n144 XThR.TBN 14.3365
R17033 XThR.TBN.n132 XThR.TBN 14.3365
R17034 XThR.TBN.n120 XThR.TBN 14.3365
R17035 XThR.TBN.n108 XThR.TBN 14.3365
R17036 XThR.TBN.n96 XThR.TBN 14.3365
R17037 XThR.TBN.n85 XThR.TBN 14.3365
R17038 XThR.TBN XThR.TBN.n182 13.5685
R17039 XThR.TBN.n177 XThR.TBN.n176 12.2885
R17040 XThR.TBN XThR.TBN.n181 10.7525
R17041 XThR.TBN.n156 XThR.TBN 9.2165
R17042 XThR.TBN.n144 XThR.TBN 9.2165
R17043 XThR.TBN.n132 XThR.TBN 9.2165
R17044 XThR.TBN.n120 XThR.TBN 9.2165
R17045 XThR.TBN.n108 XThR.TBN 9.2165
R17046 XThR.TBN.n96 XThR.TBN 9.2165
R17047 XThR.TBN.n85 XThR.TBN 9.2165
R17048 XThR.TBN.n160 XThR.TBN 7.1685
R17049 XThR.TBN.n148 XThR.TBN 7.1685
R17050 XThR.TBN.n136 XThR.TBN 7.1685
R17051 XThR.TBN.n124 XThR.TBN 7.1685
R17052 XThR.TBN.n112 XThR.TBN 7.1685
R17053 XThR.TBN.n100 XThR.TBN 7.1685
R17054 XThR.TBN.n89 XThR.TBN 7.1685
R17055 XThR.TBN.n177 XThR.TBN 6.9125
R17056 XThR.TBN.n181 XThR.TBN 6.6565
R17057 XThR.TBN.n6 XThR.TBN.n2 6.57323
R17058 XThR.TBN.n17 XThR.TBN.n13 6.57323
R17059 XThR.TBN.n29 XThR.TBN.n25 6.57323
R17060 XThR.TBN.n41 XThR.TBN.n37 6.57323
R17061 XThR.TBN.n53 XThR.TBN.n49 6.57323
R17062 XThR.TBN.n65 XThR.TBN.n61 6.57323
R17063 XThR.TBN.n77 XThR.TBN.n73 6.57323
R17064 XThR.TBN.n172 XThR.TBN 6.4005
R17065 XThR.TBN.n171 XThR.TBN 6.4005
R17066 XThR.TBN.n179 XThR.TBN.n178 5.74665
R17067 XThR.TBN.n178 XThR.TBN.n166 5.74569
R17068 XThR.TBN.n161 XThR.TBN 5.1205
R17069 XThR.TBN.n149 XThR.TBN 5.1205
R17070 XThR.TBN.n137 XThR.TBN 5.1205
R17071 XThR.TBN.n125 XThR.TBN 5.1205
R17072 XThR.TBN.n113 XThR.TBN 5.1205
R17073 XThR.TBN.n101 XThR.TBN 5.1205
R17074 XThR.TBN.n90 XThR.TBN 5.1205
R17075 XThR.TBN.n8 XThR.TBN.n7 5.11262
R17076 XThR.TBN.n19 XThR.TBN.n18 5.11262
R17077 XThR.TBN.n31 XThR.TBN.n30 5.11262
R17078 XThR.TBN.n43 XThR.TBN.n42 5.11262
R17079 XThR.TBN.n55 XThR.TBN.n54 5.11262
R17080 XThR.TBN.n67 XThR.TBN.n66 5.11262
R17081 XThR.TBN.n79 XThR.TBN.n78 5.11262
R17082 XThR.TBN.n182 XThR.TBN.n179 5.06717
R17083 XThR.TBN.n181 XThR.TBN 5.04292
R17084 XThR.TBN.n178 XThR.TBN.n177 4.6505
R17085 XThR.TBN.n176 XThR.TBN 4.3525
R17086 XThR.TBN XThR.TBN.n0 4.1605
R17087 XThR.TBN XThR.TBN.n11 4.1605
R17088 XThR.TBN XThR.TBN.n23 4.1605
R17089 XThR.TBN XThR.TBN.n35 4.1605
R17090 XThR.TBN XThR.TBN.n47 4.1605
R17091 XThR.TBN XThR.TBN.n59 4.1605
R17092 XThR.TBN XThR.TBN.n71 4.1605
R17093 XThR.TBN.n182 XThR.TBN 3.8405
R17094 XThR.TBN.n184 XThR.TBN 2.5605
R17095 XThR.TBN.n164 XThR.TBN 2.3045
R17096 XThR.TBN.n152 XThR.TBN 2.3045
R17097 XThR.TBN.n140 XThR.TBN 2.3045
R17098 XThR.TBN.n128 XThR.TBN 2.3045
R17099 XThR.TBN.n116 XThR.TBN 2.3045
R17100 XThR.TBN.n104 XThR.TBN 2.3045
R17101 XThR.TBN.n93 XThR.TBN 2.3045
R17102 XThR.TBN XThR.TBN.n184 1.93989
R17103 XThR.TBN.n166 XThR.TBN.n82 1.53415
R17104 XThR.TBN.n34 XThR.TBN.n22 1.49088
R17105 XThR.TBN.n58 XThR.TBN.n46 1.49088
R17106 XThR.TBN.n82 XThR.TBN.n70 1.48608
R17107 XThR.TBN.n153 XThR.TBN.n141 1.46204
R17108 XThR.TBN.n129 XThR.TBN.n117 1.46204
R17109 XThR.TBN.n165 XThR.TBN.n153 1.15435
R17110 XThR.TBN.n141 XThR.TBN.n129 1.15435
R17111 XThR.TBN.n117 XThR.TBN.n105 1.15435
R17112 XThR.TBN XThR.TBN.n165 1.14473
R17113 XThR.TBN.n70 XThR.TBN.n58 1.13031
R17114 XThR.TBN.n46 XThR.TBN.n34 1.1255
R17115 XThR.TBN.n166 XThR.TBN 0.063
R17116 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R17117 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R17118 XThR.Tn[6] XThR.Tn[6].n82 161.363
R17119 XThR.Tn[6] XThR.Tn[6].n77 161.363
R17120 XThR.Tn[6] XThR.Tn[6].n72 161.363
R17121 XThR.Tn[6] XThR.Tn[6].n67 161.363
R17122 XThR.Tn[6] XThR.Tn[6].n62 161.363
R17123 XThR.Tn[6] XThR.Tn[6].n57 161.363
R17124 XThR.Tn[6] XThR.Tn[6].n52 161.363
R17125 XThR.Tn[6] XThR.Tn[6].n47 161.363
R17126 XThR.Tn[6] XThR.Tn[6].n42 161.363
R17127 XThR.Tn[6] XThR.Tn[6].n37 161.363
R17128 XThR.Tn[6] XThR.Tn[6].n32 161.363
R17129 XThR.Tn[6] XThR.Tn[6].n27 161.363
R17130 XThR.Tn[6] XThR.Tn[6].n22 161.363
R17131 XThR.Tn[6] XThR.Tn[6].n17 161.363
R17132 XThR.Tn[6] XThR.Tn[6].n12 161.363
R17133 XThR.Tn[6] XThR.Tn[6].n10 161.363
R17134 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R17135 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R17136 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R17137 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R17138 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R17139 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R17140 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R17141 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R17142 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R17143 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R17144 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R17145 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R17146 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R17147 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R17148 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R17149 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R17150 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R17151 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R17152 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R17153 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R17154 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R17155 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R17156 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R17157 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R17158 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R17159 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R17160 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R17161 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R17162 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R17163 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R17164 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R17165 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R17166 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R17167 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R17168 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R17169 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R17170 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R17171 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R17172 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R17173 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R17174 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R17175 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R17176 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R17177 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R17178 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R17179 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R17180 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R17181 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R17182 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R17183 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R17184 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R17185 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R17186 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R17187 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R17188 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R17189 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R17190 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R17191 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R17192 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R17193 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R17194 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R17195 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R17196 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R17197 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R17198 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R17199 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R17200 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R17201 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R17202 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R17203 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R17204 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R17205 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R17206 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R17207 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R17208 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R17209 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R17210 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R17211 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R17212 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R17213 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R17214 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R17215 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R17216 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R17217 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R17218 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R17219 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R17220 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R17221 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R17222 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R17223 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R17224 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R17225 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R17226 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R17227 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R17228 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R17229 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R17230 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R17231 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R17232 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R17233 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R17234 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R17235 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R17236 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R17237 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R17238 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R17239 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R17240 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R17241 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R17242 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R17243 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R17244 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R17245 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R17246 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R17247 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R17248 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R17249 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R17250 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R17251 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R17252 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R17253 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R17254 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R17255 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R17256 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R17257 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R17258 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R17259 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R17260 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R17261 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R17262 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R17263 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R17264 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R17265 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R17266 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R17267 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R17268 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R17269 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R17270 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R17271 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R17272 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R17273 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R17274 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R17275 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R17276 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R17277 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R17278 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R17279 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R17280 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R17281 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R17282 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R17283 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R17284 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R17285 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R17286 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R17287 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R17288 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R17289 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R17290 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R17291 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R17292 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R17293 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R17294 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R17295 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R17296 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R17297 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R17298 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R17299 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R17300 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R17301 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R17302 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R17303 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R17304 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R17305 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R17306 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R17307 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R17308 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R17309 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R17310 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R17311 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R17312 XThR.Tn[6] XThR.Tn[6].n87 0.038
R17313 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R17314 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R17315 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R17316 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R17317 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R17318 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R17319 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R17320 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R17321 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R17322 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R17323 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R17324 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R17325 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R17326 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R17327 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R17328 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R17329 XThR.Tn[14].n5 XThR.Tn[14].n4 256.103
R17330 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R17331 XThR.Tn[14].n88 XThR.Tn[14].n87 241.847
R17332 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R17333 XThR.Tn[14].n5 XThR.Tn[14].n3 202.095
R17334 XThR.Tn[14].n88 XThR.Tn[14].n86 185
R17335 XThR.Tn[14] XThR.Tn[14].n79 161.363
R17336 XThR.Tn[14] XThR.Tn[14].n74 161.363
R17337 XThR.Tn[14] XThR.Tn[14].n69 161.363
R17338 XThR.Tn[14] XThR.Tn[14].n64 161.363
R17339 XThR.Tn[14] XThR.Tn[14].n59 161.363
R17340 XThR.Tn[14] XThR.Tn[14].n54 161.363
R17341 XThR.Tn[14] XThR.Tn[14].n49 161.363
R17342 XThR.Tn[14] XThR.Tn[14].n44 161.363
R17343 XThR.Tn[14] XThR.Tn[14].n39 161.363
R17344 XThR.Tn[14] XThR.Tn[14].n34 161.363
R17345 XThR.Tn[14] XThR.Tn[14].n29 161.363
R17346 XThR.Tn[14] XThR.Tn[14].n24 161.363
R17347 XThR.Tn[14] XThR.Tn[14].n19 161.363
R17348 XThR.Tn[14] XThR.Tn[14].n14 161.363
R17349 XThR.Tn[14] XThR.Tn[14].n9 161.363
R17350 XThR.Tn[14] XThR.Tn[14].n7 161.363
R17351 XThR.Tn[14].n81 XThR.Tn[14].n80 161.3
R17352 XThR.Tn[14].n76 XThR.Tn[14].n75 161.3
R17353 XThR.Tn[14].n71 XThR.Tn[14].n70 161.3
R17354 XThR.Tn[14].n66 XThR.Tn[14].n65 161.3
R17355 XThR.Tn[14].n61 XThR.Tn[14].n60 161.3
R17356 XThR.Tn[14].n56 XThR.Tn[14].n55 161.3
R17357 XThR.Tn[14].n51 XThR.Tn[14].n50 161.3
R17358 XThR.Tn[14].n46 XThR.Tn[14].n45 161.3
R17359 XThR.Tn[14].n41 XThR.Tn[14].n40 161.3
R17360 XThR.Tn[14].n36 XThR.Tn[14].n35 161.3
R17361 XThR.Tn[14].n31 XThR.Tn[14].n30 161.3
R17362 XThR.Tn[14].n26 XThR.Tn[14].n25 161.3
R17363 XThR.Tn[14].n21 XThR.Tn[14].n20 161.3
R17364 XThR.Tn[14].n16 XThR.Tn[14].n15 161.3
R17365 XThR.Tn[14].n11 XThR.Tn[14].n10 161.3
R17366 XThR.Tn[14].n79 XThR.Tn[14].t51 161.106
R17367 XThR.Tn[14].n74 XThR.Tn[14].t58 161.106
R17368 XThR.Tn[14].n69 XThR.Tn[14].t39 161.106
R17369 XThR.Tn[14].n64 XThR.Tn[14].t22 161.106
R17370 XThR.Tn[14].n59 XThR.Tn[14].t49 161.106
R17371 XThR.Tn[14].n54 XThR.Tn[14].t12 161.106
R17372 XThR.Tn[14].n49 XThR.Tn[14].t56 161.106
R17373 XThR.Tn[14].n44 XThR.Tn[14].t36 161.106
R17374 XThR.Tn[14].n39 XThR.Tn[14].t19 161.106
R17375 XThR.Tn[14].n34 XThR.Tn[14].t25 161.106
R17376 XThR.Tn[14].n29 XThR.Tn[14].t73 161.106
R17377 XThR.Tn[14].n24 XThR.Tn[14].t38 161.106
R17378 XThR.Tn[14].n19 XThR.Tn[14].t72 161.106
R17379 XThR.Tn[14].n14 XThR.Tn[14].t54 161.106
R17380 XThR.Tn[14].n9 XThR.Tn[14].t13 161.106
R17381 XThR.Tn[14].n7 XThR.Tn[14].t62 161.106
R17382 XThR.Tn[14].n80 XThR.Tn[14].t32 159.978
R17383 XThR.Tn[14].n75 XThR.Tn[14].t37 159.978
R17384 XThR.Tn[14].n70 XThR.Tn[14].t20 159.978
R17385 XThR.Tn[14].n65 XThR.Tn[14].t68 159.978
R17386 XThR.Tn[14].n60 XThR.Tn[14].t30 159.978
R17387 XThR.Tn[14].n55 XThR.Tn[14].t55 159.978
R17388 XThR.Tn[14].n50 XThR.Tn[14].t35 159.978
R17389 XThR.Tn[14].n45 XThR.Tn[14].t16 159.978
R17390 XThR.Tn[14].n40 XThR.Tn[14].t66 159.978
R17391 XThR.Tn[14].n35 XThR.Tn[14].t71 159.978
R17392 XThR.Tn[14].n30 XThR.Tn[14].t53 159.978
R17393 XThR.Tn[14].n25 XThR.Tn[14].t18 159.978
R17394 XThR.Tn[14].n20 XThR.Tn[14].t52 159.978
R17395 XThR.Tn[14].n15 XThR.Tn[14].t34 159.978
R17396 XThR.Tn[14].n10 XThR.Tn[14].t60 159.978
R17397 XThR.Tn[14].n79 XThR.Tn[14].t41 145.038
R17398 XThR.Tn[14].n74 XThR.Tn[14].t65 145.038
R17399 XThR.Tn[14].n69 XThR.Tn[14].t45 145.038
R17400 XThR.Tn[14].n64 XThR.Tn[14].t26 145.038
R17401 XThR.Tn[14].n59 XThR.Tn[14].t59 145.038
R17402 XThR.Tn[14].n54 XThR.Tn[14].t40 145.038
R17403 XThR.Tn[14].n49 XThR.Tn[14].t46 145.038
R17404 XThR.Tn[14].n44 XThR.Tn[14].t27 145.038
R17405 XThR.Tn[14].n39 XThR.Tn[14].t23 145.038
R17406 XThR.Tn[14].n34 XThR.Tn[14].t57 145.038
R17407 XThR.Tn[14].n29 XThR.Tn[14].t15 145.038
R17408 XThR.Tn[14].n24 XThR.Tn[14].t44 145.038
R17409 XThR.Tn[14].n19 XThR.Tn[14].t14 145.038
R17410 XThR.Tn[14].n14 XThR.Tn[14].t64 145.038
R17411 XThR.Tn[14].n9 XThR.Tn[14].t24 145.038
R17412 XThR.Tn[14].n7 XThR.Tn[14].t69 145.038
R17413 XThR.Tn[14].n80 XThR.Tn[14].t43 143.911
R17414 XThR.Tn[14].n75 XThR.Tn[14].t70 143.911
R17415 XThR.Tn[14].n70 XThR.Tn[14].t48 143.911
R17416 XThR.Tn[14].n65 XThR.Tn[14].t31 143.911
R17417 XThR.Tn[14].n60 XThR.Tn[14].t63 143.911
R17418 XThR.Tn[14].n55 XThR.Tn[14].t42 143.911
R17419 XThR.Tn[14].n50 XThR.Tn[14].t50 143.911
R17420 XThR.Tn[14].n45 XThR.Tn[14].t33 143.911
R17421 XThR.Tn[14].n40 XThR.Tn[14].t29 143.911
R17422 XThR.Tn[14].n35 XThR.Tn[14].t61 143.911
R17423 XThR.Tn[14].n30 XThR.Tn[14].t21 143.911
R17424 XThR.Tn[14].n25 XThR.Tn[14].t47 143.911
R17425 XThR.Tn[14].n20 XThR.Tn[14].t17 143.911
R17426 XThR.Tn[14].n15 XThR.Tn[14].t67 143.911
R17427 XThR.Tn[14].n10 XThR.Tn[14].t28 143.911
R17428 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17429 XThR.Tn[14].n3 XThR.Tn[14].t6 26.5955
R17430 XThR.Tn[14].n3 XThR.Tn[14].t7 26.5955
R17431 XThR.Tn[14].n4 XThR.Tn[14].t4 26.5955
R17432 XThR.Tn[14].n4 XThR.Tn[14].t5 26.5955
R17433 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R17434 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R17435 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R17436 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R17437 XThR.Tn[14].n86 XThR.Tn[14].t0 24.9236
R17438 XThR.Tn[14].n86 XThR.Tn[14].t1 24.9236
R17439 XThR.Tn[14].n87 XThR.Tn[14].t2 24.9236
R17440 XThR.Tn[14].n87 XThR.Tn[14].t3 24.9236
R17441 XThR.Tn[14] XThR.Tn[14].n88 18.8943
R17442 XThR.Tn[14].n6 XThR.Tn[14].n5 13.5534
R17443 XThR.Tn[14].n85 XThR.Tn[14] 8.47191
R17444 XThR.Tn[14] XThR.Tn[14].n85 6.34069
R17445 XThR.Tn[14] XThR.Tn[14].n8 5.34038
R17446 XThR.Tn[14].n13 XThR.Tn[14].n12 4.5005
R17447 XThR.Tn[14].n18 XThR.Tn[14].n17 4.5005
R17448 XThR.Tn[14].n23 XThR.Tn[14].n22 4.5005
R17449 XThR.Tn[14].n28 XThR.Tn[14].n27 4.5005
R17450 XThR.Tn[14].n33 XThR.Tn[14].n32 4.5005
R17451 XThR.Tn[14].n38 XThR.Tn[14].n37 4.5005
R17452 XThR.Tn[14].n43 XThR.Tn[14].n42 4.5005
R17453 XThR.Tn[14].n48 XThR.Tn[14].n47 4.5005
R17454 XThR.Tn[14].n53 XThR.Tn[14].n52 4.5005
R17455 XThR.Tn[14].n58 XThR.Tn[14].n57 4.5005
R17456 XThR.Tn[14].n63 XThR.Tn[14].n62 4.5005
R17457 XThR.Tn[14].n68 XThR.Tn[14].n67 4.5005
R17458 XThR.Tn[14].n73 XThR.Tn[14].n72 4.5005
R17459 XThR.Tn[14].n78 XThR.Tn[14].n77 4.5005
R17460 XThR.Tn[14].n83 XThR.Tn[14].n82 4.5005
R17461 XThR.Tn[14].n84 XThR.Tn[14] 3.70586
R17462 XThR.Tn[14].n13 XThR.Tn[14] 2.52282
R17463 XThR.Tn[14].n18 XThR.Tn[14] 2.52282
R17464 XThR.Tn[14].n23 XThR.Tn[14] 2.52282
R17465 XThR.Tn[14].n28 XThR.Tn[14] 2.52282
R17466 XThR.Tn[14].n33 XThR.Tn[14] 2.52282
R17467 XThR.Tn[14].n38 XThR.Tn[14] 2.52282
R17468 XThR.Tn[14].n43 XThR.Tn[14] 2.52282
R17469 XThR.Tn[14].n48 XThR.Tn[14] 2.52282
R17470 XThR.Tn[14].n53 XThR.Tn[14] 2.52282
R17471 XThR.Tn[14].n58 XThR.Tn[14] 2.52282
R17472 XThR.Tn[14].n63 XThR.Tn[14] 2.52282
R17473 XThR.Tn[14].n68 XThR.Tn[14] 2.52282
R17474 XThR.Tn[14].n73 XThR.Tn[14] 2.52282
R17475 XThR.Tn[14].n78 XThR.Tn[14] 2.52282
R17476 XThR.Tn[14].n83 XThR.Tn[14] 2.52282
R17477 XThR.Tn[14].n85 XThR.Tn[14] 1.79489
R17478 XThR.Tn[14].n6 XThR.Tn[14] 1.50638
R17479 XThR.Tn[14] XThR.Tn[14].n6 1.19676
R17480 XThR.Tn[14].n81 XThR.Tn[14] 1.08677
R17481 XThR.Tn[14].n76 XThR.Tn[14] 1.08677
R17482 XThR.Tn[14].n71 XThR.Tn[14] 1.08677
R17483 XThR.Tn[14].n66 XThR.Tn[14] 1.08677
R17484 XThR.Tn[14].n61 XThR.Tn[14] 1.08677
R17485 XThR.Tn[14].n56 XThR.Tn[14] 1.08677
R17486 XThR.Tn[14].n51 XThR.Tn[14] 1.08677
R17487 XThR.Tn[14].n46 XThR.Tn[14] 1.08677
R17488 XThR.Tn[14].n41 XThR.Tn[14] 1.08677
R17489 XThR.Tn[14].n36 XThR.Tn[14] 1.08677
R17490 XThR.Tn[14].n31 XThR.Tn[14] 1.08677
R17491 XThR.Tn[14].n26 XThR.Tn[14] 1.08677
R17492 XThR.Tn[14].n21 XThR.Tn[14] 1.08677
R17493 XThR.Tn[14].n16 XThR.Tn[14] 1.08677
R17494 XThR.Tn[14].n11 XThR.Tn[14] 1.08677
R17495 XThR.Tn[14] XThR.Tn[14].n13 0.839786
R17496 XThR.Tn[14] XThR.Tn[14].n18 0.839786
R17497 XThR.Tn[14] XThR.Tn[14].n23 0.839786
R17498 XThR.Tn[14] XThR.Tn[14].n28 0.839786
R17499 XThR.Tn[14] XThR.Tn[14].n33 0.839786
R17500 XThR.Tn[14] XThR.Tn[14].n38 0.839786
R17501 XThR.Tn[14] XThR.Tn[14].n43 0.839786
R17502 XThR.Tn[14] XThR.Tn[14].n48 0.839786
R17503 XThR.Tn[14] XThR.Tn[14].n53 0.839786
R17504 XThR.Tn[14] XThR.Tn[14].n58 0.839786
R17505 XThR.Tn[14] XThR.Tn[14].n63 0.839786
R17506 XThR.Tn[14] XThR.Tn[14].n68 0.839786
R17507 XThR.Tn[14] XThR.Tn[14].n73 0.839786
R17508 XThR.Tn[14] XThR.Tn[14].n78 0.839786
R17509 XThR.Tn[14] XThR.Tn[14].n83 0.839786
R17510 XThR.Tn[14].n8 XThR.Tn[14] 0.499542
R17511 XThR.Tn[14].n82 XThR.Tn[14] 0.063
R17512 XThR.Tn[14].n77 XThR.Tn[14] 0.063
R17513 XThR.Tn[14].n72 XThR.Tn[14] 0.063
R17514 XThR.Tn[14].n67 XThR.Tn[14] 0.063
R17515 XThR.Tn[14].n62 XThR.Tn[14] 0.063
R17516 XThR.Tn[14].n57 XThR.Tn[14] 0.063
R17517 XThR.Tn[14].n52 XThR.Tn[14] 0.063
R17518 XThR.Tn[14].n47 XThR.Tn[14] 0.063
R17519 XThR.Tn[14].n42 XThR.Tn[14] 0.063
R17520 XThR.Tn[14].n37 XThR.Tn[14] 0.063
R17521 XThR.Tn[14].n32 XThR.Tn[14] 0.063
R17522 XThR.Tn[14].n27 XThR.Tn[14] 0.063
R17523 XThR.Tn[14].n22 XThR.Tn[14] 0.063
R17524 XThR.Tn[14].n17 XThR.Tn[14] 0.063
R17525 XThR.Tn[14].n12 XThR.Tn[14] 0.063
R17526 XThR.Tn[14].n84 XThR.Tn[14] 0.0540714
R17527 XThR.Tn[14] XThR.Tn[14].n84 0.038
R17528 XThR.Tn[14].n8 XThR.Tn[14] 0.0143889
R17529 XThR.Tn[14].n82 XThR.Tn[14].n81 0.00771154
R17530 XThR.Tn[14].n77 XThR.Tn[14].n76 0.00771154
R17531 XThR.Tn[14].n72 XThR.Tn[14].n71 0.00771154
R17532 XThR.Tn[14].n67 XThR.Tn[14].n66 0.00771154
R17533 XThR.Tn[14].n62 XThR.Tn[14].n61 0.00771154
R17534 XThR.Tn[14].n57 XThR.Tn[14].n56 0.00771154
R17535 XThR.Tn[14].n52 XThR.Tn[14].n51 0.00771154
R17536 XThR.Tn[14].n47 XThR.Tn[14].n46 0.00771154
R17537 XThR.Tn[14].n42 XThR.Tn[14].n41 0.00771154
R17538 XThR.Tn[14].n37 XThR.Tn[14].n36 0.00771154
R17539 XThR.Tn[14].n32 XThR.Tn[14].n31 0.00771154
R17540 XThR.Tn[14].n27 XThR.Tn[14].n26 0.00771154
R17541 XThR.Tn[14].n22 XThR.Tn[14].n21 0.00771154
R17542 XThR.Tn[14].n17 XThR.Tn[14].n16 0.00771154
R17543 XThR.Tn[14].n12 XThR.Tn[14].n11 0.00771154
R17544 XThR.Tn[12].n5 XThR.Tn[12].n4 256.103
R17545 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R17546 XThR.Tn[12].n88 XThR.Tn[12].n87 241.847
R17547 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R17548 XThR.Tn[12].n5 XThR.Tn[12].n3 202.095
R17549 XThR.Tn[12].n88 XThR.Tn[12].n86 185
R17550 XThR.Tn[12] XThR.Tn[12].n79 161.363
R17551 XThR.Tn[12] XThR.Tn[12].n74 161.363
R17552 XThR.Tn[12] XThR.Tn[12].n69 161.363
R17553 XThR.Tn[12] XThR.Tn[12].n64 161.363
R17554 XThR.Tn[12] XThR.Tn[12].n59 161.363
R17555 XThR.Tn[12] XThR.Tn[12].n54 161.363
R17556 XThR.Tn[12] XThR.Tn[12].n49 161.363
R17557 XThR.Tn[12] XThR.Tn[12].n44 161.363
R17558 XThR.Tn[12] XThR.Tn[12].n39 161.363
R17559 XThR.Tn[12] XThR.Tn[12].n34 161.363
R17560 XThR.Tn[12] XThR.Tn[12].n29 161.363
R17561 XThR.Tn[12] XThR.Tn[12].n24 161.363
R17562 XThR.Tn[12] XThR.Tn[12].n19 161.363
R17563 XThR.Tn[12] XThR.Tn[12].n14 161.363
R17564 XThR.Tn[12] XThR.Tn[12].n9 161.363
R17565 XThR.Tn[12] XThR.Tn[12].n7 161.363
R17566 XThR.Tn[12].n81 XThR.Tn[12].n80 161.3
R17567 XThR.Tn[12].n76 XThR.Tn[12].n75 161.3
R17568 XThR.Tn[12].n71 XThR.Tn[12].n70 161.3
R17569 XThR.Tn[12].n66 XThR.Tn[12].n65 161.3
R17570 XThR.Tn[12].n61 XThR.Tn[12].n60 161.3
R17571 XThR.Tn[12].n56 XThR.Tn[12].n55 161.3
R17572 XThR.Tn[12].n51 XThR.Tn[12].n50 161.3
R17573 XThR.Tn[12].n46 XThR.Tn[12].n45 161.3
R17574 XThR.Tn[12].n41 XThR.Tn[12].n40 161.3
R17575 XThR.Tn[12].n36 XThR.Tn[12].n35 161.3
R17576 XThR.Tn[12].n31 XThR.Tn[12].n30 161.3
R17577 XThR.Tn[12].n26 XThR.Tn[12].n25 161.3
R17578 XThR.Tn[12].n21 XThR.Tn[12].n20 161.3
R17579 XThR.Tn[12].n16 XThR.Tn[12].n15 161.3
R17580 XThR.Tn[12].n11 XThR.Tn[12].n10 161.3
R17581 XThR.Tn[12].n79 XThR.Tn[12].t18 161.106
R17582 XThR.Tn[12].n74 XThR.Tn[12].t24 161.106
R17583 XThR.Tn[12].n69 XThR.Tn[12].t67 161.106
R17584 XThR.Tn[12].n64 XThR.Tn[12].t52 161.106
R17585 XThR.Tn[12].n59 XThR.Tn[12].t16 161.106
R17586 XThR.Tn[12].n54 XThR.Tn[12].t40 161.106
R17587 XThR.Tn[12].n49 XThR.Tn[12].t22 161.106
R17588 XThR.Tn[12].n44 XThR.Tn[12].t65 161.106
R17589 XThR.Tn[12].n39 XThR.Tn[12].t51 161.106
R17590 XThR.Tn[12].n34 XThR.Tn[12].t56 161.106
R17591 XThR.Tn[12].n29 XThR.Tn[12].t39 161.106
R17592 XThR.Tn[12].n24 XThR.Tn[12].t66 161.106
R17593 XThR.Tn[12].n19 XThR.Tn[12].t38 161.106
R17594 XThR.Tn[12].n14 XThR.Tn[12].t20 161.106
R17595 XThR.Tn[12].n9 XThR.Tn[12].t43 161.106
R17596 XThR.Tn[12].n7 XThR.Tn[12].t28 161.106
R17597 XThR.Tn[12].n80 XThR.Tn[12].t58 159.978
R17598 XThR.Tn[12].n75 XThR.Tn[12].t62 159.978
R17599 XThR.Tn[12].n70 XThR.Tn[12].t47 159.978
R17600 XThR.Tn[12].n65 XThR.Tn[12].t31 159.978
R17601 XThR.Tn[12].n60 XThR.Tn[12].t55 159.978
R17602 XThR.Tn[12].n55 XThR.Tn[12].t19 159.978
R17603 XThR.Tn[12].n50 XThR.Tn[12].t61 159.978
R17604 XThR.Tn[12].n45 XThR.Tn[12].t44 159.978
R17605 XThR.Tn[12].n40 XThR.Tn[12].t29 159.978
R17606 XThR.Tn[12].n35 XThR.Tn[12].t37 159.978
R17607 XThR.Tn[12].n30 XThR.Tn[12].t17 159.978
R17608 XThR.Tn[12].n25 XThR.Tn[12].t46 159.978
R17609 XThR.Tn[12].n20 XThR.Tn[12].t15 159.978
R17610 XThR.Tn[12].n15 XThR.Tn[12].t60 159.978
R17611 XThR.Tn[12].n10 XThR.Tn[12].t21 159.978
R17612 XThR.Tn[12].n79 XThR.Tn[12].t69 145.038
R17613 XThR.Tn[12].n74 XThR.Tn[12].t32 145.038
R17614 XThR.Tn[12].n69 XThR.Tn[12].t73 145.038
R17615 XThR.Tn[12].n64 XThR.Tn[12].t57 145.038
R17616 XThR.Tn[12].n59 XThR.Tn[12].t25 145.038
R17617 XThR.Tn[12].n54 XThR.Tn[12].t68 145.038
R17618 XThR.Tn[12].n49 XThR.Tn[12].t12 145.038
R17619 XThR.Tn[12].n44 XThR.Tn[12].t59 145.038
R17620 XThR.Tn[12].n39 XThR.Tn[12].t54 145.038
R17621 XThR.Tn[12].n34 XThR.Tn[12].t23 145.038
R17622 XThR.Tn[12].n29 XThR.Tn[12].t48 145.038
R17623 XThR.Tn[12].n24 XThR.Tn[12].t70 145.038
R17624 XThR.Tn[12].n19 XThR.Tn[12].t45 145.038
R17625 XThR.Tn[12].n14 XThR.Tn[12].t30 145.038
R17626 XThR.Tn[12].n9 XThR.Tn[12].t53 145.038
R17627 XThR.Tn[12].n7 XThR.Tn[12].t36 145.038
R17628 XThR.Tn[12].n80 XThR.Tn[12].t27 143.911
R17629 XThR.Tn[12].n75 XThR.Tn[12].t50 143.911
R17630 XThR.Tn[12].n70 XThR.Tn[12].t34 143.911
R17631 XThR.Tn[12].n65 XThR.Tn[12].t13 143.911
R17632 XThR.Tn[12].n60 XThR.Tn[12].t42 143.911
R17633 XThR.Tn[12].n55 XThR.Tn[12].t26 143.911
R17634 XThR.Tn[12].n50 XThR.Tn[12].t35 143.911
R17635 XThR.Tn[12].n45 XThR.Tn[12].t14 143.911
R17636 XThR.Tn[12].n40 XThR.Tn[12].t72 143.911
R17637 XThR.Tn[12].n35 XThR.Tn[12].t41 143.911
R17638 XThR.Tn[12].n30 XThR.Tn[12].t64 143.911
R17639 XThR.Tn[12].n25 XThR.Tn[12].t33 143.911
R17640 XThR.Tn[12].n20 XThR.Tn[12].t63 143.911
R17641 XThR.Tn[12].n15 XThR.Tn[12].t49 143.911
R17642 XThR.Tn[12].n10 XThR.Tn[12].t71 143.911
R17643 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17644 XThR.Tn[12].n3 XThR.Tn[12].t6 26.5955
R17645 XThR.Tn[12].n3 XThR.Tn[12].t4 26.5955
R17646 XThR.Tn[12].n4 XThR.Tn[12].t7 26.5955
R17647 XThR.Tn[12].n4 XThR.Tn[12].t5 26.5955
R17648 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R17649 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R17650 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R17651 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R17652 XThR.Tn[12].n86 XThR.Tn[12].t2 24.9236
R17653 XThR.Tn[12].n86 XThR.Tn[12].t0 24.9236
R17654 XThR.Tn[12].n87 XThR.Tn[12].t3 24.9236
R17655 XThR.Tn[12].n87 XThR.Tn[12].t1 24.9236
R17656 XThR.Tn[12] XThR.Tn[12].n88 18.8943
R17657 XThR.Tn[12].n6 XThR.Tn[12].n5 13.5534
R17658 XThR.Tn[12].n85 XThR.Tn[12] 8.18715
R17659 XThR.Tn[12] XThR.Tn[12].n85 6.34069
R17660 XThR.Tn[12] XThR.Tn[12].n8 5.34038
R17661 XThR.Tn[12].n13 XThR.Tn[12].n12 4.5005
R17662 XThR.Tn[12].n18 XThR.Tn[12].n17 4.5005
R17663 XThR.Tn[12].n23 XThR.Tn[12].n22 4.5005
R17664 XThR.Tn[12].n28 XThR.Tn[12].n27 4.5005
R17665 XThR.Tn[12].n33 XThR.Tn[12].n32 4.5005
R17666 XThR.Tn[12].n38 XThR.Tn[12].n37 4.5005
R17667 XThR.Tn[12].n43 XThR.Tn[12].n42 4.5005
R17668 XThR.Tn[12].n48 XThR.Tn[12].n47 4.5005
R17669 XThR.Tn[12].n53 XThR.Tn[12].n52 4.5005
R17670 XThR.Tn[12].n58 XThR.Tn[12].n57 4.5005
R17671 XThR.Tn[12].n63 XThR.Tn[12].n62 4.5005
R17672 XThR.Tn[12].n68 XThR.Tn[12].n67 4.5005
R17673 XThR.Tn[12].n73 XThR.Tn[12].n72 4.5005
R17674 XThR.Tn[12].n78 XThR.Tn[12].n77 4.5005
R17675 XThR.Tn[12].n83 XThR.Tn[12].n82 4.5005
R17676 XThR.Tn[12].n84 XThR.Tn[12] 3.70586
R17677 XThR.Tn[12].n13 XThR.Tn[12] 2.52282
R17678 XThR.Tn[12].n18 XThR.Tn[12] 2.52282
R17679 XThR.Tn[12].n23 XThR.Tn[12] 2.52282
R17680 XThR.Tn[12].n28 XThR.Tn[12] 2.52282
R17681 XThR.Tn[12].n33 XThR.Tn[12] 2.52282
R17682 XThR.Tn[12].n38 XThR.Tn[12] 2.52282
R17683 XThR.Tn[12].n43 XThR.Tn[12] 2.52282
R17684 XThR.Tn[12].n48 XThR.Tn[12] 2.52282
R17685 XThR.Tn[12].n53 XThR.Tn[12] 2.52282
R17686 XThR.Tn[12].n58 XThR.Tn[12] 2.52282
R17687 XThR.Tn[12].n63 XThR.Tn[12] 2.52282
R17688 XThR.Tn[12].n68 XThR.Tn[12] 2.52282
R17689 XThR.Tn[12].n73 XThR.Tn[12] 2.52282
R17690 XThR.Tn[12].n78 XThR.Tn[12] 2.52282
R17691 XThR.Tn[12].n83 XThR.Tn[12] 2.52282
R17692 XThR.Tn[12].n85 XThR.Tn[12] 1.79489
R17693 XThR.Tn[12].n6 XThR.Tn[12] 1.50638
R17694 XThR.Tn[12] XThR.Tn[12].n6 1.19676
R17695 XThR.Tn[12].n81 XThR.Tn[12] 1.08677
R17696 XThR.Tn[12].n76 XThR.Tn[12] 1.08677
R17697 XThR.Tn[12].n71 XThR.Tn[12] 1.08677
R17698 XThR.Tn[12].n66 XThR.Tn[12] 1.08677
R17699 XThR.Tn[12].n61 XThR.Tn[12] 1.08677
R17700 XThR.Tn[12].n56 XThR.Tn[12] 1.08677
R17701 XThR.Tn[12].n51 XThR.Tn[12] 1.08677
R17702 XThR.Tn[12].n46 XThR.Tn[12] 1.08677
R17703 XThR.Tn[12].n41 XThR.Tn[12] 1.08677
R17704 XThR.Tn[12].n36 XThR.Tn[12] 1.08677
R17705 XThR.Tn[12].n31 XThR.Tn[12] 1.08677
R17706 XThR.Tn[12].n26 XThR.Tn[12] 1.08677
R17707 XThR.Tn[12].n21 XThR.Tn[12] 1.08677
R17708 XThR.Tn[12].n16 XThR.Tn[12] 1.08677
R17709 XThR.Tn[12].n11 XThR.Tn[12] 1.08677
R17710 XThR.Tn[12] XThR.Tn[12].n13 0.839786
R17711 XThR.Tn[12] XThR.Tn[12].n18 0.839786
R17712 XThR.Tn[12] XThR.Tn[12].n23 0.839786
R17713 XThR.Tn[12] XThR.Tn[12].n28 0.839786
R17714 XThR.Tn[12] XThR.Tn[12].n33 0.839786
R17715 XThR.Tn[12] XThR.Tn[12].n38 0.839786
R17716 XThR.Tn[12] XThR.Tn[12].n43 0.839786
R17717 XThR.Tn[12] XThR.Tn[12].n48 0.839786
R17718 XThR.Tn[12] XThR.Tn[12].n53 0.839786
R17719 XThR.Tn[12] XThR.Tn[12].n58 0.839786
R17720 XThR.Tn[12] XThR.Tn[12].n63 0.839786
R17721 XThR.Tn[12] XThR.Tn[12].n68 0.839786
R17722 XThR.Tn[12] XThR.Tn[12].n73 0.839786
R17723 XThR.Tn[12] XThR.Tn[12].n78 0.839786
R17724 XThR.Tn[12] XThR.Tn[12].n83 0.839786
R17725 XThR.Tn[12].n8 XThR.Tn[12] 0.499542
R17726 XThR.Tn[12].n82 XThR.Tn[12] 0.063
R17727 XThR.Tn[12].n77 XThR.Tn[12] 0.063
R17728 XThR.Tn[12].n72 XThR.Tn[12] 0.063
R17729 XThR.Tn[12].n67 XThR.Tn[12] 0.063
R17730 XThR.Tn[12].n62 XThR.Tn[12] 0.063
R17731 XThR.Tn[12].n57 XThR.Tn[12] 0.063
R17732 XThR.Tn[12].n52 XThR.Tn[12] 0.063
R17733 XThR.Tn[12].n47 XThR.Tn[12] 0.063
R17734 XThR.Tn[12].n42 XThR.Tn[12] 0.063
R17735 XThR.Tn[12].n37 XThR.Tn[12] 0.063
R17736 XThR.Tn[12].n32 XThR.Tn[12] 0.063
R17737 XThR.Tn[12].n27 XThR.Tn[12] 0.063
R17738 XThR.Tn[12].n22 XThR.Tn[12] 0.063
R17739 XThR.Tn[12].n17 XThR.Tn[12] 0.063
R17740 XThR.Tn[12].n12 XThR.Tn[12] 0.063
R17741 XThR.Tn[12].n84 XThR.Tn[12] 0.0540714
R17742 XThR.Tn[12] XThR.Tn[12].n84 0.038
R17743 XThR.Tn[12].n8 XThR.Tn[12] 0.0143889
R17744 XThR.Tn[12].n82 XThR.Tn[12].n81 0.00771154
R17745 XThR.Tn[12].n77 XThR.Tn[12].n76 0.00771154
R17746 XThR.Tn[12].n72 XThR.Tn[12].n71 0.00771154
R17747 XThR.Tn[12].n67 XThR.Tn[12].n66 0.00771154
R17748 XThR.Tn[12].n62 XThR.Tn[12].n61 0.00771154
R17749 XThR.Tn[12].n57 XThR.Tn[12].n56 0.00771154
R17750 XThR.Tn[12].n52 XThR.Tn[12].n51 0.00771154
R17751 XThR.Tn[12].n47 XThR.Tn[12].n46 0.00771154
R17752 XThR.Tn[12].n42 XThR.Tn[12].n41 0.00771154
R17753 XThR.Tn[12].n37 XThR.Tn[12].n36 0.00771154
R17754 XThR.Tn[12].n32 XThR.Tn[12].n31 0.00771154
R17755 XThR.Tn[12].n27 XThR.Tn[12].n26 0.00771154
R17756 XThR.Tn[12].n22 XThR.Tn[12].n21 0.00771154
R17757 XThR.Tn[12].n17 XThR.Tn[12].n16 0.00771154
R17758 XThR.Tn[12].n12 XThR.Tn[12].n11 0.00771154
R17759 XThC.TBN.n183 XThC.TBN.t9 212.081
R17760 XThC.TBN.n182 XThC.TBN.t75 212.081
R17761 XThC.TBN.n176 XThC.TBN.t33 212.081
R17762 XThC.TBN.n177 XThC.TBN.t27 212.081
R17763 XThC.TBN.n87 XThC.TBN.t25 212.081
R17764 XThC.TBN.n78 XThC.TBN.t100 212.081
R17765 XThC.TBN.n82 XThC.TBN.t93 212.081
R17766 XThC.TBN.n80 XThC.TBN.t90 212.081
R17767 XThC.TBN.n61 XThC.TBN.t47 212.081
R17768 XThC.TBN.n52 XThC.TBN.t17 212.081
R17769 XThC.TBN.n56 XThC.TBN.t116 212.081
R17770 XThC.TBN.n54 XThC.TBN.t111 212.081
R17771 XThC.TBN.n35 XThC.TBN.t106 212.081
R17772 XThC.TBN.n26 XThC.TBN.t70 212.081
R17773 XThC.TBN.n30 XThC.TBN.t56 212.081
R17774 XThC.TBN.n28 XThC.TBN.t48 212.081
R17775 XThC.TBN.n10 XThC.TBN.t50 212.081
R17776 XThC.TBN.n1 XThC.TBN.t18 212.081
R17777 XThC.TBN.n5 XThC.TBN.t120 212.081
R17778 XThC.TBN.n3 XThC.TBN.t114 212.081
R17779 XThC.TBN.n74 XThC.TBN.t101 212.081
R17780 XThC.TBN.n65 XThC.TBN.t63 212.081
R17781 XThC.TBN.n69 XThC.TBN.t52 212.081
R17782 XThC.TBN.n67 XThC.TBN.t44 212.081
R17783 XThC.TBN.n48 XThC.TBN.t39 212.081
R17784 XThC.TBN.n39 XThC.TBN.t122 212.081
R17785 XThC.TBN.n43 XThC.TBN.t109 212.081
R17786 XThC.TBN.n41 XThC.TBN.t102 212.081
R17787 XThC.TBN.n22 XThC.TBN.t79 212.081
R17788 XThC.TBN.n13 XThC.TBN.t36 212.081
R17789 XThC.TBN.n17 XThC.TBN.t26 212.081
R17790 XThC.TBN.n15 XThC.TBN.t21 212.081
R17791 XThC.TBN.n100 XThC.TBN.t54 212.081
R17792 XThC.TBN.n99 XThC.TBN.t46 212.081
R17793 XThC.TBN.n94 XThC.TBN.t12 212.081
R17794 XThC.TBN.n93 XThC.TBN.t6 212.081
R17795 XThC.TBN.n123 XThC.TBN.t34 212.081
R17796 XThC.TBN.n122 XThC.TBN.t30 212.081
R17797 XThC.TBN.n117 XThC.TBN.t103 212.081
R17798 XThC.TBN.n116 XThC.TBN.t98 212.081
R17799 XThC.TBN.n147 XThC.TBN.t91 212.081
R17800 XThC.TBN.n146 XThC.TBN.t88 212.081
R17801 XThC.TBN.n141 XThC.TBN.t40 212.081
R17802 XThC.TBN.n140 XThC.TBN.t37 212.081
R17803 XThC.TBN.n171 XThC.TBN.t28 212.081
R17804 XThC.TBN.n170 XThC.TBN.t23 212.081
R17805 XThC.TBN.n165 XThC.TBN.t97 212.081
R17806 XThC.TBN.n164 XThC.TBN.t95 212.081
R17807 XThC.TBN.n111 XThC.TBN.t42 212.081
R17808 XThC.TBN.n110 XThC.TBN.t38 212.081
R17809 XThC.TBN.n105 XThC.TBN.t119 212.081
R17810 XThC.TBN.n104 XThC.TBN.t113 212.081
R17811 XThC.TBN.n135 XThC.TBN.t99 212.081
R17812 XThC.TBN.n134 XThC.TBN.t96 212.081
R17813 XThC.TBN.n129 XThC.TBN.t58 212.081
R17814 XThC.TBN.n128 XThC.TBN.t51 212.081
R17815 XThC.TBN.n159 XThC.TBN.t13 212.081
R17816 XThC.TBN.n158 XThC.TBN.t7 212.081
R17817 XThC.TBN.n153 XThC.TBN.t86 212.081
R17818 XThC.TBN.n152 XThC.TBN.t81 212.081
R17819 XThC.TBN.n190 XThC.TBN.n189 208.965
R17820 XThC.TBN.n177 XThC.TBN.n0 188.516
R17821 XThC.TBN.n88 XThC.TBN.n87 180.482
R17822 XThC.TBN.n62 XThC.TBN.n61 180.482
R17823 XThC.TBN.n36 XThC.TBN.n35 180.482
R17824 XThC.TBN.n11 XThC.TBN.n10 180.482
R17825 XThC.TBN.n75 XThC.TBN.n74 180.482
R17826 XThC.TBN.n49 XThC.TBN.n48 180.482
R17827 XThC.TBN.n23 XThC.TBN.n22 180.482
R17828 XThC.TBN.n96 XThC.TBN.n95 173.761
R17829 XThC.TBN.n119 XThC.TBN.n118 173.761
R17830 XThC.TBN.n143 XThC.TBN.n142 173.761
R17831 XThC.TBN.n167 XThC.TBN.n166 173.761
R17832 XThC.TBN.n107 XThC.TBN.n106 173.761
R17833 XThC.TBN.n131 XThC.TBN.n130 173.761
R17834 XThC.TBN.n155 XThC.TBN.n154 173.761
R17835 XThC.TBN.n81 XThC.TBN.n79 152
R17836 XThC.TBN.n84 XThC.TBN.n83 152
R17837 XThC.TBN.n86 XThC.TBN.n85 152
R17838 XThC.TBN.n55 XThC.TBN.n53 152
R17839 XThC.TBN.n58 XThC.TBN.n57 152
R17840 XThC.TBN.n60 XThC.TBN.n59 152
R17841 XThC.TBN.n29 XThC.TBN.n27 152
R17842 XThC.TBN.n32 XThC.TBN.n31 152
R17843 XThC.TBN.n34 XThC.TBN.n33 152
R17844 XThC.TBN.n4 XThC.TBN.n2 152
R17845 XThC.TBN.n7 XThC.TBN.n6 152
R17846 XThC.TBN.n9 XThC.TBN.n8 152
R17847 XThC.TBN.n68 XThC.TBN.n66 152
R17848 XThC.TBN.n71 XThC.TBN.n70 152
R17849 XThC.TBN.n73 XThC.TBN.n72 152
R17850 XThC.TBN.n42 XThC.TBN.n40 152
R17851 XThC.TBN.n45 XThC.TBN.n44 152
R17852 XThC.TBN.n47 XThC.TBN.n46 152
R17853 XThC.TBN.n16 XThC.TBN.n14 152
R17854 XThC.TBN.n19 XThC.TBN.n18 152
R17855 XThC.TBN.n21 XThC.TBN.n20 152
R17856 XThC.TBN.n96 XThC.TBN.n92 152
R17857 XThC.TBN.n98 XThC.TBN.n97 152
R17858 XThC.TBN.n102 XThC.TBN.n101 152
R17859 XThC.TBN.n119 XThC.TBN.n115 152
R17860 XThC.TBN.n121 XThC.TBN.n120 152
R17861 XThC.TBN.n125 XThC.TBN.n124 152
R17862 XThC.TBN.n143 XThC.TBN.n139 152
R17863 XThC.TBN.n145 XThC.TBN.n144 152
R17864 XThC.TBN.n149 XThC.TBN.n148 152
R17865 XThC.TBN.n167 XThC.TBN.n163 152
R17866 XThC.TBN.n169 XThC.TBN.n168 152
R17867 XThC.TBN.n173 XThC.TBN.n172 152
R17868 XThC.TBN.n107 XThC.TBN.n103 152
R17869 XThC.TBN.n109 XThC.TBN.n108 152
R17870 XThC.TBN.n113 XThC.TBN.n112 152
R17871 XThC.TBN.n131 XThC.TBN.n127 152
R17872 XThC.TBN.n133 XThC.TBN.n132 152
R17873 XThC.TBN.n137 XThC.TBN.n136 152
R17874 XThC.TBN.n155 XThC.TBN.n151 152
R17875 XThC.TBN.n157 XThC.TBN.n156 152
R17876 XThC.TBN.n161 XThC.TBN.n160 152
R17877 XThC.TBN.n179 XThC.TBN.n178 152
R17878 XThC.TBN.n181 XThC.TBN.n180 152
R17879 XThC.TBN.n185 XThC.TBN.n184 152
R17880 XThC.TBN.n183 XThC.TBN.t14 139.78
R17881 XThC.TBN.n182 XThC.TBN.t105 139.78
R17882 XThC.TBN.n176 XThC.TBN.t69 139.78
R17883 XThC.TBN.n177 XThC.TBN.t61 139.78
R17884 XThC.TBN.n87 XThC.TBN.t123 139.78
R17885 XThC.TBN.n78 XThC.TBN.t85 139.78
R17886 XThC.TBN.n82 XThC.TBN.t74 139.78
R17887 XThC.TBN.n80 XThC.TBN.t65 139.78
R17888 XThC.TBN.n61 XThC.TBN.t31 139.78
R17889 XThC.TBN.n52 XThC.TBN.t104 139.78
R17890 XThC.TBN.n56 XThC.TBN.t94 139.78
R17891 XThC.TBN.n54 XThC.TBN.t92 139.78
R17892 XThC.TBN.n35 XThC.TBN.t89 139.78
R17893 XThC.TBN.n26 XThC.TBN.t41 139.78
R17894 XThC.TBN.n30 XThC.TBN.t35 139.78
R17895 XThC.TBN.n28 XThC.TBN.t32 139.78
R17896 XThC.TBN.n10 XThC.TBN.t118 139.78
R17897 XThC.TBN.n1 XThC.TBN.t83 139.78
R17898 XThC.TBN.n5 XThC.TBN.t71 139.78
R17899 XThC.TBN.n3 XThC.TBN.t62 139.78
R17900 XThC.TBN.n74 XThC.TBN.t107 139.78
R17901 XThC.TBN.n65 XThC.TBN.t72 139.78
R17902 XThC.TBN.n69 XThC.TBN.t57 139.78
R17903 XThC.TBN.n67 XThC.TBN.t49 139.78
R17904 XThC.TBN.n48 XThC.TBN.t43 139.78
R17905 XThC.TBN.n39 XThC.TBN.t10 139.78
R17906 XThC.TBN.n43 XThC.TBN.t112 139.78
R17907 XThC.TBN.n41 XThC.TBN.t108 139.78
R17908 XThC.TBN.n22 XThC.TBN.t121 139.78
R17909 XThC.TBN.n13 XThC.TBN.t84 139.78
R17910 XThC.TBN.n17 XThC.TBN.t73 139.78
R17911 XThC.TBN.n15 XThC.TBN.t64 139.78
R17912 XThC.TBN.n100 XThC.TBN.t76 139.78
R17913 XThC.TBN.n99 XThC.TBN.t67 139.78
R17914 XThC.TBN.n94 XThC.TBN.t29 139.78
R17915 XThC.TBN.n93 XThC.TBN.t24 139.78
R17916 XThC.TBN.n123 XThC.TBN.t15 139.78
R17917 XThC.TBN.n122 XThC.TBN.t8 139.78
R17918 XThC.TBN.n117 XThC.TBN.t87 139.78
R17919 XThC.TBN.n116 XThC.TBN.t82 139.78
R17920 XThC.TBN.n147 XThC.TBN.t66 139.78
R17921 XThC.TBN.n146 XThC.TBN.t60 139.78
R17922 XThC.TBN.n141 XThC.TBN.t22 139.78
R17923 XThC.TBN.n140 XThC.TBN.t20 139.78
R17924 XThC.TBN.n171 XThC.TBN.t4 139.78
R17925 XThC.TBN.n170 XThC.TBN.t117 139.78
R17926 XThC.TBN.n165 XThC.TBN.t80 139.78
R17927 XThC.TBN.n164 XThC.TBN.t78 139.78
R17928 XThC.TBN.n111 XThC.TBN.t59 139.78
R17929 XThC.TBN.n110 XThC.TBN.t55 139.78
R17930 XThC.TBN.n105 XThC.TBN.t19 139.78
R17931 XThC.TBN.n104 XThC.TBN.t16 139.78
R17932 XThC.TBN.n135 XThC.TBN.t115 139.78
R17933 XThC.TBN.n134 XThC.TBN.t110 139.78
R17934 XThC.TBN.n129 XThC.TBN.t77 139.78
R17935 XThC.TBN.n128 XThC.TBN.t68 139.78
R17936 XThC.TBN.n159 XThC.TBN.t53 139.78
R17937 XThC.TBN.n158 XThC.TBN.t45 139.78
R17938 XThC.TBN.n153 XThC.TBN.t11 139.78
R17939 XThC.TBN.n152 XThC.TBN.t5 139.78
R17940 XThC.TBN XThC.TBN.n193 96.8352
R17941 XThC.TBN.n188 XThC.TBN.n0 64.6909
R17942 XThC.TBN.n98 XThC.TBN.n92 49.6611
R17943 XThC.TBN.n121 XThC.TBN.n115 49.6611
R17944 XThC.TBN.n145 XThC.TBN.n139 49.6611
R17945 XThC.TBN.n169 XThC.TBN.n163 49.6611
R17946 XThC.TBN.n109 XThC.TBN.n103 49.6611
R17947 XThC.TBN.n133 XThC.TBN.n127 49.6611
R17948 XThC.TBN.n157 XThC.TBN.n151 49.6611
R17949 XThC.TBN.n101 XThC.TBN.n99 44.549
R17950 XThC.TBN.n124 XThC.TBN.n122 44.549
R17951 XThC.TBN.n148 XThC.TBN.n146 44.549
R17952 XThC.TBN.n172 XThC.TBN.n170 44.549
R17953 XThC.TBN.n112 XThC.TBN.n110 44.549
R17954 XThC.TBN.n136 XThC.TBN.n134 44.549
R17955 XThC.TBN.n160 XThC.TBN.n158 44.549
R17956 XThC.TBN.n95 XThC.TBN.n94 43.0884
R17957 XThC.TBN.n118 XThC.TBN.n117 43.0884
R17958 XThC.TBN.n142 XThC.TBN.n141 43.0884
R17959 XThC.TBN.n166 XThC.TBN.n165 43.0884
R17960 XThC.TBN.n106 XThC.TBN.n105 43.0884
R17961 XThC.TBN.n130 XThC.TBN.n129 43.0884
R17962 XThC.TBN.n154 XThC.TBN.n153 43.0884
R17963 XThC.TBN.n178 XThC.TBN.n177 30.6732
R17964 XThC.TBN.n178 XThC.TBN.n176 30.6732
R17965 XThC.TBN.n181 XThC.TBN.n176 30.6732
R17966 XThC.TBN.n182 XThC.TBN.n181 30.6732
R17967 XThC.TBN.n184 XThC.TBN.n182 30.6732
R17968 XThC.TBN.n184 XThC.TBN.n183 30.6732
R17969 XThC.TBN.n81 XThC.TBN.n80 30.6732
R17970 XThC.TBN.n82 XThC.TBN.n81 30.6732
R17971 XThC.TBN.n83 XThC.TBN.n82 30.6732
R17972 XThC.TBN.n83 XThC.TBN.n78 30.6732
R17973 XThC.TBN.n86 XThC.TBN.n78 30.6732
R17974 XThC.TBN.n87 XThC.TBN.n86 30.6732
R17975 XThC.TBN.n55 XThC.TBN.n54 30.6732
R17976 XThC.TBN.n56 XThC.TBN.n55 30.6732
R17977 XThC.TBN.n57 XThC.TBN.n56 30.6732
R17978 XThC.TBN.n57 XThC.TBN.n52 30.6732
R17979 XThC.TBN.n60 XThC.TBN.n52 30.6732
R17980 XThC.TBN.n61 XThC.TBN.n60 30.6732
R17981 XThC.TBN.n29 XThC.TBN.n28 30.6732
R17982 XThC.TBN.n30 XThC.TBN.n29 30.6732
R17983 XThC.TBN.n31 XThC.TBN.n30 30.6732
R17984 XThC.TBN.n31 XThC.TBN.n26 30.6732
R17985 XThC.TBN.n34 XThC.TBN.n26 30.6732
R17986 XThC.TBN.n35 XThC.TBN.n34 30.6732
R17987 XThC.TBN.n4 XThC.TBN.n3 30.6732
R17988 XThC.TBN.n5 XThC.TBN.n4 30.6732
R17989 XThC.TBN.n6 XThC.TBN.n5 30.6732
R17990 XThC.TBN.n6 XThC.TBN.n1 30.6732
R17991 XThC.TBN.n9 XThC.TBN.n1 30.6732
R17992 XThC.TBN.n10 XThC.TBN.n9 30.6732
R17993 XThC.TBN.n68 XThC.TBN.n67 30.6732
R17994 XThC.TBN.n69 XThC.TBN.n68 30.6732
R17995 XThC.TBN.n70 XThC.TBN.n69 30.6732
R17996 XThC.TBN.n70 XThC.TBN.n65 30.6732
R17997 XThC.TBN.n73 XThC.TBN.n65 30.6732
R17998 XThC.TBN.n74 XThC.TBN.n73 30.6732
R17999 XThC.TBN.n42 XThC.TBN.n41 30.6732
R18000 XThC.TBN.n43 XThC.TBN.n42 30.6732
R18001 XThC.TBN.n44 XThC.TBN.n43 30.6732
R18002 XThC.TBN.n44 XThC.TBN.n39 30.6732
R18003 XThC.TBN.n47 XThC.TBN.n39 30.6732
R18004 XThC.TBN.n48 XThC.TBN.n47 30.6732
R18005 XThC.TBN.n16 XThC.TBN.n15 30.6732
R18006 XThC.TBN.n17 XThC.TBN.n16 30.6732
R18007 XThC.TBN.n18 XThC.TBN.n17 30.6732
R18008 XThC.TBN.n18 XThC.TBN.n13 30.6732
R18009 XThC.TBN.n21 XThC.TBN.n13 30.6732
R18010 XThC.TBN.n22 XThC.TBN.n21 30.6732
R18011 XThC.TBN.n189 XThC.TBN.t2 26.5955
R18012 XThC.TBN.n189 XThC.TBN.t3 26.5955
R18013 XThC.TBN.n193 XThC.TBN.t1 24.9236
R18014 XThC.TBN.n193 XThC.TBN.t0 24.9236
R18015 XThC.TBN.n97 XThC.TBN.n96 21.7605
R18016 XThC.TBN.n120 XThC.TBN.n119 21.7605
R18017 XThC.TBN.n144 XThC.TBN.n143 21.7605
R18018 XThC.TBN.n168 XThC.TBN.n167 21.7605
R18019 XThC.TBN.n108 XThC.TBN.n107 21.7605
R18020 XThC.TBN.n132 XThC.TBN.n131 21.7605
R18021 XThC.TBN.n156 XThC.TBN.n155 21.7605
R18022 XThC.TBN.n84 XThC.TBN.n79 21.5045
R18023 XThC.TBN.n58 XThC.TBN.n53 21.5045
R18024 XThC.TBN.n32 XThC.TBN.n27 21.5045
R18025 XThC.TBN.n7 XThC.TBN.n2 21.5045
R18026 XThC.TBN.n71 XThC.TBN.n66 21.5045
R18027 XThC.TBN.n45 XThC.TBN.n40 21.5045
R18028 XThC.TBN.n19 XThC.TBN.n14 21.5045
R18029 XThC.TBN.n179 XThC.TBN 21.2485
R18030 XThC.TBN.n85 XThC.TBN 19.9685
R18031 XThC.TBN.n59 XThC.TBN 19.9685
R18032 XThC.TBN.n33 XThC.TBN 19.9685
R18033 XThC.TBN.n8 XThC.TBN 19.9685
R18034 XThC.TBN.n72 XThC.TBN 19.9685
R18035 XThC.TBN.n46 XThC.TBN 19.9685
R18036 XThC.TBN.n20 XThC.TBN 19.9685
R18037 XThC.TBN.n180 XThC.TBN 19.2005
R18038 XThC.TBN.n95 XThC.TBN.n93 18.2581
R18039 XThC.TBN.n118 XThC.TBN.n116 18.2581
R18040 XThC.TBN.n142 XThC.TBN.n140 18.2581
R18041 XThC.TBN.n166 XThC.TBN.n164 18.2581
R18042 XThC.TBN.n106 XThC.TBN.n104 18.2581
R18043 XThC.TBN.n130 XThC.TBN.n128 18.2581
R18044 XThC.TBN.n154 XThC.TBN.n152 18.2581
R18045 XThC.TBN.n114 XThC.TBN.n102 17.1655
R18046 XThC.TBN.n88 XThC.TBN 17.1525
R18047 XThC.TBN.n62 XThC.TBN 17.1525
R18048 XThC.TBN.n36 XThC.TBN 17.1525
R18049 XThC.TBN.n11 XThC.TBN 17.1525
R18050 XThC.TBN.n75 XThC.TBN 17.1525
R18051 XThC.TBN.n49 XThC.TBN 17.1525
R18052 XThC.TBN.n23 XThC.TBN 17.1525
R18053 XThC.TBN.n101 XThC.TBN.n100 16.7975
R18054 XThC.TBN.n124 XThC.TBN.n123 16.7975
R18055 XThC.TBN.n148 XThC.TBN.n147 16.7975
R18056 XThC.TBN.n172 XThC.TBN.n171 16.7975
R18057 XThC.TBN.n112 XThC.TBN.n111 16.7975
R18058 XThC.TBN.n136 XThC.TBN.n135 16.7975
R18059 XThC.TBN.n160 XThC.TBN.n159 16.7975
R18060 XThC.TBN.n126 XThC.TBN.n125 16.0405
R18061 XThC.TBN.n150 XThC.TBN.n149 16.0405
R18062 XThC.TBN.n174 XThC.TBN.n173 16.0405
R18063 XThC.TBN.n114 XThC.TBN.n113 16.0405
R18064 XThC.TBN.n138 XThC.TBN.n137 16.0405
R18065 XThC.TBN.n162 XThC.TBN.n161 16.0405
R18066 XThC.TBN.n25 XThC.TBN.n12 15.262
R18067 XThC.TBN.n102 XThC.TBN 15.0405
R18068 XThC.TBN.n125 XThC.TBN 15.0405
R18069 XThC.TBN.n149 XThC.TBN 15.0405
R18070 XThC.TBN.n173 XThC.TBN 15.0405
R18071 XThC.TBN.n113 XThC.TBN 15.0405
R18072 XThC.TBN.n137 XThC.TBN 15.0405
R18073 XThC.TBN.n161 XThC.TBN 15.0405
R18074 XThC.TBN.n90 XThC.TBN.n89 13.8005
R18075 XThC.TBN.n64 XThC.TBN.n63 13.8005
R18076 XThC.TBN.n38 XThC.TBN.n37 13.8005
R18077 XThC.TBN.n77 XThC.TBN.n76 13.8005
R18078 XThC.TBN.n51 XThC.TBN.n50 13.8005
R18079 XThC.TBN.n25 XThC.TBN.n24 13.8005
R18080 XThC.TBN.n191 XThC.TBN 12.5445
R18081 XThC.TBN.n192 XThC.TBN 11.2645
R18082 XThC.TBN.n186 XThC.TBN.n185 9.2165
R18083 XThC.TBN.n186 XThC.TBN 7.9365
R18084 XThC.TBN.n97 XThC.TBN 6.7205
R18085 XThC.TBN.n120 XThC.TBN 6.7205
R18086 XThC.TBN.n144 XThC.TBN 6.7205
R18087 XThC.TBN.n168 XThC.TBN 6.7205
R18088 XThC.TBN.n108 XThC.TBN 6.7205
R18089 XThC.TBN.n132 XThC.TBN 6.7205
R18090 XThC.TBN.n156 XThC.TBN 6.7205
R18091 XThC.TBN.n94 XThC.TBN.n92 6.57323
R18092 XThC.TBN.n117 XThC.TBN.n115 6.57323
R18093 XThC.TBN.n141 XThC.TBN.n139 6.57323
R18094 XThC.TBN.n165 XThC.TBN.n163 6.57323
R18095 XThC.TBN.n105 XThC.TBN.n103 6.57323
R18096 XThC.TBN.n129 XThC.TBN.n127 6.57323
R18097 XThC.TBN.n153 XThC.TBN.n151 6.57323
R18098 XThC.TBN.n185 XThC.TBN 6.4005
R18099 XThC.TBN.n192 XThC.TBN 6.1445
R18100 XThC.TBN.n188 XThC.TBN.n187 5.74665
R18101 XThC.TBN.n187 XThC.TBN.n175 5.68319
R18102 XThC.TBN.n99 XThC.TBN.n98 5.11262
R18103 XThC.TBN.n122 XThC.TBN.n121 5.11262
R18104 XThC.TBN.n146 XThC.TBN.n145 5.11262
R18105 XThC.TBN.n170 XThC.TBN.n169 5.11262
R18106 XThC.TBN.n110 XThC.TBN.n109 5.11262
R18107 XThC.TBN.n134 XThC.TBN.n133 5.11262
R18108 XThC.TBN.n158 XThC.TBN.n157 5.11262
R18109 XThC.TBN.n191 XThC.TBN.n188 5.06717
R18110 XThC.TBN XThC.TBN.n191 4.8645
R18111 XThC.TBN XThC.TBN.n192 4.65505
R18112 XThC.TBN.n187 XThC.TBN.n186 4.6505
R18113 XThC.TBN.n89 XThC.TBN 4.6085
R18114 XThC.TBN.n63 XThC.TBN 4.6085
R18115 XThC.TBN.n37 XThC.TBN 4.6085
R18116 XThC.TBN.n12 XThC.TBN 4.6085
R18117 XThC.TBN.n76 XThC.TBN 4.6085
R18118 XThC.TBN.n50 XThC.TBN 4.6085
R18119 XThC.TBN.n24 XThC.TBN 4.6085
R18120 XThC.TBN.n180 XThC.TBN 4.3525
R18121 XThC.TBN.n85 XThC.TBN 3.5845
R18122 XThC.TBN.n59 XThC.TBN 3.5845
R18123 XThC.TBN.n33 XThC.TBN 3.5845
R18124 XThC.TBN.n8 XThC.TBN 3.5845
R18125 XThC.TBN.n72 XThC.TBN 3.5845
R18126 XThC.TBN.n46 XThC.TBN 3.5845
R18127 XThC.TBN.n20 XThC.TBN 3.5845
R18128 XThC.TBN XThC.TBN.n0 2.3045
R18129 XThC.TBN XThC.TBN.n179 2.3045
R18130 XThC.TBN XThC.TBN.n190 2.0485
R18131 XThC.TBN.n89 XThC.TBN.n88 1.7925
R18132 XThC.TBN.n63 XThC.TBN.n62 1.7925
R18133 XThC.TBN.n37 XThC.TBN.n36 1.7925
R18134 XThC.TBN.n12 XThC.TBN.n11 1.7925
R18135 XThC.TBN.n76 XThC.TBN.n75 1.7925
R18136 XThC.TBN.n50 XThC.TBN.n49 1.7925
R18137 XThC.TBN.n24 XThC.TBN.n23 1.7925
R18138 XThC.TBN.n175 XThC.TBN.n174 1.59665
R18139 XThC.TBN.n190 XThC.TBN 1.55202
R18140 XThC.TBN XThC.TBN.n84 1.5365
R18141 XThC.TBN XThC.TBN.n58 1.5365
R18142 XThC.TBN XThC.TBN.n32 1.5365
R18143 XThC.TBN XThC.TBN.n7 1.5365
R18144 XThC.TBN XThC.TBN.n71 1.5365
R18145 XThC.TBN XThC.TBN.n45 1.5365
R18146 XThC.TBN XThC.TBN.n19 1.5365
R18147 XThC.TBN.n150 XThC.TBN.n138 1.49088
R18148 XThC.TBN.n126 XThC.TBN.n114 1.49088
R18149 XThC.TBN.n174 XThC.TBN.n162 1.48608
R18150 XThC.TBN.n51 XThC.TBN.n38 1.46204
R18151 XThC.TBN.n77 XThC.TBN.n64 1.46204
R18152 XThC.TBN.n38 XThC.TBN.n25 1.15435
R18153 XThC.TBN.n64 XThC.TBN.n51 1.15435
R18154 XThC.TBN.n90 XThC.TBN.n77 1.15435
R18155 XThC.TBN.n162 XThC.TBN.n150 1.13031
R18156 XThC.TBN.n138 XThC.TBN.n126 1.1255
R18157 XThC.TBN.n91 XThC.TBN.n90 1.00531
R18158 XThC.TBN.n79 XThC.TBN 0.5125
R18159 XThC.TBN.n53 XThC.TBN 0.5125
R18160 XThC.TBN.n27 XThC.TBN 0.5125
R18161 XThC.TBN.n2 XThC.TBN 0.5125
R18162 XThC.TBN.n66 XThC.TBN 0.5125
R18163 XThC.TBN.n40 XThC.TBN 0.5125
R18164 XThC.TBN.n14 XThC.TBN 0.5125
R18165 XThC.TBN.n175 XThC.TBN.n91 0.139923
R18166 XThC.TBN.n91 XThC.TBN 0.1255
R18167 XThC.TBN.n91 XThC.TBN 0.063
R18168 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R18169 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R18170 XThC.Tn[6].n71 XThC.Tn[6].n69 161.365
R18171 XThC.Tn[6].n67 XThC.Tn[6].n65 161.365
R18172 XThC.Tn[6].n63 XThC.Tn[6].n61 161.365
R18173 XThC.Tn[6].n59 XThC.Tn[6].n57 161.365
R18174 XThC.Tn[6].n55 XThC.Tn[6].n53 161.365
R18175 XThC.Tn[6].n51 XThC.Tn[6].n49 161.365
R18176 XThC.Tn[6].n47 XThC.Tn[6].n45 161.365
R18177 XThC.Tn[6].n43 XThC.Tn[6].n41 161.365
R18178 XThC.Tn[6].n39 XThC.Tn[6].n37 161.365
R18179 XThC.Tn[6].n35 XThC.Tn[6].n33 161.365
R18180 XThC.Tn[6].n31 XThC.Tn[6].n29 161.365
R18181 XThC.Tn[6].n27 XThC.Tn[6].n25 161.365
R18182 XThC.Tn[6].n23 XThC.Tn[6].n21 161.365
R18183 XThC.Tn[6].n19 XThC.Tn[6].n17 161.365
R18184 XThC.Tn[6].n15 XThC.Tn[6].n13 161.365
R18185 XThC.Tn[6].n12 XThC.Tn[6].n10 161.365
R18186 XThC.Tn[6].n69 XThC.Tn[6].t34 161.202
R18187 XThC.Tn[6].n65 XThC.Tn[6].t24 161.202
R18188 XThC.Tn[6].n61 XThC.Tn[6].t43 161.202
R18189 XThC.Tn[6].n57 XThC.Tn[6].t41 161.202
R18190 XThC.Tn[6].n53 XThC.Tn[6].t32 161.202
R18191 XThC.Tn[6].n49 XThC.Tn[6].t21 161.202
R18192 XThC.Tn[6].n45 XThC.Tn[6].t19 161.202
R18193 XThC.Tn[6].n41 XThC.Tn[6].t31 161.202
R18194 XThC.Tn[6].n37 XThC.Tn[6].t29 161.202
R18195 XThC.Tn[6].n33 XThC.Tn[6].t22 161.202
R18196 XThC.Tn[6].n29 XThC.Tn[6].t38 161.202
R18197 XThC.Tn[6].n25 XThC.Tn[6].t37 161.202
R18198 XThC.Tn[6].n21 XThC.Tn[6].t18 161.202
R18199 XThC.Tn[6].n17 XThC.Tn[6].t17 161.202
R18200 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R18201 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R18202 XThC.Tn[6].n69 XThC.Tn[6].t30 145.137
R18203 XThC.Tn[6].n65 XThC.Tn[6].t20 145.137
R18204 XThC.Tn[6].n61 XThC.Tn[6].t39 145.137
R18205 XThC.Tn[6].n57 XThC.Tn[6].t36 145.137
R18206 XThC.Tn[6].n53 XThC.Tn[6].t28 145.137
R18207 XThC.Tn[6].n49 XThC.Tn[6].t15 145.137
R18208 XThC.Tn[6].n45 XThC.Tn[6].t14 145.137
R18209 XThC.Tn[6].n41 XThC.Tn[6].t27 145.137
R18210 XThC.Tn[6].n37 XThC.Tn[6].t25 145.137
R18211 XThC.Tn[6].n33 XThC.Tn[6].t16 145.137
R18212 XThC.Tn[6].n29 XThC.Tn[6].t35 145.137
R18213 XThC.Tn[6].n25 XThC.Tn[6].t33 145.137
R18214 XThC.Tn[6].n21 XThC.Tn[6].t12 145.137
R18215 XThC.Tn[6].n17 XThC.Tn[6].t42 145.137
R18216 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R18217 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R18218 XThC.Tn[6].n7 XThC.Tn[6].n6 135.248
R18219 XThC.Tn[6].n9 XThC.Tn[6].n3 98.982
R18220 XThC.Tn[6].n8 XThC.Tn[6].n4 98.982
R18221 XThC.Tn[6].n7 XThC.Tn[6].n5 98.982
R18222 XThC.Tn[6].n9 XThC.Tn[6].n8 36.2672
R18223 XThC.Tn[6].n8 XThC.Tn[6].n7 36.2672
R18224 XThC.Tn[6].n73 XThC.Tn[6].n9 32.6405
R18225 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R18226 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R18227 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R18228 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R18229 XThC.Tn[6].n3 XThC.Tn[6].t8 24.9236
R18230 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R18231 XThC.Tn[6].n4 XThC.Tn[6].t10 24.9236
R18232 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R18233 XThC.Tn[6].n5 XThC.Tn[6].t1 24.9236
R18234 XThC.Tn[6].n5 XThC.Tn[6].t0 24.9236
R18235 XThC.Tn[6].n6 XThC.Tn[6].t3 24.9236
R18236 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R18237 XThC.Tn[6].n74 XThC.Tn[6].n2 18.5605
R18238 XThC.Tn[6].n74 XThC.Tn[6].n73 11.5205
R18239 XThC.Tn[6] XThC.Tn[6].n12 8.0245
R18240 XThC.Tn[6].n72 XThC.Tn[6].n71 7.9105
R18241 XThC.Tn[6].n68 XThC.Tn[6].n67 7.9105
R18242 XThC.Tn[6].n64 XThC.Tn[6].n63 7.9105
R18243 XThC.Tn[6].n60 XThC.Tn[6].n59 7.9105
R18244 XThC.Tn[6].n56 XThC.Tn[6].n55 7.9105
R18245 XThC.Tn[6].n52 XThC.Tn[6].n51 7.9105
R18246 XThC.Tn[6].n48 XThC.Tn[6].n47 7.9105
R18247 XThC.Tn[6].n44 XThC.Tn[6].n43 7.9105
R18248 XThC.Tn[6].n40 XThC.Tn[6].n39 7.9105
R18249 XThC.Tn[6].n36 XThC.Tn[6].n35 7.9105
R18250 XThC.Tn[6].n32 XThC.Tn[6].n31 7.9105
R18251 XThC.Tn[6].n28 XThC.Tn[6].n27 7.9105
R18252 XThC.Tn[6].n24 XThC.Tn[6].n23 7.9105
R18253 XThC.Tn[6].n20 XThC.Tn[6].n19 7.9105
R18254 XThC.Tn[6].n16 XThC.Tn[6].n15 7.9105
R18255 XThC.Tn[6].n73 XThC.Tn[6] 5.42203
R18256 XThC.Tn[6] XThC.Tn[6].n74 0.6405
R18257 XThC.Tn[6].n16 XThC.Tn[6] 0.235138
R18258 XThC.Tn[6].n20 XThC.Tn[6] 0.235138
R18259 XThC.Tn[6].n24 XThC.Tn[6] 0.235138
R18260 XThC.Tn[6].n28 XThC.Tn[6] 0.235138
R18261 XThC.Tn[6].n32 XThC.Tn[6] 0.235138
R18262 XThC.Tn[6].n36 XThC.Tn[6] 0.235138
R18263 XThC.Tn[6].n40 XThC.Tn[6] 0.235138
R18264 XThC.Tn[6].n44 XThC.Tn[6] 0.235138
R18265 XThC.Tn[6].n48 XThC.Tn[6] 0.235138
R18266 XThC.Tn[6].n52 XThC.Tn[6] 0.235138
R18267 XThC.Tn[6].n56 XThC.Tn[6] 0.235138
R18268 XThC.Tn[6].n60 XThC.Tn[6] 0.235138
R18269 XThC.Tn[6].n64 XThC.Tn[6] 0.235138
R18270 XThC.Tn[6].n68 XThC.Tn[6] 0.235138
R18271 XThC.Tn[6].n72 XThC.Tn[6] 0.235138
R18272 XThC.Tn[6] XThC.Tn[6].n16 0.114505
R18273 XThC.Tn[6] XThC.Tn[6].n20 0.114505
R18274 XThC.Tn[6] XThC.Tn[6].n24 0.114505
R18275 XThC.Tn[6] XThC.Tn[6].n28 0.114505
R18276 XThC.Tn[6] XThC.Tn[6].n32 0.114505
R18277 XThC.Tn[6] XThC.Tn[6].n36 0.114505
R18278 XThC.Tn[6] XThC.Tn[6].n40 0.114505
R18279 XThC.Tn[6] XThC.Tn[6].n44 0.114505
R18280 XThC.Tn[6] XThC.Tn[6].n48 0.114505
R18281 XThC.Tn[6] XThC.Tn[6].n52 0.114505
R18282 XThC.Tn[6] XThC.Tn[6].n56 0.114505
R18283 XThC.Tn[6] XThC.Tn[6].n60 0.114505
R18284 XThC.Tn[6] XThC.Tn[6].n64 0.114505
R18285 XThC.Tn[6] XThC.Tn[6].n68 0.114505
R18286 XThC.Tn[6] XThC.Tn[6].n72 0.114505
R18287 XThC.Tn[6].n71 XThC.Tn[6].n70 0.0599512
R18288 XThC.Tn[6].n67 XThC.Tn[6].n66 0.0599512
R18289 XThC.Tn[6].n63 XThC.Tn[6].n62 0.0599512
R18290 XThC.Tn[6].n59 XThC.Tn[6].n58 0.0599512
R18291 XThC.Tn[6].n55 XThC.Tn[6].n54 0.0599512
R18292 XThC.Tn[6].n51 XThC.Tn[6].n50 0.0599512
R18293 XThC.Tn[6].n47 XThC.Tn[6].n46 0.0599512
R18294 XThC.Tn[6].n43 XThC.Tn[6].n42 0.0599512
R18295 XThC.Tn[6].n39 XThC.Tn[6].n38 0.0599512
R18296 XThC.Tn[6].n35 XThC.Tn[6].n34 0.0599512
R18297 XThC.Tn[6].n31 XThC.Tn[6].n30 0.0599512
R18298 XThC.Tn[6].n27 XThC.Tn[6].n26 0.0599512
R18299 XThC.Tn[6].n23 XThC.Tn[6].n22 0.0599512
R18300 XThC.Tn[6].n19 XThC.Tn[6].n18 0.0599512
R18301 XThC.Tn[6].n15 XThC.Tn[6].n14 0.0599512
R18302 XThC.Tn[6].n12 XThC.Tn[6].n11 0.0599512
R18303 XThC.Tn[6].n70 XThC.Tn[6] 0.0469286
R18304 XThC.Tn[6].n66 XThC.Tn[6] 0.0469286
R18305 XThC.Tn[6].n62 XThC.Tn[6] 0.0469286
R18306 XThC.Tn[6].n58 XThC.Tn[6] 0.0469286
R18307 XThC.Tn[6].n54 XThC.Tn[6] 0.0469286
R18308 XThC.Tn[6].n50 XThC.Tn[6] 0.0469286
R18309 XThC.Tn[6].n46 XThC.Tn[6] 0.0469286
R18310 XThC.Tn[6].n42 XThC.Tn[6] 0.0469286
R18311 XThC.Tn[6].n38 XThC.Tn[6] 0.0469286
R18312 XThC.Tn[6].n34 XThC.Tn[6] 0.0469286
R18313 XThC.Tn[6].n30 XThC.Tn[6] 0.0469286
R18314 XThC.Tn[6].n26 XThC.Tn[6] 0.0469286
R18315 XThC.Tn[6].n22 XThC.Tn[6] 0.0469286
R18316 XThC.Tn[6].n18 XThC.Tn[6] 0.0469286
R18317 XThC.Tn[6].n14 XThC.Tn[6] 0.0469286
R18318 XThC.Tn[6].n11 XThC.Tn[6] 0.0469286
R18319 XThC.Tn[6].n70 XThC.Tn[6] 0.0401341
R18320 XThC.Tn[6].n66 XThC.Tn[6] 0.0401341
R18321 XThC.Tn[6].n62 XThC.Tn[6] 0.0401341
R18322 XThC.Tn[6].n58 XThC.Tn[6] 0.0401341
R18323 XThC.Tn[6].n54 XThC.Tn[6] 0.0401341
R18324 XThC.Tn[6].n50 XThC.Tn[6] 0.0401341
R18325 XThC.Tn[6].n46 XThC.Tn[6] 0.0401341
R18326 XThC.Tn[6].n42 XThC.Tn[6] 0.0401341
R18327 XThC.Tn[6].n38 XThC.Tn[6] 0.0401341
R18328 XThC.Tn[6].n34 XThC.Tn[6] 0.0401341
R18329 XThC.Tn[6].n30 XThC.Tn[6] 0.0401341
R18330 XThC.Tn[6].n26 XThC.Tn[6] 0.0401341
R18331 XThC.Tn[6].n22 XThC.Tn[6] 0.0401341
R18332 XThC.Tn[6].n18 XThC.Tn[6] 0.0401341
R18333 XThC.Tn[6].n14 XThC.Tn[6] 0.0401341
R18334 XThC.Tn[6].n11 XThC.Tn[6] 0.0401341
R18335 XThR.Tn[9].n87 XThR.Tn[9].n86 256.104
R18336 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R18337 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R18338 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R18339 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R18340 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R18341 XThR.Tn[9] XThR.Tn[9].n78 161.363
R18342 XThR.Tn[9] XThR.Tn[9].n73 161.363
R18343 XThR.Tn[9] XThR.Tn[9].n68 161.363
R18344 XThR.Tn[9] XThR.Tn[9].n63 161.363
R18345 XThR.Tn[9] XThR.Tn[9].n58 161.363
R18346 XThR.Tn[9] XThR.Tn[9].n53 161.363
R18347 XThR.Tn[9] XThR.Tn[9].n48 161.363
R18348 XThR.Tn[9] XThR.Tn[9].n43 161.363
R18349 XThR.Tn[9] XThR.Tn[9].n38 161.363
R18350 XThR.Tn[9] XThR.Tn[9].n33 161.363
R18351 XThR.Tn[9] XThR.Tn[9].n28 161.363
R18352 XThR.Tn[9] XThR.Tn[9].n23 161.363
R18353 XThR.Tn[9] XThR.Tn[9].n18 161.363
R18354 XThR.Tn[9] XThR.Tn[9].n13 161.363
R18355 XThR.Tn[9] XThR.Tn[9].n8 161.363
R18356 XThR.Tn[9] XThR.Tn[9].n6 161.363
R18357 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R18358 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R18359 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R18360 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R18361 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R18362 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R18363 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R18364 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R18365 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R18366 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R18367 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R18368 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R18369 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R18370 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R18371 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R18372 XThR.Tn[9].n78 XThR.Tn[9].t63 161.106
R18373 XThR.Tn[9].n73 XThR.Tn[9].t69 161.106
R18374 XThR.Tn[9].n68 XThR.Tn[9].t47 161.106
R18375 XThR.Tn[9].n63 XThR.Tn[9].t34 161.106
R18376 XThR.Tn[9].n58 XThR.Tn[9].t62 161.106
R18377 XThR.Tn[9].n53 XThR.Tn[9].t24 161.106
R18378 XThR.Tn[9].n48 XThR.Tn[9].t66 161.106
R18379 XThR.Tn[9].n43 XThR.Tn[9].t45 161.106
R18380 XThR.Tn[9].n38 XThR.Tn[9].t32 161.106
R18381 XThR.Tn[9].n33 XThR.Tn[9].t37 161.106
R18382 XThR.Tn[9].n28 XThR.Tn[9].t23 161.106
R18383 XThR.Tn[9].n23 XThR.Tn[9].t46 161.106
R18384 XThR.Tn[9].n18 XThR.Tn[9].t21 161.106
R18385 XThR.Tn[9].n13 XThR.Tn[9].t64 161.106
R18386 XThR.Tn[9].n8 XThR.Tn[9].t28 161.106
R18387 XThR.Tn[9].n6 XThR.Tn[9].t71 161.106
R18388 XThR.Tn[9].n79 XThR.Tn[9].t54 159.978
R18389 XThR.Tn[9].n74 XThR.Tn[9].t61 159.978
R18390 XThR.Tn[9].n69 XThR.Tn[9].t43 159.978
R18391 XThR.Tn[9].n64 XThR.Tn[9].t27 159.978
R18392 XThR.Tn[9].n59 XThR.Tn[9].t52 159.978
R18393 XThR.Tn[9].n54 XThR.Tn[9].t18 159.978
R18394 XThR.Tn[9].n49 XThR.Tn[9].t60 159.978
R18395 XThR.Tn[9].n44 XThR.Tn[9].t40 159.978
R18396 XThR.Tn[9].n39 XThR.Tn[9].t25 159.978
R18397 XThR.Tn[9].n34 XThR.Tn[9].t33 159.978
R18398 XThR.Tn[9].n29 XThR.Tn[9].t16 159.978
R18399 XThR.Tn[9].n24 XThR.Tn[9].t42 159.978
R18400 XThR.Tn[9].n19 XThR.Tn[9].t15 159.978
R18401 XThR.Tn[9].n14 XThR.Tn[9].t59 159.978
R18402 XThR.Tn[9].n9 XThR.Tn[9].t19 159.978
R18403 XThR.Tn[9].n78 XThR.Tn[9].t49 145.038
R18404 XThR.Tn[9].n73 XThR.Tn[9].t14 145.038
R18405 XThR.Tn[9].n68 XThR.Tn[9].t57 145.038
R18406 XThR.Tn[9].n63 XThR.Tn[9].t38 145.038
R18407 XThR.Tn[9].n58 XThR.Tn[9].t70 145.038
R18408 XThR.Tn[9].n53 XThR.Tn[9].t48 145.038
R18409 XThR.Tn[9].n48 XThR.Tn[9].t58 145.038
R18410 XThR.Tn[9].n43 XThR.Tn[9].t39 145.038
R18411 XThR.Tn[9].n38 XThR.Tn[9].t36 145.038
R18412 XThR.Tn[9].n33 XThR.Tn[9].t67 145.038
R18413 XThR.Tn[9].n28 XThR.Tn[9].t31 145.038
R18414 XThR.Tn[9].n23 XThR.Tn[9].t56 145.038
R18415 XThR.Tn[9].n18 XThR.Tn[9].t29 145.038
R18416 XThR.Tn[9].n13 XThR.Tn[9].t72 145.038
R18417 XThR.Tn[9].n8 XThR.Tn[9].t35 145.038
R18418 XThR.Tn[9].n6 XThR.Tn[9].t17 145.038
R18419 XThR.Tn[9].n79 XThR.Tn[9].t68 143.911
R18420 XThR.Tn[9].n74 XThR.Tn[9].t30 143.911
R18421 XThR.Tn[9].n69 XThR.Tn[9].t12 143.911
R18422 XThR.Tn[9].n64 XThR.Tn[9].t53 143.911
R18423 XThR.Tn[9].n59 XThR.Tn[9].t22 143.911
R18424 XThR.Tn[9].n54 XThR.Tn[9].t65 143.911
R18425 XThR.Tn[9].n49 XThR.Tn[9].t13 143.911
R18426 XThR.Tn[9].n44 XThR.Tn[9].t55 143.911
R18427 XThR.Tn[9].n39 XThR.Tn[9].t51 143.911
R18428 XThR.Tn[9].n34 XThR.Tn[9].t20 143.911
R18429 XThR.Tn[9].n29 XThR.Tn[9].t44 143.911
R18430 XThR.Tn[9].n24 XThR.Tn[9].t73 143.911
R18431 XThR.Tn[9].n19 XThR.Tn[9].t41 143.911
R18432 XThR.Tn[9].n14 XThR.Tn[9].t26 143.911
R18433 XThR.Tn[9].n9 XThR.Tn[9].t50 143.911
R18434 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R18435 XThR.Tn[9].n0 XThR.Tn[9].t2 26.5955
R18436 XThR.Tn[9].n0 XThR.Tn[9].t0 26.5955
R18437 XThR.Tn[9].n85 XThR.Tn[9].t10 26.5955
R18438 XThR.Tn[9].n85 XThR.Tn[9].t8 26.5955
R18439 XThR.Tn[9].n86 XThR.Tn[9].t11 26.5955
R18440 XThR.Tn[9].n86 XThR.Tn[9].t9 26.5955
R18441 XThR.Tn[9].n1 XThR.Tn[9].t3 26.5955
R18442 XThR.Tn[9].n1 XThR.Tn[9].t1 26.5955
R18443 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R18444 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R18445 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R18446 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R18447 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R18448 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R18449 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R18450 XThR.Tn[9] XThR.Tn[9].n7 5.34038
R18451 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R18452 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R18453 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R18454 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R18455 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R18456 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R18457 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R18458 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R18459 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R18460 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R18461 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R18462 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R18463 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R18464 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R18465 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R18466 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R18467 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R18468 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R18469 XThR.Tn[9].n12 XThR.Tn[9] 2.52282
R18470 XThR.Tn[9].n17 XThR.Tn[9] 2.52282
R18471 XThR.Tn[9].n22 XThR.Tn[9] 2.52282
R18472 XThR.Tn[9].n27 XThR.Tn[9] 2.52282
R18473 XThR.Tn[9].n32 XThR.Tn[9] 2.52282
R18474 XThR.Tn[9].n37 XThR.Tn[9] 2.52282
R18475 XThR.Tn[9].n42 XThR.Tn[9] 2.52282
R18476 XThR.Tn[9].n47 XThR.Tn[9] 2.52282
R18477 XThR.Tn[9].n52 XThR.Tn[9] 2.52282
R18478 XThR.Tn[9].n57 XThR.Tn[9] 2.52282
R18479 XThR.Tn[9].n62 XThR.Tn[9] 2.52282
R18480 XThR.Tn[9].n67 XThR.Tn[9] 2.52282
R18481 XThR.Tn[9].n72 XThR.Tn[9] 2.52282
R18482 XThR.Tn[9].n77 XThR.Tn[9] 2.52282
R18483 XThR.Tn[9].n82 XThR.Tn[9] 2.52282
R18484 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R18485 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R18486 XThR.Tn[9].n80 XThR.Tn[9] 1.08677
R18487 XThR.Tn[9].n75 XThR.Tn[9] 1.08677
R18488 XThR.Tn[9].n70 XThR.Tn[9] 1.08677
R18489 XThR.Tn[9].n65 XThR.Tn[9] 1.08677
R18490 XThR.Tn[9].n60 XThR.Tn[9] 1.08677
R18491 XThR.Tn[9].n55 XThR.Tn[9] 1.08677
R18492 XThR.Tn[9].n50 XThR.Tn[9] 1.08677
R18493 XThR.Tn[9].n45 XThR.Tn[9] 1.08677
R18494 XThR.Tn[9].n40 XThR.Tn[9] 1.08677
R18495 XThR.Tn[9].n35 XThR.Tn[9] 1.08677
R18496 XThR.Tn[9].n30 XThR.Tn[9] 1.08677
R18497 XThR.Tn[9].n25 XThR.Tn[9] 1.08677
R18498 XThR.Tn[9].n20 XThR.Tn[9] 1.08677
R18499 XThR.Tn[9].n15 XThR.Tn[9] 1.08677
R18500 XThR.Tn[9].n10 XThR.Tn[9] 1.08677
R18501 XThR.Tn[9] XThR.Tn[9].n12 0.839786
R18502 XThR.Tn[9] XThR.Tn[9].n17 0.839786
R18503 XThR.Tn[9] XThR.Tn[9].n22 0.839786
R18504 XThR.Tn[9] XThR.Tn[9].n27 0.839786
R18505 XThR.Tn[9] XThR.Tn[9].n32 0.839786
R18506 XThR.Tn[9] XThR.Tn[9].n37 0.839786
R18507 XThR.Tn[9] XThR.Tn[9].n42 0.839786
R18508 XThR.Tn[9] XThR.Tn[9].n47 0.839786
R18509 XThR.Tn[9] XThR.Tn[9].n52 0.839786
R18510 XThR.Tn[9] XThR.Tn[9].n57 0.839786
R18511 XThR.Tn[9] XThR.Tn[9].n62 0.839786
R18512 XThR.Tn[9] XThR.Tn[9].n67 0.839786
R18513 XThR.Tn[9] XThR.Tn[9].n72 0.839786
R18514 XThR.Tn[9] XThR.Tn[9].n77 0.839786
R18515 XThR.Tn[9] XThR.Tn[9].n82 0.839786
R18516 XThR.Tn[9].n7 XThR.Tn[9] 0.499542
R18517 XThR.Tn[9].n81 XThR.Tn[9] 0.063
R18518 XThR.Tn[9].n76 XThR.Tn[9] 0.063
R18519 XThR.Tn[9].n71 XThR.Tn[9] 0.063
R18520 XThR.Tn[9].n66 XThR.Tn[9] 0.063
R18521 XThR.Tn[9].n61 XThR.Tn[9] 0.063
R18522 XThR.Tn[9].n56 XThR.Tn[9] 0.063
R18523 XThR.Tn[9].n51 XThR.Tn[9] 0.063
R18524 XThR.Tn[9].n46 XThR.Tn[9] 0.063
R18525 XThR.Tn[9].n41 XThR.Tn[9] 0.063
R18526 XThR.Tn[9].n36 XThR.Tn[9] 0.063
R18527 XThR.Tn[9].n31 XThR.Tn[9] 0.063
R18528 XThR.Tn[9].n26 XThR.Tn[9] 0.063
R18529 XThR.Tn[9].n21 XThR.Tn[9] 0.063
R18530 XThR.Tn[9].n16 XThR.Tn[9] 0.063
R18531 XThR.Tn[9].n11 XThR.Tn[9] 0.063
R18532 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R18533 XThR.Tn[9] XThR.Tn[9].n83 0.038
R18534 XThR.Tn[9].n7 XThR.Tn[9] 0.0143889
R18535 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00771154
R18536 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00771154
R18537 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00771154
R18538 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00771154
R18539 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00771154
R18540 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00771154
R18541 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00771154
R18542 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00771154
R18543 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00771154
R18544 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00771154
R18545 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00771154
R18546 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00771154
R18547 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00771154
R18548 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00771154
R18549 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00771154
R18550 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18551 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18552 XThC.Tn[5].n71 XThC.Tn[5].n69 161.365
R18553 XThC.Tn[5].n67 XThC.Tn[5].n65 161.365
R18554 XThC.Tn[5].n63 XThC.Tn[5].n61 161.365
R18555 XThC.Tn[5].n59 XThC.Tn[5].n57 161.365
R18556 XThC.Tn[5].n55 XThC.Tn[5].n53 161.365
R18557 XThC.Tn[5].n51 XThC.Tn[5].n49 161.365
R18558 XThC.Tn[5].n47 XThC.Tn[5].n45 161.365
R18559 XThC.Tn[5].n43 XThC.Tn[5].n41 161.365
R18560 XThC.Tn[5].n39 XThC.Tn[5].n37 161.365
R18561 XThC.Tn[5].n35 XThC.Tn[5].n33 161.365
R18562 XThC.Tn[5].n31 XThC.Tn[5].n29 161.365
R18563 XThC.Tn[5].n27 XThC.Tn[5].n25 161.365
R18564 XThC.Tn[5].n23 XThC.Tn[5].n21 161.365
R18565 XThC.Tn[5].n19 XThC.Tn[5].n17 161.365
R18566 XThC.Tn[5].n15 XThC.Tn[5].n13 161.365
R18567 XThC.Tn[5].n12 XThC.Tn[5].n10 161.365
R18568 XThC.Tn[5].n69 XThC.Tn[5].t41 161.202
R18569 XThC.Tn[5].n65 XThC.Tn[5].t30 161.202
R18570 XThC.Tn[5].n61 XThC.Tn[5].t18 161.202
R18571 XThC.Tn[5].n57 XThC.Tn[5].t16 161.202
R18572 XThC.Tn[5].n53 XThC.Tn[5].t39 161.202
R18573 XThC.Tn[5].n49 XThC.Tn[5].t26 161.202
R18574 XThC.Tn[5].n45 XThC.Tn[5].t25 161.202
R18575 XThC.Tn[5].n41 XThC.Tn[5].t37 161.202
R18576 XThC.Tn[5].n37 XThC.Tn[5].t35 161.202
R18577 XThC.Tn[5].n33 XThC.Tn[5].t27 161.202
R18578 XThC.Tn[5].n29 XThC.Tn[5].t14 161.202
R18579 XThC.Tn[5].n25 XThC.Tn[5].t13 161.202
R18580 XThC.Tn[5].n21 XThC.Tn[5].t24 161.202
R18581 XThC.Tn[5].n17 XThC.Tn[5].t23 161.202
R18582 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18583 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18584 XThC.Tn[5].n69 XThC.Tn[5].t22 145.137
R18585 XThC.Tn[5].n65 XThC.Tn[5].t12 145.137
R18586 XThC.Tn[5].n61 XThC.Tn[5].t32 145.137
R18587 XThC.Tn[5].n57 XThC.Tn[5].t31 145.137
R18588 XThC.Tn[5].n53 XThC.Tn[5].t21 145.137
R18589 XThC.Tn[5].n49 XThC.Tn[5].t42 145.137
R18590 XThC.Tn[5].n45 XThC.Tn[5].t40 145.137
R18591 XThC.Tn[5].n41 XThC.Tn[5].t20 145.137
R18592 XThC.Tn[5].n37 XThC.Tn[5].t17 145.137
R18593 XThC.Tn[5].n33 XThC.Tn[5].t43 145.137
R18594 XThC.Tn[5].n29 XThC.Tn[5].t29 145.137
R18595 XThC.Tn[5].n25 XThC.Tn[5].t28 145.137
R18596 XThC.Tn[5].n21 XThC.Tn[5].t38 145.137
R18597 XThC.Tn[5].n17 XThC.Tn[5].t36 145.137
R18598 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18599 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18600 XThC.Tn[5].n7 XThC.Tn[5].n6 135.249
R18601 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18602 XThC.Tn[5].n8 XThC.Tn[5].n4 98.981
R18603 XThC.Tn[5].n7 XThC.Tn[5].n5 98.981
R18604 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18605 XThC.Tn[5].n8 XThC.Tn[5].n7 36.2672
R18606 XThC.Tn[5].n73 XThC.Tn[5].n9 32.6405
R18607 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R18608 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R18609 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R18610 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R18611 XThC.Tn[5].n3 XThC.Tn[5].t9 24.9236
R18612 XThC.Tn[5].n3 XThC.Tn[5].t8 24.9236
R18613 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R18614 XThC.Tn[5].n4 XThC.Tn[5].t10 24.9236
R18615 XThC.Tn[5].n5 XThC.Tn[5].t2 24.9236
R18616 XThC.Tn[5].n5 XThC.Tn[5].t1 24.9236
R18617 XThC.Tn[5].n6 XThC.Tn[5].t0 24.9236
R18618 XThC.Tn[5].n6 XThC.Tn[5].t3 24.9236
R18619 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18620 XThC.Tn[5] XThC.Tn[5].n12 8.0245
R18621 XThC.Tn[5].n72 XThC.Tn[5].n71 7.9105
R18622 XThC.Tn[5].n68 XThC.Tn[5].n67 7.9105
R18623 XThC.Tn[5].n64 XThC.Tn[5].n63 7.9105
R18624 XThC.Tn[5].n60 XThC.Tn[5].n59 7.9105
R18625 XThC.Tn[5].n56 XThC.Tn[5].n55 7.9105
R18626 XThC.Tn[5].n52 XThC.Tn[5].n51 7.9105
R18627 XThC.Tn[5].n48 XThC.Tn[5].n47 7.9105
R18628 XThC.Tn[5].n44 XThC.Tn[5].n43 7.9105
R18629 XThC.Tn[5].n40 XThC.Tn[5].n39 7.9105
R18630 XThC.Tn[5].n36 XThC.Tn[5].n35 7.9105
R18631 XThC.Tn[5].n32 XThC.Tn[5].n31 7.9105
R18632 XThC.Tn[5].n28 XThC.Tn[5].n27 7.9105
R18633 XThC.Tn[5].n24 XThC.Tn[5].n23 7.9105
R18634 XThC.Tn[5].n20 XThC.Tn[5].n19 7.9105
R18635 XThC.Tn[5].n16 XThC.Tn[5].n15 7.9105
R18636 XThC.Tn[5] XThC.Tn[5].n73 6.7205
R18637 XThC.Tn[5].n73 XThC.Tn[5] 5.69842
R18638 XThC.Tn[5].n16 XThC.Tn[5] 0.235138
R18639 XThC.Tn[5].n20 XThC.Tn[5] 0.235138
R18640 XThC.Tn[5].n24 XThC.Tn[5] 0.235138
R18641 XThC.Tn[5].n28 XThC.Tn[5] 0.235138
R18642 XThC.Tn[5].n32 XThC.Tn[5] 0.235138
R18643 XThC.Tn[5].n36 XThC.Tn[5] 0.235138
R18644 XThC.Tn[5].n40 XThC.Tn[5] 0.235138
R18645 XThC.Tn[5].n44 XThC.Tn[5] 0.235138
R18646 XThC.Tn[5].n48 XThC.Tn[5] 0.235138
R18647 XThC.Tn[5].n52 XThC.Tn[5] 0.235138
R18648 XThC.Tn[5].n56 XThC.Tn[5] 0.235138
R18649 XThC.Tn[5].n60 XThC.Tn[5] 0.235138
R18650 XThC.Tn[5].n64 XThC.Tn[5] 0.235138
R18651 XThC.Tn[5].n68 XThC.Tn[5] 0.235138
R18652 XThC.Tn[5].n72 XThC.Tn[5] 0.235138
R18653 XThC.Tn[5] XThC.Tn[5].n16 0.114505
R18654 XThC.Tn[5] XThC.Tn[5].n20 0.114505
R18655 XThC.Tn[5] XThC.Tn[5].n24 0.114505
R18656 XThC.Tn[5] XThC.Tn[5].n28 0.114505
R18657 XThC.Tn[5] XThC.Tn[5].n32 0.114505
R18658 XThC.Tn[5] XThC.Tn[5].n36 0.114505
R18659 XThC.Tn[5] XThC.Tn[5].n40 0.114505
R18660 XThC.Tn[5] XThC.Tn[5].n44 0.114505
R18661 XThC.Tn[5] XThC.Tn[5].n48 0.114505
R18662 XThC.Tn[5] XThC.Tn[5].n52 0.114505
R18663 XThC.Tn[5] XThC.Tn[5].n56 0.114505
R18664 XThC.Tn[5] XThC.Tn[5].n60 0.114505
R18665 XThC.Tn[5] XThC.Tn[5].n64 0.114505
R18666 XThC.Tn[5] XThC.Tn[5].n68 0.114505
R18667 XThC.Tn[5] XThC.Tn[5].n72 0.114505
R18668 XThC.Tn[5].n71 XThC.Tn[5].n70 0.0599512
R18669 XThC.Tn[5].n67 XThC.Tn[5].n66 0.0599512
R18670 XThC.Tn[5].n63 XThC.Tn[5].n62 0.0599512
R18671 XThC.Tn[5].n59 XThC.Tn[5].n58 0.0599512
R18672 XThC.Tn[5].n55 XThC.Tn[5].n54 0.0599512
R18673 XThC.Tn[5].n51 XThC.Tn[5].n50 0.0599512
R18674 XThC.Tn[5].n47 XThC.Tn[5].n46 0.0599512
R18675 XThC.Tn[5].n43 XThC.Tn[5].n42 0.0599512
R18676 XThC.Tn[5].n39 XThC.Tn[5].n38 0.0599512
R18677 XThC.Tn[5].n35 XThC.Tn[5].n34 0.0599512
R18678 XThC.Tn[5].n31 XThC.Tn[5].n30 0.0599512
R18679 XThC.Tn[5].n27 XThC.Tn[5].n26 0.0599512
R18680 XThC.Tn[5].n23 XThC.Tn[5].n22 0.0599512
R18681 XThC.Tn[5].n19 XThC.Tn[5].n18 0.0599512
R18682 XThC.Tn[5].n15 XThC.Tn[5].n14 0.0599512
R18683 XThC.Tn[5].n12 XThC.Tn[5].n11 0.0599512
R18684 XThC.Tn[5].n70 XThC.Tn[5] 0.0469286
R18685 XThC.Tn[5].n66 XThC.Tn[5] 0.0469286
R18686 XThC.Tn[5].n62 XThC.Tn[5] 0.0469286
R18687 XThC.Tn[5].n58 XThC.Tn[5] 0.0469286
R18688 XThC.Tn[5].n54 XThC.Tn[5] 0.0469286
R18689 XThC.Tn[5].n50 XThC.Tn[5] 0.0469286
R18690 XThC.Tn[5].n46 XThC.Tn[5] 0.0469286
R18691 XThC.Tn[5].n42 XThC.Tn[5] 0.0469286
R18692 XThC.Tn[5].n38 XThC.Tn[5] 0.0469286
R18693 XThC.Tn[5].n34 XThC.Tn[5] 0.0469286
R18694 XThC.Tn[5].n30 XThC.Tn[5] 0.0469286
R18695 XThC.Tn[5].n26 XThC.Tn[5] 0.0469286
R18696 XThC.Tn[5].n22 XThC.Tn[5] 0.0469286
R18697 XThC.Tn[5].n18 XThC.Tn[5] 0.0469286
R18698 XThC.Tn[5].n14 XThC.Tn[5] 0.0469286
R18699 XThC.Tn[5].n11 XThC.Tn[5] 0.0469286
R18700 XThC.Tn[5].n70 XThC.Tn[5] 0.0401341
R18701 XThC.Tn[5].n66 XThC.Tn[5] 0.0401341
R18702 XThC.Tn[5].n62 XThC.Tn[5] 0.0401341
R18703 XThC.Tn[5].n58 XThC.Tn[5] 0.0401341
R18704 XThC.Tn[5].n54 XThC.Tn[5] 0.0401341
R18705 XThC.Tn[5].n50 XThC.Tn[5] 0.0401341
R18706 XThC.Tn[5].n46 XThC.Tn[5] 0.0401341
R18707 XThC.Tn[5].n42 XThC.Tn[5] 0.0401341
R18708 XThC.Tn[5].n38 XThC.Tn[5] 0.0401341
R18709 XThC.Tn[5].n34 XThC.Tn[5] 0.0401341
R18710 XThC.Tn[5].n30 XThC.Tn[5] 0.0401341
R18711 XThC.Tn[5].n26 XThC.Tn[5] 0.0401341
R18712 XThC.Tn[5].n22 XThC.Tn[5] 0.0401341
R18713 XThC.Tn[5].n18 XThC.Tn[5] 0.0401341
R18714 XThC.Tn[5].n14 XThC.Tn[5] 0.0401341
R18715 XThC.Tn[5].n11 XThC.Tn[5] 0.0401341
R18716 XThC.Tn[9].n2 XThC.Tn[9].n1 265.341
R18717 XThC.Tn[9].n5 XThC.Tn[9].n3 243.68
R18718 XThC.Tn[9].n74 XThC.Tn[9].n72 241.847
R18719 XThC.Tn[9].n5 XThC.Tn[9].n4 205.28
R18720 XThC.Tn[9].n2 XThC.Tn[9].n0 202.094
R18721 XThC.Tn[9].n74 XThC.Tn[9].n73 185
R18722 XThC.Tn[9].n68 XThC.Tn[9].n66 161.365
R18723 XThC.Tn[9].n64 XThC.Tn[9].n62 161.365
R18724 XThC.Tn[9].n60 XThC.Tn[9].n58 161.365
R18725 XThC.Tn[9].n56 XThC.Tn[9].n54 161.365
R18726 XThC.Tn[9].n52 XThC.Tn[9].n50 161.365
R18727 XThC.Tn[9].n48 XThC.Tn[9].n46 161.365
R18728 XThC.Tn[9].n44 XThC.Tn[9].n42 161.365
R18729 XThC.Tn[9].n40 XThC.Tn[9].n38 161.365
R18730 XThC.Tn[9].n36 XThC.Tn[9].n34 161.365
R18731 XThC.Tn[9].n32 XThC.Tn[9].n30 161.365
R18732 XThC.Tn[9].n28 XThC.Tn[9].n26 161.365
R18733 XThC.Tn[9].n24 XThC.Tn[9].n22 161.365
R18734 XThC.Tn[9].n20 XThC.Tn[9].n18 161.365
R18735 XThC.Tn[9].n16 XThC.Tn[9].n14 161.365
R18736 XThC.Tn[9].n12 XThC.Tn[9].n10 161.365
R18737 XThC.Tn[9].n9 XThC.Tn[9].n7 161.365
R18738 XThC.Tn[9].n66 XThC.Tn[9].t20 161.202
R18739 XThC.Tn[9].n62 XThC.Tn[9].t41 161.202
R18740 XThC.Tn[9].n58 XThC.Tn[9].t29 161.202
R18741 XThC.Tn[9].n54 XThC.Tn[9].t27 161.202
R18742 XThC.Tn[9].n50 XThC.Tn[9].t18 161.202
R18743 XThC.Tn[9].n46 XThC.Tn[9].t37 161.202
R18744 XThC.Tn[9].n42 XThC.Tn[9].t36 161.202
R18745 XThC.Tn[9].n38 XThC.Tn[9].t16 161.202
R18746 XThC.Tn[9].n34 XThC.Tn[9].t14 161.202
R18747 XThC.Tn[9].n30 XThC.Tn[9].t38 161.202
R18748 XThC.Tn[9].n26 XThC.Tn[9].t25 161.202
R18749 XThC.Tn[9].n22 XThC.Tn[9].t24 161.202
R18750 XThC.Tn[9].n18 XThC.Tn[9].t35 161.202
R18751 XThC.Tn[9].n14 XThC.Tn[9].t34 161.202
R18752 XThC.Tn[9].n10 XThC.Tn[9].t30 161.202
R18753 XThC.Tn[9].n7 XThC.Tn[9].t12 161.202
R18754 XThC.Tn[9].n66 XThC.Tn[9].t33 145.137
R18755 XThC.Tn[9].n62 XThC.Tn[9].t23 145.137
R18756 XThC.Tn[9].n58 XThC.Tn[9].t43 145.137
R18757 XThC.Tn[9].n54 XThC.Tn[9].t42 145.137
R18758 XThC.Tn[9].n50 XThC.Tn[9].t32 145.137
R18759 XThC.Tn[9].n46 XThC.Tn[9].t21 145.137
R18760 XThC.Tn[9].n42 XThC.Tn[9].t19 145.137
R18761 XThC.Tn[9].n38 XThC.Tn[9].t31 145.137
R18762 XThC.Tn[9].n34 XThC.Tn[9].t28 145.137
R18763 XThC.Tn[9].n30 XThC.Tn[9].t22 145.137
R18764 XThC.Tn[9].n26 XThC.Tn[9].t40 145.137
R18765 XThC.Tn[9].n22 XThC.Tn[9].t39 145.137
R18766 XThC.Tn[9].n18 XThC.Tn[9].t17 145.137
R18767 XThC.Tn[9].n14 XThC.Tn[9].t15 145.137
R18768 XThC.Tn[9].n10 XThC.Tn[9].t13 145.137
R18769 XThC.Tn[9].n7 XThC.Tn[9].t26 145.137
R18770 XThC.Tn[9].n1 XThC.Tn[9].t6 26.5955
R18771 XThC.Tn[9].n1 XThC.Tn[9].t5 26.5955
R18772 XThC.Tn[9].n0 XThC.Tn[9].t4 26.5955
R18773 XThC.Tn[9].n0 XThC.Tn[9].t7 26.5955
R18774 XThC.Tn[9].n3 XThC.Tn[9].t9 26.5955
R18775 XThC.Tn[9].n3 XThC.Tn[9].t8 26.5955
R18776 XThC.Tn[9].n4 XThC.Tn[9].t11 26.5955
R18777 XThC.Tn[9].n4 XThC.Tn[9].t10 26.5955
R18778 XThC.Tn[9].n72 XThC.Tn[9].t1 24.9236
R18779 XThC.Tn[9].n72 XThC.Tn[9].t0 24.9236
R18780 XThC.Tn[9].n73 XThC.Tn[9].t2 24.9236
R18781 XThC.Tn[9].n73 XThC.Tn[9].t3 24.9236
R18782 XThC.Tn[9] XThC.Tn[9].n5 22.9652
R18783 XThC.Tn[9] XThC.Tn[9].n74 18.8943
R18784 XThC.Tn[9].n6 XThC.Tn[9].n2 13.9299
R18785 XThC.Tn[9].n6 XThC.Tn[9] 13.9299
R18786 XThC.Tn[9] XThC.Tn[9].n9 8.0245
R18787 XThC.Tn[9].n69 XThC.Tn[9].n68 7.9105
R18788 XThC.Tn[9].n65 XThC.Tn[9].n64 7.9105
R18789 XThC.Tn[9].n61 XThC.Tn[9].n60 7.9105
R18790 XThC.Tn[9].n57 XThC.Tn[9].n56 7.9105
R18791 XThC.Tn[9].n53 XThC.Tn[9].n52 7.9105
R18792 XThC.Tn[9].n49 XThC.Tn[9].n48 7.9105
R18793 XThC.Tn[9].n45 XThC.Tn[9].n44 7.9105
R18794 XThC.Tn[9].n41 XThC.Tn[9].n40 7.9105
R18795 XThC.Tn[9].n37 XThC.Tn[9].n36 7.9105
R18796 XThC.Tn[9].n33 XThC.Tn[9].n32 7.9105
R18797 XThC.Tn[9].n29 XThC.Tn[9].n28 7.9105
R18798 XThC.Tn[9].n25 XThC.Tn[9].n24 7.9105
R18799 XThC.Tn[9].n21 XThC.Tn[9].n20 7.9105
R18800 XThC.Tn[9].n17 XThC.Tn[9].n16 7.9105
R18801 XThC.Tn[9].n13 XThC.Tn[9].n12 7.9105
R18802 XThC.Tn[9].n71 XThC.Tn[9].n70 7.44831
R18803 XThC.Tn[9] XThC.Tn[9].n71 6.34069
R18804 XThC.Tn[9].n70 XThC.Tn[9] 4.25199
R18805 XThC.Tn[9].n71 XThC.Tn[9] 1.79489
R18806 XThC.Tn[9] XThC.Tn[9].n6 1.19676
R18807 XThC.Tn[9].n70 XThC.Tn[9] 0.657022
R18808 XThC.Tn[9].n13 XThC.Tn[9] 0.235138
R18809 XThC.Tn[9].n17 XThC.Tn[9] 0.235138
R18810 XThC.Tn[9].n21 XThC.Tn[9] 0.235138
R18811 XThC.Tn[9].n25 XThC.Tn[9] 0.235138
R18812 XThC.Tn[9].n29 XThC.Tn[9] 0.235138
R18813 XThC.Tn[9].n33 XThC.Tn[9] 0.235138
R18814 XThC.Tn[9].n37 XThC.Tn[9] 0.235138
R18815 XThC.Tn[9].n41 XThC.Tn[9] 0.235138
R18816 XThC.Tn[9].n45 XThC.Tn[9] 0.235138
R18817 XThC.Tn[9].n49 XThC.Tn[9] 0.235138
R18818 XThC.Tn[9].n53 XThC.Tn[9] 0.235138
R18819 XThC.Tn[9].n57 XThC.Tn[9] 0.235138
R18820 XThC.Tn[9].n61 XThC.Tn[9] 0.235138
R18821 XThC.Tn[9].n65 XThC.Tn[9] 0.235138
R18822 XThC.Tn[9].n69 XThC.Tn[9] 0.235138
R18823 XThC.Tn[9] XThC.Tn[9].n13 0.114505
R18824 XThC.Tn[9] XThC.Tn[9].n17 0.114505
R18825 XThC.Tn[9] XThC.Tn[9].n21 0.114505
R18826 XThC.Tn[9] XThC.Tn[9].n25 0.114505
R18827 XThC.Tn[9] XThC.Tn[9].n29 0.114505
R18828 XThC.Tn[9] XThC.Tn[9].n33 0.114505
R18829 XThC.Tn[9] XThC.Tn[9].n37 0.114505
R18830 XThC.Tn[9] XThC.Tn[9].n41 0.114505
R18831 XThC.Tn[9] XThC.Tn[9].n45 0.114505
R18832 XThC.Tn[9] XThC.Tn[9].n49 0.114505
R18833 XThC.Tn[9] XThC.Tn[9].n53 0.114505
R18834 XThC.Tn[9] XThC.Tn[9].n57 0.114505
R18835 XThC.Tn[9] XThC.Tn[9].n61 0.114505
R18836 XThC.Tn[9] XThC.Tn[9].n65 0.114505
R18837 XThC.Tn[9] XThC.Tn[9].n69 0.114505
R18838 XThC.Tn[9].n68 XThC.Tn[9].n67 0.0599512
R18839 XThC.Tn[9].n64 XThC.Tn[9].n63 0.0599512
R18840 XThC.Tn[9].n60 XThC.Tn[9].n59 0.0599512
R18841 XThC.Tn[9].n56 XThC.Tn[9].n55 0.0599512
R18842 XThC.Tn[9].n52 XThC.Tn[9].n51 0.0599512
R18843 XThC.Tn[9].n48 XThC.Tn[9].n47 0.0599512
R18844 XThC.Tn[9].n44 XThC.Tn[9].n43 0.0599512
R18845 XThC.Tn[9].n40 XThC.Tn[9].n39 0.0599512
R18846 XThC.Tn[9].n36 XThC.Tn[9].n35 0.0599512
R18847 XThC.Tn[9].n32 XThC.Tn[9].n31 0.0599512
R18848 XThC.Tn[9].n28 XThC.Tn[9].n27 0.0599512
R18849 XThC.Tn[9].n24 XThC.Tn[9].n23 0.0599512
R18850 XThC.Tn[9].n20 XThC.Tn[9].n19 0.0599512
R18851 XThC.Tn[9].n16 XThC.Tn[9].n15 0.0599512
R18852 XThC.Tn[9].n12 XThC.Tn[9].n11 0.0599512
R18853 XThC.Tn[9].n9 XThC.Tn[9].n8 0.0599512
R18854 XThC.Tn[9].n67 XThC.Tn[9] 0.0469286
R18855 XThC.Tn[9].n63 XThC.Tn[9] 0.0469286
R18856 XThC.Tn[9].n59 XThC.Tn[9] 0.0469286
R18857 XThC.Tn[9].n55 XThC.Tn[9] 0.0469286
R18858 XThC.Tn[9].n51 XThC.Tn[9] 0.0469286
R18859 XThC.Tn[9].n47 XThC.Tn[9] 0.0469286
R18860 XThC.Tn[9].n43 XThC.Tn[9] 0.0469286
R18861 XThC.Tn[9].n39 XThC.Tn[9] 0.0469286
R18862 XThC.Tn[9].n35 XThC.Tn[9] 0.0469286
R18863 XThC.Tn[9].n31 XThC.Tn[9] 0.0469286
R18864 XThC.Tn[9].n27 XThC.Tn[9] 0.0469286
R18865 XThC.Tn[9].n23 XThC.Tn[9] 0.0469286
R18866 XThC.Tn[9].n19 XThC.Tn[9] 0.0469286
R18867 XThC.Tn[9].n15 XThC.Tn[9] 0.0469286
R18868 XThC.Tn[9].n11 XThC.Tn[9] 0.0469286
R18869 XThC.Tn[9].n8 XThC.Tn[9] 0.0469286
R18870 XThC.Tn[9].n67 XThC.Tn[9] 0.0401341
R18871 XThC.Tn[9].n63 XThC.Tn[9] 0.0401341
R18872 XThC.Tn[9].n59 XThC.Tn[9] 0.0401341
R18873 XThC.Tn[9].n55 XThC.Tn[9] 0.0401341
R18874 XThC.Tn[9].n51 XThC.Tn[9] 0.0401341
R18875 XThC.Tn[9].n47 XThC.Tn[9] 0.0401341
R18876 XThC.Tn[9].n43 XThC.Tn[9] 0.0401341
R18877 XThC.Tn[9].n39 XThC.Tn[9] 0.0401341
R18878 XThC.Tn[9].n35 XThC.Tn[9] 0.0401341
R18879 XThC.Tn[9].n31 XThC.Tn[9] 0.0401341
R18880 XThC.Tn[9].n27 XThC.Tn[9] 0.0401341
R18881 XThC.Tn[9].n23 XThC.Tn[9] 0.0401341
R18882 XThC.Tn[9].n19 XThC.Tn[9] 0.0401341
R18883 XThC.Tn[9].n15 XThC.Tn[9] 0.0401341
R18884 XThC.Tn[9].n11 XThC.Tn[9] 0.0401341
R18885 XThC.Tn[9].n8 XThC.Tn[9] 0.0401341
R18886 XThC.Tn[11].n70 XThC.Tn[11].n69 265.341
R18887 XThC.Tn[11].n74 XThC.Tn[11].n72 243.68
R18888 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R18889 XThC.Tn[11].n74 XThC.Tn[11].n73 205.28
R18890 XThC.Tn[11].n70 XThC.Tn[11].n68 202.094
R18891 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R18892 XThC.Tn[11].n64 XThC.Tn[11].n62 161.365
R18893 XThC.Tn[11].n60 XThC.Tn[11].n58 161.365
R18894 XThC.Tn[11].n56 XThC.Tn[11].n54 161.365
R18895 XThC.Tn[11].n52 XThC.Tn[11].n50 161.365
R18896 XThC.Tn[11].n48 XThC.Tn[11].n46 161.365
R18897 XThC.Tn[11].n44 XThC.Tn[11].n42 161.365
R18898 XThC.Tn[11].n40 XThC.Tn[11].n38 161.365
R18899 XThC.Tn[11].n36 XThC.Tn[11].n34 161.365
R18900 XThC.Tn[11].n32 XThC.Tn[11].n30 161.365
R18901 XThC.Tn[11].n28 XThC.Tn[11].n26 161.365
R18902 XThC.Tn[11].n24 XThC.Tn[11].n22 161.365
R18903 XThC.Tn[11].n20 XThC.Tn[11].n18 161.365
R18904 XThC.Tn[11].n16 XThC.Tn[11].n14 161.365
R18905 XThC.Tn[11].n12 XThC.Tn[11].n10 161.365
R18906 XThC.Tn[11].n8 XThC.Tn[11].n6 161.365
R18907 XThC.Tn[11].n5 XThC.Tn[11].n3 161.365
R18908 XThC.Tn[11].n62 XThC.Tn[11].t24 161.202
R18909 XThC.Tn[11].n58 XThC.Tn[11].t14 161.202
R18910 XThC.Tn[11].n54 XThC.Tn[11].t33 161.202
R18911 XThC.Tn[11].n50 XThC.Tn[11].t30 161.202
R18912 XThC.Tn[11].n46 XThC.Tn[11].t22 161.202
R18913 XThC.Tn[11].n42 XThC.Tn[11].t41 161.202
R18914 XThC.Tn[11].n38 XThC.Tn[11].t40 161.202
R18915 XThC.Tn[11].n34 XThC.Tn[11].t21 161.202
R18916 XThC.Tn[11].n30 XThC.Tn[11].t19 161.202
R18917 XThC.Tn[11].n26 XThC.Tn[11].t42 161.202
R18918 XThC.Tn[11].n22 XThC.Tn[11].t29 161.202
R18919 XThC.Tn[11].n18 XThC.Tn[11].t28 161.202
R18920 XThC.Tn[11].n14 XThC.Tn[11].t39 161.202
R18921 XThC.Tn[11].n10 XThC.Tn[11].t37 161.202
R18922 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R18923 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R18924 XThC.Tn[11].n62 XThC.Tn[11].t27 145.137
R18925 XThC.Tn[11].n58 XThC.Tn[11].t17 145.137
R18926 XThC.Tn[11].n54 XThC.Tn[11].t36 145.137
R18927 XThC.Tn[11].n50 XThC.Tn[11].t34 145.137
R18928 XThC.Tn[11].n46 XThC.Tn[11].t26 145.137
R18929 XThC.Tn[11].n42 XThC.Tn[11].t15 145.137
R18930 XThC.Tn[11].n38 XThC.Tn[11].t13 145.137
R18931 XThC.Tn[11].n34 XThC.Tn[11].t25 145.137
R18932 XThC.Tn[11].n30 XThC.Tn[11].t23 145.137
R18933 XThC.Tn[11].n26 XThC.Tn[11].t16 145.137
R18934 XThC.Tn[11].n22 XThC.Tn[11].t32 145.137
R18935 XThC.Tn[11].n18 XThC.Tn[11].t31 145.137
R18936 XThC.Tn[11].n14 XThC.Tn[11].t12 145.137
R18937 XThC.Tn[11].n10 XThC.Tn[11].t43 145.137
R18938 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R18939 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R18940 XThC.Tn[11].n68 XThC.Tn[11].t4 26.5955
R18941 XThC.Tn[11].n68 XThC.Tn[11].t1 26.5955
R18942 XThC.Tn[11].n72 XThC.Tn[11].t7 26.5955
R18943 XThC.Tn[11].n72 XThC.Tn[11].t10 26.5955
R18944 XThC.Tn[11].n73 XThC.Tn[11].t9 26.5955
R18945 XThC.Tn[11].n73 XThC.Tn[11].t8 26.5955
R18946 XThC.Tn[11].n69 XThC.Tn[11].t6 26.5955
R18947 XThC.Tn[11].n69 XThC.Tn[11].t0 26.5955
R18948 XThC.Tn[11].n1 XThC.Tn[11].t5 24.9236
R18949 XThC.Tn[11].n1 XThC.Tn[11].t3 24.9236
R18950 XThC.Tn[11].n0 XThC.Tn[11].t11 24.9236
R18951 XThC.Tn[11].n0 XThC.Tn[11].t2 24.9236
R18952 XThC.Tn[11] XThC.Tn[11].n74 22.9652
R18953 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R18954 XThC.Tn[11].n71 XThC.Tn[11].n70 13.9299
R18955 XThC.Tn[11] XThC.Tn[11].n71 13.9299
R18956 XThC.Tn[11] XThC.Tn[11].n5 8.0245
R18957 XThC.Tn[11].n65 XThC.Tn[11].n64 7.9105
R18958 XThC.Tn[11].n61 XThC.Tn[11].n60 7.9105
R18959 XThC.Tn[11].n57 XThC.Tn[11].n56 7.9105
R18960 XThC.Tn[11].n53 XThC.Tn[11].n52 7.9105
R18961 XThC.Tn[11].n49 XThC.Tn[11].n48 7.9105
R18962 XThC.Tn[11].n45 XThC.Tn[11].n44 7.9105
R18963 XThC.Tn[11].n41 XThC.Tn[11].n40 7.9105
R18964 XThC.Tn[11].n37 XThC.Tn[11].n36 7.9105
R18965 XThC.Tn[11].n33 XThC.Tn[11].n32 7.9105
R18966 XThC.Tn[11].n29 XThC.Tn[11].n28 7.9105
R18967 XThC.Tn[11].n25 XThC.Tn[11].n24 7.9105
R18968 XThC.Tn[11].n21 XThC.Tn[11].n20 7.9105
R18969 XThC.Tn[11].n17 XThC.Tn[11].n16 7.9105
R18970 XThC.Tn[11].n13 XThC.Tn[11].n12 7.9105
R18971 XThC.Tn[11].n9 XThC.Tn[11].n8 7.9105
R18972 XThC.Tn[11].n67 XThC.Tn[11].n66 7.44831
R18973 XThC.Tn[11].n67 XThC.Tn[11] 6.34069
R18974 XThC.Tn[11].n66 XThC.Tn[11] 4.37928
R18975 XThC.Tn[11] XThC.Tn[11].n67 1.79489
R18976 XThC.Tn[11].n71 XThC.Tn[11] 1.19676
R18977 XThC.Tn[11].n66 XThC.Tn[11] 1.0918
R18978 XThC.Tn[11].n9 XThC.Tn[11] 0.235138
R18979 XThC.Tn[11].n13 XThC.Tn[11] 0.235138
R18980 XThC.Tn[11].n17 XThC.Tn[11] 0.235138
R18981 XThC.Tn[11].n21 XThC.Tn[11] 0.235138
R18982 XThC.Tn[11].n25 XThC.Tn[11] 0.235138
R18983 XThC.Tn[11].n29 XThC.Tn[11] 0.235138
R18984 XThC.Tn[11].n33 XThC.Tn[11] 0.235138
R18985 XThC.Tn[11].n37 XThC.Tn[11] 0.235138
R18986 XThC.Tn[11].n41 XThC.Tn[11] 0.235138
R18987 XThC.Tn[11].n45 XThC.Tn[11] 0.235138
R18988 XThC.Tn[11].n49 XThC.Tn[11] 0.235138
R18989 XThC.Tn[11].n53 XThC.Tn[11] 0.235138
R18990 XThC.Tn[11].n57 XThC.Tn[11] 0.235138
R18991 XThC.Tn[11].n61 XThC.Tn[11] 0.235138
R18992 XThC.Tn[11].n65 XThC.Tn[11] 0.235138
R18993 XThC.Tn[11] XThC.Tn[11].n9 0.114505
R18994 XThC.Tn[11] XThC.Tn[11].n13 0.114505
R18995 XThC.Tn[11] XThC.Tn[11].n17 0.114505
R18996 XThC.Tn[11] XThC.Tn[11].n21 0.114505
R18997 XThC.Tn[11] XThC.Tn[11].n25 0.114505
R18998 XThC.Tn[11] XThC.Tn[11].n29 0.114505
R18999 XThC.Tn[11] XThC.Tn[11].n33 0.114505
R19000 XThC.Tn[11] XThC.Tn[11].n37 0.114505
R19001 XThC.Tn[11] XThC.Tn[11].n41 0.114505
R19002 XThC.Tn[11] XThC.Tn[11].n45 0.114505
R19003 XThC.Tn[11] XThC.Tn[11].n49 0.114505
R19004 XThC.Tn[11] XThC.Tn[11].n53 0.114505
R19005 XThC.Tn[11] XThC.Tn[11].n57 0.114505
R19006 XThC.Tn[11] XThC.Tn[11].n61 0.114505
R19007 XThC.Tn[11] XThC.Tn[11].n65 0.114505
R19008 XThC.Tn[11].n64 XThC.Tn[11].n63 0.0599512
R19009 XThC.Tn[11].n60 XThC.Tn[11].n59 0.0599512
R19010 XThC.Tn[11].n56 XThC.Tn[11].n55 0.0599512
R19011 XThC.Tn[11].n52 XThC.Tn[11].n51 0.0599512
R19012 XThC.Tn[11].n48 XThC.Tn[11].n47 0.0599512
R19013 XThC.Tn[11].n44 XThC.Tn[11].n43 0.0599512
R19014 XThC.Tn[11].n40 XThC.Tn[11].n39 0.0599512
R19015 XThC.Tn[11].n36 XThC.Tn[11].n35 0.0599512
R19016 XThC.Tn[11].n32 XThC.Tn[11].n31 0.0599512
R19017 XThC.Tn[11].n28 XThC.Tn[11].n27 0.0599512
R19018 XThC.Tn[11].n24 XThC.Tn[11].n23 0.0599512
R19019 XThC.Tn[11].n20 XThC.Tn[11].n19 0.0599512
R19020 XThC.Tn[11].n16 XThC.Tn[11].n15 0.0599512
R19021 XThC.Tn[11].n12 XThC.Tn[11].n11 0.0599512
R19022 XThC.Tn[11].n8 XThC.Tn[11].n7 0.0599512
R19023 XThC.Tn[11].n5 XThC.Tn[11].n4 0.0599512
R19024 XThC.Tn[11].n63 XThC.Tn[11] 0.0469286
R19025 XThC.Tn[11].n59 XThC.Tn[11] 0.0469286
R19026 XThC.Tn[11].n55 XThC.Tn[11] 0.0469286
R19027 XThC.Tn[11].n51 XThC.Tn[11] 0.0469286
R19028 XThC.Tn[11].n47 XThC.Tn[11] 0.0469286
R19029 XThC.Tn[11].n43 XThC.Tn[11] 0.0469286
R19030 XThC.Tn[11].n39 XThC.Tn[11] 0.0469286
R19031 XThC.Tn[11].n35 XThC.Tn[11] 0.0469286
R19032 XThC.Tn[11].n31 XThC.Tn[11] 0.0469286
R19033 XThC.Tn[11].n27 XThC.Tn[11] 0.0469286
R19034 XThC.Tn[11].n23 XThC.Tn[11] 0.0469286
R19035 XThC.Tn[11].n19 XThC.Tn[11] 0.0469286
R19036 XThC.Tn[11].n15 XThC.Tn[11] 0.0469286
R19037 XThC.Tn[11].n11 XThC.Tn[11] 0.0469286
R19038 XThC.Tn[11].n7 XThC.Tn[11] 0.0469286
R19039 XThC.Tn[11].n4 XThC.Tn[11] 0.0469286
R19040 XThC.Tn[11].n63 XThC.Tn[11] 0.0401341
R19041 XThC.Tn[11].n59 XThC.Tn[11] 0.0401341
R19042 XThC.Tn[11].n55 XThC.Tn[11] 0.0401341
R19043 XThC.Tn[11].n51 XThC.Tn[11] 0.0401341
R19044 XThC.Tn[11].n47 XThC.Tn[11] 0.0401341
R19045 XThC.Tn[11].n43 XThC.Tn[11] 0.0401341
R19046 XThC.Tn[11].n39 XThC.Tn[11] 0.0401341
R19047 XThC.Tn[11].n35 XThC.Tn[11] 0.0401341
R19048 XThC.Tn[11].n31 XThC.Tn[11] 0.0401341
R19049 XThC.Tn[11].n27 XThC.Tn[11] 0.0401341
R19050 XThC.Tn[11].n23 XThC.Tn[11] 0.0401341
R19051 XThC.Tn[11].n19 XThC.Tn[11] 0.0401341
R19052 XThC.Tn[11].n15 XThC.Tn[11] 0.0401341
R19053 XThC.Tn[11].n11 XThC.Tn[11] 0.0401341
R19054 XThC.Tn[11].n7 XThC.Tn[11] 0.0401341
R19055 XThC.Tn[11].n4 XThC.Tn[11] 0.0401341
R19056 XThC.Tn[12].n70 XThC.Tn[12].n69 256.104
R19057 XThC.Tn[12].n74 XThC.Tn[12].n72 243.68
R19058 XThC.Tn[12].n2 XThC.Tn[12].n0 241.847
R19059 XThC.Tn[12].n74 XThC.Tn[12].n73 205.28
R19060 XThC.Tn[12].n70 XThC.Tn[12].n68 202.095
R19061 XThC.Tn[12].n2 XThC.Tn[12].n1 185
R19062 XThC.Tn[12].n64 XThC.Tn[12].n62 161.365
R19063 XThC.Tn[12].n60 XThC.Tn[12].n58 161.365
R19064 XThC.Tn[12].n56 XThC.Tn[12].n54 161.365
R19065 XThC.Tn[12].n52 XThC.Tn[12].n50 161.365
R19066 XThC.Tn[12].n48 XThC.Tn[12].n46 161.365
R19067 XThC.Tn[12].n44 XThC.Tn[12].n42 161.365
R19068 XThC.Tn[12].n40 XThC.Tn[12].n38 161.365
R19069 XThC.Tn[12].n36 XThC.Tn[12].n34 161.365
R19070 XThC.Tn[12].n32 XThC.Tn[12].n30 161.365
R19071 XThC.Tn[12].n28 XThC.Tn[12].n26 161.365
R19072 XThC.Tn[12].n24 XThC.Tn[12].n22 161.365
R19073 XThC.Tn[12].n20 XThC.Tn[12].n18 161.365
R19074 XThC.Tn[12].n16 XThC.Tn[12].n14 161.365
R19075 XThC.Tn[12].n12 XThC.Tn[12].n10 161.365
R19076 XThC.Tn[12].n8 XThC.Tn[12].n6 161.365
R19077 XThC.Tn[12].n5 XThC.Tn[12].n3 161.365
R19078 XThC.Tn[12].n62 XThC.Tn[12].t41 161.202
R19079 XThC.Tn[12].n58 XThC.Tn[12].t31 161.202
R19080 XThC.Tn[12].n54 XThC.Tn[12].t18 161.202
R19081 XThC.Tn[12].n50 XThC.Tn[12].t15 161.202
R19082 XThC.Tn[12].n46 XThC.Tn[12].t39 161.202
R19083 XThC.Tn[12].n42 XThC.Tn[12].t26 161.202
R19084 XThC.Tn[12].n38 XThC.Tn[12].t25 161.202
R19085 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R19086 XThC.Tn[12].n30 XThC.Tn[12].t36 161.202
R19087 XThC.Tn[12].n26 XThC.Tn[12].t27 161.202
R19088 XThC.Tn[12].n22 XThC.Tn[12].t14 161.202
R19089 XThC.Tn[12].n18 XThC.Tn[12].t13 161.202
R19090 XThC.Tn[12].n14 XThC.Tn[12].t24 161.202
R19091 XThC.Tn[12].n10 XThC.Tn[12].t22 161.202
R19092 XThC.Tn[12].n6 XThC.Tn[12].t20 161.202
R19093 XThC.Tn[12].n3 XThC.Tn[12].t35 161.202
R19094 XThC.Tn[12].n62 XThC.Tn[12].t12 145.137
R19095 XThC.Tn[12].n58 XThC.Tn[12].t34 145.137
R19096 XThC.Tn[12].n54 XThC.Tn[12].t21 145.137
R19097 XThC.Tn[12].n50 XThC.Tn[12].t19 145.137
R19098 XThC.Tn[12].n46 XThC.Tn[12].t43 145.137
R19099 XThC.Tn[12].n42 XThC.Tn[12].t32 145.137
R19100 XThC.Tn[12].n38 XThC.Tn[12].t30 145.137
R19101 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R19102 XThC.Tn[12].n30 XThC.Tn[12].t40 145.137
R19103 XThC.Tn[12].n26 XThC.Tn[12].t33 145.137
R19104 XThC.Tn[12].n22 XThC.Tn[12].t17 145.137
R19105 XThC.Tn[12].n18 XThC.Tn[12].t16 145.137
R19106 XThC.Tn[12].n14 XThC.Tn[12].t29 145.137
R19107 XThC.Tn[12].n10 XThC.Tn[12].t28 145.137
R19108 XThC.Tn[12].n6 XThC.Tn[12].t23 145.137
R19109 XThC.Tn[12].n3 XThC.Tn[12].t37 145.137
R19110 XThC.Tn[12].n72 XThC.Tn[12].t1 26.5955
R19111 XThC.Tn[12].n72 XThC.Tn[12].t0 26.5955
R19112 XThC.Tn[12].n68 XThC.Tn[12].t9 26.5955
R19113 XThC.Tn[12].n68 XThC.Tn[12].t10 26.5955
R19114 XThC.Tn[12].n69 XThC.Tn[12].t8 26.5955
R19115 XThC.Tn[12].n69 XThC.Tn[12].t11 26.5955
R19116 XThC.Tn[12].n73 XThC.Tn[12].t3 26.5955
R19117 XThC.Tn[12].n73 XThC.Tn[12].t2 26.5955
R19118 XThC.Tn[12].n1 XThC.Tn[12].t5 24.9236
R19119 XThC.Tn[12].n1 XThC.Tn[12].t4 24.9236
R19120 XThC.Tn[12].n0 XThC.Tn[12].t7 24.9236
R19121 XThC.Tn[12].n0 XThC.Tn[12].t6 24.9236
R19122 XThC.Tn[12] XThC.Tn[12].n74 22.9652
R19123 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R19124 XThC.Tn[12].n71 XThC.Tn[12].n70 13.9299
R19125 XThC.Tn[12] XThC.Tn[12].n71 13.9299
R19126 XThC.Tn[12] XThC.Tn[12].n5 8.0245
R19127 XThC.Tn[12].n65 XThC.Tn[12].n64 7.9105
R19128 XThC.Tn[12].n61 XThC.Tn[12].n60 7.9105
R19129 XThC.Tn[12].n57 XThC.Tn[12].n56 7.9105
R19130 XThC.Tn[12].n53 XThC.Tn[12].n52 7.9105
R19131 XThC.Tn[12].n49 XThC.Tn[12].n48 7.9105
R19132 XThC.Tn[12].n45 XThC.Tn[12].n44 7.9105
R19133 XThC.Tn[12].n41 XThC.Tn[12].n40 7.9105
R19134 XThC.Tn[12].n37 XThC.Tn[12].n36 7.9105
R19135 XThC.Tn[12].n33 XThC.Tn[12].n32 7.9105
R19136 XThC.Tn[12].n29 XThC.Tn[12].n28 7.9105
R19137 XThC.Tn[12].n25 XThC.Tn[12].n24 7.9105
R19138 XThC.Tn[12].n21 XThC.Tn[12].n20 7.9105
R19139 XThC.Tn[12].n17 XThC.Tn[12].n16 7.9105
R19140 XThC.Tn[12].n13 XThC.Tn[12].n12 7.9105
R19141 XThC.Tn[12].n9 XThC.Tn[12].n8 7.9105
R19142 XThC.Tn[12].n67 XThC.Tn[12].n66 7.4309
R19143 XThC.Tn[12].n66 XThC.Tn[12] 4.71945
R19144 XThC.Tn[12].n71 XThC.Tn[12].n67 2.99115
R19145 XThC.Tn[12].n71 XThC.Tn[12] 2.87153
R19146 XThC.Tn[12].n67 XThC.Tn[12] 2.2734
R19147 XThC.Tn[12].n66 XThC.Tn[12] 0.88175
R19148 XThC.Tn[12].n9 XThC.Tn[12] 0.235138
R19149 XThC.Tn[12].n13 XThC.Tn[12] 0.235138
R19150 XThC.Tn[12].n17 XThC.Tn[12] 0.235138
R19151 XThC.Tn[12].n21 XThC.Tn[12] 0.235138
R19152 XThC.Tn[12].n25 XThC.Tn[12] 0.235138
R19153 XThC.Tn[12].n29 XThC.Tn[12] 0.235138
R19154 XThC.Tn[12].n33 XThC.Tn[12] 0.235138
R19155 XThC.Tn[12].n37 XThC.Tn[12] 0.235138
R19156 XThC.Tn[12].n41 XThC.Tn[12] 0.235138
R19157 XThC.Tn[12].n45 XThC.Tn[12] 0.235138
R19158 XThC.Tn[12].n49 XThC.Tn[12] 0.235138
R19159 XThC.Tn[12].n53 XThC.Tn[12] 0.235138
R19160 XThC.Tn[12].n57 XThC.Tn[12] 0.235138
R19161 XThC.Tn[12].n61 XThC.Tn[12] 0.235138
R19162 XThC.Tn[12].n65 XThC.Tn[12] 0.235138
R19163 XThC.Tn[12] XThC.Tn[12].n9 0.114505
R19164 XThC.Tn[12] XThC.Tn[12].n13 0.114505
R19165 XThC.Tn[12] XThC.Tn[12].n17 0.114505
R19166 XThC.Tn[12] XThC.Tn[12].n21 0.114505
R19167 XThC.Tn[12] XThC.Tn[12].n25 0.114505
R19168 XThC.Tn[12] XThC.Tn[12].n29 0.114505
R19169 XThC.Tn[12] XThC.Tn[12].n33 0.114505
R19170 XThC.Tn[12] XThC.Tn[12].n37 0.114505
R19171 XThC.Tn[12] XThC.Tn[12].n41 0.114505
R19172 XThC.Tn[12] XThC.Tn[12].n45 0.114505
R19173 XThC.Tn[12] XThC.Tn[12].n49 0.114505
R19174 XThC.Tn[12] XThC.Tn[12].n53 0.114505
R19175 XThC.Tn[12] XThC.Tn[12].n57 0.114505
R19176 XThC.Tn[12] XThC.Tn[12].n61 0.114505
R19177 XThC.Tn[12] XThC.Tn[12].n65 0.114505
R19178 XThC.Tn[12].n64 XThC.Tn[12].n63 0.0599512
R19179 XThC.Tn[12].n60 XThC.Tn[12].n59 0.0599512
R19180 XThC.Tn[12].n56 XThC.Tn[12].n55 0.0599512
R19181 XThC.Tn[12].n52 XThC.Tn[12].n51 0.0599512
R19182 XThC.Tn[12].n48 XThC.Tn[12].n47 0.0599512
R19183 XThC.Tn[12].n44 XThC.Tn[12].n43 0.0599512
R19184 XThC.Tn[12].n40 XThC.Tn[12].n39 0.0599512
R19185 XThC.Tn[12].n36 XThC.Tn[12].n35 0.0599512
R19186 XThC.Tn[12].n32 XThC.Tn[12].n31 0.0599512
R19187 XThC.Tn[12].n28 XThC.Tn[12].n27 0.0599512
R19188 XThC.Tn[12].n24 XThC.Tn[12].n23 0.0599512
R19189 XThC.Tn[12].n20 XThC.Tn[12].n19 0.0599512
R19190 XThC.Tn[12].n16 XThC.Tn[12].n15 0.0599512
R19191 XThC.Tn[12].n12 XThC.Tn[12].n11 0.0599512
R19192 XThC.Tn[12].n8 XThC.Tn[12].n7 0.0599512
R19193 XThC.Tn[12].n5 XThC.Tn[12].n4 0.0599512
R19194 XThC.Tn[12].n63 XThC.Tn[12] 0.0469286
R19195 XThC.Tn[12].n59 XThC.Tn[12] 0.0469286
R19196 XThC.Tn[12].n55 XThC.Tn[12] 0.0469286
R19197 XThC.Tn[12].n51 XThC.Tn[12] 0.0469286
R19198 XThC.Tn[12].n47 XThC.Tn[12] 0.0469286
R19199 XThC.Tn[12].n43 XThC.Tn[12] 0.0469286
R19200 XThC.Tn[12].n39 XThC.Tn[12] 0.0469286
R19201 XThC.Tn[12].n35 XThC.Tn[12] 0.0469286
R19202 XThC.Tn[12].n31 XThC.Tn[12] 0.0469286
R19203 XThC.Tn[12].n27 XThC.Tn[12] 0.0469286
R19204 XThC.Tn[12].n23 XThC.Tn[12] 0.0469286
R19205 XThC.Tn[12].n19 XThC.Tn[12] 0.0469286
R19206 XThC.Tn[12].n15 XThC.Tn[12] 0.0469286
R19207 XThC.Tn[12].n11 XThC.Tn[12] 0.0469286
R19208 XThC.Tn[12].n7 XThC.Tn[12] 0.0469286
R19209 XThC.Tn[12].n4 XThC.Tn[12] 0.0469286
R19210 XThC.Tn[12].n63 XThC.Tn[12] 0.0401341
R19211 XThC.Tn[12].n59 XThC.Tn[12] 0.0401341
R19212 XThC.Tn[12].n55 XThC.Tn[12] 0.0401341
R19213 XThC.Tn[12].n51 XThC.Tn[12] 0.0401341
R19214 XThC.Tn[12].n47 XThC.Tn[12] 0.0401341
R19215 XThC.Tn[12].n43 XThC.Tn[12] 0.0401341
R19216 XThC.Tn[12].n39 XThC.Tn[12] 0.0401341
R19217 XThC.Tn[12].n35 XThC.Tn[12] 0.0401341
R19218 XThC.Tn[12].n31 XThC.Tn[12] 0.0401341
R19219 XThC.Tn[12].n27 XThC.Tn[12] 0.0401341
R19220 XThC.Tn[12].n23 XThC.Tn[12] 0.0401341
R19221 XThC.Tn[12].n19 XThC.Tn[12] 0.0401341
R19222 XThC.Tn[12].n15 XThC.Tn[12] 0.0401341
R19223 XThC.Tn[12].n11 XThC.Tn[12] 0.0401341
R19224 XThC.Tn[12].n7 XThC.Tn[12] 0.0401341
R19225 XThC.Tn[12].n4 XThC.Tn[12] 0.0401341
R19226 XThC.Tn[13].n2 XThC.Tn[13].n1 265.341
R19227 XThC.Tn[13].n5 XThC.Tn[13].n3 243.68
R19228 XThC.Tn[13].n74 XThC.Tn[13].n73 241.847
R19229 XThC.Tn[13].n5 XThC.Tn[13].n4 205.28
R19230 XThC.Tn[13].n2 XThC.Tn[13].n0 202.094
R19231 XThC.Tn[13].n74 XThC.Tn[13].n72 185
R19232 XThC.Tn[13].n68 XThC.Tn[13].n66 161.365
R19233 XThC.Tn[13].n64 XThC.Tn[13].n62 161.365
R19234 XThC.Tn[13].n60 XThC.Tn[13].n58 161.365
R19235 XThC.Tn[13].n56 XThC.Tn[13].n54 161.365
R19236 XThC.Tn[13].n52 XThC.Tn[13].n50 161.365
R19237 XThC.Tn[13].n48 XThC.Tn[13].n46 161.365
R19238 XThC.Tn[13].n44 XThC.Tn[13].n42 161.365
R19239 XThC.Tn[13].n40 XThC.Tn[13].n38 161.365
R19240 XThC.Tn[13].n36 XThC.Tn[13].n34 161.365
R19241 XThC.Tn[13].n32 XThC.Tn[13].n30 161.365
R19242 XThC.Tn[13].n28 XThC.Tn[13].n26 161.365
R19243 XThC.Tn[13].n24 XThC.Tn[13].n22 161.365
R19244 XThC.Tn[13].n20 XThC.Tn[13].n18 161.365
R19245 XThC.Tn[13].n16 XThC.Tn[13].n14 161.365
R19246 XThC.Tn[13].n12 XThC.Tn[13].n10 161.365
R19247 XThC.Tn[13].n9 XThC.Tn[13].n7 161.365
R19248 XThC.Tn[13].n66 XThC.Tn[13].t33 161.202
R19249 XThC.Tn[13].n62 XThC.Tn[13].t23 161.202
R19250 XThC.Tn[13].n58 XThC.Tn[13].t42 161.202
R19251 XThC.Tn[13].n54 XThC.Tn[13].t39 161.202
R19252 XThC.Tn[13].n50 XThC.Tn[13].t31 161.202
R19253 XThC.Tn[13].n46 XThC.Tn[13].t18 161.202
R19254 XThC.Tn[13].n42 XThC.Tn[13].t17 161.202
R19255 XThC.Tn[13].n38 XThC.Tn[13].t30 161.202
R19256 XThC.Tn[13].n34 XThC.Tn[13].t28 161.202
R19257 XThC.Tn[13].n30 XThC.Tn[13].t19 161.202
R19258 XThC.Tn[13].n26 XThC.Tn[13].t38 161.202
R19259 XThC.Tn[13].n22 XThC.Tn[13].t37 161.202
R19260 XThC.Tn[13].n18 XThC.Tn[13].t16 161.202
R19261 XThC.Tn[13].n14 XThC.Tn[13].t14 161.202
R19262 XThC.Tn[13].n10 XThC.Tn[13].t12 161.202
R19263 XThC.Tn[13].n7 XThC.Tn[13].t27 161.202
R19264 XThC.Tn[13].n66 XThC.Tn[13].t36 145.137
R19265 XThC.Tn[13].n62 XThC.Tn[13].t26 145.137
R19266 XThC.Tn[13].n58 XThC.Tn[13].t13 145.137
R19267 XThC.Tn[13].n54 XThC.Tn[13].t43 145.137
R19268 XThC.Tn[13].n50 XThC.Tn[13].t35 145.137
R19269 XThC.Tn[13].n46 XThC.Tn[13].t24 145.137
R19270 XThC.Tn[13].n42 XThC.Tn[13].t22 145.137
R19271 XThC.Tn[13].n38 XThC.Tn[13].t34 145.137
R19272 XThC.Tn[13].n34 XThC.Tn[13].t32 145.137
R19273 XThC.Tn[13].n30 XThC.Tn[13].t25 145.137
R19274 XThC.Tn[13].n26 XThC.Tn[13].t41 145.137
R19275 XThC.Tn[13].n22 XThC.Tn[13].t40 145.137
R19276 XThC.Tn[13].n18 XThC.Tn[13].t21 145.137
R19277 XThC.Tn[13].n14 XThC.Tn[13].t20 145.137
R19278 XThC.Tn[13].n10 XThC.Tn[13].t15 145.137
R19279 XThC.Tn[13].n7 XThC.Tn[13].t29 145.137
R19280 XThC.Tn[13].n1 XThC.Tn[13].t4 26.5955
R19281 XThC.Tn[13].n1 XThC.Tn[13].t7 26.5955
R19282 XThC.Tn[13].n0 XThC.Tn[13].t6 26.5955
R19283 XThC.Tn[13].n0 XThC.Tn[13].t5 26.5955
R19284 XThC.Tn[13].n3 XThC.Tn[13].t9 26.5955
R19285 XThC.Tn[13].n3 XThC.Tn[13].t8 26.5955
R19286 XThC.Tn[13].n4 XThC.Tn[13].t11 26.5955
R19287 XThC.Tn[13].n4 XThC.Tn[13].t10 26.5955
R19288 XThC.Tn[13].n72 XThC.Tn[13].t0 24.9236
R19289 XThC.Tn[13].n72 XThC.Tn[13].t2 24.9236
R19290 XThC.Tn[13].n73 XThC.Tn[13].t3 24.9236
R19291 XThC.Tn[13].n73 XThC.Tn[13].t1 24.9236
R19292 XThC.Tn[13] XThC.Tn[13].n5 22.9652
R19293 XThC.Tn[13] XThC.Tn[13].n74 18.8943
R19294 XThC.Tn[13].n6 XThC.Tn[13].n2 13.9299
R19295 XThC.Tn[13].n6 XThC.Tn[13] 13.9299
R19296 XThC.Tn[13] XThC.Tn[13].n9 8.0245
R19297 XThC.Tn[13].n69 XThC.Tn[13].n68 7.9105
R19298 XThC.Tn[13].n65 XThC.Tn[13].n64 7.9105
R19299 XThC.Tn[13].n61 XThC.Tn[13].n60 7.9105
R19300 XThC.Tn[13].n57 XThC.Tn[13].n56 7.9105
R19301 XThC.Tn[13].n53 XThC.Tn[13].n52 7.9105
R19302 XThC.Tn[13].n49 XThC.Tn[13].n48 7.9105
R19303 XThC.Tn[13].n45 XThC.Tn[13].n44 7.9105
R19304 XThC.Tn[13].n41 XThC.Tn[13].n40 7.9105
R19305 XThC.Tn[13].n37 XThC.Tn[13].n36 7.9105
R19306 XThC.Tn[13].n33 XThC.Tn[13].n32 7.9105
R19307 XThC.Tn[13].n29 XThC.Tn[13].n28 7.9105
R19308 XThC.Tn[13].n25 XThC.Tn[13].n24 7.9105
R19309 XThC.Tn[13].n21 XThC.Tn[13].n20 7.9105
R19310 XThC.Tn[13].n17 XThC.Tn[13].n16 7.9105
R19311 XThC.Tn[13].n13 XThC.Tn[13].n12 7.9105
R19312 XThC.Tn[13].n71 XThC.Tn[13].n70 7.46054
R19313 XThC.Tn[13] XThC.Tn[13].n71 6.34069
R19314 XThC.Tn[13].n70 XThC.Tn[13] 4.78838
R19315 XThC.Tn[13].n71 XThC.Tn[13] 1.79489
R19316 XThC.Tn[13].n70 XThC.Tn[13] 1.51436
R19317 XThC.Tn[13] XThC.Tn[13].n6 1.19676
R19318 XThC.Tn[13].n13 XThC.Tn[13] 0.235138
R19319 XThC.Tn[13].n17 XThC.Tn[13] 0.235138
R19320 XThC.Tn[13].n21 XThC.Tn[13] 0.235138
R19321 XThC.Tn[13].n25 XThC.Tn[13] 0.235138
R19322 XThC.Tn[13].n29 XThC.Tn[13] 0.235138
R19323 XThC.Tn[13].n33 XThC.Tn[13] 0.235138
R19324 XThC.Tn[13].n37 XThC.Tn[13] 0.235138
R19325 XThC.Tn[13].n41 XThC.Tn[13] 0.235138
R19326 XThC.Tn[13].n45 XThC.Tn[13] 0.235138
R19327 XThC.Tn[13].n49 XThC.Tn[13] 0.235138
R19328 XThC.Tn[13].n53 XThC.Tn[13] 0.235138
R19329 XThC.Tn[13].n57 XThC.Tn[13] 0.235138
R19330 XThC.Tn[13].n61 XThC.Tn[13] 0.235138
R19331 XThC.Tn[13].n65 XThC.Tn[13] 0.235138
R19332 XThC.Tn[13].n69 XThC.Tn[13] 0.235138
R19333 XThC.Tn[13] XThC.Tn[13].n13 0.114505
R19334 XThC.Tn[13] XThC.Tn[13].n17 0.114505
R19335 XThC.Tn[13] XThC.Tn[13].n21 0.114505
R19336 XThC.Tn[13] XThC.Tn[13].n25 0.114505
R19337 XThC.Tn[13] XThC.Tn[13].n29 0.114505
R19338 XThC.Tn[13] XThC.Tn[13].n33 0.114505
R19339 XThC.Tn[13] XThC.Tn[13].n37 0.114505
R19340 XThC.Tn[13] XThC.Tn[13].n41 0.114505
R19341 XThC.Tn[13] XThC.Tn[13].n45 0.114505
R19342 XThC.Tn[13] XThC.Tn[13].n49 0.114505
R19343 XThC.Tn[13] XThC.Tn[13].n53 0.114505
R19344 XThC.Tn[13] XThC.Tn[13].n57 0.114505
R19345 XThC.Tn[13] XThC.Tn[13].n61 0.114505
R19346 XThC.Tn[13] XThC.Tn[13].n65 0.114505
R19347 XThC.Tn[13] XThC.Tn[13].n69 0.114505
R19348 XThC.Tn[13].n68 XThC.Tn[13].n67 0.0599512
R19349 XThC.Tn[13].n64 XThC.Tn[13].n63 0.0599512
R19350 XThC.Tn[13].n60 XThC.Tn[13].n59 0.0599512
R19351 XThC.Tn[13].n56 XThC.Tn[13].n55 0.0599512
R19352 XThC.Tn[13].n52 XThC.Tn[13].n51 0.0599512
R19353 XThC.Tn[13].n48 XThC.Tn[13].n47 0.0599512
R19354 XThC.Tn[13].n44 XThC.Tn[13].n43 0.0599512
R19355 XThC.Tn[13].n40 XThC.Tn[13].n39 0.0599512
R19356 XThC.Tn[13].n36 XThC.Tn[13].n35 0.0599512
R19357 XThC.Tn[13].n32 XThC.Tn[13].n31 0.0599512
R19358 XThC.Tn[13].n28 XThC.Tn[13].n27 0.0599512
R19359 XThC.Tn[13].n24 XThC.Tn[13].n23 0.0599512
R19360 XThC.Tn[13].n20 XThC.Tn[13].n19 0.0599512
R19361 XThC.Tn[13].n16 XThC.Tn[13].n15 0.0599512
R19362 XThC.Tn[13].n12 XThC.Tn[13].n11 0.0599512
R19363 XThC.Tn[13].n9 XThC.Tn[13].n8 0.0599512
R19364 XThC.Tn[13].n67 XThC.Tn[13] 0.0469286
R19365 XThC.Tn[13].n63 XThC.Tn[13] 0.0469286
R19366 XThC.Tn[13].n59 XThC.Tn[13] 0.0469286
R19367 XThC.Tn[13].n55 XThC.Tn[13] 0.0469286
R19368 XThC.Tn[13].n51 XThC.Tn[13] 0.0469286
R19369 XThC.Tn[13].n47 XThC.Tn[13] 0.0469286
R19370 XThC.Tn[13].n43 XThC.Tn[13] 0.0469286
R19371 XThC.Tn[13].n39 XThC.Tn[13] 0.0469286
R19372 XThC.Tn[13].n35 XThC.Tn[13] 0.0469286
R19373 XThC.Tn[13].n31 XThC.Tn[13] 0.0469286
R19374 XThC.Tn[13].n27 XThC.Tn[13] 0.0469286
R19375 XThC.Tn[13].n23 XThC.Tn[13] 0.0469286
R19376 XThC.Tn[13].n19 XThC.Tn[13] 0.0469286
R19377 XThC.Tn[13].n15 XThC.Tn[13] 0.0469286
R19378 XThC.Tn[13].n11 XThC.Tn[13] 0.0469286
R19379 XThC.Tn[13].n8 XThC.Tn[13] 0.0469286
R19380 XThC.Tn[13].n67 XThC.Tn[13] 0.0401341
R19381 XThC.Tn[13].n63 XThC.Tn[13] 0.0401341
R19382 XThC.Tn[13].n59 XThC.Tn[13] 0.0401341
R19383 XThC.Tn[13].n55 XThC.Tn[13] 0.0401341
R19384 XThC.Tn[13].n51 XThC.Tn[13] 0.0401341
R19385 XThC.Tn[13].n47 XThC.Tn[13] 0.0401341
R19386 XThC.Tn[13].n43 XThC.Tn[13] 0.0401341
R19387 XThC.Tn[13].n39 XThC.Tn[13] 0.0401341
R19388 XThC.Tn[13].n35 XThC.Tn[13] 0.0401341
R19389 XThC.Tn[13].n31 XThC.Tn[13] 0.0401341
R19390 XThC.Tn[13].n27 XThC.Tn[13] 0.0401341
R19391 XThC.Tn[13].n23 XThC.Tn[13] 0.0401341
R19392 XThC.Tn[13].n19 XThC.Tn[13] 0.0401341
R19393 XThC.Tn[13].n15 XThC.Tn[13] 0.0401341
R19394 XThC.Tn[13].n11 XThC.Tn[13] 0.0401341
R19395 XThC.Tn[13].n8 XThC.Tn[13] 0.0401341
R19396 XThC.Tn[0].n2 XThC.Tn[0].n1 332.332
R19397 XThC.Tn[0].n2 XThC.Tn[0].n0 296.493
R19398 XThC.Tn[0].n71 XThC.Tn[0].n69 161.365
R19399 XThC.Tn[0].n67 XThC.Tn[0].n65 161.365
R19400 XThC.Tn[0].n63 XThC.Tn[0].n61 161.365
R19401 XThC.Tn[0].n59 XThC.Tn[0].n57 161.365
R19402 XThC.Tn[0].n55 XThC.Tn[0].n53 161.365
R19403 XThC.Tn[0].n51 XThC.Tn[0].n49 161.365
R19404 XThC.Tn[0].n47 XThC.Tn[0].n45 161.365
R19405 XThC.Tn[0].n43 XThC.Tn[0].n41 161.365
R19406 XThC.Tn[0].n39 XThC.Tn[0].n37 161.365
R19407 XThC.Tn[0].n35 XThC.Tn[0].n33 161.365
R19408 XThC.Tn[0].n31 XThC.Tn[0].n29 161.365
R19409 XThC.Tn[0].n27 XThC.Tn[0].n25 161.365
R19410 XThC.Tn[0].n23 XThC.Tn[0].n21 161.365
R19411 XThC.Tn[0].n19 XThC.Tn[0].n17 161.365
R19412 XThC.Tn[0].n15 XThC.Tn[0].n13 161.365
R19413 XThC.Tn[0].n12 XThC.Tn[0].n10 161.365
R19414 XThC.Tn[0].n69 XThC.Tn[0].t29 161.202
R19415 XThC.Tn[0].n65 XThC.Tn[0].t19 161.202
R19416 XThC.Tn[0].n61 XThC.Tn[0].t38 161.202
R19417 XThC.Tn[0].n57 XThC.Tn[0].t36 161.202
R19418 XThC.Tn[0].n53 XThC.Tn[0].t27 161.202
R19419 XThC.Tn[0].n49 XThC.Tn[0].t16 161.202
R19420 XThC.Tn[0].n45 XThC.Tn[0].t15 161.202
R19421 XThC.Tn[0].n41 XThC.Tn[0].t26 161.202
R19422 XThC.Tn[0].n37 XThC.Tn[0].t25 161.202
R19423 XThC.Tn[0].n33 XThC.Tn[0].t17 161.202
R19424 XThC.Tn[0].n29 XThC.Tn[0].t34 161.202
R19425 XThC.Tn[0].n25 XThC.Tn[0].t32 161.202
R19426 XThC.Tn[0].n21 XThC.Tn[0].t13 161.202
R19427 XThC.Tn[0].n17 XThC.Tn[0].t12 161.202
R19428 XThC.Tn[0].n13 XThC.Tn[0].t41 161.202
R19429 XThC.Tn[0].n10 XThC.Tn[0].t22 161.202
R19430 XThC.Tn[0].n69 XThC.Tn[0].t24 145.137
R19431 XThC.Tn[0].n65 XThC.Tn[0].t14 145.137
R19432 XThC.Tn[0].n61 XThC.Tn[0].t33 145.137
R19433 XThC.Tn[0].n57 XThC.Tn[0].t31 145.137
R19434 XThC.Tn[0].n53 XThC.Tn[0].t23 145.137
R19435 XThC.Tn[0].n49 XThC.Tn[0].t42 145.137
R19436 XThC.Tn[0].n45 XThC.Tn[0].t40 145.137
R19437 XThC.Tn[0].n41 XThC.Tn[0].t21 145.137
R19438 XThC.Tn[0].n37 XThC.Tn[0].t20 145.137
R19439 XThC.Tn[0].n33 XThC.Tn[0].t43 145.137
R19440 XThC.Tn[0].n29 XThC.Tn[0].t30 145.137
R19441 XThC.Tn[0].n25 XThC.Tn[0].t28 145.137
R19442 XThC.Tn[0].n21 XThC.Tn[0].t39 145.137
R19443 XThC.Tn[0].n17 XThC.Tn[0].t37 145.137
R19444 XThC.Tn[0].n13 XThC.Tn[0].t35 145.137
R19445 XThC.Tn[0].n10 XThC.Tn[0].t18 145.137
R19446 XThC.Tn[0].n7 XThC.Tn[0].n6 135.248
R19447 XThC.Tn[0].n9 XThC.Tn[0].n3 98.982
R19448 XThC.Tn[0].n8 XThC.Tn[0].n4 98.982
R19449 XThC.Tn[0].n7 XThC.Tn[0].n5 98.982
R19450 XThC.Tn[0].n9 XThC.Tn[0].n8 36.2672
R19451 XThC.Tn[0].n8 XThC.Tn[0].n7 36.2672
R19452 XThC.Tn[0].n74 XThC.Tn[0].n9 32.6405
R19453 XThC.Tn[0].n1 XThC.Tn[0].t4 26.5955
R19454 XThC.Tn[0].n1 XThC.Tn[0].t3 26.5955
R19455 XThC.Tn[0].n0 XThC.Tn[0].t2 26.5955
R19456 XThC.Tn[0].n0 XThC.Tn[0].t1 26.5955
R19457 XThC.Tn[0].n3 XThC.Tn[0].t6 24.9236
R19458 XThC.Tn[0].n3 XThC.Tn[0].t5 24.9236
R19459 XThC.Tn[0].n4 XThC.Tn[0].t8 24.9236
R19460 XThC.Tn[0].n4 XThC.Tn[0].t7 24.9236
R19461 XThC.Tn[0].n5 XThC.Tn[0].t10 24.9236
R19462 XThC.Tn[0].n5 XThC.Tn[0].t11 24.9236
R19463 XThC.Tn[0].n6 XThC.Tn[0].t0 24.9236
R19464 XThC.Tn[0].n6 XThC.Tn[0].t9 24.9236
R19465 XThC.Tn[0].n75 XThC.Tn[0].n2 18.5605
R19466 XThC.Tn[0].n75 XThC.Tn[0].n74 11.5205
R19467 XThC.Tn[0] XThC.Tn[0].n12 8.0245
R19468 XThC.Tn[0].n72 XThC.Tn[0].n71 7.9105
R19469 XThC.Tn[0].n68 XThC.Tn[0].n67 7.9105
R19470 XThC.Tn[0].n64 XThC.Tn[0].n63 7.9105
R19471 XThC.Tn[0].n60 XThC.Tn[0].n59 7.9105
R19472 XThC.Tn[0].n56 XThC.Tn[0].n55 7.9105
R19473 XThC.Tn[0].n52 XThC.Tn[0].n51 7.9105
R19474 XThC.Tn[0].n48 XThC.Tn[0].n47 7.9105
R19475 XThC.Tn[0].n44 XThC.Tn[0].n43 7.9105
R19476 XThC.Tn[0].n40 XThC.Tn[0].n39 7.9105
R19477 XThC.Tn[0].n36 XThC.Tn[0].n35 7.9105
R19478 XThC.Tn[0].n32 XThC.Tn[0].n31 7.9105
R19479 XThC.Tn[0].n28 XThC.Tn[0].n27 7.9105
R19480 XThC.Tn[0].n24 XThC.Tn[0].n23 7.9105
R19481 XThC.Tn[0].n20 XThC.Tn[0].n19 7.9105
R19482 XThC.Tn[0].n16 XThC.Tn[0].n15 7.9105
R19483 XThC.Tn[0].n73 XThC.Tn[0] 5.95611
R19484 XThC.Tn[0].n74 XThC.Tn[0].n73 4.6005
R19485 XThC.Tn[0].n73 XThC.Tn[0] 1.89022
R19486 XThC.Tn[0] XThC.Tn[0].n75 0.6405
R19487 XThC.Tn[0].n16 XThC.Tn[0] 0.235138
R19488 XThC.Tn[0].n20 XThC.Tn[0] 0.235138
R19489 XThC.Tn[0].n24 XThC.Tn[0] 0.235138
R19490 XThC.Tn[0].n28 XThC.Tn[0] 0.235138
R19491 XThC.Tn[0].n32 XThC.Tn[0] 0.235138
R19492 XThC.Tn[0].n36 XThC.Tn[0] 0.235138
R19493 XThC.Tn[0].n40 XThC.Tn[0] 0.235138
R19494 XThC.Tn[0].n44 XThC.Tn[0] 0.235138
R19495 XThC.Tn[0].n48 XThC.Tn[0] 0.235138
R19496 XThC.Tn[0].n52 XThC.Tn[0] 0.235138
R19497 XThC.Tn[0].n56 XThC.Tn[0] 0.235138
R19498 XThC.Tn[0].n60 XThC.Tn[0] 0.235138
R19499 XThC.Tn[0].n64 XThC.Tn[0] 0.235138
R19500 XThC.Tn[0].n68 XThC.Tn[0] 0.235138
R19501 XThC.Tn[0].n72 XThC.Tn[0] 0.235138
R19502 XThC.Tn[0] XThC.Tn[0].n16 0.114505
R19503 XThC.Tn[0] XThC.Tn[0].n20 0.114505
R19504 XThC.Tn[0] XThC.Tn[0].n24 0.114505
R19505 XThC.Tn[0] XThC.Tn[0].n28 0.114505
R19506 XThC.Tn[0] XThC.Tn[0].n32 0.114505
R19507 XThC.Tn[0] XThC.Tn[0].n36 0.114505
R19508 XThC.Tn[0] XThC.Tn[0].n40 0.114505
R19509 XThC.Tn[0] XThC.Tn[0].n44 0.114505
R19510 XThC.Tn[0] XThC.Tn[0].n48 0.114505
R19511 XThC.Tn[0] XThC.Tn[0].n52 0.114505
R19512 XThC.Tn[0] XThC.Tn[0].n56 0.114505
R19513 XThC.Tn[0] XThC.Tn[0].n60 0.114505
R19514 XThC.Tn[0] XThC.Tn[0].n64 0.114505
R19515 XThC.Tn[0] XThC.Tn[0].n68 0.114505
R19516 XThC.Tn[0] XThC.Tn[0].n72 0.114505
R19517 XThC.Tn[0].n71 XThC.Tn[0].n70 0.0599512
R19518 XThC.Tn[0].n67 XThC.Tn[0].n66 0.0599512
R19519 XThC.Tn[0].n63 XThC.Tn[0].n62 0.0599512
R19520 XThC.Tn[0].n59 XThC.Tn[0].n58 0.0599512
R19521 XThC.Tn[0].n55 XThC.Tn[0].n54 0.0599512
R19522 XThC.Tn[0].n51 XThC.Tn[0].n50 0.0599512
R19523 XThC.Tn[0].n47 XThC.Tn[0].n46 0.0599512
R19524 XThC.Tn[0].n43 XThC.Tn[0].n42 0.0599512
R19525 XThC.Tn[0].n39 XThC.Tn[0].n38 0.0599512
R19526 XThC.Tn[0].n35 XThC.Tn[0].n34 0.0599512
R19527 XThC.Tn[0].n31 XThC.Tn[0].n30 0.0599512
R19528 XThC.Tn[0].n27 XThC.Tn[0].n26 0.0599512
R19529 XThC.Tn[0].n23 XThC.Tn[0].n22 0.0599512
R19530 XThC.Tn[0].n19 XThC.Tn[0].n18 0.0599512
R19531 XThC.Tn[0].n15 XThC.Tn[0].n14 0.0599512
R19532 XThC.Tn[0].n12 XThC.Tn[0].n11 0.0599512
R19533 XThC.Tn[0].n70 XThC.Tn[0] 0.0469286
R19534 XThC.Tn[0].n66 XThC.Tn[0] 0.0469286
R19535 XThC.Tn[0].n62 XThC.Tn[0] 0.0469286
R19536 XThC.Tn[0].n58 XThC.Tn[0] 0.0469286
R19537 XThC.Tn[0].n54 XThC.Tn[0] 0.0469286
R19538 XThC.Tn[0].n50 XThC.Tn[0] 0.0469286
R19539 XThC.Tn[0].n46 XThC.Tn[0] 0.0469286
R19540 XThC.Tn[0].n42 XThC.Tn[0] 0.0469286
R19541 XThC.Tn[0].n38 XThC.Tn[0] 0.0469286
R19542 XThC.Tn[0].n34 XThC.Tn[0] 0.0469286
R19543 XThC.Tn[0].n30 XThC.Tn[0] 0.0469286
R19544 XThC.Tn[0].n26 XThC.Tn[0] 0.0469286
R19545 XThC.Tn[0].n22 XThC.Tn[0] 0.0469286
R19546 XThC.Tn[0].n18 XThC.Tn[0] 0.0469286
R19547 XThC.Tn[0].n14 XThC.Tn[0] 0.0469286
R19548 XThC.Tn[0].n11 XThC.Tn[0] 0.0469286
R19549 XThC.Tn[0].n70 XThC.Tn[0] 0.0401341
R19550 XThC.Tn[0].n66 XThC.Tn[0] 0.0401341
R19551 XThC.Tn[0].n62 XThC.Tn[0] 0.0401341
R19552 XThC.Tn[0].n58 XThC.Tn[0] 0.0401341
R19553 XThC.Tn[0].n54 XThC.Tn[0] 0.0401341
R19554 XThC.Tn[0].n50 XThC.Tn[0] 0.0401341
R19555 XThC.Tn[0].n46 XThC.Tn[0] 0.0401341
R19556 XThC.Tn[0].n42 XThC.Tn[0] 0.0401341
R19557 XThC.Tn[0].n38 XThC.Tn[0] 0.0401341
R19558 XThC.Tn[0].n34 XThC.Tn[0] 0.0401341
R19559 XThC.Tn[0].n30 XThC.Tn[0] 0.0401341
R19560 XThC.Tn[0].n26 XThC.Tn[0] 0.0401341
R19561 XThC.Tn[0].n22 XThC.Tn[0] 0.0401341
R19562 XThC.Tn[0].n18 XThC.Tn[0] 0.0401341
R19563 XThC.Tn[0].n14 XThC.Tn[0] 0.0401341
R19564 XThC.Tn[0].n11 XThC.Tn[0] 0.0401341
R19565 XThC.TB4.t0 XThC.TB4.n21 268.738
R19566 XThC.TB4.n22 XThC.TB4.t0 268.077
R19567 XThC.TB4.n0 XThC.TB4.t1 235.56
R19568 XThC.TB4.n4 XThC.TB4.t3 212.081
R19569 XThC.TB4.n3 XThC.TB4.t2 212.081
R19570 XThC.TB4.n9 XThC.TB4.t17 212.081
R19571 XThC.TB4.n1 XThC.TB4.t13 212.081
R19572 XThC.TB4.n13 XThC.TB4.t8 212.081
R19573 XThC.TB4.n14 XThC.TB4.t12 212.081
R19574 XThC.TB4.n16 XThC.TB4.t6 212.081
R19575 XThC.TB4.n12 XThC.TB4.t16 212.081
R19576 XThC.TB4.n6 XThC.TB4.n5 173.761
R19577 XThC.TB4.n15 XThC.TB4 158.656
R19578 XThC.TB4.n8 XThC.TB4.n7 152
R19579 XThC.TB4.n6 XThC.TB4.n2 152
R19580 XThC.TB4.n11 XThC.TB4.n10 152
R19581 XThC.TB4.n18 XThC.TB4.n17 152
R19582 XThC.TB4.n4 XThC.TB4.t14 139.78
R19583 XThC.TB4.n3 XThC.TB4.t10 139.78
R19584 XThC.TB4.n9 XThC.TB4.t7 139.78
R19585 XThC.TB4.n1 XThC.TB4.t4 139.78
R19586 XThC.TB4.n13 XThC.TB4.t11 139.78
R19587 XThC.TB4.n14 XThC.TB4.t15 139.78
R19588 XThC.TB4.n16 XThC.TB4.t9 139.78
R19589 XThC.TB4.n12 XThC.TB4.t5 139.78
R19590 XThC.TB4.n20 XThC.TB4.n11 72.9296
R19591 XThC.TB4.n14 XThC.TB4.n13 61.346
R19592 XThC.TB4.n8 XThC.TB4.n2 49.6611
R19593 XThC.TB4.n10 XThC.TB4.n9 45.2793
R19594 XThC.TB4.n5 XThC.TB4.n3 42.3581
R19595 XThC.TB4 XThC.TB4.n19 32.9276
R19596 XThC.TB4.n17 XThC.TB4.n12 30.6732
R19597 XThC.TB4.n17 XThC.TB4.n16 30.6732
R19598 XThC.TB4.n16 XThC.TB4.n15 30.6732
R19599 XThC.TB4.n15 XThC.TB4.n14 30.6732
R19600 XThC.TB4.n7 XThC.TB4.n6 21.7605
R19601 XThC.TB4.n5 XThC.TB4.n4 18.9884
R19602 XThC.TB4 XThC.TB4.n22 17.8682
R19603 XThC.TB4.n10 XThC.TB4.n1 16.0672
R19604 XThC.TB4.n18 XThC.TB4 14.7905
R19605 XThC.TB4.n11 XThC.TB4 11.5205
R19606 XThC.TB4.n21 XThC.TB4.n20 10.353
R19607 XThC.TB4.n7 XThC.TB4 10.2405
R19608 XThC.TB4.n3 XThC.TB4.n2 7.30353
R19609 XThC.TB4.n19 XThC.TB4.n18 7.24578
R19610 XThC.TB4.n20 XThC.TB4 5.25834
R19611 XThC.TB4.n9 XThC.TB4.n8 4.38232
R19612 XThC.TB4.n22 XThC.TB4.n21 3.29747
R19613 XThC.TB4 XThC.TB4.n0 2.22659
R19614 XThC.TB4.n0 XThC.TB4 1.55202
R19615 XThC.TB4.n19 XThC.TB4 0.966538
R19616 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19617 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19618 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19619 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19620 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19621 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19622 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19623 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19624 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19625 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19626 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19627 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19628 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19629 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19630 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19631 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19632 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19633 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19634 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19635 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19636 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19637 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19638 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19639 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19640 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19641 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19642 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19643 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19644 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19645 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19646 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19647 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19648 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19649 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19650 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19651 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19652 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19653 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19654 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19655 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19656 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19657 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19658 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19659 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19660 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19661 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19662 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19663 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19664 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19665 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19666 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19667 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19668 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19669 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19670 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19671 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19672 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19673 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19674 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19675 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19676 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19677 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19678 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19679 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19680 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19681 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19682 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19683 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19684 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19685 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19686 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19687 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19688 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19689 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19690 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19691 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19692 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19693 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19694 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19695 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19696 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19697 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19698 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19699 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19700 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19701 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19702 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19703 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19704 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19705 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19706 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19707 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19708 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19709 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19710 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19711 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R19712 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19713 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19714 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R19715 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19716 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19717 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19718 XThR.Tn[3].n1 XThR.Tn[3].t4 26.5955
R19719 XThR.Tn[3].n1 XThR.Tn[3].t7 26.5955
R19720 XThR.Tn[3].n0 XThR.Tn[3].t5 26.5955
R19721 XThR.Tn[3].n0 XThR.Tn[3].t6 26.5955
R19722 XThR.Tn[3].n3 XThR.Tn[3].t11 24.9236
R19723 XThR.Tn[3].n3 XThR.Tn[3].t8 24.9236
R19724 XThR.Tn[3].n4 XThR.Tn[3].t10 24.9236
R19725 XThR.Tn[3].n4 XThR.Tn[3].t9 24.9236
R19726 XThR.Tn[3].n5 XThR.Tn[3].t0 24.9236
R19727 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19728 XThR.Tn[3].n6 XThR.Tn[3].t3 24.9236
R19729 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19730 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19731 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19732 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19733 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19734 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19735 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19736 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19737 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19738 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19739 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19740 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19741 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19742 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19743 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19744 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19745 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19746 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19747 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19748 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19749 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19750 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19751 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19752 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19753 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19754 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19755 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19756 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19757 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19758 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19759 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19760 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19761 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19762 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19763 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19764 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19765 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19766 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19767 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19768 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19769 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19770 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19771 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19772 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19773 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19774 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19775 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19776 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19777 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19778 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19779 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19780 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19781 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19782 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19783 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19784 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19785 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19786 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19787 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19788 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19789 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19790 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19791 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19792 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19793 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19794 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19795 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19796 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19797 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19798 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19799 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19800 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19801 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19802 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19803 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19804 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19805 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19806 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19807 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19808 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19809 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19810 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19811 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19812 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19813 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19814 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19815 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19816 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19817 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19818 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19819 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19820 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19821 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19822 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19823 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19824 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19825 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19826 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19827 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19828 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19829 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19830 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19831 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19832 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19833 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19834 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19835 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19836 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19837 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19838 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19839 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19840 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19841 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19842 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19843 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19844 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19845 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19846 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19847 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19848 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19849 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19850 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19851 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19852 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19853 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19854 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19855 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19856 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19857 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19858 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19859 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19860 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19861 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19862 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19863 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19864 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19865 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19866 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19867 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19868 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19869 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19870 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19871 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19872 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19873 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19874 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19875 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19876 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19877 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19878 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19879 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19880 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19881 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19882 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19883 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19884 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19885 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19886 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19887 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19888 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19889 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19890 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19891 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19892 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19893 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19894 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19895 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19896 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19897 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19898 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19899 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19900 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19901 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19902 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19903 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19904 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19905 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19906 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19907 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19908 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19909 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19910 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19911 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19912 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19913 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19914 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19915 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19916 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19917 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19918 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19919 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19920 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19921 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19922 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19923 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19924 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19925 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19926 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19927 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19928 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19929 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19930 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19931 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19932 XThR.Tn[5].n1 XThR.Tn[5].t5 26.5955
R19933 XThR.Tn[5].n1 XThR.Tn[5].t4 26.5955
R19934 XThR.Tn[5].n0 XThR.Tn[5].t6 26.5955
R19935 XThR.Tn[5].n0 XThR.Tn[5].t7 26.5955
R19936 XThR.Tn[5].n3 XThR.Tn[5].t11 24.9236
R19937 XThR.Tn[5].n3 XThR.Tn[5].t8 24.9236
R19938 XThR.Tn[5].n4 XThR.Tn[5].t10 24.9236
R19939 XThR.Tn[5].n4 XThR.Tn[5].t9 24.9236
R19940 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19941 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19942 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19943 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19944 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19945 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19946 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19947 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19948 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19949 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19950 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19951 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19952 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19953 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19954 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19955 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19956 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19957 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19958 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19959 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19960 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19961 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19962 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19963 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19964 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19965 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19966 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19967 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19968 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19969 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19970 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19971 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19972 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19973 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19974 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19975 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19976 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19977 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19978 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19979 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19980 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19981 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19982 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19983 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19984 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19985 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19986 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19987 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19988 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19989 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19990 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19991 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19992 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19993 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19994 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19995 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19996 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19997 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19998 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19999 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R20000 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R20001 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R20002 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R20003 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R20004 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R20005 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R20006 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R20007 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R20008 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R20009 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R20010 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R20011 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R20012 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R20013 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R20014 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R20015 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R20016 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R20017 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R20018 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R20019 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R20020 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R20021 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R20022 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R20023 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R20024 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R20025 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R20026 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R20027 XThR.Tn[5] XThR.Tn[5].n87 0.038
R20028 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R20029 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R20030 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R20031 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R20032 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R20033 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R20034 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R20035 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R20036 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R20037 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R20038 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R20039 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R20040 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R20041 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R20042 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R20043 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R20044 XThC.Tn[4].n73 XThC.Tn[4].n72 332.332
R20045 XThC.Tn[4].n73 XThC.Tn[4].n71 296.493
R20046 XThC.Tn[4].n68 XThC.Tn[4].n66 161.365
R20047 XThC.Tn[4].n64 XThC.Tn[4].n62 161.365
R20048 XThC.Tn[4].n60 XThC.Tn[4].n58 161.365
R20049 XThC.Tn[4].n56 XThC.Tn[4].n54 161.365
R20050 XThC.Tn[4].n52 XThC.Tn[4].n50 161.365
R20051 XThC.Tn[4].n48 XThC.Tn[4].n46 161.365
R20052 XThC.Tn[4].n44 XThC.Tn[4].n42 161.365
R20053 XThC.Tn[4].n40 XThC.Tn[4].n38 161.365
R20054 XThC.Tn[4].n36 XThC.Tn[4].n34 161.365
R20055 XThC.Tn[4].n32 XThC.Tn[4].n30 161.365
R20056 XThC.Tn[4].n28 XThC.Tn[4].n26 161.365
R20057 XThC.Tn[4].n24 XThC.Tn[4].n22 161.365
R20058 XThC.Tn[4].n20 XThC.Tn[4].n18 161.365
R20059 XThC.Tn[4].n16 XThC.Tn[4].n14 161.365
R20060 XThC.Tn[4].n12 XThC.Tn[4].n10 161.365
R20061 XThC.Tn[4].n9 XThC.Tn[4].n7 161.365
R20062 XThC.Tn[4].n66 XThC.Tn[4].t32 161.202
R20063 XThC.Tn[4].n62 XThC.Tn[4].t22 161.202
R20064 XThC.Tn[4].n58 XThC.Tn[4].t41 161.202
R20065 XThC.Tn[4].n54 XThC.Tn[4].t38 161.202
R20066 XThC.Tn[4].n50 XThC.Tn[4].t30 161.202
R20067 XThC.Tn[4].n46 XThC.Tn[4].t17 161.202
R20068 XThC.Tn[4].n42 XThC.Tn[4].t16 161.202
R20069 XThC.Tn[4].n38 XThC.Tn[4].t29 161.202
R20070 XThC.Tn[4].n34 XThC.Tn[4].t27 161.202
R20071 XThC.Tn[4].n30 XThC.Tn[4].t18 161.202
R20072 XThC.Tn[4].n26 XThC.Tn[4].t37 161.202
R20073 XThC.Tn[4].n22 XThC.Tn[4].t36 161.202
R20074 XThC.Tn[4].n18 XThC.Tn[4].t15 161.202
R20075 XThC.Tn[4].n14 XThC.Tn[4].t13 161.202
R20076 XThC.Tn[4].n10 XThC.Tn[4].t43 161.202
R20077 XThC.Tn[4].n7 XThC.Tn[4].t26 161.202
R20078 XThC.Tn[4].n66 XThC.Tn[4].t35 145.137
R20079 XThC.Tn[4].n62 XThC.Tn[4].t25 145.137
R20080 XThC.Tn[4].n58 XThC.Tn[4].t12 145.137
R20081 XThC.Tn[4].n54 XThC.Tn[4].t42 145.137
R20082 XThC.Tn[4].n50 XThC.Tn[4].t34 145.137
R20083 XThC.Tn[4].n46 XThC.Tn[4].t23 145.137
R20084 XThC.Tn[4].n42 XThC.Tn[4].t21 145.137
R20085 XThC.Tn[4].n38 XThC.Tn[4].t33 145.137
R20086 XThC.Tn[4].n34 XThC.Tn[4].t31 145.137
R20087 XThC.Tn[4].n30 XThC.Tn[4].t24 145.137
R20088 XThC.Tn[4].n26 XThC.Tn[4].t40 145.137
R20089 XThC.Tn[4].n22 XThC.Tn[4].t39 145.137
R20090 XThC.Tn[4].n18 XThC.Tn[4].t20 145.137
R20091 XThC.Tn[4].n14 XThC.Tn[4].t19 145.137
R20092 XThC.Tn[4].n10 XThC.Tn[4].t14 145.137
R20093 XThC.Tn[4].n7 XThC.Tn[4].t28 145.137
R20094 XThC.Tn[4].n2 XThC.Tn[4].n0 135.248
R20095 XThC.Tn[4].n2 XThC.Tn[4].n1 98.982
R20096 XThC.Tn[4].n4 XThC.Tn[4].n3 98.982
R20097 XThC.Tn[4].n6 XThC.Tn[4].n5 98.982
R20098 XThC.Tn[4].n4 XThC.Tn[4].n2 36.2672
R20099 XThC.Tn[4].n6 XThC.Tn[4].n4 36.2672
R20100 XThC.Tn[4].n70 XThC.Tn[4].n6 32.6405
R20101 XThC.Tn[4].n71 XThC.Tn[4].t1 26.5955
R20102 XThC.Tn[4].n71 XThC.Tn[4].t0 26.5955
R20103 XThC.Tn[4].n72 XThC.Tn[4].t3 26.5955
R20104 XThC.Tn[4].n72 XThC.Tn[4].t2 26.5955
R20105 XThC.Tn[4].n0 XThC.Tn[4].t8 24.9236
R20106 XThC.Tn[4].n0 XThC.Tn[4].t11 24.9236
R20107 XThC.Tn[4].n1 XThC.Tn[4].t10 24.9236
R20108 XThC.Tn[4].n1 XThC.Tn[4].t9 24.9236
R20109 XThC.Tn[4].n3 XThC.Tn[4].t7 24.9236
R20110 XThC.Tn[4].n3 XThC.Tn[4].t6 24.9236
R20111 XThC.Tn[4].n5 XThC.Tn[4].t5 24.9236
R20112 XThC.Tn[4].n5 XThC.Tn[4].t4 24.9236
R20113 XThC.Tn[4].n74 XThC.Tn[4].n73 18.5605
R20114 XThC.Tn[4].n74 XThC.Tn[4].n70 11.5205
R20115 XThC.Tn[4] XThC.Tn[4].n9 8.0245
R20116 XThC.Tn[4].n69 XThC.Tn[4].n68 7.9105
R20117 XThC.Tn[4].n65 XThC.Tn[4].n64 7.9105
R20118 XThC.Tn[4].n61 XThC.Tn[4].n60 7.9105
R20119 XThC.Tn[4].n57 XThC.Tn[4].n56 7.9105
R20120 XThC.Tn[4].n53 XThC.Tn[4].n52 7.9105
R20121 XThC.Tn[4].n49 XThC.Tn[4].n48 7.9105
R20122 XThC.Tn[4].n45 XThC.Tn[4].n44 7.9105
R20123 XThC.Tn[4].n41 XThC.Tn[4].n40 7.9105
R20124 XThC.Tn[4].n37 XThC.Tn[4].n36 7.9105
R20125 XThC.Tn[4].n33 XThC.Tn[4].n32 7.9105
R20126 XThC.Tn[4].n29 XThC.Tn[4].n28 7.9105
R20127 XThC.Tn[4].n25 XThC.Tn[4].n24 7.9105
R20128 XThC.Tn[4].n21 XThC.Tn[4].n20 7.9105
R20129 XThC.Tn[4].n17 XThC.Tn[4].n16 7.9105
R20130 XThC.Tn[4].n13 XThC.Tn[4].n12 7.9105
R20131 XThC.Tn[4].n70 XThC.Tn[4] 5.77342
R20132 XThC.Tn[4] XThC.Tn[4].n74 0.6405
R20133 XThC.Tn[4].n13 XThC.Tn[4] 0.235138
R20134 XThC.Tn[4].n17 XThC.Tn[4] 0.235138
R20135 XThC.Tn[4].n21 XThC.Tn[4] 0.235138
R20136 XThC.Tn[4].n25 XThC.Tn[4] 0.235138
R20137 XThC.Tn[4].n29 XThC.Tn[4] 0.235138
R20138 XThC.Tn[4].n33 XThC.Tn[4] 0.235138
R20139 XThC.Tn[4].n37 XThC.Tn[4] 0.235138
R20140 XThC.Tn[4].n41 XThC.Tn[4] 0.235138
R20141 XThC.Tn[4].n45 XThC.Tn[4] 0.235138
R20142 XThC.Tn[4].n49 XThC.Tn[4] 0.235138
R20143 XThC.Tn[4].n53 XThC.Tn[4] 0.235138
R20144 XThC.Tn[4].n57 XThC.Tn[4] 0.235138
R20145 XThC.Tn[4].n61 XThC.Tn[4] 0.235138
R20146 XThC.Tn[4].n65 XThC.Tn[4] 0.235138
R20147 XThC.Tn[4].n69 XThC.Tn[4] 0.235138
R20148 XThC.Tn[4] XThC.Tn[4].n13 0.114505
R20149 XThC.Tn[4] XThC.Tn[4].n17 0.114505
R20150 XThC.Tn[4] XThC.Tn[4].n21 0.114505
R20151 XThC.Tn[4] XThC.Tn[4].n25 0.114505
R20152 XThC.Tn[4] XThC.Tn[4].n29 0.114505
R20153 XThC.Tn[4] XThC.Tn[4].n33 0.114505
R20154 XThC.Tn[4] XThC.Tn[4].n37 0.114505
R20155 XThC.Tn[4] XThC.Tn[4].n41 0.114505
R20156 XThC.Tn[4] XThC.Tn[4].n45 0.114505
R20157 XThC.Tn[4] XThC.Tn[4].n49 0.114505
R20158 XThC.Tn[4] XThC.Tn[4].n53 0.114505
R20159 XThC.Tn[4] XThC.Tn[4].n57 0.114505
R20160 XThC.Tn[4] XThC.Tn[4].n61 0.114505
R20161 XThC.Tn[4] XThC.Tn[4].n65 0.114505
R20162 XThC.Tn[4] XThC.Tn[4].n69 0.114505
R20163 XThC.Tn[4].n68 XThC.Tn[4].n67 0.0599512
R20164 XThC.Tn[4].n64 XThC.Tn[4].n63 0.0599512
R20165 XThC.Tn[4].n60 XThC.Tn[4].n59 0.0599512
R20166 XThC.Tn[4].n56 XThC.Tn[4].n55 0.0599512
R20167 XThC.Tn[4].n52 XThC.Tn[4].n51 0.0599512
R20168 XThC.Tn[4].n48 XThC.Tn[4].n47 0.0599512
R20169 XThC.Tn[4].n44 XThC.Tn[4].n43 0.0599512
R20170 XThC.Tn[4].n40 XThC.Tn[4].n39 0.0599512
R20171 XThC.Tn[4].n36 XThC.Tn[4].n35 0.0599512
R20172 XThC.Tn[4].n32 XThC.Tn[4].n31 0.0599512
R20173 XThC.Tn[4].n28 XThC.Tn[4].n27 0.0599512
R20174 XThC.Tn[4].n24 XThC.Tn[4].n23 0.0599512
R20175 XThC.Tn[4].n20 XThC.Tn[4].n19 0.0599512
R20176 XThC.Tn[4].n16 XThC.Tn[4].n15 0.0599512
R20177 XThC.Tn[4].n12 XThC.Tn[4].n11 0.0599512
R20178 XThC.Tn[4].n9 XThC.Tn[4].n8 0.0599512
R20179 XThC.Tn[4].n67 XThC.Tn[4] 0.0469286
R20180 XThC.Tn[4].n63 XThC.Tn[4] 0.0469286
R20181 XThC.Tn[4].n59 XThC.Tn[4] 0.0469286
R20182 XThC.Tn[4].n55 XThC.Tn[4] 0.0469286
R20183 XThC.Tn[4].n51 XThC.Tn[4] 0.0469286
R20184 XThC.Tn[4].n47 XThC.Tn[4] 0.0469286
R20185 XThC.Tn[4].n43 XThC.Tn[4] 0.0469286
R20186 XThC.Tn[4].n39 XThC.Tn[4] 0.0469286
R20187 XThC.Tn[4].n35 XThC.Tn[4] 0.0469286
R20188 XThC.Tn[4].n31 XThC.Tn[4] 0.0469286
R20189 XThC.Tn[4].n27 XThC.Tn[4] 0.0469286
R20190 XThC.Tn[4].n23 XThC.Tn[4] 0.0469286
R20191 XThC.Tn[4].n19 XThC.Tn[4] 0.0469286
R20192 XThC.Tn[4].n15 XThC.Tn[4] 0.0469286
R20193 XThC.Tn[4].n11 XThC.Tn[4] 0.0469286
R20194 XThC.Tn[4].n8 XThC.Tn[4] 0.0469286
R20195 XThC.Tn[4].n67 XThC.Tn[4] 0.0401341
R20196 XThC.Tn[4].n63 XThC.Tn[4] 0.0401341
R20197 XThC.Tn[4].n59 XThC.Tn[4] 0.0401341
R20198 XThC.Tn[4].n55 XThC.Tn[4] 0.0401341
R20199 XThC.Tn[4].n51 XThC.Tn[4] 0.0401341
R20200 XThC.Tn[4].n47 XThC.Tn[4] 0.0401341
R20201 XThC.Tn[4].n43 XThC.Tn[4] 0.0401341
R20202 XThC.Tn[4].n39 XThC.Tn[4] 0.0401341
R20203 XThC.Tn[4].n35 XThC.Tn[4] 0.0401341
R20204 XThC.Tn[4].n31 XThC.Tn[4] 0.0401341
R20205 XThC.Tn[4].n27 XThC.Tn[4] 0.0401341
R20206 XThC.Tn[4].n23 XThC.Tn[4] 0.0401341
R20207 XThC.Tn[4].n19 XThC.Tn[4] 0.0401341
R20208 XThC.Tn[4].n15 XThC.Tn[4] 0.0401341
R20209 XThC.Tn[4].n11 XThC.Tn[4] 0.0401341
R20210 XThC.Tn[4].n8 XThC.Tn[4] 0.0401341
R20211 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R20212 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R20213 XThC.Tn[2].n71 XThC.Tn[2].n69 161.365
R20214 XThC.Tn[2].n67 XThC.Tn[2].n65 161.365
R20215 XThC.Tn[2].n63 XThC.Tn[2].n61 161.365
R20216 XThC.Tn[2].n59 XThC.Tn[2].n57 161.365
R20217 XThC.Tn[2].n55 XThC.Tn[2].n53 161.365
R20218 XThC.Tn[2].n51 XThC.Tn[2].n49 161.365
R20219 XThC.Tn[2].n47 XThC.Tn[2].n45 161.365
R20220 XThC.Tn[2].n43 XThC.Tn[2].n41 161.365
R20221 XThC.Tn[2].n39 XThC.Tn[2].n37 161.365
R20222 XThC.Tn[2].n35 XThC.Tn[2].n33 161.365
R20223 XThC.Tn[2].n31 XThC.Tn[2].n29 161.365
R20224 XThC.Tn[2].n27 XThC.Tn[2].n25 161.365
R20225 XThC.Tn[2].n23 XThC.Tn[2].n21 161.365
R20226 XThC.Tn[2].n19 XThC.Tn[2].n17 161.365
R20227 XThC.Tn[2].n15 XThC.Tn[2].n13 161.365
R20228 XThC.Tn[2].n12 XThC.Tn[2].n10 161.365
R20229 XThC.Tn[2].n69 XThC.Tn[2].t24 161.202
R20230 XThC.Tn[2].n65 XThC.Tn[2].t14 161.202
R20231 XThC.Tn[2].n61 XThC.Tn[2].t33 161.202
R20232 XThC.Tn[2].n57 XThC.Tn[2].t30 161.202
R20233 XThC.Tn[2].n53 XThC.Tn[2].t22 161.202
R20234 XThC.Tn[2].n49 XThC.Tn[2].t41 161.202
R20235 XThC.Tn[2].n45 XThC.Tn[2].t40 161.202
R20236 XThC.Tn[2].n41 XThC.Tn[2].t21 161.202
R20237 XThC.Tn[2].n37 XThC.Tn[2].t19 161.202
R20238 XThC.Tn[2].n33 XThC.Tn[2].t42 161.202
R20239 XThC.Tn[2].n29 XThC.Tn[2].t29 161.202
R20240 XThC.Tn[2].n25 XThC.Tn[2].t28 161.202
R20241 XThC.Tn[2].n21 XThC.Tn[2].t39 161.202
R20242 XThC.Tn[2].n17 XThC.Tn[2].t37 161.202
R20243 XThC.Tn[2].n13 XThC.Tn[2].t35 161.202
R20244 XThC.Tn[2].n10 XThC.Tn[2].t18 161.202
R20245 XThC.Tn[2].n69 XThC.Tn[2].t27 145.137
R20246 XThC.Tn[2].n65 XThC.Tn[2].t17 145.137
R20247 XThC.Tn[2].n61 XThC.Tn[2].t36 145.137
R20248 XThC.Tn[2].n57 XThC.Tn[2].t34 145.137
R20249 XThC.Tn[2].n53 XThC.Tn[2].t26 145.137
R20250 XThC.Tn[2].n49 XThC.Tn[2].t15 145.137
R20251 XThC.Tn[2].n45 XThC.Tn[2].t13 145.137
R20252 XThC.Tn[2].n41 XThC.Tn[2].t25 145.137
R20253 XThC.Tn[2].n37 XThC.Tn[2].t23 145.137
R20254 XThC.Tn[2].n33 XThC.Tn[2].t16 145.137
R20255 XThC.Tn[2].n29 XThC.Tn[2].t32 145.137
R20256 XThC.Tn[2].n25 XThC.Tn[2].t31 145.137
R20257 XThC.Tn[2].n21 XThC.Tn[2].t12 145.137
R20258 XThC.Tn[2].n17 XThC.Tn[2].t43 145.137
R20259 XThC.Tn[2].n13 XThC.Tn[2].t38 145.137
R20260 XThC.Tn[2].n10 XThC.Tn[2].t20 145.137
R20261 XThC.Tn[2].n7 XThC.Tn[2].n6 135.248
R20262 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R20263 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R20264 XThC.Tn[2].n7 XThC.Tn[2].n5 98.982
R20265 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R20266 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R20267 XThC.Tn[2].n74 XThC.Tn[2].n9 32.6405
R20268 XThC.Tn[2].n1 XThC.Tn[2].t5 26.5955
R20269 XThC.Tn[2].n1 XThC.Tn[2].t4 26.5955
R20270 XThC.Tn[2].n0 XThC.Tn[2].t7 26.5955
R20271 XThC.Tn[2].n0 XThC.Tn[2].t6 26.5955
R20272 XThC.Tn[2].n3 XThC.Tn[2].t11 24.9236
R20273 XThC.Tn[2].n3 XThC.Tn[2].t10 24.9236
R20274 XThC.Tn[2].n4 XThC.Tn[2].t9 24.9236
R20275 XThC.Tn[2].n4 XThC.Tn[2].t8 24.9236
R20276 XThC.Tn[2].n5 XThC.Tn[2].t1 24.9236
R20277 XThC.Tn[2].n5 XThC.Tn[2].t2 24.9236
R20278 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R20279 XThC.Tn[2].n6 XThC.Tn[2].t3 24.9236
R20280 XThC.Tn[2].n75 XThC.Tn[2].n2 18.5605
R20281 XThC.Tn[2].n75 XThC.Tn[2].n74 11.5205
R20282 XThC.Tn[2] XThC.Tn[2].n12 8.0245
R20283 XThC.Tn[2].n72 XThC.Tn[2].n71 7.9105
R20284 XThC.Tn[2].n68 XThC.Tn[2].n67 7.9105
R20285 XThC.Tn[2].n64 XThC.Tn[2].n63 7.9105
R20286 XThC.Tn[2].n60 XThC.Tn[2].n59 7.9105
R20287 XThC.Tn[2].n56 XThC.Tn[2].n55 7.9105
R20288 XThC.Tn[2].n52 XThC.Tn[2].n51 7.9105
R20289 XThC.Tn[2].n48 XThC.Tn[2].n47 7.9105
R20290 XThC.Tn[2].n44 XThC.Tn[2].n43 7.9105
R20291 XThC.Tn[2].n40 XThC.Tn[2].n39 7.9105
R20292 XThC.Tn[2].n36 XThC.Tn[2].n35 7.9105
R20293 XThC.Tn[2].n32 XThC.Tn[2].n31 7.9105
R20294 XThC.Tn[2].n28 XThC.Tn[2].n27 7.9105
R20295 XThC.Tn[2].n24 XThC.Tn[2].n23 7.9105
R20296 XThC.Tn[2].n20 XThC.Tn[2].n19 7.9105
R20297 XThC.Tn[2].n16 XThC.Tn[2].n15 7.9105
R20298 XThC.Tn[2].n73 XThC.Tn[2] 5.58686
R20299 XThC.Tn[2].n74 XThC.Tn[2].n73 4.6005
R20300 XThC.Tn[2].n73 XThC.Tn[2] 1.83383
R20301 XThC.Tn[2] XThC.Tn[2].n75 0.6405
R20302 XThC.Tn[2].n16 XThC.Tn[2] 0.235138
R20303 XThC.Tn[2].n20 XThC.Tn[2] 0.235138
R20304 XThC.Tn[2].n24 XThC.Tn[2] 0.235138
R20305 XThC.Tn[2].n28 XThC.Tn[2] 0.235138
R20306 XThC.Tn[2].n32 XThC.Tn[2] 0.235138
R20307 XThC.Tn[2].n36 XThC.Tn[2] 0.235138
R20308 XThC.Tn[2].n40 XThC.Tn[2] 0.235138
R20309 XThC.Tn[2].n44 XThC.Tn[2] 0.235138
R20310 XThC.Tn[2].n48 XThC.Tn[2] 0.235138
R20311 XThC.Tn[2].n52 XThC.Tn[2] 0.235138
R20312 XThC.Tn[2].n56 XThC.Tn[2] 0.235138
R20313 XThC.Tn[2].n60 XThC.Tn[2] 0.235138
R20314 XThC.Tn[2].n64 XThC.Tn[2] 0.235138
R20315 XThC.Tn[2].n68 XThC.Tn[2] 0.235138
R20316 XThC.Tn[2].n72 XThC.Tn[2] 0.235138
R20317 XThC.Tn[2] XThC.Tn[2].n16 0.114505
R20318 XThC.Tn[2] XThC.Tn[2].n20 0.114505
R20319 XThC.Tn[2] XThC.Tn[2].n24 0.114505
R20320 XThC.Tn[2] XThC.Tn[2].n28 0.114505
R20321 XThC.Tn[2] XThC.Tn[2].n32 0.114505
R20322 XThC.Tn[2] XThC.Tn[2].n36 0.114505
R20323 XThC.Tn[2] XThC.Tn[2].n40 0.114505
R20324 XThC.Tn[2] XThC.Tn[2].n44 0.114505
R20325 XThC.Tn[2] XThC.Tn[2].n48 0.114505
R20326 XThC.Tn[2] XThC.Tn[2].n52 0.114505
R20327 XThC.Tn[2] XThC.Tn[2].n56 0.114505
R20328 XThC.Tn[2] XThC.Tn[2].n60 0.114505
R20329 XThC.Tn[2] XThC.Tn[2].n64 0.114505
R20330 XThC.Tn[2] XThC.Tn[2].n68 0.114505
R20331 XThC.Tn[2] XThC.Tn[2].n72 0.114505
R20332 XThC.Tn[2].n71 XThC.Tn[2].n70 0.0599512
R20333 XThC.Tn[2].n67 XThC.Tn[2].n66 0.0599512
R20334 XThC.Tn[2].n63 XThC.Tn[2].n62 0.0599512
R20335 XThC.Tn[2].n59 XThC.Tn[2].n58 0.0599512
R20336 XThC.Tn[2].n55 XThC.Tn[2].n54 0.0599512
R20337 XThC.Tn[2].n51 XThC.Tn[2].n50 0.0599512
R20338 XThC.Tn[2].n47 XThC.Tn[2].n46 0.0599512
R20339 XThC.Tn[2].n43 XThC.Tn[2].n42 0.0599512
R20340 XThC.Tn[2].n39 XThC.Tn[2].n38 0.0599512
R20341 XThC.Tn[2].n35 XThC.Tn[2].n34 0.0599512
R20342 XThC.Tn[2].n31 XThC.Tn[2].n30 0.0599512
R20343 XThC.Tn[2].n27 XThC.Tn[2].n26 0.0599512
R20344 XThC.Tn[2].n23 XThC.Tn[2].n22 0.0599512
R20345 XThC.Tn[2].n19 XThC.Tn[2].n18 0.0599512
R20346 XThC.Tn[2].n15 XThC.Tn[2].n14 0.0599512
R20347 XThC.Tn[2].n12 XThC.Tn[2].n11 0.0599512
R20348 XThC.Tn[2].n70 XThC.Tn[2] 0.0469286
R20349 XThC.Tn[2].n66 XThC.Tn[2] 0.0469286
R20350 XThC.Tn[2].n62 XThC.Tn[2] 0.0469286
R20351 XThC.Tn[2].n58 XThC.Tn[2] 0.0469286
R20352 XThC.Tn[2].n54 XThC.Tn[2] 0.0469286
R20353 XThC.Tn[2].n50 XThC.Tn[2] 0.0469286
R20354 XThC.Tn[2].n46 XThC.Tn[2] 0.0469286
R20355 XThC.Tn[2].n42 XThC.Tn[2] 0.0469286
R20356 XThC.Tn[2].n38 XThC.Tn[2] 0.0469286
R20357 XThC.Tn[2].n34 XThC.Tn[2] 0.0469286
R20358 XThC.Tn[2].n30 XThC.Tn[2] 0.0469286
R20359 XThC.Tn[2].n26 XThC.Tn[2] 0.0469286
R20360 XThC.Tn[2].n22 XThC.Tn[2] 0.0469286
R20361 XThC.Tn[2].n18 XThC.Tn[2] 0.0469286
R20362 XThC.Tn[2].n14 XThC.Tn[2] 0.0469286
R20363 XThC.Tn[2].n11 XThC.Tn[2] 0.0469286
R20364 XThC.Tn[2].n70 XThC.Tn[2] 0.0401341
R20365 XThC.Tn[2].n66 XThC.Tn[2] 0.0401341
R20366 XThC.Tn[2].n62 XThC.Tn[2] 0.0401341
R20367 XThC.Tn[2].n58 XThC.Tn[2] 0.0401341
R20368 XThC.Tn[2].n54 XThC.Tn[2] 0.0401341
R20369 XThC.Tn[2].n50 XThC.Tn[2] 0.0401341
R20370 XThC.Tn[2].n46 XThC.Tn[2] 0.0401341
R20371 XThC.Tn[2].n42 XThC.Tn[2] 0.0401341
R20372 XThC.Tn[2].n38 XThC.Tn[2] 0.0401341
R20373 XThC.Tn[2].n34 XThC.Tn[2] 0.0401341
R20374 XThC.Tn[2].n30 XThC.Tn[2] 0.0401341
R20375 XThC.Tn[2].n26 XThC.Tn[2] 0.0401341
R20376 XThC.Tn[2].n22 XThC.Tn[2] 0.0401341
R20377 XThC.Tn[2].n18 XThC.Tn[2] 0.0401341
R20378 XThC.Tn[2].n14 XThC.Tn[2] 0.0401341
R20379 XThC.Tn[2].n11 XThC.Tn[2] 0.0401341
R20380 Vbias.n1 Vbias.t5 651.571
R20381 Vbias.n1 Vbias.t3 651.571
R20382 Vbias.n2 Vbias.t0 651.571
R20383 Vbias.n2 Vbias.t4 651.571
R20384 Vbias.n337 Vbias.t261 119.309
R20385 Vbias.n383 Vbias.t194 119.309
R20386 Vbias.n384 Vbias.t61 119.309
R20387 Vbias.n334 Vbias.t215 119.309
R20388 Vbias.n292 Vbias.t86 119.309
R20389 Vbias.n284 Vbias.t186 119.309
R20390 Vbias.n288 Vbias.t109 119.309
R20391 Vbias.n280 Vbias.t189 119.309
R20392 Vbias.n194 Vbias.t64 119.309
R20393 Vbias.n149 Vbias.t82 119.309
R20394 Vbias.n189 Vbias.t105 119.309
R20395 Vbias.n145 Vbias.t121 119.309
R20396 Vbias.n679 Vbias.t255 119.309
R20397 Vbias.n102 Vbias.t16 119.309
R20398 Vbias.n10 Vbias.t146 119.309
R20399 Vbias.n57 Vbias.t57 119.309
R20400 Vbias.n58 Vbias.t129 119.309
R20401 Vbias.n54 Vbias.t201 119.309
R20402 Vbias.n441 Vbias.t79 119.309
R20403 Vbias.n343 Vbias.t216 119.309
R20404 Vbias.n333 Vbias.t31 119.309
R20405 Vbias.n331 Vbias.t100 119.309
R20406 Vbias.n578 Vbias.t6 119.309
R20407 Vbias.n278 Vbias.t128 119.309
R20408 Vbias.n276 Vbias.t10 119.309
R20409 Vbias.n197 Vbias.t83 119.309
R20410 Vbias.n150 Vbias.t154 119.309
R20411 Vbias.n152 Vbias.t122 119.309
R20412 Vbias.n790 Vbias.t195 119.309
R20413 Vbias.n105 Vbias.t17 119.309
R20414 Vbias.n103 Vbias.t88 119.309
R20415 Vbias.n97 Vbias.t160 119.309
R20416 Vbias.n56 Vbias.t130 119.309
R20417 Vbias.n53 Vbias.t41 119.309
R20418 Vbias.n438 Vbias.t174 119.309
R20419 Vbias.n346 Vbias.t59 119.309
R20420 Vbias.n326 Vbias.t132 119.309
R20421 Vbias.n328 Vbias.t203 119.309
R20422 Vbias.n575 Vbias.t103 119.309
R20423 Vbias.n273 Vbias.t226 119.309
R20424 Vbias.n275 Vbias.t108 119.309
R20425 Vbias.n200 Vbias.t180 119.309
R20426 Vbias.n155 Vbias.t257 119.309
R20427 Vbias.n153 Vbias.t222 119.309
R20428 Vbias.n793 Vbias.t37 119.309
R20429 Vbias.n106 Vbias.t113 119.309
R20430 Vbias.n108 Vbias.t185 119.309
R20431 Vbias.n94 Vbias.t262 119.309
R20432 Vbias.n51 Vbias.t229 119.309
R20433 Vbias.n48 Vbias.t56 119.309
R20434 Vbias.n435 Vbias.t182 119.309
R20435 Vbias.n349 Vbias.t67 119.309
R20436 Vbias.n325 Vbias.t139 119.309
R20437 Vbias.n323 Vbias.t214 119.309
R20438 Vbias.n572 Vbias.t115 119.309
R20439 Vbias.n272 Vbias.t241 119.309
R20440 Vbias.n270 Vbias.t117 119.309
R20441 Vbias.n203 Vbias.t188 119.309
R20442 Vbias.n156 Vbias.t8 119.309
R20443 Vbias.n158 Vbias.t235 119.309
R20444 Vbias.n796 Vbias.t48 119.309
R20445 Vbias.n111 Vbias.t124 119.309
R20446 Vbias.n109 Vbias.t196 119.309
R20447 Vbias.n91 Vbias.t14 119.309
R20448 Vbias.n50 Vbias.t242 119.309
R20449 Vbias.n47 Vbias.t141 119.309
R20450 Vbias.n432 Vbias.t15 119.309
R20451 Vbias.n352 Vbias.t152 119.309
R20452 Vbias.n320 Vbias.t224 119.309
R20453 Vbias.n322 Vbias.t38 119.309
R20454 Vbias.n569 Vbias.t206 119.309
R20455 Vbias.n267 Vbias.t66 119.309
R20456 Vbias.n269 Vbias.t208 119.309
R20457 Vbias.n206 Vbias.t23 119.309
R20458 Vbias.n161 Vbias.t93 119.309
R20459 Vbias.n159 Vbias.t63 119.309
R20460 Vbias.n799 Vbias.t135 119.309
R20461 Vbias.n112 Vbias.t213 119.309
R20462 Vbias.n114 Vbias.t29 119.309
R20463 Vbias.n88 Vbias.t99 119.309
R20464 Vbias.n45 Vbias.t69 119.309
R20465 Vbias.n42 Vbias.t227 119.309
R20466 Vbias.n429 Vbias.t101 119.309
R20467 Vbias.n355 Vbias.t245 119.309
R20468 Vbias.n319 Vbias.t58 119.309
R20469 Vbias.n317 Vbias.t131 119.309
R20470 Vbias.n566 Vbias.t34 119.309
R20471 Vbias.n266 Vbias.t155 119.309
R20472 Vbias.n264 Vbias.t36 119.309
R20473 Vbias.n209 Vbias.t107 119.309
R20474 Vbias.n162 Vbias.t179 119.309
R20475 Vbias.n164 Vbias.t150 119.309
R20476 Vbias.n802 Vbias.t221 119.309
R20477 Vbias.n117 Vbias.t40 119.309
R20478 Vbias.n115 Vbias.t112 119.309
R20479 Vbias.n85 Vbias.t183 119.309
R20480 Vbias.n44 Vbias.t156 119.309
R20481 Vbias.n41 Vbias.t60 119.309
R20482 Vbias.n426 Vbias.t184 119.309
R20483 Vbias.n358 Vbias.t72 119.309
R20484 Vbias.n314 Vbias.t145 119.309
R20485 Vbias.n316 Vbias.t218 119.309
R20486 Vbias.n563 Vbias.t116 119.309
R20487 Vbias.n261 Vbias.t244 119.309
R20488 Vbias.n263 Vbias.t120 119.309
R20489 Vbias.n212 Vbias.t192 119.309
R20490 Vbias.n167 Vbias.t11 119.309
R20491 Vbias.n165 Vbias.t237 119.309
R20492 Vbias.n805 Vbias.t50 119.309
R20493 Vbias.n118 Vbias.t127 119.309
R20494 Vbias.n120 Vbias.t200 119.309
R20495 Vbias.n82 Vbias.t18 119.309
R20496 Vbias.n39 Vbias.t247 119.309
R20497 Vbias.n36 Vbias.t147 119.309
R20498 Vbias.n423 Vbias.t19 119.309
R20499 Vbias.n361 Vbias.t158 119.309
R20500 Vbias.n313 Vbias.t230 119.309
R20501 Vbias.n311 Vbias.t42 119.309
R20502 Vbias.n560 Vbias.t209 119.309
R20503 Vbias.n260 Vbias.t74 119.309
R20504 Vbias.n258 Vbias.t212 119.309
R20505 Vbias.n215 Vbias.t28 119.309
R20506 Vbias.n168 Vbias.t98 119.309
R20507 Vbias.n170 Vbias.t68 119.309
R20508 Vbias.n808 Vbias.t138 119.309
R20509 Vbias.n123 Vbias.t219 119.309
R20510 Vbias.n121 Vbias.t33 119.309
R20511 Vbias.n79 Vbias.t102 119.309
R20512 Vbias.n38 Vbias.t76 119.309
R20513 Vbias.n35 Vbias.t169 119.309
R20514 Vbias.n420 Vbias.t39 119.309
R20515 Vbias.n364 Vbias.t178 119.309
R20516 Vbias.n308 Vbias.t253 119.309
R20517 Vbias.n310 Vbias.t70 119.309
R20518 Vbias.n557 Vbias.t231 119.309
R20519 Vbias.n255 Vbias.t94 119.309
R20520 Vbias.n257 Vbias.t234 119.309
R20521 Vbias.n218 Vbias.t45 119.309
R20522 Vbias.n173 Vbias.t118 119.309
R20523 Vbias.n171 Vbias.t91 119.309
R20524 Vbias.n811 Vbias.t163 119.309
R20525 Vbias.n124 Vbias.t240 119.309
R20526 Vbias.n126 Vbias.t53 119.309
R20527 Vbias.n76 Vbias.t125 119.309
R20528 Vbias.n33 Vbias.t96 119.309
R20529 Vbias.n30 Vbias.t246 119.309
R20530 Vbias.n417 Vbias.t111 119.309
R20531 Vbias.n367 Vbias.t254 119.309
R20532 Vbias.n307 Vbias.t71 119.309
R20533 Vbias.n305 Vbias.t143 119.309
R20534 Vbias.n554 Vbias.t43 119.309
R20535 Vbias.n254 Vbias.t167 119.309
R20536 Vbias.n252 Vbias.t46 119.309
R20537 Vbias.n221 Vbias.t119 119.309
R20538 Vbias.n174 Vbias.t190 119.309
R20539 Vbias.n176 Vbias.t164 119.309
R20540 Vbias.n814 Vbias.t236 119.309
R20541 Vbias.n129 Vbias.t54 119.309
R20542 Vbias.n127 Vbias.t126 119.309
R20543 Vbias.n73 Vbias.t199 119.309
R20544 Vbias.n32 Vbias.t171 119.309
R20545 Vbias.n29 Vbias.t75 119.309
R20546 Vbias.n414 Vbias.t202 119.309
R20547 Vbias.n370 Vbias.t84 119.309
R20548 Vbias.n302 Vbias.t157 119.309
R20549 Vbias.n304 Vbias.t228 119.309
R20550 Vbias.n551 Vbias.t134 119.309
R20551 Vbias.n249 Vbias.t256 119.309
R20552 Vbias.n251 Vbias.t136 119.309
R20553 Vbias.n224 Vbias.t211 119.309
R20554 Vbias.n179 Vbias.t27 119.309
R20555 Vbias.n177 Vbias.t251 119.309
R20556 Vbias.n817 Vbias.t65 119.309
R20557 Vbias.n130 Vbias.t144 119.309
R20558 Vbias.n132 Vbias.t217 119.309
R20559 Vbias.n70 Vbias.t32 119.309
R20560 Vbias.n27 Vbias.t258 119.309
R20561 Vbias.n24 Vbias.t95 119.309
R20562 Vbias.n411 Vbias.t223 119.309
R20563 Vbias.n373 Vbias.t106 119.309
R20564 Vbias.n301 Vbias.t177 119.309
R20565 Vbias.n299 Vbias.t252 119.309
R20566 Vbias.n548 Vbias.t159 119.309
R20567 Vbias.n248 Vbias.t22 119.309
R20568 Vbias.n246 Vbias.t162 119.309
R20569 Vbias.n227 Vbias.t233 119.309
R20570 Vbias.n180 Vbias.t44 119.309
R20571 Vbias.n182 Vbias.t21 119.309
R20572 Vbias.n820 Vbias.t90 119.309
R20573 Vbias.n135 Vbias.t166 119.309
R20574 Vbias.n133 Vbias.t239 119.309
R20575 Vbias.n67 Vbias.t52 119.309
R20576 Vbias.n26 Vbias.t25 119.309
R20577 Vbias.n23 Vbias.t248 119.309
R20578 Vbias.n408 Vbias.t114 119.309
R20579 Vbias.n376 Vbias.t259 119.309
R20580 Vbias.n296 Vbias.t77 119.309
R20581 Vbias.n298 Vbias.t148 119.309
R20582 Vbias.n545 Vbias.t47 119.309
R20583 Vbias.n243 Vbias.t172 119.309
R20584 Vbias.n245 Vbias.t51 119.309
R20585 Vbias.n230 Vbias.t123 119.309
R20586 Vbias.n185 Vbias.t197 119.309
R20587 Vbias.n183 Vbias.t168 119.309
R20588 Vbias.n823 Vbias.t243 119.309
R20589 Vbias.n136 Vbias.t62 119.309
R20590 Vbias.n138 Vbias.t133 119.309
R20591 Vbias.n64 Vbias.t205 119.309
R20592 Vbias.n21 Vbias.t173 119.309
R20593 Vbias.n16 Vbias.t12 119.309
R20594 Vbias.n405 Vbias.t142 119.309
R20595 Vbias.n379 Vbias.t26 119.309
R20596 Vbias.n295 Vbias.t97 119.309
R20597 Vbias.n293 Vbias.t170 119.309
R20598 Vbias.n542 Vbias.t78 119.309
R20599 Vbias.n242 Vbias.t191 119.309
R20600 Vbias.n240 Vbias.t80 119.309
R20601 Vbias.n233 Vbias.t149 119.309
R20602 Vbias.n186 Vbias.t220 119.309
R20603 Vbias.n188 Vbias.t187 119.309
R20604 Vbias.n826 Vbias.t7 119.309
R20605 Vbias.n141 Vbias.t81 119.309
R20606 Vbias.n139 Vbias.t153 119.309
R20607 Vbias.n61 Vbias.t225 119.309
R20608 Vbias.n18 Vbias.t193 119.309
R20609 Vbias.n15 Vbias.t24 119.309
R20610 Vbias.n338 Vbias.t151 119.309
R20611 Vbias.n339 Vbias.t35 119.309
R20612 Vbias.n341 Vbias.t104 119.309
R20613 Vbias.n526 Vbias.t175 119.309
R20614 Vbias.n285 Vbias.t85 119.309
R20615 Vbias.n287 Vbias.t207 119.309
R20616 Vbias.n663 Vbias.t89 119.309
R20617 Vbias.n236 Vbias.t161 119.309
R20618 Vbias.n238 Vbias.t232 119.309
R20619 Vbias.n704 Vbias.t204 119.309
R20620 Vbias.n144 Vbias.t20 119.309
R20621 Vbias.n142 Vbias.t92 119.309
R20622 Vbias.n672 Vbias.t165 119.309
R20623 Vbias.n11 Vbias.t238 119.309
R20624 Vbias.n13 Vbias.t210 119.309
R20625 Vbias.n6 Vbias.t181 119.309
R20626 Vbias.n7 Vbias.t110 119.309
R20627 Vbias.n60 Vbias.t87 119.309
R20628 Vbias.n675 Vbias.t73 119.309
R20629 Vbias.n907 Vbias.t198 119.309
R20630 Vbias.n684 Vbias.t176 119.309
R20631 Vbias.n146 Vbias.t49 119.309
R20632 Vbias.n191 Vbias.t137 119.309
R20633 Vbias.n195 Vbias.t9 119.309
R20634 Vbias.n666 Vbias.t250 119.309
R20635 Vbias.n279 Vbias.t55 119.309
R20636 Vbias.n289 Vbias.t249 119.309
R20637 Vbias.n329 Vbias.t30 119.309
R20638 Vbias.n396 Vbias.t13 119.309
R20639 Vbias.n335 Vbias.t140 119.309
R20640 Vbias.n0 Vbias.t1 77.1834
R20641 Vbias.n0 Vbias.t2 34.3787
R20642 Vbias.n3 Vbias.n1 4.78773
R20643 Vbias.n3 Vbias.n2 4.78773
R20644 Vbias.n387 Vbias.n384 4.5005
R20645 Vbias.n442 Vbias.n441 4.5005
R20646 Vbias.n344 Vbias.n343 4.5005
R20647 Vbias.n449 Vbias.n333 4.5005
R20648 Vbias.n452 Vbias.n331 4.5005
R20649 Vbias.n579 Vbias.n578 4.5005
R20650 Vbias.n586 Vbias.n278 4.5005
R20651 Vbias.n589 Vbias.n276 4.5005
R20652 Vbias.n198 Vbias.n197 4.5005
R20653 Vbias.n783 Vbias.n150 4.5005
R20654 Vbias.n780 Vbias.n152 4.5005
R20655 Vbias.n791 Vbias.n790 4.5005
R20656 Vbias.n910 Vbias.n105 4.5005
R20657 Vbias.n913 Vbias.n103 4.5005
R20658 Vbias.n98 Vbias.n97 4.5005
R20659 Vbias.n921 Vbias.n56 4.5005
R20660 Vbias.n923 Vbias.n54 4.5005
R20661 Vbias.n439 Vbias.n438 4.5005
R20662 Vbias.n347 Vbias.n346 4.5005
R20663 Vbias.n458 Vbias.n326 4.5005
R20664 Vbias.n455 Vbias.n328 4.5005
R20665 Vbias.n576 Vbias.n575 4.5005
R20666 Vbias.n595 Vbias.n273 4.5005
R20667 Vbias.n592 Vbias.n275 4.5005
R20668 Vbias.n201 Vbias.n200 4.5005
R20669 Vbias.n774 Vbias.n155 4.5005
R20670 Vbias.n777 Vbias.n153 4.5005
R20671 Vbias.n794 Vbias.n793 4.5005
R20672 Vbias.n905 Vbias.n106 4.5005
R20673 Vbias.n902 Vbias.n108 4.5005
R20674 Vbias.n95 Vbias.n94 4.5005
R20675 Vbias.n928 Vbias.n51 4.5005
R20676 Vbias.n926 Vbias.n53 4.5005
R20677 Vbias.n436 Vbias.n435 4.5005
R20678 Vbias.n350 Vbias.n349 4.5005
R20679 Vbias.n461 Vbias.n325 4.5005
R20680 Vbias.n464 Vbias.n323 4.5005
R20681 Vbias.n573 Vbias.n572 4.5005
R20682 Vbias.n598 Vbias.n272 4.5005
R20683 Vbias.n601 Vbias.n270 4.5005
R20684 Vbias.n204 Vbias.n203 4.5005
R20685 Vbias.n771 Vbias.n156 4.5005
R20686 Vbias.n768 Vbias.n158 4.5005
R20687 Vbias.n797 Vbias.n796 4.5005
R20688 Vbias.n896 Vbias.n111 4.5005
R20689 Vbias.n899 Vbias.n109 4.5005
R20690 Vbias.n92 Vbias.n91 4.5005
R20691 Vbias.n931 Vbias.n50 4.5005
R20692 Vbias.n933 Vbias.n48 4.5005
R20693 Vbias.n433 Vbias.n432 4.5005
R20694 Vbias.n353 Vbias.n352 4.5005
R20695 Vbias.n470 Vbias.n320 4.5005
R20696 Vbias.n467 Vbias.n322 4.5005
R20697 Vbias.n570 Vbias.n569 4.5005
R20698 Vbias.n607 Vbias.n267 4.5005
R20699 Vbias.n604 Vbias.n269 4.5005
R20700 Vbias.n207 Vbias.n206 4.5005
R20701 Vbias.n762 Vbias.n161 4.5005
R20702 Vbias.n765 Vbias.n159 4.5005
R20703 Vbias.n800 Vbias.n799 4.5005
R20704 Vbias.n893 Vbias.n112 4.5005
R20705 Vbias.n890 Vbias.n114 4.5005
R20706 Vbias.n89 Vbias.n88 4.5005
R20707 Vbias.n938 Vbias.n45 4.5005
R20708 Vbias.n936 Vbias.n47 4.5005
R20709 Vbias.n430 Vbias.n429 4.5005
R20710 Vbias.n356 Vbias.n355 4.5005
R20711 Vbias.n473 Vbias.n319 4.5005
R20712 Vbias.n476 Vbias.n317 4.5005
R20713 Vbias.n567 Vbias.n566 4.5005
R20714 Vbias.n610 Vbias.n266 4.5005
R20715 Vbias.n613 Vbias.n264 4.5005
R20716 Vbias.n210 Vbias.n209 4.5005
R20717 Vbias.n759 Vbias.n162 4.5005
R20718 Vbias.n756 Vbias.n164 4.5005
R20719 Vbias.n803 Vbias.n802 4.5005
R20720 Vbias.n884 Vbias.n117 4.5005
R20721 Vbias.n887 Vbias.n115 4.5005
R20722 Vbias.n86 Vbias.n85 4.5005
R20723 Vbias.n941 Vbias.n44 4.5005
R20724 Vbias.n943 Vbias.n42 4.5005
R20725 Vbias.n427 Vbias.n426 4.5005
R20726 Vbias.n359 Vbias.n358 4.5005
R20727 Vbias.n482 Vbias.n314 4.5005
R20728 Vbias.n479 Vbias.n316 4.5005
R20729 Vbias.n564 Vbias.n563 4.5005
R20730 Vbias.n619 Vbias.n261 4.5005
R20731 Vbias.n616 Vbias.n263 4.5005
R20732 Vbias.n213 Vbias.n212 4.5005
R20733 Vbias.n750 Vbias.n167 4.5005
R20734 Vbias.n753 Vbias.n165 4.5005
R20735 Vbias.n806 Vbias.n805 4.5005
R20736 Vbias.n881 Vbias.n118 4.5005
R20737 Vbias.n878 Vbias.n120 4.5005
R20738 Vbias.n83 Vbias.n82 4.5005
R20739 Vbias.n948 Vbias.n39 4.5005
R20740 Vbias.n946 Vbias.n41 4.5005
R20741 Vbias.n424 Vbias.n423 4.5005
R20742 Vbias.n362 Vbias.n361 4.5005
R20743 Vbias.n485 Vbias.n313 4.5005
R20744 Vbias.n488 Vbias.n311 4.5005
R20745 Vbias.n561 Vbias.n560 4.5005
R20746 Vbias.n622 Vbias.n260 4.5005
R20747 Vbias.n625 Vbias.n258 4.5005
R20748 Vbias.n216 Vbias.n215 4.5005
R20749 Vbias.n747 Vbias.n168 4.5005
R20750 Vbias.n744 Vbias.n170 4.5005
R20751 Vbias.n809 Vbias.n808 4.5005
R20752 Vbias.n872 Vbias.n123 4.5005
R20753 Vbias.n875 Vbias.n121 4.5005
R20754 Vbias.n80 Vbias.n79 4.5005
R20755 Vbias.n951 Vbias.n38 4.5005
R20756 Vbias.n953 Vbias.n36 4.5005
R20757 Vbias.n421 Vbias.n420 4.5005
R20758 Vbias.n365 Vbias.n364 4.5005
R20759 Vbias.n494 Vbias.n308 4.5005
R20760 Vbias.n491 Vbias.n310 4.5005
R20761 Vbias.n558 Vbias.n557 4.5005
R20762 Vbias.n631 Vbias.n255 4.5005
R20763 Vbias.n628 Vbias.n257 4.5005
R20764 Vbias.n219 Vbias.n218 4.5005
R20765 Vbias.n738 Vbias.n173 4.5005
R20766 Vbias.n741 Vbias.n171 4.5005
R20767 Vbias.n812 Vbias.n811 4.5005
R20768 Vbias.n869 Vbias.n124 4.5005
R20769 Vbias.n866 Vbias.n126 4.5005
R20770 Vbias.n77 Vbias.n76 4.5005
R20771 Vbias.n958 Vbias.n33 4.5005
R20772 Vbias.n956 Vbias.n35 4.5005
R20773 Vbias.n418 Vbias.n417 4.5005
R20774 Vbias.n368 Vbias.n367 4.5005
R20775 Vbias.n497 Vbias.n307 4.5005
R20776 Vbias.n500 Vbias.n305 4.5005
R20777 Vbias.n555 Vbias.n554 4.5005
R20778 Vbias.n634 Vbias.n254 4.5005
R20779 Vbias.n637 Vbias.n252 4.5005
R20780 Vbias.n222 Vbias.n221 4.5005
R20781 Vbias.n735 Vbias.n174 4.5005
R20782 Vbias.n732 Vbias.n176 4.5005
R20783 Vbias.n815 Vbias.n814 4.5005
R20784 Vbias.n860 Vbias.n129 4.5005
R20785 Vbias.n863 Vbias.n127 4.5005
R20786 Vbias.n74 Vbias.n73 4.5005
R20787 Vbias.n961 Vbias.n32 4.5005
R20788 Vbias.n963 Vbias.n30 4.5005
R20789 Vbias.n415 Vbias.n414 4.5005
R20790 Vbias.n371 Vbias.n370 4.5005
R20791 Vbias.n506 Vbias.n302 4.5005
R20792 Vbias.n503 Vbias.n304 4.5005
R20793 Vbias.n552 Vbias.n551 4.5005
R20794 Vbias.n643 Vbias.n249 4.5005
R20795 Vbias.n640 Vbias.n251 4.5005
R20796 Vbias.n225 Vbias.n224 4.5005
R20797 Vbias.n726 Vbias.n179 4.5005
R20798 Vbias.n729 Vbias.n177 4.5005
R20799 Vbias.n818 Vbias.n817 4.5005
R20800 Vbias.n857 Vbias.n130 4.5005
R20801 Vbias.n854 Vbias.n132 4.5005
R20802 Vbias.n71 Vbias.n70 4.5005
R20803 Vbias.n968 Vbias.n27 4.5005
R20804 Vbias.n966 Vbias.n29 4.5005
R20805 Vbias.n412 Vbias.n411 4.5005
R20806 Vbias.n374 Vbias.n373 4.5005
R20807 Vbias.n509 Vbias.n301 4.5005
R20808 Vbias.n512 Vbias.n299 4.5005
R20809 Vbias.n549 Vbias.n548 4.5005
R20810 Vbias.n646 Vbias.n248 4.5005
R20811 Vbias.n649 Vbias.n246 4.5005
R20812 Vbias.n228 Vbias.n227 4.5005
R20813 Vbias.n723 Vbias.n180 4.5005
R20814 Vbias.n720 Vbias.n182 4.5005
R20815 Vbias.n821 Vbias.n820 4.5005
R20816 Vbias.n848 Vbias.n135 4.5005
R20817 Vbias.n851 Vbias.n133 4.5005
R20818 Vbias.n68 Vbias.n67 4.5005
R20819 Vbias.n971 Vbias.n26 4.5005
R20820 Vbias.n973 Vbias.n24 4.5005
R20821 Vbias.n409 Vbias.n408 4.5005
R20822 Vbias.n377 Vbias.n376 4.5005
R20823 Vbias.n518 Vbias.n296 4.5005
R20824 Vbias.n515 Vbias.n298 4.5005
R20825 Vbias.n546 Vbias.n545 4.5005
R20826 Vbias.n655 Vbias.n243 4.5005
R20827 Vbias.n652 Vbias.n245 4.5005
R20828 Vbias.n231 Vbias.n230 4.5005
R20829 Vbias.n714 Vbias.n185 4.5005
R20830 Vbias.n717 Vbias.n183 4.5005
R20831 Vbias.n824 Vbias.n823 4.5005
R20832 Vbias.n845 Vbias.n136 4.5005
R20833 Vbias.n842 Vbias.n138 4.5005
R20834 Vbias.n65 Vbias.n64 4.5005
R20835 Vbias.n978 Vbias.n21 4.5005
R20836 Vbias.n976 Vbias.n23 4.5005
R20837 Vbias.n406 Vbias.n405 4.5005
R20838 Vbias.n380 Vbias.n379 4.5005
R20839 Vbias.n521 Vbias.n295 4.5005
R20840 Vbias.n524 Vbias.n293 4.5005
R20841 Vbias.n543 Vbias.n542 4.5005
R20842 Vbias.n658 Vbias.n242 4.5005
R20843 Vbias.n661 Vbias.n240 4.5005
R20844 Vbias.n234 Vbias.n233 4.5005
R20845 Vbias.n711 Vbias.n186 4.5005
R20846 Vbias.n708 Vbias.n188 4.5005
R20847 Vbias.n827 Vbias.n826 4.5005
R20848 Vbias.n836 Vbias.n141 4.5005
R20849 Vbias.n839 Vbias.n139 4.5005
R20850 Vbias.n62 Vbias.n61 4.5005
R20851 Vbias.n981 Vbias.n18 4.5005
R20852 Vbias.n983 Vbias.n16 4.5005
R20853 Vbias.n403 Vbias.n338 4.5005
R20854 Vbias.n340 Vbias.n339 4.5005
R20855 Vbias.n400 Vbias.n341 4.5005
R20856 Vbias.n527 Vbias.n526 4.5005
R20857 Vbias.n540 Vbias.n285 4.5005
R20858 Vbias.n537 Vbias.n287 4.5005
R20859 Vbias.n664 Vbias.n663 4.5005
R20860 Vbias.n695 Vbias.n236 4.5005
R20861 Vbias.n692 Vbias.n238 4.5005
R20862 Vbias.n705 Vbias.n704 4.5005
R20863 Vbias.n830 Vbias.n144 4.5005
R20864 Vbias.n833 Vbias.n142 4.5005
R20865 Vbias.n673 Vbias.n672 4.5005
R20866 Vbias.n989 Vbias.n11 4.5005
R20867 Vbias.n14 Vbias.n13 4.5005
R20868 Vbias.n986 Vbias.n15 4.5005
R20869 Vbias.n995 Vbias.n6 4.5005
R20870 Vbias.n59 Vbias.n58 4.5005
R20871 Vbias.n919 Vbias.n57 4.5005
R20872 Vbias.n8 Vbias.n7 4.5005
R20873 Vbias.n992 Vbias.n10 4.5005
R20874 Vbias.n100 Vbias.n60 4.5005
R20875 Vbias.n915 Vbias.n102 4.5005
R20876 Vbias.n676 Vbias.n675 4.5005
R20877 Vbias.n681 Vbias.n679 4.5005
R20878 Vbias.n908 Vbias.n907 4.5005
R20879 Vbias.n789 Vbias.n145 4.5005
R20880 Vbias.n685 Vbias.n684 4.5005
R20881 Vbias.n702 Vbias.n189 4.5005
R20882 Vbias.n147 Vbias.n146 4.5005
R20883 Vbias.n785 Vbias.n149 4.5005
R20884 Vbias.n192 Vbias.n191 4.5005
R20885 Vbias.n698 Vbias.n194 4.5005
R20886 Vbias.n196 Vbias.n195 4.5005
R20887 Vbias.n281 Vbias.n280 4.5005
R20888 Vbias.n667 Vbias.n666 4.5005
R20889 Vbias.n534 Vbias.n288 4.5005
R20890 Vbias.n584 Vbias.n279 4.5005
R20891 Vbias.n581 Vbias.n284 4.5005
R20892 Vbias.n290 Vbias.n289 4.5005
R20893 Vbias.n530 Vbias.n292 4.5005
R20894 Vbias.n330 Vbias.n329 4.5005
R20895 Vbias.n447 Vbias.n334 4.5005
R20896 Vbias.n397 Vbias.n396 4.5005
R20897 Vbias.n389 Vbias.n383 4.5005
R20898 Vbias.n336 Vbias.n335 4.5005
R20899 Vbias.n444 Vbias.n337 4.5005
R20900 Vbias.n59 Vbias 3.50727
R20901 Vbias Vbias.n919 3.50727
R20902 Vbias.n100 Vbias 3.50727
R20903 Vbias.n915 Vbias 3.50727
R20904 Vbias Vbias.n908 3.50727
R20905 Vbias Vbias.n789 3.50727
R20906 Vbias Vbias.n147 3.50727
R20907 Vbias.n785 Vbias 3.50727
R20908 Vbias Vbias.n196 3.50727
R20909 Vbias.n281 Vbias 3.50727
R20910 Vbias Vbias.n584 3.50727
R20911 Vbias.n581 Vbias 3.50727
R20912 Vbias Vbias.n330 3.50727
R20913 Vbias Vbias.n447 3.50727
R20914 Vbias Vbias.n336 3.50727
R20915 Vbias.n444 Vbias 3.50727
R20916 Vbias.n996 Vbias.n995 3.4105
R20917 Vbias.n986 Vbias.n985 3.4105
R20918 Vbias.n984 Vbias.n983 3.4105
R20919 Vbias.n976 Vbias.n975 3.4105
R20920 Vbias.n974 Vbias.n973 3.4105
R20921 Vbias.n966 Vbias.n965 3.4105
R20922 Vbias.n964 Vbias.n963 3.4105
R20923 Vbias.n956 Vbias.n955 3.4105
R20924 Vbias.n954 Vbias.n953 3.4105
R20925 Vbias.n946 Vbias.n945 3.4105
R20926 Vbias.n944 Vbias.n943 3.4105
R20927 Vbias.n936 Vbias.n935 3.4105
R20928 Vbias.n934 Vbias.n933 3.4105
R20929 Vbias.n926 Vbias.n925 3.4105
R20930 Vbias.n924 Vbias.n923 3.4105
R20931 Vbias.n921 Vbias.n920 3.4105
R20932 Vbias.n929 Vbias.n928 3.4105
R20933 Vbias.n931 Vbias.n930 3.4105
R20934 Vbias.n939 Vbias.n938 3.4105
R20935 Vbias.n941 Vbias.n940 3.4105
R20936 Vbias.n949 Vbias.n948 3.4105
R20937 Vbias.n951 Vbias.n950 3.4105
R20938 Vbias.n959 Vbias.n958 3.4105
R20939 Vbias.n961 Vbias.n960 3.4105
R20940 Vbias.n969 Vbias.n968 3.4105
R20941 Vbias.n971 Vbias.n970 3.4105
R20942 Vbias.n979 Vbias.n978 3.4105
R20943 Vbias.n981 Vbias.n980 3.4105
R20944 Vbias.n20 Vbias.n14 3.4105
R20945 Vbias.n19 Vbias.n8 3.4105
R20946 Vbias.n992 Vbias.n991 3.4105
R20947 Vbias.n990 Vbias.n989 3.4105
R20948 Vbias.n63 Vbias.n62 3.4105
R20949 Vbias.n66 Vbias.n65 3.4105
R20950 Vbias.n69 Vbias.n68 3.4105
R20951 Vbias.n72 Vbias.n71 3.4105
R20952 Vbias.n75 Vbias.n74 3.4105
R20953 Vbias.n78 Vbias.n77 3.4105
R20954 Vbias.n81 Vbias.n80 3.4105
R20955 Vbias.n84 Vbias.n83 3.4105
R20956 Vbias.n87 Vbias.n86 3.4105
R20957 Vbias.n90 Vbias.n89 3.4105
R20958 Vbias.n93 Vbias.n92 3.4105
R20959 Vbias.n96 Vbias.n95 3.4105
R20960 Vbias.n99 Vbias.n98 3.4105
R20961 Vbias.n914 Vbias.n913 3.4105
R20962 Vbias.n902 Vbias.n901 3.4105
R20963 Vbias.n900 Vbias.n899 3.4105
R20964 Vbias.n890 Vbias.n889 3.4105
R20965 Vbias.n888 Vbias.n887 3.4105
R20966 Vbias.n878 Vbias.n877 3.4105
R20967 Vbias.n876 Vbias.n875 3.4105
R20968 Vbias.n866 Vbias.n865 3.4105
R20969 Vbias.n864 Vbias.n863 3.4105
R20970 Vbias.n854 Vbias.n853 3.4105
R20971 Vbias.n852 Vbias.n851 3.4105
R20972 Vbias.n842 Vbias.n841 3.4105
R20973 Vbias.n840 Vbias.n839 3.4105
R20974 Vbias.n674 Vbias.n673 3.4105
R20975 Vbias.n677 Vbias.n676 3.4105
R20976 Vbias.n682 Vbias.n681 3.4105
R20977 Vbias.n834 Vbias.n833 3.4105
R20978 Vbias.n836 Vbias.n835 3.4105
R20979 Vbias.n846 Vbias.n845 3.4105
R20980 Vbias.n848 Vbias.n847 3.4105
R20981 Vbias.n858 Vbias.n857 3.4105
R20982 Vbias.n860 Vbias.n859 3.4105
R20983 Vbias.n870 Vbias.n869 3.4105
R20984 Vbias.n872 Vbias.n871 3.4105
R20985 Vbias.n882 Vbias.n881 3.4105
R20986 Vbias.n884 Vbias.n883 3.4105
R20987 Vbias.n894 Vbias.n893 3.4105
R20988 Vbias.n896 Vbias.n895 3.4105
R20989 Vbias.n906 Vbias.n905 3.4105
R20990 Vbias.n910 Vbias.n909 3.4105
R20991 Vbias.n792 Vbias.n791 3.4105
R20992 Vbias.n795 Vbias.n794 3.4105
R20993 Vbias.n798 Vbias.n797 3.4105
R20994 Vbias.n801 Vbias.n800 3.4105
R20995 Vbias.n804 Vbias.n803 3.4105
R20996 Vbias.n807 Vbias.n806 3.4105
R20997 Vbias.n810 Vbias.n809 3.4105
R20998 Vbias.n813 Vbias.n812 3.4105
R20999 Vbias.n816 Vbias.n815 3.4105
R21000 Vbias.n819 Vbias.n818 3.4105
R21001 Vbias.n822 Vbias.n821 3.4105
R21002 Vbias.n825 Vbias.n824 3.4105
R21003 Vbias.n828 Vbias.n827 3.4105
R21004 Vbias.n830 Vbias.n829 3.4105
R21005 Vbias.n686 Vbias.n685 3.4105
R21006 Vbias.n703 Vbias.n702 3.4105
R21007 Vbias.n706 Vbias.n705 3.4105
R21008 Vbias.n708 Vbias.n707 3.4105
R21009 Vbias.n718 Vbias.n717 3.4105
R21010 Vbias.n720 Vbias.n719 3.4105
R21011 Vbias.n730 Vbias.n729 3.4105
R21012 Vbias.n732 Vbias.n731 3.4105
R21013 Vbias.n742 Vbias.n741 3.4105
R21014 Vbias.n744 Vbias.n743 3.4105
R21015 Vbias.n754 Vbias.n753 3.4105
R21016 Vbias.n756 Vbias.n755 3.4105
R21017 Vbias.n766 Vbias.n765 3.4105
R21018 Vbias.n768 Vbias.n767 3.4105
R21019 Vbias.n778 Vbias.n777 3.4105
R21020 Vbias.n780 Vbias.n779 3.4105
R21021 Vbias.n784 Vbias.n783 3.4105
R21022 Vbias.n774 Vbias.n773 3.4105
R21023 Vbias.n772 Vbias.n771 3.4105
R21024 Vbias.n762 Vbias.n761 3.4105
R21025 Vbias.n760 Vbias.n759 3.4105
R21026 Vbias.n750 Vbias.n749 3.4105
R21027 Vbias.n748 Vbias.n747 3.4105
R21028 Vbias.n738 Vbias.n737 3.4105
R21029 Vbias.n736 Vbias.n735 3.4105
R21030 Vbias.n726 Vbias.n725 3.4105
R21031 Vbias.n724 Vbias.n723 3.4105
R21032 Vbias.n714 Vbias.n713 3.4105
R21033 Vbias.n712 Vbias.n711 3.4105
R21034 Vbias.n692 Vbias.n691 3.4105
R21035 Vbias.n690 Vbias.n192 3.4105
R21036 Vbias.n698 Vbias.n697 3.4105
R21037 Vbias.n696 Vbias.n695 3.4105
R21038 Vbias.n235 Vbias.n234 3.4105
R21039 Vbias.n232 Vbias.n231 3.4105
R21040 Vbias.n229 Vbias.n228 3.4105
R21041 Vbias.n226 Vbias.n225 3.4105
R21042 Vbias.n223 Vbias.n222 3.4105
R21043 Vbias.n220 Vbias.n219 3.4105
R21044 Vbias.n217 Vbias.n216 3.4105
R21045 Vbias.n214 Vbias.n213 3.4105
R21046 Vbias.n211 Vbias.n210 3.4105
R21047 Vbias.n208 Vbias.n207 3.4105
R21048 Vbias.n205 Vbias.n204 3.4105
R21049 Vbias.n202 Vbias.n201 3.4105
R21050 Vbias.n199 Vbias.n198 3.4105
R21051 Vbias.n590 Vbias.n589 3.4105
R21052 Vbias.n592 Vbias.n591 3.4105
R21053 Vbias.n602 Vbias.n601 3.4105
R21054 Vbias.n604 Vbias.n603 3.4105
R21055 Vbias.n614 Vbias.n613 3.4105
R21056 Vbias.n616 Vbias.n615 3.4105
R21057 Vbias.n626 Vbias.n625 3.4105
R21058 Vbias.n628 Vbias.n627 3.4105
R21059 Vbias.n638 Vbias.n637 3.4105
R21060 Vbias.n640 Vbias.n639 3.4105
R21061 Vbias.n650 Vbias.n649 3.4105
R21062 Vbias.n652 Vbias.n651 3.4105
R21063 Vbias.n662 Vbias.n661 3.4105
R21064 Vbias.n665 Vbias.n664 3.4105
R21065 Vbias.n668 Vbias.n667 3.4105
R21066 Vbias.n535 Vbias.n534 3.4105
R21067 Vbias.n537 Vbias.n536 3.4105
R21068 Vbias.n658 Vbias.n657 3.4105
R21069 Vbias.n656 Vbias.n655 3.4105
R21070 Vbias.n646 Vbias.n645 3.4105
R21071 Vbias.n644 Vbias.n643 3.4105
R21072 Vbias.n634 Vbias.n633 3.4105
R21073 Vbias.n632 Vbias.n631 3.4105
R21074 Vbias.n622 Vbias.n621 3.4105
R21075 Vbias.n620 Vbias.n619 3.4105
R21076 Vbias.n610 Vbias.n609 3.4105
R21077 Vbias.n608 Vbias.n607 3.4105
R21078 Vbias.n598 Vbias.n597 3.4105
R21079 Vbias.n596 Vbias.n595 3.4105
R21080 Vbias.n586 Vbias.n585 3.4105
R21081 Vbias.n580 Vbias.n579 3.4105
R21082 Vbias.n577 Vbias.n576 3.4105
R21083 Vbias.n574 Vbias.n573 3.4105
R21084 Vbias.n571 Vbias.n570 3.4105
R21085 Vbias.n568 Vbias.n567 3.4105
R21086 Vbias.n565 Vbias.n564 3.4105
R21087 Vbias.n562 Vbias.n561 3.4105
R21088 Vbias.n559 Vbias.n558 3.4105
R21089 Vbias.n556 Vbias.n555 3.4105
R21090 Vbias.n553 Vbias.n552 3.4105
R21091 Vbias.n550 Vbias.n549 3.4105
R21092 Vbias.n547 Vbias.n546 3.4105
R21093 Vbias.n544 Vbias.n543 3.4105
R21094 Vbias.n541 Vbias.n540 3.4105
R21095 Vbias.n392 Vbias.n290 3.4105
R21096 Vbias.n530 Vbias.n529 3.4105
R21097 Vbias.n528 Vbias.n527 3.4105
R21098 Vbias.n525 Vbias.n524 3.4105
R21099 Vbias.n515 Vbias.n514 3.4105
R21100 Vbias.n513 Vbias.n512 3.4105
R21101 Vbias.n503 Vbias.n502 3.4105
R21102 Vbias.n501 Vbias.n500 3.4105
R21103 Vbias.n491 Vbias.n490 3.4105
R21104 Vbias.n489 Vbias.n488 3.4105
R21105 Vbias.n479 Vbias.n478 3.4105
R21106 Vbias.n477 Vbias.n476 3.4105
R21107 Vbias.n467 Vbias.n466 3.4105
R21108 Vbias.n465 Vbias.n464 3.4105
R21109 Vbias.n455 Vbias.n454 3.4105
R21110 Vbias.n453 Vbias.n452 3.4105
R21111 Vbias.n449 Vbias.n448 3.4105
R21112 Vbias.n459 Vbias.n458 3.4105
R21113 Vbias.n461 Vbias.n460 3.4105
R21114 Vbias.n471 Vbias.n470 3.4105
R21115 Vbias.n473 Vbias.n472 3.4105
R21116 Vbias.n483 Vbias.n482 3.4105
R21117 Vbias.n485 Vbias.n484 3.4105
R21118 Vbias.n495 Vbias.n494 3.4105
R21119 Vbias.n497 Vbias.n496 3.4105
R21120 Vbias.n507 Vbias.n506 3.4105
R21121 Vbias.n509 Vbias.n508 3.4105
R21122 Vbias.n519 Vbias.n518 3.4105
R21123 Vbias.n521 Vbias.n520 3.4105
R21124 Vbias.n400 Vbias.n399 3.4105
R21125 Vbias.n398 Vbias.n397 3.4105
R21126 Vbias.n390 Vbias.n389 3.4105
R21127 Vbias.n382 Vbias.n340 3.4105
R21128 Vbias.n381 Vbias.n380 3.4105
R21129 Vbias.n378 Vbias.n377 3.4105
R21130 Vbias.n375 Vbias.n374 3.4105
R21131 Vbias.n372 Vbias.n371 3.4105
R21132 Vbias.n369 Vbias.n368 3.4105
R21133 Vbias.n366 Vbias.n365 3.4105
R21134 Vbias.n363 Vbias.n362 3.4105
R21135 Vbias.n360 Vbias.n359 3.4105
R21136 Vbias.n357 Vbias.n356 3.4105
R21137 Vbias.n354 Vbias.n353 3.4105
R21138 Vbias.n351 Vbias.n350 3.4105
R21139 Vbias.n348 Vbias.n347 3.4105
R21140 Vbias.n345 Vbias.n344 3.4105
R21141 Vbias.n443 Vbias.n442 3.4105
R21142 Vbias.n440 Vbias.n439 3.4105
R21143 Vbias.n437 Vbias.n436 3.4105
R21144 Vbias.n434 Vbias.n433 3.4105
R21145 Vbias.n431 Vbias.n430 3.4105
R21146 Vbias.n428 Vbias.n427 3.4105
R21147 Vbias.n425 Vbias.n424 3.4105
R21148 Vbias.n422 Vbias.n421 3.4105
R21149 Vbias.n419 Vbias.n418 3.4105
R21150 Vbias.n416 Vbias.n415 3.4105
R21151 Vbias.n413 Vbias.n412 3.4105
R21152 Vbias.n410 Vbias.n409 3.4105
R21153 Vbias.n407 Vbias.n406 3.4105
R21154 Vbias.n404 Vbias.n403 3.4105
R21155 Vbias.n387 Vbias.n386 3.4105
R21156 Vbias.n388 Vbias.n387 2.9408
R21157 Vbias.n442 Vbias.n332 2.9408
R21158 Vbias.n923 Vbias.n922 2.9408
R21159 Vbias.n439 Vbias.n327 2.9408
R21160 Vbias.n927 Vbias.n926 2.9408
R21161 Vbias.n436 Vbias.n324 2.9408
R21162 Vbias.n933 Vbias.n932 2.9408
R21163 Vbias.n433 Vbias.n321 2.9408
R21164 Vbias.n937 Vbias.n936 2.9408
R21165 Vbias.n430 Vbias.n318 2.9408
R21166 Vbias.n943 Vbias.n942 2.9408
R21167 Vbias.n427 Vbias.n315 2.9408
R21168 Vbias.n947 Vbias.n946 2.9408
R21169 Vbias.n424 Vbias.n312 2.9408
R21170 Vbias.n953 Vbias.n952 2.9408
R21171 Vbias.n421 Vbias.n309 2.9408
R21172 Vbias.n957 Vbias.n956 2.9408
R21173 Vbias.n418 Vbias.n306 2.9408
R21174 Vbias.n963 Vbias.n962 2.9408
R21175 Vbias.n415 Vbias.n303 2.9408
R21176 Vbias.n967 Vbias.n966 2.9408
R21177 Vbias.n412 Vbias.n300 2.9408
R21178 Vbias.n973 Vbias.n972 2.9408
R21179 Vbias.n409 Vbias.n297 2.9408
R21180 Vbias.n977 Vbias.n976 2.9408
R21181 Vbias.n406 Vbias.n294 2.9408
R21182 Vbias.n983 Vbias.n982 2.9408
R21183 Vbias.n403 Vbias.n402 2.9408
R21184 Vbias.n987 Vbias.n986 2.9408
R21185 Vbias.n995 Vbias.n994 2.9408
R21186 Vbias.n918 Vbias.n59 2.9408
R21187 Vbias.n445 Vbias.n444 2.9408
R21188 Vbias.n450 Vbias.n332 2.76612
R21189 Vbias.n451 Vbias.n450 2.76612
R21190 Vbias.n451 Vbias.n277 2.76612
R21191 Vbias.n587 Vbias.n277 2.76612
R21192 Vbias.n588 Vbias.n587 2.76612
R21193 Vbias.n588 Vbias.n151 2.76612
R21194 Vbias.n782 Vbias.n151 2.76612
R21195 Vbias.n782 Vbias.n781 2.76612
R21196 Vbias.n781 Vbias.n104 2.76612
R21197 Vbias.n911 Vbias.n104 2.76612
R21198 Vbias.n912 Vbias.n911 2.76612
R21199 Vbias.n912 Vbias.n55 2.76612
R21200 Vbias.n922 Vbias.n55 2.76612
R21201 Vbias.n457 Vbias.n327 2.76612
R21202 Vbias.n457 Vbias.n456 2.76612
R21203 Vbias.n456 Vbias.n274 2.76612
R21204 Vbias.n594 Vbias.n274 2.76612
R21205 Vbias.n594 Vbias.n593 2.76612
R21206 Vbias.n593 Vbias.n154 2.76612
R21207 Vbias.n775 Vbias.n154 2.76612
R21208 Vbias.n776 Vbias.n775 2.76612
R21209 Vbias.n776 Vbias.n107 2.76612
R21210 Vbias.n904 Vbias.n107 2.76612
R21211 Vbias.n904 Vbias.n903 2.76612
R21212 Vbias.n903 Vbias.n52 2.76612
R21213 Vbias.n927 Vbias.n52 2.76612
R21214 Vbias.n462 Vbias.n324 2.76612
R21215 Vbias.n463 Vbias.n462 2.76612
R21216 Vbias.n463 Vbias.n271 2.76612
R21217 Vbias.n599 Vbias.n271 2.76612
R21218 Vbias.n600 Vbias.n599 2.76612
R21219 Vbias.n600 Vbias.n157 2.76612
R21220 Vbias.n770 Vbias.n157 2.76612
R21221 Vbias.n770 Vbias.n769 2.76612
R21222 Vbias.n769 Vbias.n110 2.76612
R21223 Vbias.n897 Vbias.n110 2.76612
R21224 Vbias.n898 Vbias.n897 2.76612
R21225 Vbias.n898 Vbias.n49 2.76612
R21226 Vbias.n932 Vbias.n49 2.76612
R21227 Vbias.n469 Vbias.n321 2.76612
R21228 Vbias.n469 Vbias.n468 2.76612
R21229 Vbias.n468 Vbias.n268 2.76612
R21230 Vbias.n606 Vbias.n268 2.76612
R21231 Vbias.n606 Vbias.n605 2.76612
R21232 Vbias.n605 Vbias.n160 2.76612
R21233 Vbias.n763 Vbias.n160 2.76612
R21234 Vbias.n764 Vbias.n763 2.76612
R21235 Vbias.n764 Vbias.n113 2.76612
R21236 Vbias.n892 Vbias.n113 2.76612
R21237 Vbias.n892 Vbias.n891 2.76612
R21238 Vbias.n891 Vbias.n46 2.76612
R21239 Vbias.n937 Vbias.n46 2.76612
R21240 Vbias.n474 Vbias.n318 2.76612
R21241 Vbias.n475 Vbias.n474 2.76612
R21242 Vbias.n475 Vbias.n265 2.76612
R21243 Vbias.n611 Vbias.n265 2.76612
R21244 Vbias.n612 Vbias.n611 2.76612
R21245 Vbias.n612 Vbias.n163 2.76612
R21246 Vbias.n758 Vbias.n163 2.76612
R21247 Vbias.n758 Vbias.n757 2.76612
R21248 Vbias.n757 Vbias.n116 2.76612
R21249 Vbias.n885 Vbias.n116 2.76612
R21250 Vbias.n886 Vbias.n885 2.76612
R21251 Vbias.n886 Vbias.n43 2.76612
R21252 Vbias.n942 Vbias.n43 2.76612
R21253 Vbias.n481 Vbias.n315 2.76612
R21254 Vbias.n481 Vbias.n480 2.76612
R21255 Vbias.n480 Vbias.n262 2.76612
R21256 Vbias.n618 Vbias.n262 2.76612
R21257 Vbias.n618 Vbias.n617 2.76612
R21258 Vbias.n617 Vbias.n166 2.76612
R21259 Vbias.n751 Vbias.n166 2.76612
R21260 Vbias.n752 Vbias.n751 2.76612
R21261 Vbias.n752 Vbias.n119 2.76612
R21262 Vbias.n880 Vbias.n119 2.76612
R21263 Vbias.n880 Vbias.n879 2.76612
R21264 Vbias.n879 Vbias.n40 2.76612
R21265 Vbias.n947 Vbias.n40 2.76612
R21266 Vbias.n486 Vbias.n312 2.76612
R21267 Vbias.n487 Vbias.n486 2.76612
R21268 Vbias.n487 Vbias.n259 2.76612
R21269 Vbias.n623 Vbias.n259 2.76612
R21270 Vbias.n624 Vbias.n623 2.76612
R21271 Vbias.n624 Vbias.n169 2.76612
R21272 Vbias.n746 Vbias.n169 2.76612
R21273 Vbias.n746 Vbias.n745 2.76612
R21274 Vbias.n745 Vbias.n122 2.76612
R21275 Vbias.n873 Vbias.n122 2.76612
R21276 Vbias.n874 Vbias.n873 2.76612
R21277 Vbias.n874 Vbias.n37 2.76612
R21278 Vbias.n952 Vbias.n37 2.76612
R21279 Vbias.n493 Vbias.n309 2.76612
R21280 Vbias.n493 Vbias.n492 2.76612
R21281 Vbias.n492 Vbias.n256 2.76612
R21282 Vbias.n630 Vbias.n256 2.76612
R21283 Vbias.n630 Vbias.n629 2.76612
R21284 Vbias.n629 Vbias.n172 2.76612
R21285 Vbias.n739 Vbias.n172 2.76612
R21286 Vbias.n740 Vbias.n739 2.76612
R21287 Vbias.n740 Vbias.n125 2.76612
R21288 Vbias.n868 Vbias.n125 2.76612
R21289 Vbias.n868 Vbias.n867 2.76612
R21290 Vbias.n867 Vbias.n34 2.76612
R21291 Vbias.n957 Vbias.n34 2.76612
R21292 Vbias.n498 Vbias.n306 2.76612
R21293 Vbias.n499 Vbias.n498 2.76612
R21294 Vbias.n499 Vbias.n253 2.76612
R21295 Vbias.n635 Vbias.n253 2.76612
R21296 Vbias.n636 Vbias.n635 2.76612
R21297 Vbias.n636 Vbias.n175 2.76612
R21298 Vbias.n734 Vbias.n175 2.76612
R21299 Vbias.n734 Vbias.n733 2.76612
R21300 Vbias.n733 Vbias.n128 2.76612
R21301 Vbias.n861 Vbias.n128 2.76612
R21302 Vbias.n862 Vbias.n861 2.76612
R21303 Vbias.n862 Vbias.n31 2.76612
R21304 Vbias.n962 Vbias.n31 2.76612
R21305 Vbias.n505 Vbias.n303 2.76612
R21306 Vbias.n505 Vbias.n504 2.76612
R21307 Vbias.n504 Vbias.n250 2.76612
R21308 Vbias.n642 Vbias.n250 2.76612
R21309 Vbias.n642 Vbias.n641 2.76612
R21310 Vbias.n641 Vbias.n178 2.76612
R21311 Vbias.n727 Vbias.n178 2.76612
R21312 Vbias.n728 Vbias.n727 2.76612
R21313 Vbias.n728 Vbias.n131 2.76612
R21314 Vbias.n856 Vbias.n131 2.76612
R21315 Vbias.n856 Vbias.n855 2.76612
R21316 Vbias.n855 Vbias.n28 2.76612
R21317 Vbias.n967 Vbias.n28 2.76612
R21318 Vbias.n510 Vbias.n300 2.76612
R21319 Vbias.n511 Vbias.n510 2.76612
R21320 Vbias.n511 Vbias.n247 2.76612
R21321 Vbias.n647 Vbias.n247 2.76612
R21322 Vbias.n648 Vbias.n647 2.76612
R21323 Vbias.n648 Vbias.n181 2.76612
R21324 Vbias.n722 Vbias.n181 2.76612
R21325 Vbias.n722 Vbias.n721 2.76612
R21326 Vbias.n721 Vbias.n134 2.76612
R21327 Vbias.n849 Vbias.n134 2.76612
R21328 Vbias.n850 Vbias.n849 2.76612
R21329 Vbias.n850 Vbias.n25 2.76612
R21330 Vbias.n972 Vbias.n25 2.76612
R21331 Vbias.n517 Vbias.n297 2.76612
R21332 Vbias.n517 Vbias.n516 2.76612
R21333 Vbias.n516 Vbias.n244 2.76612
R21334 Vbias.n654 Vbias.n244 2.76612
R21335 Vbias.n654 Vbias.n653 2.76612
R21336 Vbias.n653 Vbias.n184 2.76612
R21337 Vbias.n715 Vbias.n184 2.76612
R21338 Vbias.n716 Vbias.n715 2.76612
R21339 Vbias.n716 Vbias.n137 2.76612
R21340 Vbias.n844 Vbias.n137 2.76612
R21341 Vbias.n844 Vbias.n843 2.76612
R21342 Vbias.n843 Vbias.n22 2.76612
R21343 Vbias.n977 Vbias.n22 2.76612
R21344 Vbias.n522 Vbias.n294 2.76612
R21345 Vbias.n523 Vbias.n522 2.76612
R21346 Vbias.n523 Vbias.n241 2.76612
R21347 Vbias.n659 Vbias.n241 2.76612
R21348 Vbias.n660 Vbias.n659 2.76612
R21349 Vbias.n660 Vbias.n187 2.76612
R21350 Vbias.n710 Vbias.n187 2.76612
R21351 Vbias.n710 Vbias.n709 2.76612
R21352 Vbias.n709 Vbias.n140 2.76612
R21353 Vbias.n837 Vbias.n140 2.76612
R21354 Vbias.n838 Vbias.n837 2.76612
R21355 Vbias.n838 Vbias.n17 2.76612
R21356 Vbias.n982 Vbias.n17 2.76612
R21357 Vbias.n402 Vbias.n401 2.76612
R21358 Vbias.n401 Vbias.n286 2.76612
R21359 Vbias.n539 Vbias.n286 2.76612
R21360 Vbias.n539 Vbias.n538 2.76612
R21361 Vbias.n538 Vbias.n237 2.76612
R21362 Vbias.n694 Vbias.n237 2.76612
R21363 Vbias.n694 Vbias.n693 2.76612
R21364 Vbias.n693 Vbias.n143 2.76612
R21365 Vbias.n831 Vbias.n143 2.76612
R21366 Vbias.n832 Vbias.n831 2.76612
R21367 Vbias.n832 Vbias.n12 2.76612
R21368 Vbias.n988 Vbias.n12 2.76612
R21369 Vbias.n988 Vbias.n987 2.76612
R21370 Vbias.n918 Vbias.n917 2.76612
R21371 Vbias.n994 Vbias.n993 2.76612
R21372 Vbias.n993 Vbias.n9 2.76612
R21373 Vbias.n917 Vbias.n916 2.76612
R21374 Vbias.n916 Vbias.n101 2.76612
R21375 Vbias.n680 Vbias.n9 2.76612
R21376 Vbias.n680 Vbias.n190 2.76612
R21377 Vbias.n788 Vbias.n101 2.76612
R21378 Vbias.n788 Vbias.n787 2.76612
R21379 Vbias.n701 Vbias.n190 2.76612
R21380 Vbias.n701 Vbias.n700 2.76612
R21381 Vbias.n787 Vbias.n786 2.76612
R21382 Vbias.n786 Vbias.n148 2.76612
R21383 Vbias.n700 Vbias.n699 2.76612
R21384 Vbias.n699 Vbias.n193 2.76612
R21385 Vbias.n282 Vbias.n148 2.76612
R21386 Vbias.n583 Vbias.n282 2.76612
R21387 Vbias.n533 Vbias.n193 2.76612
R21388 Vbias.n533 Vbias.n532 2.76612
R21389 Vbias.n583 Vbias.n582 2.76612
R21390 Vbias.n582 Vbias.n283 2.76612
R21391 Vbias.n532 Vbias.n531 2.76612
R21392 Vbias.n531 Vbias.n291 2.76612
R21393 Vbias.n446 Vbias.n283 2.76612
R21394 Vbias.n446 Vbias.n445 2.76612
R21395 Vbias.n388 Vbias.n291 2.76612
R21396 Vbias.n4 Vbias.n3 2.06591
R21397 Vbias Vbias.n385 1.6647
R21398 Vbias Vbias.n395 1.6647
R21399 Vbias.n393 Vbias 1.6647
R21400 Vbias.n669 Vbias 1.6647
R21401 Vbias Vbias.n689 1.6647
R21402 Vbias.n687 Vbias 1.6647
R21403 Vbias.n678 Vbias 1.6647
R21404 Vbias Vbias.n5 1.6647
R21405 Vbias.n997 Vbias 1.6647
R21406 Vbias.n671 Vbias 1.6647
R21407 Vbias.n683 Vbias 1.6647
R21408 Vbias.n688 Vbias 1.6647
R21409 Vbias.n670 Vbias 1.6647
R21410 Vbias Vbias.n239 1.6647
R21411 Vbias.n394 Vbias 1.6647
R21412 Vbias.n391 Vbias 1.6647
R21413 Vbias Vbias.n998 1.57836
R21414 Vbias.n4 Vbias.n0 1.13456
R21415 Vbias Vbias.n4 0.782551
R21416 Vbias.n998 Vbias 0.412011
R21417 Vbias.n395 Vbias.n391 0.410967
R21418 Vbias.n395 Vbias.n394 0.410967
R21419 Vbias.n394 Vbias.n393 0.410967
R21420 Vbias.n393 Vbias.n239 0.410967
R21421 Vbias.n669 Vbias.n239 0.410967
R21422 Vbias.n670 Vbias.n669 0.410967
R21423 Vbias.n689 Vbias.n670 0.410967
R21424 Vbias.n689 Vbias.n688 0.410967
R21425 Vbias.n688 Vbias.n687 0.410967
R21426 Vbias.n687 Vbias.n683 0.410967
R21427 Vbias.n683 Vbias.n678 0.410967
R21428 Vbias.n678 Vbias.n671 0.410967
R21429 Vbias.n671 Vbias.n5 0.410967
R21430 Vbias.n997 Vbias.n5 0.410967
R21431 Vbias.n385 Vbias 0.383811
R21432 Vbias.n998 Vbias.n997 0.332633
R21433 Vbias.n342 Vbias.t260 0.322387
R21434 Vbias.n996 Vbias 0.252372
R21435 Vbias.n985 Vbias 0.252372
R21436 Vbias.n984 Vbias 0.252372
R21437 Vbias.n975 Vbias 0.252372
R21438 Vbias.n974 Vbias 0.252372
R21439 Vbias.n965 Vbias 0.252372
R21440 Vbias.n964 Vbias 0.252372
R21441 Vbias.n955 Vbias 0.252372
R21442 Vbias.n954 Vbias 0.252372
R21443 Vbias.n945 Vbias 0.252372
R21444 Vbias.n944 Vbias 0.252372
R21445 Vbias.n935 Vbias 0.252372
R21446 Vbias.n934 Vbias 0.252372
R21447 Vbias.n925 Vbias 0.252372
R21448 Vbias.n924 Vbias 0.252372
R21449 Vbias.n920 Vbias 0.252372
R21450 Vbias.n929 Vbias 0.252372
R21451 Vbias.n930 Vbias 0.252372
R21452 Vbias.n939 Vbias 0.252372
R21453 Vbias.n940 Vbias 0.252372
R21454 Vbias.n949 Vbias 0.252372
R21455 Vbias.n950 Vbias 0.252372
R21456 Vbias.n959 Vbias 0.252372
R21457 Vbias.n960 Vbias 0.252372
R21458 Vbias.n969 Vbias 0.252372
R21459 Vbias.n970 Vbias 0.252372
R21460 Vbias.n979 Vbias 0.252372
R21461 Vbias.n980 Vbias 0.252372
R21462 Vbias Vbias.n20 0.252372
R21463 Vbias Vbias.n19 0.252372
R21464 Vbias.n991 Vbias 0.252372
R21465 Vbias.n990 Vbias 0.252372
R21466 Vbias Vbias.n63 0.252372
R21467 Vbias Vbias.n66 0.252372
R21468 Vbias Vbias.n69 0.252372
R21469 Vbias Vbias.n72 0.252372
R21470 Vbias Vbias.n75 0.252372
R21471 Vbias Vbias.n78 0.252372
R21472 Vbias Vbias.n81 0.252372
R21473 Vbias Vbias.n84 0.252372
R21474 Vbias Vbias.n87 0.252372
R21475 Vbias Vbias.n90 0.252372
R21476 Vbias Vbias.n93 0.252372
R21477 Vbias Vbias.n96 0.252372
R21478 Vbias Vbias.n99 0.252372
R21479 Vbias Vbias.n914 0.252372
R21480 Vbias.n901 Vbias 0.252372
R21481 Vbias Vbias.n900 0.252372
R21482 Vbias.n889 Vbias 0.252372
R21483 Vbias Vbias.n888 0.252372
R21484 Vbias.n877 Vbias 0.252372
R21485 Vbias Vbias.n876 0.252372
R21486 Vbias.n865 Vbias 0.252372
R21487 Vbias Vbias.n864 0.252372
R21488 Vbias.n853 Vbias 0.252372
R21489 Vbias Vbias.n852 0.252372
R21490 Vbias.n841 Vbias 0.252372
R21491 Vbias Vbias.n840 0.252372
R21492 Vbias.n674 Vbias 0.252372
R21493 Vbias.n677 Vbias 0.252372
R21494 Vbias.n682 Vbias 0.252372
R21495 Vbias Vbias.n834 0.252372
R21496 Vbias.n835 Vbias 0.252372
R21497 Vbias Vbias.n846 0.252372
R21498 Vbias.n847 Vbias 0.252372
R21499 Vbias Vbias.n858 0.252372
R21500 Vbias.n859 Vbias 0.252372
R21501 Vbias Vbias.n870 0.252372
R21502 Vbias.n871 Vbias 0.252372
R21503 Vbias Vbias.n882 0.252372
R21504 Vbias.n883 Vbias 0.252372
R21505 Vbias Vbias.n894 0.252372
R21506 Vbias.n895 Vbias 0.252372
R21507 Vbias Vbias.n906 0.252372
R21508 Vbias.n909 Vbias 0.252372
R21509 Vbias.n792 Vbias 0.252372
R21510 Vbias.n795 Vbias 0.252372
R21511 Vbias.n798 Vbias 0.252372
R21512 Vbias.n801 Vbias 0.252372
R21513 Vbias.n804 Vbias 0.252372
R21514 Vbias.n807 Vbias 0.252372
R21515 Vbias.n810 Vbias 0.252372
R21516 Vbias.n813 Vbias 0.252372
R21517 Vbias.n816 Vbias 0.252372
R21518 Vbias.n819 Vbias 0.252372
R21519 Vbias.n822 Vbias 0.252372
R21520 Vbias.n825 Vbias 0.252372
R21521 Vbias.n828 Vbias 0.252372
R21522 Vbias.n829 Vbias 0.252372
R21523 Vbias.n686 Vbias 0.252372
R21524 Vbias Vbias.n703 0.252372
R21525 Vbias Vbias.n706 0.252372
R21526 Vbias.n707 Vbias 0.252372
R21527 Vbias Vbias.n718 0.252372
R21528 Vbias.n719 Vbias 0.252372
R21529 Vbias Vbias.n730 0.252372
R21530 Vbias.n731 Vbias 0.252372
R21531 Vbias Vbias.n742 0.252372
R21532 Vbias.n743 Vbias 0.252372
R21533 Vbias Vbias.n754 0.252372
R21534 Vbias.n755 Vbias 0.252372
R21535 Vbias Vbias.n766 0.252372
R21536 Vbias.n767 Vbias 0.252372
R21537 Vbias Vbias.n778 0.252372
R21538 Vbias.n779 Vbias 0.252372
R21539 Vbias Vbias.n784 0.252372
R21540 Vbias.n773 Vbias 0.252372
R21541 Vbias Vbias.n772 0.252372
R21542 Vbias.n761 Vbias 0.252372
R21543 Vbias Vbias.n760 0.252372
R21544 Vbias.n749 Vbias 0.252372
R21545 Vbias Vbias.n748 0.252372
R21546 Vbias.n737 Vbias 0.252372
R21547 Vbias Vbias.n736 0.252372
R21548 Vbias.n725 Vbias 0.252372
R21549 Vbias Vbias.n724 0.252372
R21550 Vbias.n713 Vbias 0.252372
R21551 Vbias Vbias.n712 0.252372
R21552 Vbias.n691 Vbias 0.252372
R21553 Vbias Vbias.n690 0.252372
R21554 Vbias.n697 Vbias 0.252372
R21555 Vbias.n696 Vbias 0.252372
R21556 Vbias.n235 Vbias 0.252372
R21557 Vbias.n232 Vbias 0.252372
R21558 Vbias.n229 Vbias 0.252372
R21559 Vbias.n226 Vbias 0.252372
R21560 Vbias.n223 Vbias 0.252372
R21561 Vbias.n220 Vbias 0.252372
R21562 Vbias.n217 Vbias 0.252372
R21563 Vbias.n214 Vbias 0.252372
R21564 Vbias.n211 Vbias 0.252372
R21565 Vbias.n208 Vbias 0.252372
R21566 Vbias.n205 Vbias 0.252372
R21567 Vbias.n202 Vbias 0.252372
R21568 Vbias.n199 Vbias 0.252372
R21569 Vbias.n590 Vbias 0.252372
R21570 Vbias.n591 Vbias 0.252372
R21571 Vbias.n602 Vbias 0.252372
R21572 Vbias.n603 Vbias 0.252372
R21573 Vbias.n614 Vbias 0.252372
R21574 Vbias.n615 Vbias 0.252372
R21575 Vbias.n626 Vbias 0.252372
R21576 Vbias.n627 Vbias 0.252372
R21577 Vbias.n638 Vbias 0.252372
R21578 Vbias.n639 Vbias 0.252372
R21579 Vbias.n650 Vbias 0.252372
R21580 Vbias.n651 Vbias 0.252372
R21581 Vbias.n662 Vbias 0.252372
R21582 Vbias.n665 Vbias 0.252372
R21583 Vbias.n668 Vbias 0.252372
R21584 Vbias Vbias.n535 0.252372
R21585 Vbias.n536 Vbias 0.252372
R21586 Vbias.n657 Vbias 0.252372
R21587 Vbias.n656 Vbias 0.252372
R21588 Vbias.n645 Vbias 0.252372
R21589 Vbias.n644 Vbias 0.252372
R21590 Vbias.n633 Vbias 0.252372
R21591 Vbias.n632 Vbias 0.252372
R21592 Vbias.n621 Vbias 0.252372
R21593 Vbias.n620 Vbias 0.252372
R21594 Vbias.n609 Vbias 0.252372
R21595 Vbias.n608 Vbias 0.252372
R21596 Vbias.n597 Vbias 0.252372
R21597 Vbias.n596 Vbias 0.252372
R21598 Vbias.n585 Vbias 0.252372
R21599 Vbias Vbias.n580 0.252372
R21600 Vbias Vbias.n577 0.252372
R21601 Vbias Vbias.n574 0.252372
R21602 Vbias Vbias.n571 0.252372
R21603 Vbias Vbias.n568 0.252372
R21604 Vbias Vbias.n565 0.252372
R21605 Vbias Vbias.n562 0.252372
R21606 Vbias Vbias.n559 0.252372
R21607 Vbias Vbias.n556 0.252372
R21608 Vbias Vbias.n553 0.252372
R21609 Vbias Vbias.n550 0.252372
R21610 Vbias Vbias.n547 0.252372
R21611 Vbias Vbias.n544 0.252372
R21612 Vbias Vbias.n541 0.252372
R21613 Vbias.n392 Vbias 0.252372
R21614 Vbias.n529 Vbias 0.252372
R21615 Vbias.n528 Vbias 0.252372
R21616 Vbias.n525 Vbias 0.252372
R21617 Vbias.n514 Vbias 0.252372
R21618 Vbias.n513 Vbias 0.252372
R21619 Vbias.n502 Vbias 0.252372
R21620 Vbias.n501 Vbias 0.252372
R21621 Vbias.n490 Vbias 0.252372
R21622 Vbias.n489 Vbias 0.252372
R21623 Vbias.n478 Vbias 0.252372
R21624 Vbias.n477 Vbias 0.252372
R21625 Vbias.n466 Vbias 0.252372
R21626 Vbias.n465 Vbias 0.252372
R21627 Vbias.n454 Vbias 0.252372
R21628 Vbias.n453 Vbias 0.252372
R21629 Vbias.n448 Vbias 0.252372
R21630 Vbias.n459 Vbias 0.252372
R21631 Vbias.n460 Vbias 0.252372
R21632 Vbias.n471 Vbias 0.252372
R21633 Vbias.n472 Vbias 0.252372
R21634 Vbias.n483 Vbias 0.252372
R21635 Vbias.n484 Vbias 0.252372
R21636 Vbias.n495 Vbias 0.252372
R21637 Vbias.n496 Vbias 0.252372
R21638 Vbias.n507 Vbias 0.252372
R21639 Vbias.n508 Vbias 0.252372
R21640 Vbias.n519 Vbias 0.252372
R21641 Vbias.n520 Vbias 0.252372
R21642 Vbias.n399 Vbias 0.252372
R21643 Vbias Vbias.n398 0.252372
R21644 Vbias.n390 Vbias 0.252372
R21645 Vbias.n382 Vbias 0.252372
R21646 Vbias.n381 Vbias 0.252372
R21647 Vbias.n378 Vbias 0.252372
R21648 Vbias.n375 Vbias 0.252372
R21649 Vbias.n372 Vbias 0.252372
R21650 Vbias.n369 Vbias 0.252372
R21651 Vbias.n366 Vbias 0.252372
R21652 Vbias.n363 Vbias 0.252372
R21653 Vbias.n360 Vbias 0.252372
R21654 Vbias.n357 Vbias 0.252372
R21655 Vbias.n354 Vbias 0.252372
R21656 Vbias.n351 Vbias 0.252372
R21657 Vbias.n348 Vbias 0.252372
R21658 Vbias.n345 Vbias 0.252372
R21659 Vbias Vbias.n443 0.252372
R21660 Vbias Vbias.n440 0.252372
R21661 Vbias Vbias.n437 0.252372
R21662 Vbias Vbias.n434 0.252372
R21663 Vbias Vbias.n431 0.252372
R21664 Vbias Vbias.n428 0.252372
R21665 Vbias Vbias.n425 0.252372
R21666 Vbias Vbias.n422 0.252372
R21667 Vbias Vbias.n419 0.252372
R21668 Vbias Vbias.n416 0.252372
R21669 Vbias Vbias.n413 0.252372
R21670 Vbias Vbias.n410 0.252372
R21671 Vbias Vbias.n407 0.252372
R21672 Vbias Vbias.n404 0.252372
R21673 Vbias.n386 Vbias 0.252372
R21674 Vbias.n385 Vbias.n342 0.227144
R21675 Vbias.n391 Vbias.n342 0.184322
R21676 Vbias.n344 Vbias.n332 0.175179
R21677 Vbias.n450 Vbias.n449 0.175179
R21678 Vbias.n452 Vbias.n451 0.175179
R21679 Vbias.n579 Vbias.n277 0.175179
R21680 Vbias.n587 Vbias.n586 0.175179
R21681 Vbias.n589 Vbias.n588 0.175179
R21682 Vbias.n198 Vbias.n151 0.175179
R21683 Vbias.n783 Vbias.n782 0.175179
R21684 Vbias.n781 Vbias.n780 0.175179
R21685 Vbias.n791 Vbias.n104 0.175179
R21686 Vbias.n911 Vbias.n910 0.175179
R21687 Vbias.n913 Vbias.n912 0.175179
R21688 Vbias.n98 Vbias.n55 0.175179
R21689 Vbias.n922 Vbias.n921 0.175179
R21690 Vbias.n347 Vbias.n327 0.175179
R21691 Vbias.n458 Vbias.n457 0.175179
R21692 Vbias.n456 Vbias.n455 0.175179
R21693 Vbias.n576 Vbias.n274 0.175179
R21694 Vbias.n595 Vbias.n594 0.175179
R21695 Vbias.n593 Vbias.n592 0.175179
R21696 Vbias.n201 Vbias.n154 0.175179
R21697 Vbias.n775 Vbias.n774 0.175179
R21698 Vbias.n777 Vbias.n776 0.175179
R21699 Vbias.n794 Vbias.n107 0.175179
R21700 Vbias.n905 Vbias.n904 0.175179
R21701 Vbias.n903 Vbias.n902 0.175179
R21702 Vbias.n95 Vbias.n52 0.175179
R21703 Vbias.n928 Vbias.n927 0.175179
R21704 Vbias.n350 Vbias.n324 0.175179
R21705 Vbias.n462 Vbias.n461 0.175179
R21706 Vbias.n464 Vbias.n463 0.175179
R21707 Vbias.n573 Vbias.n271 0.175179
R21708 Vbias.n599 Vbias.n598 0.175179
R21709 Vbias.n601 Vbias.n600 0.175179
R21710 Vbias.n204 Vbias.n157 0.175179
R21711 Vbias.n771 Vbias.n770 0.175179
R21712 Vbias.n769 Vbias.n768 0.175179
R21713 Vbias.n797 Vbias.n110 0.175179
R21714 Vbias.n897 Vbias.n896 0.175179
R21715 Vbias.n899 Vbias.n898 0.175179
R21716 Vbias.n92 Vbias.n49 0.175179
R21717 Vbias.n932 Vbias.n931 0.175179
R21718 Vbias.n353 Vbias.n321 0.175179
R21719 Vbias.n470 Vbias.n469 0.175179
R21720 Vbias.n468 Vbias.n467 0.175179
R21721 Vbias.n570 Vbias.n268 0.175179
R21722 Vbias.n607 Vbias.n606 0.175179
R21723 Vbias.n605 Vbias.n604 0.175179
R21724 Vbias.n207 Vbias.n160 0.175179
R21725 Vbias.n763 Vbias.n762 0.175179
R21726 Vbias.n765 Vbias.n764 0.175179
R21727 Vbias.n800 Vbias.n113 0.175179
R21728 Vbias.n893 Vbias.n892 0.175179
R21729 Vbias.n891 Vbias.n890 0.175179
R21730 Vbias.n89 Vbias.n46 0.175179
R21731 Vbias.n938 Vbias.n937 0.175179
R21732 Vbias.n356 Vbias.n318 0.175179
R21733 Vbias.n474 Vbias.n473 0.175179
R21734 Vbias.n476 Vbias.n475 0.175179
R21735 Vbias.n567 Vbias.n265 0.175179
R21736 Vbias.n611 Vbias.n610 0.175179
R21737 Vbias.n613 Vbias.n612 0.175179
R21738 Vbias.n210 Vbias.n163 0.175179
R21739 Vbias.n759 Vbias.n758 0.175179
R21740 Vbias.n757 Vbias.n756 0.175179
R21741 Vbias.n803 Vbias.n116 0.175179
R21742 Vbias.n885 Vbias.n884 0.175179
R21743 Vbias.n887 Vbias.n886 0.175179
R21744 Vbias.n86 Vbias.n43 0.175179
R21745 Vbias.n942 Vbias.n941 0.175179
R21746 Vbias.n359 Vbias.n315 0.175179
R21747 Vbias.n482 Vbias.n481 0.175179
R21748 Vbias.n480 Vbias.n479 0.175179
R21749 Vbias.n564 Vbias.n262 0.175179
R21750 Vbias.n619 Vbias.n618 0.175179
R21751 Vbias.n617 Vbias.n616 0.175179
R21752 Vbias.n213 Vbias.n166 0.175179
R21753 Vbias.n751 Vbias.n750 0.175179
R21754 Vbias.n753 Vbias.n752 0.175179
R21755 Vbias.n806 Vbias.n119 0.175179
R21756 Vbias.n881 Vbias.n880 0.175179
R21757 Vbias.n879 Vbias.n878 0.175179
R21758 Vbias.n83 Vbias.n40 0.175179
R21759 Vbias.n948 Vbias.n947 0.175179
R21760 Vbias.n362 Vbias.n312 0.175179
R21761 Vbias.n486 Vbias.n485 0.175179
R21762 Vbias.n488 Vbias.n487 0.175179
R21763 Vbias.n561 Vbias.n259 0.175179
R21764 Vbias.n623 Vbias.n622 0.175179
R21765 Vbias.n625 Vbias.n624 0.175179
R21766 Vbias.n216 Vbias.n169 0.175179
R21767 Vbias.n747 Vbias.n746 0.175179
R21768 Vbias.n745 Vbias.n744 0.175179
R21769 Vbias.n809 Vbias.n122 0.175179
R21770 Vbias.n873 Vbias.n872 0.175179
R21771 Vbias.n875 Vbias.n874 0.175179
R21772 Vbias.n80 Vbias.n37 0.175179
R21773 Vbias.n952 Vbias.n951 0.175179
R21774 Vbias.n365 Vbias.n309 0.175179
R21775 Vbias.n494 Vbias.n493 0.175179
R21776 Vbias.n492 Vbias.n491 0.175179
R21777 Vbias.n558 Vbias.n256 0.175179
R21778 Vbias.n631 Vbias.n630 0.175179
R21779 Vbias.n629 Vbias.n628 0.175179
R21780 Vbias.n219 Vbias.n172 0.175179
R21781 Vbias.n739 Vbias.n738 0.175179
R21782 Vbias.n741 Vbias.n740 0.175179
R21783 Vbias.n812 Vbias.n125 0.175179
R21784 Vbias.n869 Vbias.n868 0.175179
R21785 Vbias.n867 Vbias.n866 0.175179
R21786 Vbias.n77 Vbias.n34 0.175179
R21787 Vbias.n958 Vbias.n957 0.175179
R21788 Vbias.n368 Vbias.n306 0.175179
R21789 Vbias.n498 Vbias.n497 0.175179
R21790 Vbias.n500 Vbias.n499 0.175179
R21791 Vbias.n555 Vbias.n253 0.175179
R21792 Vbias.n635 Vbias.n634 0.175179
R21793 Vbias.n637 Vbias.n636 0.175179
R21794 Vbias.n222 Vbias.n175 0.175179
R21795 Vbias.n735 Vbias.n734 0.175179
R21796 Vbias.n733 Vbias.n732 0.175179
R21797 Vbias.n815 Vbias.n128 0.175179
R21798 Vbias.n861 Vbias.n860 0.175179
R21799 Vbias.n863 Vbias.n862 0.175179
R21800 Vbias.n74 Vbias.n31 0.175179
R21801 Vbias.n962 Vbias.n961 0.175179
R21802 Vbias.n371 Vbias.n303 0.175179
R21803 Vbias.n506 Vbias.n505 0.175179
R21804 Vbias.n504 Vbias.n503 0.175179
R21805 Vbias.n552 Vbias.n250 0.175179
R21806 Vbias.n643 Vbias.n642 0.175179
R21807 Vbias.n641 Vbias.n640 0.175179
R21808 Vbias.n225 Vbias.n178 0.175179
R21809 Vbias.n727 Vbias.n726 0.175179
R21810 Vbias.n729 Vbias.n728 0.175179
R21811 Vbias.n818 Vbias.n131 0.175179
R21812 Vbias.n857 Vbias.n856 0.175179
R21813 Vbias.n855 Vbias.n854 0.175179
R21814 Vbias.n71 Vbias.n28 0.175179
R21815 Vbias.n968 Vbias.n967 0.175179
R21816 Vbias.n374 Vbias.n300 0.175179
R21817 Vbias.n510 Vbias.n509 0.175179
R21818 Vbias.n512 Vbias.n511 0.175179
R21819 Vbias.n549 Vbias.n247 0.175179
R21820 Vbias.n647 Vbias.n646 0.175179
R21821 Vbias.n649 Vbias.n648 0.175179
R21822 Vbias.n228 Vbias.n181 0.175179
R21823 Vbias.n723 Vbias.n722 0.175179
R21824 Vbias.n721 Vbias.n720 0.175179
R21825 Vbias.n821 Vbias.n134 0.175179
R21826 Vbias.n849 Vbias.n848 0.175179
R21827 Vbias.n851 Vbias.n850 0.175179
R21828 Vbias.n68 Vbias.n25 0.175179
R21829 Vbias.n972 Vbias.n971 0.175179
R21830 Vbias.n377 Vbias.n297 0.175179
R21831 Vbias.n518 Vbias.n517 0.175179
R21832 Vbias.n516 Vbias.n515 0.175179
R21833 Vbias.n546 Vbias.n244 0.175179
R21834 Vbias.n655 Vbias.n654 0.175179
R21835 Vbias.n653 Vbias.n652 0.175179
R21836 Vbias.n231 Vbias.n184 0.175179
R21837 Vbias.n715 Vbias.n714 0.175179
R21838 Vbias.n717 Vbias.n716 0.175179
R21839 Vbias.n824 Vbias.n137 0.175179
R21840 Vbias.n845 Vbias.n844 0.175179
R21841 Vbias.n843 Vbias.n842 0.175179
R21842 Vbias.n65 Vbias.n22 0.175179
R21843 Vbias.n978 Vbias.n977 0.175179
R21844 Vbias.n380 Vbias.n294 0.175179
R21845 Vbias.n522 Vbias.n521 0.175179
R21846 Vbias.n524 Vbias.n523 0.175179
R21847 Vbias.n543 Vbias.n241 0.175179
R21848 Vbias.n659 Vbias.n658 0.175179
R21849 Vbias.n661 Vbias.n660 0.175179
R21850 Vbias.n234 Vbias.n187 0.175179
R21851 Vbias.n711 Vbias.n710 0.175179
R21852 Vbias.n709 Vbias.n708 0.175179
R21853 Vbias.n827 Vbias.n140 0.175179
R21854 Vbias.n837 Vbias.n836 0.175179
R21855 Vbias.n839 Vbias.n838 0.175179
R21856 Vbias.n62 Vbias.n17 0.175179
R21857 Vbias.n982 Vbias.n981 0.175179
R21858 Vbias.n402 Vbias.n340 0.175179
R21859 Vbias.n401 Vbias.n400 0.175179
R21860 Vbias.n527 Vbias.n286 0.175179
R21861 Vbias.n540 Vbias.n539 0.175179
R21862 Vbias.n538 Vbias.n537 0.175179
R21863 Vbias.n664 Vbias.n237 0.175179
R21864 Vbias.n695 Vbias.n694 0.175179
R21865 Vbias.n693 Vbias.n692 0.175179
R21866 Vbias.n705 Vbias.n143 0.175179
R21867 Vbias.n831 Vbias.n830 0.175179
R21868 Vbias.n833 Vbias.n832 0.175179
R21869 Vbias.n673 Vbias.n12 0.175179
R21870 Vbias.n989 Vbias.n988 0.175179
R21871 Vbias.n987 Vbias.n14 0.175179
R21872 Vbias.n919 Vbias.n918 0.175179
R21873 Vbias.n994 Vbias.n8 0.175179
R21874 Vbias.n993 Vbias.n992 0.175179
R21875 Vbias.n917 Vbias.n100 0.175179
R21876 Vbias.n916 Vbias.n915 0.175179
R21877 Vbias.n676 Vbias.n9 0.175179
R21878 Vbias.n681 Vbias.n680 0.175179
R21879 Vbias.n908 Vbias.n101 0.175179
R21880 Vbias.n789 Vbias.n788 0.175179
R21881 Vbias.n685 Vbias.n190 0.175179
R21882 Vbias.n702 Vbias.n701 0.175179
R21883 Vbias.n787 Vbias.n147 0.175179
R21884 Vbias.n786 Vbias.n785 0.175179
R21885 Vbias.n700 Vbias.n192 0.175179
R21886 Vbias.n699 Vbias.n698 0.175179
R21887 Vbias.n196 Vbias.n148 0.175179
R21888 Vbias.n282 Vbias.n281 0.175179
R21889 Vbias.n667 Vbias.n193 0.175179
R21890 Vbias.n534 Vbias.n533 0.175179
R21891 Vbias.n584 Vbias.n583 0.175179
R21892 Vbias.n582 Vbias.n581 0.175179
R21893 Vbias.n532 Vbias.n290 0.175179
R21894 Vbias.n531 Vbias.n530 0.175179
R21895 Vbias.n330 Vbias.n283 0.175179
R21896 Vbias.n447 Vbias.n446 0.175179
R21897 Vbias.n397 Vbias.n291 0.175179
R21898 Vbias.n389 Vbias.n388 0.175179
R21899 Vbias.n445 Vbias.n336 0.175179
R21900 Vbias.n398 Vbias 0.0972718
R21901 Vbias Vbias.n392 0.0972718
R21902 Vbias Vbias.n668 0.0972718
R21903 Vbias.n690 Vbias 0.0972718
R21904 Vbias Vbias.n686 0.0972718
R21905 Vbias Vbias.n677 0.0972718
R21906 Vbias.n19 Vbias 0.0972718
R21907 Vbias Vbias.n996 0.0972718
R21908 Vbias.n985 Vbias 0.0972718
R21909 Vbias Vbias.n984 0.0972718
R21910 Vbias.n975 Vbias 0.0972718
R21911 Vbias Vbias.n974 0.0972718
R21912 Vbias.n965 Vbias 0.0972718
R21913 Vbias Vbias.n964 0.0972718
R21914 Vbias.n955 Vbias 0.0972718
R21915 Vbias Vbias.n954 0.0972718
R21916 Vbias.n945 Vbias 0.0972718
R21917 Vbias Vbias.n944 0.0972718
R21918 Vbias.n935 Vbias 0.0972718
R21919 Vbias Vbias.n934 0.0972718
R21920 Vbias.n925 Vbias 0.0972718
R21921 Vbias Vbias.n924 0.0972718
R21922 Vbias.n920 Vbias 0.0972718
R21923 Vbias Vbias.n929 0.0972718
R21924 Vbias.n930 Vbias 0.0972718
R21925 Vbias Vbias.n939 0.0972718
R21926 Vbias.n940 Vbias 0.0972718
R21927 Vbias Vbias.n949 0.0972718
R21928 Vbias.n950 Vbias 0.0972718
R21929 Vbias Vbias.n959 0.0972718
R21930 Vbias.n960 Vbias 0.0972718
R21931 Vbias Vbias.n969 0.0972718
R21932 Vbias.n970 Vbias 0.0972718
R21933 Vbias Vbias.n979 0.0972718
R21934 Vbias.n980 Vbias 0.0972718
R21935 Vbias.n20 Vbias 0.0972718
R21936 Vbias.n991 Vbias 0.0972718
R21937 Vbias Vbias.n990 0.0972718
R21938 Vbias.n63 Vbias 0.0972718
R21939 Vbias.n66 Vbias 0.0972718
R21940 Vbias.n69 Vbias 0.0972718
R21941 Vbias.n72 Vbias 0.0972718
R21942 Vbias.n75 Vbias 0.0972718
R21943 Vbias.n78 Vbias 0.0972718
R21944 Vbias.n81 Vbias 0.0972718
R21945 Vbias.n84 Vbias 0.0972718
R21946 Vbias.n87 Vbias 0.0972718
R21947 Vbias.n90 Vbias 0.0972718
R21948 Vbias.n93 Vbias 0.0972718
R21949 Vbias.n96 Vbias 0.0972718
R21950 Vbias.n99 Vbias 0.0972718
R21951 Vbias.n914 Vbias 0.0972718
R21952 Vbias.n901 Vbias 0.0972718
R21953 Vbias.n900 Vbias 0.0972718
R21954 Vbias.n889 Vbias 0.0972718
R21955 Vbias.n888 Vbias 0.0972718
R21956 Vbias.n877 Vbias 0.0972718
R21957 Vbias.n876 Vbias 0.0972718
R21958 Vbias.n865 Vbias 0.0972718
R21959 Vbias.n864 Vbias 0.0972718
R21960 Vbias.n853 Vbias 0.0972718
R21961 Vbias.n852 Vbias 0.0972718
R21962 Vbias.n841 Vbias 0.0972718
R21963 Vbias.n840 Vbias 0.0972718
R21964 Vbias Vbias.n674 0.0972718
R21965 Vbias Vbias.n682 0.0972718
R21966 Vbias.n834 Vbias 0.0972718
R21967 Vbias.n835 Vbias 0.0972718
R21968 Vbias.n846 Vbias 0.0972718
R21969 Vbias.n847 Vbias 0.0972718
R21970 Vbias.n858 Vbias 0.0972718
R21971 Vbias.n859 Vbias 0.0972718
R21972 Vbias.n870 Vbias 0.0972718
R21973 Vbias.n871 Vbias 0.0972718
R21974 Vbias.n882 Vbias 0.0972718
R21975 Vbias.n883 Vbias 0.0972718
R21976 Vbias.n894 Vbias 0.0972718
R21977 Vbias.n895 Vbias 0.0972718
R21978 Vbias.n906 Vbias 0.0972718
R21979 Vbias.n909 Vbias 0.0972718
R21980 Vbias Vbias.n792 0.0972718
R21981 Vbias Vbias.n795 0.0972718
R21982 Vbias Vbias.n798 0.0972718
R21983 Vbias Vbias.n801 0.0972718
R21984 Vbias Vbias.n804 0.0972718
R21985 Vbias Vbias.n807 0.0972718
R21986 Vbias Vbias.n810 0.0972718
R21987 Vbias Vbias.n813 0.0972718
R21988 Vbias Vbias.n816 0.0972718
R21989 Vbias Vbias.n819 0.0972718
R21990 Vbias Vbias.n822 0.0972718
R21991 Vbias Vbias.n825 0.0972718
R21992 Vbias Vbias.n828 0.0972718
R21993 Vbias.n829 Vbias 0.0972718
R21994 Vbias.n703 Vbias 0.0972718
R21995 Vbias.n706 Vbias 0.0972718
R21996 Vbias.n707 Vbias 0.0972718
R21997 Vbias.n718 Vbias 0.0972718
R21998 Vbias.n719 Vbias 0.0972718
R21999 Vbias.n730 Vbias 0.0972718
R22000 Vbias.n731 Vbias 0.0972718
R22001 Vbias.n742 Vbias 0.0972718
R22002 Vbias.n743 Vbias 0.0972718
R22003 Vbias.n754 Vbias 0.0972718
R22004 Vbias.n755 Vbias 0.0972718
R22005 Vbias.n766 Vbias 0.0972718
R22006 Vbias.n767 Vbias 0.0972718
R22007 Vbias.n778 Vbias 0.0972718
R22008 Vbias.n779 Vbias 0.0972718
R22009 Vbias.n784 Vbias 0.0972718
R22010 Vbias.n773 Vbias 0.0972718
R22011 Vbias.n772 Vbias 0.0972718
R22012 Vbias.n761 Vbias 0.0972718
R22013 Vbias.n760 Vbias 0.0972718
R22014 Vbias.n749 Vbias 0.0972718
R22015 Vbias.n748 Vbias 0.0972718
R22016 Vbias.n737 Vbias 0.0972718
R22017 Vbias.n736 Vbias 0.0972718
R22018 Vbias.n725 Vbias 0.0972718
R22019 Vbias.n724 Vbias 0.0972718
R22020 Vbias.n713 Vbias 0.0972718
R22021 Vbias.n712 Vbias 0.0972718
R22022 Vbias.n691 Vbias 0.0972718
R22023 Vbias.n697 Vbias 0.0972718
R22024 Vbias Vbias.n696 0.0972718
R22025 Vbias Vbias.n235 0.0972718
R22026 Vbias Vbias.n232 0.0972718
R22027 Vbias Vbias.n229 0.0972718
R22028 Vbias Vbias.n226 0.0972718
R22029 Vbias Vbias.n223 0.0972718
R22030 Vbias Vbias.n220 0.0972718
R22031 Vbias Vbias.n217 0.0972718
R22032 Vbias Vbias.n214 0.0972718
R22033 Vbias Vbias.n211 0.0972718
R22034 Vbias Vbias.n208 0.0972718
R22035 Vbias Vbias.n205 0.0972718
R22036 Vbias Vbias.n202 0.0972718
R22037 Vbias Vbias.n199 0.0972718
R22038 Vbias Vbias.n590 0.0972718
R22039 Vbias.n591 Vbias 0.0972718
R22040 Vbias Vbias.n602 0.0972718
R22041 Vbias.n603 Vbias 0.0972718
R22042 Vbias Vbias.n614 0.0972718
R22043 Vbias.n615 Vbias 0.0972718
R22044 Vbias Vbias.n626 0.0972718
R22045 Vbias.n627 Vbias 0.0972718
R22046 Vbias Vbias.n638 0.0972718
R22047 Vbias.n639 Vbias 0.0972718
R22048 Vbias Vbias.n650 0.0972718
R22049 Vbias.n651 Vbias 0.0972718
R22050 Vbias Vbias.n662 0.0972718
R22051 Vbias Vbias.n665 0.0972718
R22052 Vbias.n535 Vbias 0.0972718
R22053 Vbias.n536 Vbias 0.0972718
R22054 Vbias.n657 Vbias 0.0972718
R22055 Vbias Vbias.n656 0.0972718
R22056 Vbias.n645 Vbias 0.0972718
R22057 Vbias Vbias.n644 0.0972718
R22058 Vbias.n633 Vbias 0.0972718
R22059 Vbias Vbias.n632 0.0972718
R22060 Vbias.n621 Vbias 0.0972718
R22061 Vbias Vbias.n620 0.0972718
R22062 Vbias.n609 Vbias 0.0972718
R22063 Vbias Vbias.n608 0.0972718
R22064 Vbias.n597 Vbias 0.0972718
R22065 Vbias Vbias.n596 0.0972718
R22066 Vbias.n585 Vbias 0.0972718
R22067 Vbias.n580 Vbias 0.0972718
R22068 Vbias.n577 Vbias 0.0972718
R22069 Vbias.n574 Vbias 0.0972718
R22070 Vbias.n571 Vbias 0.0972718
R22071 Vbias.n568 Vbias 0.0972718
R22072 Vbias.n565 Vbias 0.0972718
R22073 Vbias.n562 Vbias 0.0972718
R22074 Vbias.n559 Vbias 0.0972718
R22075 Vbias.n556 Vbias 0.0972718
R22076 Vbias.n553 Vbias 0.0972718
R22077 Vbias.n550 Vbias 0.0972718
R22078 Vbias.n547 Vbias 0.0972718
R22079 Vbias.n544 Vbias 0.0972718
R22080 Vbias.n541 Vbias 0.0972718
R22081 Vbias.n529 Vbias 0.0972718
R22082 Vbias Vbias.n528 0.0972718
R22083 Vbias Vbias.n525 0.0972718
R22084 Vbias.n514 Vbias 0.0972718
R22085 Vbias Vbias.n513 0.0972718
R22086 Vbias.n502 Vbias 0.0972718
R22087 Vbias Vbias.n501 0.0972718
R22088 Vbias.n490 Vbias 0.0972718
R22089 Vbias Vbias.n489 0.0972718
R22090 Vbias.n478 Vbias 0.0972718
R22091 Vbias Vbias.n477 0.0972718
R22092 Vbias.n466 Vbias 0.0972718
R22093 Vbias Vbias.n465 0.0972718
R22094 Vbias.n454 Vbias 0.0972718
R22095 Vbias Vbias.n453 0.0972718
R22096 Vbias.n448 Vbias 0.0972718
R22097 Vbias Vbias.n459 0.0972718
R22098 Vbias.n460 Vbias 0.0972718
R22099 Vbias Vbias.n471 0.0972718
R22100 Vbias.n472 Vbias 0.0972718
R22101 Vbias Vbias.n483 0.0972718
R22102 Vbias.n484 Vbias 0.0972718
R22103 Vbias Vbias.n495 0.0972718
R22104 Vbias.n496 Vbias 0.0972718
R22105 Vbias Vbias.n507 0.0972718
R22106 Vbias.n508 Vbias 0.0972718
R22107 Vbias Vbias.n519 0.0972718
R22108 Vbias.n520 Vbias 0.0972718
R22109 Vbias.n399 Vbias 0.0972718
R22110 Vbias Vbias.n390 0.0972718
R22111 Vbias Vbias.n382 0.0972718
R22112 Vbias Vbias.n381 0.0972718
R22113 Vbias Vbias.n378 0.0972718
R22114 Vbias Vbias.n375 0.0972718
R22115 Vbias Vbias.n372 0.0972718
R22116 Vbias Vbias.n369 0.0972718
R22117 Vbias Vbias.n366 0.0972718
R22118 Vbias Vbias.n363 0.0972718
R22119 Vbias Vbias.n360 0.0972718
R22120 Vbias Vbias.n357 0.0972718
R22121 Vbias Vbias.n354 0.0972718
R22122 Vbias Vbias.n351 0.0972718
R22123 Vbias Vbias.n348 0.0972718
R22124 Vbias Vbias.n345 0.0972718
R22125 Vbias.n443 Vbias 0.0972718
R22126 Vbias.n440 Vbias 0.0972718
R22127 Vbias.n437 Vbias 0.0972718
R22128 Vbias.n434 Vbias 0.0972718
R22129 Vbias.n431 Vbias 0.0972718
R22130 Vbias.n428 Vbias 0.0972718
R22131 Vbias.n425 Vbias 0.0972718
R22132 Vbias.n422 Vbias 0.0972718
R22133 Vbias.n419 Vbias 0.0972718
R22134 Vbias.n416 Vbias 0.0972718
R22135 Vbias.n413 Vbias 0.0972718
R22136 Vbias.n410 Vbias 0.0972718
R22137 Vbias.n407 Vbias 0.0972718
R22138 Vbias.n404 Vbias 0.0972718
R22139 Vbias.n386 Vbias 0.0972718
R22140 Vbias.n337 Vbias 0.0489375
R22141 Vbias.n383 Vbias 0.0489375
R22142 Vbias.n384 Vbias 0.0489375
R22143 Vbias.n334 Vbias 0.0489375
R22144 Vbias.n292 Vbias 0.0489375
R22145 Vbias.n284 Vbias 0.0489375
R22146 Vbias.n288 Vbias 0.0489375
R22147 Vbias.n280 Vbias 0.0489375
R22148 Vbias.n194 Vbias 0.0489375
R22149 Vbias.n149 Vbias 0.0489375
R22150 Vbias.n189 Vbias 0.0489375
R22151 Vbias.n145 Vbias 0.0489375
R22152 Vbias.n679 Vbias 0.0489375
R22153 Vbias.n102 Vbias 0.0489375
R22154 Vbias.n10 Vbias 0.0489375
R22155 Vbias.n57 Vbias 0.0489375
R22156 Vbias.n58 Vbias 0.0489375
R22157 Vbias.n54 Vbias 0.0489375
R22158 Vbias.n441 Vbias 0.0489375
R22159 Vbias.n343 Vbias 0.0489375
R22160 Vbias.n333 Vbias 0.0489375
R22161 Vbias.n331 Vbias 0.0489375
R22162 Vbias.n578 Vbias 0.0489375
R22163 Vbias.n278 Vbias 0.0489375
R22164 Vbias.n276 Vbias 0.0489375
R22165 Vbias.n197 Vbias 0.0489375
R22166 Vbias.n150 Vbias 0.0489375
R22167 Vbias.n152 Vbias 0.0489375
R22168 Vbias.n790 Vbias 0.0489375
R22169 Vbias.n105 Vbias 0.0489375
R22170 Vbias.n103 Vbias 0.0489375
R22171 Vbias.n97 Vbias 0.0489375
R22172 Vbias.n56 Vbias 0.0489375
R22173 Vbias.n53 Vbias 0.0489375
R22174 Vbias.n438 Vbias 0.0489375
R22175 Vbias.n346 Vbias 0.0489375
R22176 Vbias.n326 Vbias 0.0489375
R22177 Vbias.n328 Vbias 0.0489375
R22178 Vbias.n575 Vbias 0.0489375
R22179 Vbias.n273 Vbias 0.0489375
R22180 Vbias.n275 Vbias 0.0489375
R22181 Vbias.n200 Vbias 0.0489375
R22182 Vbias.n155 Vbias 0.0489375
R22183 Vbias.n153 Vbias 0.0489375
R22184 Vbias.n793 Vbias 0.0489375
R22185 Vbias.n106 Vbias 0.0489375
R22186 Vbias.n108 Vbias 0.0489375
R22187 Vbias.n94 Vbias 0.0489375
R22188 Vbias.n51 Vbias 0.0489375
R22189 Vbias.n48 Vbias 0.0489375
R22190 Vbias.n435 Vbias 0.0489375
R22191 Vbias.n349 Vbias 0.0489375
R22192 Vbias.n325 Vbias 0.0489375
R22193 Vbias.n323 Vbias 0.0489375
R22194 Vbias.n572 Vbias 0.0489375
R22195 Vbias.n272 Vbias 0.0489375
R22196 Vbias.n270 Vbias 0.0489375
R22197 Vbias.n203 Vbias 0.0489375
R22198 Vbias.n156 Vbias 0.0489375
R22199 Vbias.n158 Vbias 0.0489375
R22200 Vbias.n796 Vbias 0.0489375
R22201 Vbias.n111 Vbias 0.0489375
R22202 Vbias.n109 Vbias 0.0489375
R22203 Vbias.n91 Vbias 0.0489375
R22204 Vbias.n50 Vbias 0.0489375
R22205 Vbias.n47 Vbias 0.0489375
R22206 Vbias.n432 Vbias 0.0489375
R22207 Vbias.n352 Vbias 0.0489375
R22208 Vbias.n320 Vbias 0.0489375
R22209 Vbias.n322 Vbias 0.0489375
R22210 Vbias.n569 Vbias 0.0489375
R22211 Vbias.n267 Vbias 0.0489375
R22212 Vbias.n269 Vbias 0.0489375
R22213 Vbias.n206 Vbias 0.0489375
R22214 Vbias.n161 Vbias 0.0489375
R22215 Vbias.n159 Vbias 0.0489375
R22216 Vbias.n799 Vbias 0.0489375
R22217 Vbias.n112 Vbias 0.0489375
R22218 Vbias.n114 Vbias 0.0489375
R22219 Vbias.n88 Vbias 0.0489375
R22220 Vbias.n45 Vbias 0.0489375
R22221 Vbias.n42 Vbias 0.0489375
R22222 Vbias.n429 Vbias 0.0489375
R22223 Vbias.n355 Vbias 0.0489375
R22224 Vbias.n319 Vbias 0.0489375
R22225 Vbias.n317 Vbias 0.0489375
R22226 Vbias.n566 Vbias 0.0489375
R22227 Vbias.n266 Vbias 0.0489375
R22228 Vbias.n264 Vbias 0.0489375
R22229 Vbias.n209 Vbias 0.0489375
R22230 Vbias.n162 Vbias 0.0489375
R22231 Vbias.n164 Vbias 0.0489375
R22232 Vbias.n802 Vbias 0.0489375
R22233 Vbias.n117 Vbias 0.0489375
R22234 Vbias.n115 Vbias 0.0489375
R22235 Vbias.n85 Vbias 0.0489375
R22236 Vbias.n44 Vbias 0.0489375
R22237 Vbias.n41 Vbias 0.0489375
R22238 Vbias.n426 Vbias 0.0489375
R22239 Vbias.n358 Vbias 0.0489375
R22240 Vbias.n314 Vbias 0.0489375
R22241 Vbias.n316 Vbias 0.0489375
R22242 Vbias.n563 Vbias 0.0489375
R22243 Vbias.n261 Vbias 0.0489375
R22244 Vbias.n263 Vbias 0.0489375
R22245 Vbias.n212 Vbias 0.0489375
R22246 Vbias.n167 Vbias 0.0489375
R22247 Vbias.n165 Vbias 0.0489375
R22248 Vbias.n805 Vbias 0.0489375
R22249 Vbias.n118 Vbias 0.0489375
R22250 Vbias.n120 Vbias 0.0489375
R22251 Vbias.n82 Vbias 0.0489375
R22252 Vbias.n39 Vbias 0.0489375
R22253 Vbias.n36 Vbias 0.0489375
R22254 Vbias.n423 Vbias 0.0489375
R22255 Vbias.n361 Vbias 0.0489375
R22256 Vbias.n313 Vbias 0.0489375
R22257 Vbias.n311 Vbias 0.0489375
R22258 Vbias.n560 Vbias 0.0489375
R22259 Vbias.n260 Vbias 0.0489375
R22260 Vbias.n258 Vbias 0.0489375
R22261 Vbias.n215 Vbias 0.0489375
R22262 Vbias.n168 Vbias 0.0489375
R22263 Vbias.n170 Vbias 0.0489375
R22264 Vbias.n808 Vbias 0.0489375
R22265 Vbias.n123 Vbias 0.0489375
R22266 Vbias.n121 Vbias 0.0489375
R22267 Vbias.n79 Vbias 0.0489375
R22268 Vbias.n38 Vbias 0.0489375
R22269 Vbias.n35 Vbias 0.0489375
R22270 Vbias.n420 Vbias 0.0489375
R22271 Vbias.n364 Vbias 0.0489375
R22272 Vbias.n308 Vbias 0.0489375
R22273 Vbias.n310 Vbias 0.0489375
R22274 Vbias.n557 Vbias 0.0489375
R22275 Vbias.n255 Vbias 0.0489375
R22276 Vbias.n257 Vbias 0.0489375
R22277 Vbias.n218 Vbias 0.0489375
R22278 Vbias.n173 Vbias 0.0489375
R22279 Vbias.n171 Vbias 0.0489375
R22280 Vbias.n811 Vbias 0.0489375
R22281 Vbias.n124 Vbias 0.0489375
R22282 Vbias.n126 Vbias 0.0489375
R22283 Vbias.n76 Vbias 0.0489375
R22284 Vbias.n33 Vbias 0.0489375
R22285 Vbias.n30 Vbias 0.0489375
R22286 Vbias.n417 Vbias 0.0489375
R22287 Vbias.n367 Vbias 0.0489375
R22288 Vbias.n307 Vbias 0.0489375
R22289 Vbias.n305 Vbias 0.0489375
R22290 Vbias.n554 Vbias 0.0489375
R22291 Vbias.n254 Vbias 0.0489375
R22292 Vbias.n252 Vbias 0.0489375
R22293 Vbias.n221 Vbias 0.0489375
R22294 Vbias.n174 Vbias 0.0489375
R22295 Vbias.n176 Vbias 0.0489375
R22296 Vbias.n814 Vbias 0.0489375
R22297 Vbias.n129 Vbias 0.0489375
R22298 Vbias.n127 Vbias 0.0489375
R22299 Vbias.n73 Vbias 0.0489375
R22300 Vbias.n32 Vbias 0.0489375
R22301 Vbias.n29 Vbias 0.0489375
R22302 Vbias.n414 Vbias 0.0489375
R22303 Vbias.n370 Vbias 0.0489375
R22304 Vbias.n302 Vbias 0.0489375
R22305 Vbias.n304 Vbias 0.0489375
R22306 Vbias.n551 Vbias 0.0489375
R22307 Vbias.n249 Vbias 0.0489375
R22308 Vbias.n251 Vbias 0.0489375
R22309 Vbias.n224 Vbias 0.0489375
R22310 Vbias.n179 Vbias 0.0489375
R22311 Vbias.n177 Vbias 0.0489375
R22312 Vbias.n817 Vbias 0.0489375
R22313 Vbias.n130 Vbias 0.0489375
R22314 Vbias.n132 Vbias 0.0489375
R22315 Vbias.n70 Vbias 0.0489375
R22316 Vbias.n27 Vbias 0.0489375
R22317 Vbias.n24 Vbias 0.0489375
R22318 Vbias.n411 Vbias 0.0489375
R22319 Vbias.n373 Vbias 0.0489375
R22320 Vbias.n301 Vbias 0.0489375
R22321 Vbias.n299 Vbias 0.0489375
R22322 Vbias.n548 Vbias 0.0489375
R22323 Vbias.n248 Vbias 0.0489375
R22324 Vbias.n246 Vbias 0.0489375
R22325 Vbias.n227 Vbias 0.0489375
R22326 Vbias.n180 Vbias 0.0489375
R22327 Vbias.n182 Vbias 0.0489375
R22328 Vbias.n820 Vbias 0.0489375
R22329 Vbias.n135 Vbias 0.0489375
R22330 Vbias.n133 Vbias 0.0489375
R22331 Vbias.n67 Vbias 0.0489375
R22332 Vbias.n26 Vbias 0.0489375
R22333 Vbias.n23 Vbias 0.0489375
R22334 Vbias.n408 Vbias 0.0489375
R22335 Vbias.n376 Vbias 0.0489375
R22336 Vbias.n296 Vbias 0.0489375
R22337 Vbias.n298 Vbias 0.0489375
R22338 Vbias.n545 Vbias 0.0489375
R22339 Vbias.n243 Vbias 0.0489375
R22340 Vbias.n245 Vbias 0.0489375
R22341 Vbias.n230 Vbias 0.0489375
R22342 Vbias.n185 Vbias 0.0489375
R22343 Vbias.n183 Vbias 0.0489375
R22344 Vbias.n823 Vbias 0.0489375
R22345 Vbias.n136 Vbias 0.0489375
R22346 Vbias.n138 Vbias 0.0489375
R22347 Vbias.n64 Vbias 0.0489375
R22348 Vbias.n21 Vbias 0.0489375
R22349 Vbias.n16 Vbias 0.0489375
R22350 Vbias.n405 Vbias 0.0489375
R22351 Vbias.n379 Vbias 0.0489375
R22352 Vbias.n295 Vbias 0.0489375
R22353 Vbias.n293 Vbias 0.0489375
R22354 Vbias.n542 Vbias 0.0489375
R22355 Vbias.n242 Vbias 0.0489375
R22356 Vbias.n240 Vbias 0.0489375
R22357 Vbias.n233 Vbias 0.0489375
R22358 Vbias.n186 Vbias 0.0489375
R22359 Vbias.n188 Vbias 0.0489375
R22360 Vbias.n826 Vbias 0.0489375
R22361 Vbias.n141 Vbias 0.0489375
R22362 Vbias.n139 Vbias 0.0489375
R22363 Vbias.n61 Vbias 0.0489375
R22364 Vbias.n18 Vbias 0.0489375
R22365 Vbias.n15 Vbias 0.0489375
R22366 Vbias.n338 Vbias 0.0489375
R22367 Vbias.n339 Vbias 0.0489375
R22368 Vbias.n341 Vbias 0.0489375
R22369 Vbias.n526 Vbias 0.0489375
R22370 Vbias.n285 Vbias 0.0489375
R22371 Vbias.n287 Vbias 0.0489375
R22372 Vbias.n663 Vbias 0.0489375
R22373 Vbias.n236 Vbias 0.0489375
R22374 Vbias.n238 Vbias 0.0489375
R22375 Vbias.n704 Vbias 0.0489375
R22376 Vbias.n144 Vbias 0.0489375
R22377 Vbias.n142 Vbias 0.0489375
R22378 Vbias.n672 Vbias 0.0489375
R22379 Vbias.n11 Vbias 0.0489375
R22380 Vbias.n13 Vbias 0.0489375
R22381 Vbias.n6 Vbias 0.0489375
R22382 Vbias.n7 Vbias 0.0489375
R22383 Vbias.n60 Vbias 0.0489375
R22384 Vbias.n675 Vbias 0.0489375
R22385 Vbias.n907 Vbias 0.0489375
R22386 Vbias.n684 Vbias 0.0489375
R22387 Vbias.n146 Vbias 0.0489375
R22388 Vbias.n191 Vbias 0.0489375
R22389 Vbias.n195 Vbias 0.0489375
R22390 Vbias.n666 Vbias 0.0489375
R22391 Vbias.n279 Vbias 0.0489375
R22392 Vbias.n289 Vbias 0.0489375
R22393 Vbias.n329 Vbias 0.0489375
R22394 Vbias.n396 Vbias 0.0489375
R22395 Vbias.n335 Vbias 0.0489375
R22396 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R22397 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R22398 XThC.Tn[1].n71 XThC.Tn[1].n69 161.365
R22399 XThC.Tn[1].n67 XThC.Tn[1].n65 161.365
R22400 XThC.Tn[1].n63 XThC.Tn[1].n61 161.365
R22401 XThC.Tn[1].n59 XThC.Tn[1].n57 161.365
R22402 XThC.Tn[1].n55 XThC.Tn[1].n53 161.365
R22403 XThC.Tn[1].n51 XThC.Tn[1].n49 161.365
R22404 XThC.Tn[1].n47 XThC.Tn[1].n45 161.365
R22405 XThC.Tn[1].n43 XThC.Tn[1].n41 161.365
R22406 XThC.Tn[1].n39 XThC.Tn[1].n37 161.365
R22407 XThC.Tn[1].n35 XThC.Tn[1].n33 161.365
R22408 XThC.Tn[1].n31 XThC.Tn[1].n29 161.365
R22409 XThC.Tn[1].n27 XThC.Tn[1].n25 161.365
R22410 XThC.Tn[1].n23 XThC.Tn[1].n21 161.365
R22411 XThC.Tn[1].n19 XThC.Tn[1].n17 161.365
R22412 XThC.Tn[1].n15 XThC.Tn[1].n13 161.365
R22413 XThC.Tn[1].n12 XThC.Tn[1].n10 161.365
R22414 XThC.Tn[1].n69 XThC.Tn[1].t35 161.202
R22415 XThC.Tn[1].n65 XThC.Tn[1].t25 161.202
R22416 XThC.Tn[1].n61 XThC.Tn[1].t12 161.202
R22417 XThC.Tn[1].n57 XThC.Tn[1].t41 161.202
R22418 XThC.Tn[1].n53 XThC.Tn[1].t33 161.202
R22419 XThC.Tn[1].n49 XThC.Tn[1].t20 161.202
R22420 XThC.Tn[1].n45 XThC.Tn[1].t19 161.202
R22421 XThC.Tn[1].n41 XThC.Tn[1].t32 161.202
R22422 XThC.Tn[1].n37 XThC.Tn[1].t30 161.202
R22423 XThC.Tn[1].n33 XThC.Tn[1].t21 161.202
R22424 XThC.Tn[1].n29 XThC.Tn[1].t40 161.202
R22425 XThC.Tn[1].n25 XThC.Tn[1].t39 161.202
R22426 XThC.Tn[1].n21 XThC.Tn[1].t18 161.202
R22427 XThC.Tn[1].n17 XThC.Tn[1].t16 161.202
R22428 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R22429 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R22430 XThC.Tn[1].n69 XThC.Tn[1].t38 145.137
R22431 XThC.Tn[1].n65 XThC.Tn[1].t28 145.137
R22432 XThC.Tn[1].n61 XThC.Tn[1].t15 145.137
R22433 XThC.Tn[1].n57 XThC.Tn[1].t13 145.137
R22434 XThC.Tn[1].n53 XThC.Tn[1].t37 145.137
R22435 XThC.Tn[1].n49 XThC.Tn[1].t26 145.137
R22436 XThC.Tn[1].n45 XThC.Tn[1].t24 145.137
R22437 XThC.Tn[1].n41 XThC.Tn[1].t36 145.137
R22438 XThC.Tn[1].n37 XThC.Tn[1].t34 145.137
R22439 XThC.Tn[1].n33 XThC.Tn[1].t27 145.137
R22440 XThC.Tn[1].n29 XThC.Tn[1].t43 145.137
R22441 XThC.Tn[1].n25 XThC.Tn[1].t42 145.137
R22442 XThC.Tn[1].n21 XThC.Tn[1].t23 145.137
R22443 XThC.Tn[1].n17 XThC.Tn[1].t22 145.137
R22444 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R22445 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R22446 XThC.Tn[1].n7 XThC.Tn[1].n6 135.249
R22447 XThC.Tn[1].n9 XThC.Tn[1].n3 98.981
R22448 XThC.Tn[1].n8 XThC.Tn[1].n4 98.981
R22449 XThC.Tn[1].n7 XThC.Tn[1].n5 98.981
R22450 XThC.Tn[1].n9 XThC.Tn[1].n8 36.2672
R22451 XThC.Tn[1].n8 XThC.Tn[1].n7 36.2672
R22452 XThC.Tn[1].n74 XThC.Tn[1].n9 32.6405
R22453 XThC.Tn[1].n1 XThC.Tn[1].t5 26.5955
R22454 XThC.Tn[1].n1 XThC.Tn[1].t4 26.5955
R22455 XThC.Tn[1].n0 XThC.Tn[1].t7 26.5955
R22456 XThC.Tn[1].n0 XThC.Tn[1].t6 26.5955
R22457 XThC.Tn[1].n3 XThC.Tn[1].t9 24.9236
R22458 XThC.Tn[1].n3 XThC.Tn[1].t8 24.9236
R22459 XThC.Tn[1].n4 XThC.Tn[1].t11 24.9236
R22460 XThC.Tn[1].n4 XThC.Tn[1].t10 24.9236
R22461 XThC.Tn[1].n5 XThC.Tn[1].t1 24.9236
R22462 XThC.Tn[1].n5 XThC.Tn[1].t0 24.9236
R22463 XThC.Tn[1].n6 XThC.Tn[1].t3 24.9236
R22464 XThC.Tn[1].n6 XThC.Tn[1].t2 24.9236
R22465 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R22466 XThC.Tn[1] XThC.Tn[1].n12 8.0245
R22467 XThC.Tn[1].n72 XThC.Tn[1].n71 7.9105
R22468 XThC.Tn[1].n68 XThC.Tn[1].n67 7.9105
R22469 XThC.Tn[1].n64 XThC.Tn[1].n63 7.9105
R22470 XThC.Tn[1].n60 XThC.Tn[1].n59 7.9105
R22471 XThC.Tn[1].n56 XThC.Tn[1].n55 7.9105
R22472 XThC.Tn[1].n52 XThC.Tn[1].n51 7.9105
R22473 XThC.Tn[1].n48 XThC.Tn[1].n47 7.9105
R22474 XThC.Tn[1].n44 XThC.Tn[1].n43 7.9105
R22475 XThC.Tn[1].n40 XThC.Tn[1].n39 7.9105
R22476 XThC.Tn[1].n36 XThC.Tn[1].n35 7.9105
R22477 XThC.Tn[1].n32 XThC.Tn[1].n31 7.9105
R22478 XThC.Tn[1].n28 XThC.Tn[1].n27 7.9105
R22479 XThC.Tn[1].n24 XThC.Tn[1].n23 7.9105
R22480 XThC.Tn[1].n20 XThC.Tn[1].n19 7.9105
R22481 XThC.Tn[1].n16 XThC.Tn[1].n15 7.9105
R22482 XThC.Tn[1] XThC.Tn[1].n74 6.7205
R22483 XThC.Tn[1].n73 XThC.Tn[1] 6.08068
R22484 XThC.Tn[1].n74 XThC.Tn[1].n73 4.65249
R22485 XThC.Tn[1].n73 XThC.Tn[1] 1.8942
R22486 XThC.Tn[1].n16 XThC.Tn[1] 0.235138
R22487 XThC.Tn[1].n20 XThC.Tn[1] 0.235138
R22488 XThC.Tn[1].n24 XThC.Tn[1] 0.235138
R22489 XThC.Tn[1].n28 XThC.Tn[1] 0.235138
R22490 XThC.Tn[1].n32 XThC.Tn[1] 0.235138
R22491 XThC.Tn[1].n36 XThC.Tn[1] 0.235138
R22492 XThC.Tn[1].n40 XThC.Tn[1] 0.235138
R22493 XThC.Tn[1].n44 XThC.Tn[1] 0.235138
R22494 XThC.Tn[1].n48 XThC.Tn[1] 0.235138
R22495 XThC.Tn[1].n52 XThC.Tn[1] 0.235138
R22496 XThC.Tn[1].n56 XThC.Tn[1] 0.235138
R22497 XThC.Tn[1].n60 XThC.Tn[1] 0.235138
R22498 XThC.Tn[1].n64 XThC.Tn[1] 0.235138
R22499 XThC.Tn[1].n68 XThC.Tn[1] 0.235138
R22500 XThC.Tn[1].n72 XThC.Tn[1] 0.235138
R22501 XThC.Tn[1] XThC.Tn[1].n16 0.114505
R22502 XThC.Tn[1] XThC.Tn[1].n20 0.114505
R22503 XThC.Tn[1] XThC.Tn[1].n24 0.114505
R22504 XThC.Tn[1] XThC.Tn[1].n28 0.114505
R22505 XThC.Tn[1] XThC.Tn[1].n32 0.114505
R22506 XThC.Tn[1] XThC.Tn[1].n36 0.114505
R22507 XThC.Tn[1] XThC.Tn[1].n40 0.114505
R22508 XThC.Tn[1] XThC.Tn[1].n44 0.114505
R22509 XThC.Tn[1] XThC.Tn[1].n48 0.114505
R22510 XThC.Tn[1] XThC.Tn[1].n52 0.114505
R22511 XThC.Tn[1] XThC.Tn[1].n56 0.114505
R22512 XThC.Tn[1] XThC.Tn[1].n60 0.114505
R22513 XThC.Tn[1] XThC.Tn[1].n64 0.114505
R22514 XThC.Tn[1] XThC.Tn[1].n68 0.114505
R22515 XThC.Tn[1] XThC.Tn[1].n72 0.114505
R22516 XThC.Tn[1].n71 XThC.Tn[1].n70 0.0599512
R22517 XThC.Tn[1].n67 XThC.Tn[1].n66 0.0599512
R22518 XThC.Tn[1].n63 XThC.Tn[1].n62 0.0599512
R22519 XThC.Tn[1].n59 XThC.Tn[1].n58 0.0599512
R22520 XThC.Tn[1].n55 XThC.Tn[1].n54 0.0599512
R22521 XThC.Tn[1].n51 XThC.Tn[1].n50 0.0599512
R22522 XThC.Tn[1].n47 XThC.Tn[1].n46 0.0599512
R22523 XThC.Tn[1].n43 XThC.Tn[1].n42 0.0599512
R22524 XThC.Tn[1].n39 XThC.Tn[1].n38 0.0599512
R22525 XThC.Tn[1].n35 XThC.Tn[1].n34 0.0599512
R22526 XThC.Tn[1].n31 XThC.Tn[1].n30 0.0599512
R22527 XThC.Tn[1].n27 XThC.Tn[1].n26 0.0599512
R22528 XThC.Tn[1].n23 XThC.Tn[1].n22 0.0599512
R22529 XThC.Tn[1].n19 XThC.Tn[1].n18 0.0599512
R22530 XThC.Tn[1].n15 XThC.Tn[1].n14 0.0599512
R22531 XThC.Tn[1].n12 XThC.Tn[1].n11 0.0599512
R22532 XThC.Tn[1].n70 XThC.Tn[1] 0.0469286
R22533 XThC.Tn[1].n66 XThC.Tn[1] 0.0469286
R22534 XThC.Tn[1].n62 XThC.Tn[1] 0.0469286
R22535 XThC.Tn[1].n58 XThC.Tn[1] 0.0469286
R22536 XThC.Tn[1].n54 XThC.Tn[1] 0.0469286
R22537 XThC.Tn[1].n50 XThC.Tn[1] 0.0469286
R22538 XThC.Tn[1].n46 XThC.Tn[1] 0.0469286
R22539 XThC.Tn[1].n42 XThC.Tn[1] 0.0469286
R22540 XThC.Tn[1].n38 XThC.Tn[1] 0.0469286
R22541 XThC.Tn[1].n34 XThC.Tn[1] 0.0469286
R22542 XThC.Tn[1].n30 XThC.Tn[1] 0.0469286
R22543 XThC.Tn[1].n26 XThC.Tn[1] 0.0469286
R22544 XThC.Tn[1].n22 XThC.Tn[1] 0.0469286
R22545 XThC.Tn[1].n18 XThC.Tn[1] 0.0469286
R22546 XThC.Tn[1].n14 XThC.Tn[1] 0.0469286
R22547 XThC.Tn[1].n11 XThC.Tn[1] 0.0469286
R22548 XThC.Tn[1].n70 XThC.Tn[1] 0.0401341
R22549 XThC.Tn[1].n66 XThC.Tn[1] 0.0401341
R22550 XThC.Tn[1].n62 XThC.Tn[1] 0.0401341
R22551 XThC.Tn[1].n58 XThC.Tn[1] 0.0401341
R22552 XThC.Tn[1].n54 XThC.Tn[1] 0.0401341
R22553 XThC.Tn[1].n50 XThC.Tn[1] 0.0401341
R22554 XThC.Tn[1].n46 XThC.Tn[1] 0.0401341
R22555 XThC.Tn[1].n42 XThC.Tn[1] 0.0401341
R22556 XThC.Tn[1].n38 XThC.Tn[1] 0.0401341
R22557 XThC.Tn[1].n34 XThC.Tn[1] 0.0401341
R22558 XThC.Tn[1].n30 XThC.Tn[1] 0.0401341
R22559 XThC.Tn[1].n26 XThC.Tn[1] 0.0401341
R22560 XThC.Tn[1].n22 XThC.Tn[1] 0.0401341
R22561 XThC.Tn[1].n18 XThC.Tn[1] 0.0401341
R22562 XThC.Tn[1].n14 XThC.Tn[1] 0.0401341
R22563 XThC.Tn[1].n11 XThC.Tn[1] 0.0401341
R22564 XThC.Tn[3].n2 XThC.Tn[3].n1 332.334
R22565 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R22566 XThC.Tn[3].n71 XThC.Tn[3].n69 161.365
R22567 XThC.Tn[3].n67 XThC.Tn[3].n65 161.365
R22568 XThC.Tn[3].n63 XThC.Tn[3].n61 161.365
R22569 XThC.Tn[3].n59 XThC.Tn[3].n57 161.365
R22570 XThC.Tn[3].n55 XThC.Tn[3].n53 161.365
R22571 XThC.Tn[3].n51 XThC.Tn[3].n49 161.365
R22572 XThC.Tn[3].n47 XThC.Tn[3].n45 161.365
R22573 XThC.Tn[3].n43 XThC.Tn[3].n41 161.365
R22574 XThC.Tn[3].n39 XThC.Tn[3].n37 161.365
R22575 XThC.Tn[3].n35 XThC.Tn[3].n33 161.365
R22576 XThC.Tn[3].n31 XThC.Tn[3].n29 161.365
R22577 XThC.Tn[3].n27 XThC.Tn[3].n25 161.365
R22578 XThC.Tn[3].n23 XThC.Tn[3].n21 161.365
R22579 XThC.Tn[3].n19 XThC.Tn[3].n17 161.365
R22580 XThC.Tn[3].n15 XThC.Tn[3].n13 161.365
R22581 XThC.Tn[3].n12 XThC.Tn[3].n10 161.365
R22582 XThC.Tn[3].n69 XThC.Tn[3].t16 161.202
R22583 XThC.Tn[3].n65 XThC.Tn[3].t38 161.202
R22584 XThC.Tn[3].n61 XThC.Tn[3].t25 161.202
R22585 XThC.Tn[3].n57 XThC.Tn[3].t22 161.202
R22586 XThC.Tn[3].n53 XThC.Tn[3].t14 161.202
R22587 XThC.Tn[3].n49 XThC.Tn[3].t33 161.202
R22588 XThC.Tn[3].n45 XThC.Tn[3].t32 161.202
R22589 XThC.Tn[3].n41 XThC.Tn[3].t13 161.202
R22590 XThC.Tn[3].n37 XThC.Tn[3].t43 161.202
R22591 XThC.Tn[3].n33 XThC.Tn[3].t34 161.202
R22592 XThC.Tn[3].n29 XThC.Tn[3].t21 161.202
R22593 XThC.Tn[3].n25 XThC.Tn[3].t20 161.202
R22594 XThC.Tn[3].n21 XThC.Tn[3].t31 161.202
R22595 XThC.Tn[3].n17 XThC.Tn[3].t29 161.202
R22596 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R22597 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R22598 XThC.Tn[3].n69 XThC.Tn[3].t19 145.137
R22599 XThC.Tn[3].n65 XThC.Tn[3].t41 145.137
R22600 XThC.Tn[3].n61 XThC.Tn[3].t28 145.137
R22601 XThC.Tn[3].n57 XThC.Tn[3].t26 145.137
R22602 XThC.Tn[3].n53 XThC.Tn[3].t18 145.137
R22603 XThC.Tn[3].n49 XThC.Tn[3].t39 145.137
R22604 XThC.Tn[3].n45 XThC.Tn[3].t37 145.137
R22605 XThC.Tn[3].n41 XThC.Tn[3].t17 145.137
R22606 XThC.Tn[3].n37 XThC.Tn[3].t15 145.137
R22607 XThC.Tn[3].n33 XThC.Tn[3].t40 145.137
R22608 XThC.Tn[3].n29 XThC.Tn[3].t24 145.137
R22609 XThC.Tn[3].n25 XThC.Tn[3].t23 145.137
R22610 XThC.Tn[3].n21 XThC.Tn[3].t36 145.137
R22611 XThC.Tn[3].n17 XThC.Tn[3].t35 145.137
R22612 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R22613 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R22614 XThC.Tn[3].n5 XThC.Tn[3].n3 135.249
R22615 XThC.Tn[3].n5 XThC.Tn[3].n4 98.981
R22616 XThC.Tn[3].n7 XThC.Tn[3].n6 98.981
R22617 XThC.Tn[3].n9 XThC.Tn[3].n8 98.981
R22618 XThC.Tn[3].n7 XThC.Tn[3].n5 36.2672
R22619 XThC.Tn[3].n9 XThC.Tn[3].n7 36.2672
R22620 XThC.Tn[3].n74 XThC.Tn[3].n9 32.6405
R22621 XThC.Tn[3].n0 XThC.Tn[3].t1 26.5955
R22622 XThC.Tn[3].n0 XThC.Tn[3].t0 26.5955
R22623 XThC.Tn[3].n1 XThC.Tn[3].t3 26.5955
R22624 XThC.Tn[3].n1 XThC.Tn[3].t2 26.5955
R22625 XThC.Tn[3].n3 XThC.Tn[3].t11 24.9236
R22626 XThC.Tn[3].n3 XThC.Tn[3].t10 24.9236
R22627 XThC.Tn[3].n4 XThC.Tn[3].t9 24.9236
R22628 XThC.Tn[3].n4 XThC.Tn[3].t8 24.9236
R22629 XThC.Tn[3].n6 XThC.Tn[3].t7 24.9236
R22630 XThC.Tn[3].n6 XThC.Tn[3].t6 24.9236
R22631 XThC.Tn[3].n8 XThC.Tn[3].t5 24.9236
R22632 XThC.Tn[3].n8 XThC.Tn[3].t4 24.9236
R22633 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R22634 XThC.Tn[3] XThC.Tn[3].n12 8.0245
R22635 XThC.Tn[3].n72 XThC.Tn[3].n71 7.9105
R22636 XThC.Tn[3].n68 XThC.Tn[3].n67 7.9105
R22637 XThC.Tn[3].n64 XThC.Tn[3].n63 7.9105
R22638 XThC.Tn[3].n60 XThC.Tn[3].n59 7.9105
R22639 XThC.Tn[3].n56 XThC.Tn[3].n55 7.9105
R22640 XThC.Tn[3].n52 XThC.Tn[3].n51 7.9105
R22641 XThC.Tn[3].n48 XThC.Tn[3].n47 7.9105
R22642 XThC.Tn[3].n44 XThC.Tn[3].n43 7.9105
R22643 XThC.Tn[3].n40 XThC.Tn[3].n39 7.9105
R22644 XThC.Tn[3].n36 XThC.Tn[3].n35 7.9105
R22645 XThC.Tn[3].n32 XThC.Tn[3].n31 7.9105
R22646 XThC.Tn[3].n28 XThC.Tn[3].n27 7.9105
R22647 XThC.Tn[3].n24 XThC.Tn[3].n23 7.9105
R22648 XThC.Tn[3].n20 XThC.Tn[3].n19 7.9105
R22649 XThC.Tn[3].n16 XThC.Tn[3].n15 7.9105
R22650 XThC.Tn[3].n73 XThC.Tn[3] 7.48718
R22651 XThC.Tn[3] XThC.Tn[3].n74 6.7205
R22652 XThC.Tn[3].n74 XThC.Tn[3].n73 5.06464
R22653 XThC.Tn[3].n73 XThC.Tn[3] 1.18175
R22654 XThC.Tn[3].n16 XThC.Tn[3] 0.235138
R22655 XThC.Tn[3].n20 XThC.Tn[3] 0.235138
R22656 XThC.Tn[3].n24 XThC.Tn[3] 0.235138
R22657 XThC.Tn[3].n28 XThC.Tn[3] 0.235138
R22658 XThC.Tn[3].n32 XThC.Tn[3] 0.235138
R22659 XThC.Tn[3].n36 XThC.Tn[3] 0.235138
R22660 XThC.Tn[3].n40 XThC.Tn[3] 0.235138
R22661 XThC.Tn[3].n44 XThC.Tn[3] 0.235138
R22662 XThC.Tn[3].n48 XThC.Tn[3] 0.235138
R22663 XThC.Tn[3].n52 XThC.Tn[3] 0.235138
R22664 XThC.Tn[3].n56 XThC.Tn[3] 0.235138
R22665 XThC.Tn[3].n60 XThC.Tn[3] 0.235138
R22666 XThC.Tn[3].n64 XThC.Tn[3] 0.235138
R22667 XThC.Tn[3].n68 XThC.Tn[3] 0.235138
R22668 XThC.Tn[3].n72 XThC.Tn[3] 0.235138
R22669 XThC.Tn[3] XThC.Tn[3].n16 0.114505
R22670 XThC.Tn[3] XThC.Tn[3].n20 0.114505
R22671 XThC.Tn[3] XThC.Tn[3].n24 0.114505
R22672 XThC.Tn[3] XThC.Tn[3].n28 0.114505
R22673 XThC.Tn[3] XThC.Tn[3].n32 0.114505
R22674 XThC.Tn[3] XThC.Tn[3].n36 0.114505
R22675 XThC.Tn[3] XThC.Tn[3].n40 0.114505
R22676 XThC.Tn[3] XThC.Tn[3].n44 0.114505
R22677 XThC.Tn[3] XThC.Tn[3].n48 0.114505
R22678 XThC.Tn[3] XThC.Tn[3].n52 0.114505
R22679 XThC.Tn[3] XThC.Tn[3].n56 0.114505
R22680 XThC.Tn[3] XThC.Tn[3].n60 0.114505
R22681 XThC.Tn[3] XThC.Tn[3].n64 0.114505
R22682 XThC.Tn[3] XThC.Tn[3].n68 0.114505
R22683 XThC.Tn[3] XThC.Tn[3].n72 0.114505
R22684 XThC.Tn[3].n71 XThC.Tn[3].n70 0.0599512
R22685 XThC.Tn[3].n67 XThC.Tn[3].n66 0.0599512
R22686 XThC.Tn[3].n63 XThC.Tn[3].n62 0.0599512
R22687 XThC.Tn[3].n59 XThC.Tn[3].n58 0.0599512
R22688 XThC.Tn[3].n55 XThC.Tn[3].n54 0.0599512
R22689 XThC.Tn[3].n51 XThC.Tn[3].n50 0.0599512
R22690 XThC.Tn[3].n47 XThC.Tn[3].n46 0.0599512
R22691 XThC.Tn[3].n43 XThC.Tn[3].n42 0.0599512
R22692 XThC.Tn[3].n39 XThC.Tn[3].n38 0.0599512
R22693 XThC.Tn[3].n35 XThC.Tn[3].n34 0.0599512
R22694 XThC.Tn[3].n31 XThC.Tn[3].n30 0.0599512
R22695 XThC.Tn[3].n27 XThC.Tn[3].n26 0.0599512
R22696 XThC.Tn[3].n23 XThC.Tn[3].n22 0.0599512
R22697 XThC.Tn[3].n19 XThC.Tn[3].n18 0.0599512
R22698 XThC.Tn[3].n15 XThC.Tn[3].n14 0.0599512
R22699 XThC.Tn[3].n12 XThC.Tn[3].n11 0.0599512
R22700 XThC.Tn[3].n70 XThC.Tn[3] 0.0469286
R22701 XThC.Tn[3].n66 XThC.Tn[3] 0.0469286
R22702 XThC.Tn[3].n62 XThC.Tn[3] 0.0469286
R22703 XThC.Tn[3].n58 XThC.Tn[3] 0.0469286
R22704 XThC.Tn[3].n54 XThC.Tn[3] 0.0469286
R22705 XThC.Tn[3].n50 XThC.Tn[3] 0.0469286
R22706 XThC.Tn[3].n46 XThC.Tn[3] 0.0469286
R22707 XThC.Tn[3].n42 XThC.Tn[3] 0.0469286
R22708 XThC.Tn[3].n38 XThC.Tn[3] 0.0469286
R22709 XThC.Tn[3].n34 XThC.Tn[3] 0.0469286
R22710 XThC.Tn[3].n30 XThC.Tn[3] 0.0469286
R22711 XThC.Tn[3].n26 XThC.Tn[3] 0.0469286
R22712 XThC.Tn[3].n22 XThC.Tn[3] 0.0469286
R22713 XThC.Tn[3].n18 XThC.Tn[3] 0.0469286
R22714 XThC.Tn[3].n14 XThC.Tn[3] 0.0469286
R22715 XThC.Tn[3].n11 XThC.Tn[3] 0.0469286
R22716 XThC.Tn[3].n70 XThC.Tn[3] 0.0401341
R22717 XThC.Tn[3].n66 XThC.Tn[3] 0.0401341
R22718 XThC.Tn[3].n62 XThC.Tn[3] 0.0401341
R22719 XThC.Tn[3].n58 XThC.Tn[3] 0.0401341
R22720 XThC.Tn[3].n54 XThC.Tn[3] 0.0401341
R22721 XThC.Tn[3].n50 XThC.Tn[3] 0.0401341
R22722 XThC.Tn[3].n46 XThC.Tn[3] 0.0401341
R22723 XThC.Tn[3].n42 XThC.Tn[3] 0.0401341
R22724 XThC.Tn[3].n38 XThC.Tn[3] 0.0401341
R22725 XThC.Tn[3].n34 XThC.Tn[3] 0.0401341
R22726 XThC.Tn[3].n30 XThC.Tn[3] 0.0401341
R22727 XThC.Tn[3].n26 XThC.Tn[3] 0.0401341
R22728 XThC.Tn[3].n22 XThC.Tn[3] 0.0401341
R22729 XThC.Tn[3].n18 XThC.Tn[3] 0.0401341
R22730 XThC.Tn[3].n14 XThC.Tn[3] 0.0401341
R22731 XThC.Tn[3].n11 XThC.Tn[3] 0.0401341
R22732 XThR.Tn[10].n87 XThR.Tn[10].n86 256.103
R22733 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R22734 XThR.Tn[10].n5 XThR.Tn[10].n3 241.847
R22735 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R22736 XThR.Tn[10].n87 XThR.Tn[10].n85 202.095
R22737 XThR.Tn[10].n5 XThR.Tn[10].n4 185
R22738 XThR.Tn[10] XThR.Tn[10].n78 161.363
R22739 XThR.Tn[10] XThR.Tn[10].n73 161.363
R22740 XThR.Tn[10] XThR.Tn[10].n68 161.363
R22741 XThR.Tn[10] XThR.Tn[10].n63 161.363
R22742 XThR.Tn[10] XThR.Tn[10].n58 161.363
R22743 XThR.Tn[10] XThR.Tn[10].n53 161.363
R22744 XThR.Tn[10] XThR.Tn[10].n48 161.363
R22745 XThR.Tn[10] XThR.Tn[10].n43 161.363
R22746 XThR.Tn[10] XThR.Tn[10].n38 161.363
R22747 XThR.Tn[10] XThR.Tn[10].n33 161.363
R22748 XThR.Tn[10] XThR.Tn[10].n28 161.363
R22749 XThR.Tn[10] XThR.Tn[10].n23 161.363
R22750 XThR.Tn[10] XThR.Tn[10].n18 161.363
R22751 XThR.Tn[10] XThR.Tn[10].n13 161.363
R22752 XThR.Tn[10] XThR.Tn[10].n8 161.363
R22753 XThR.Tn[10] XThR.Tn[10].n6 161.363
R22754 XThR.Tn[10].n80 XThR.Tn[10].n79 161.3
R22755 XThR.Tn[10].n75 XThR.Tn[10].n74 161.3
R22756 XThR.Tn[10].n70 XThR.Tn[10].n69 161.3
R22757 XThR.Tn[10].n65 XThR.Tn[10].n64 161.3
R22758 XThR.Tn[10].n60 XThR.Tn[10].n59 161.3
R22759 XThR.Tn[10].n55 XThR.Tn[10].n54 161.3
R22760 XThR.Tn[10].n50 XThR.Tn[10].n49 161.3
R22761 XThR.Tn[10].n45 XThR.Tn[10].n44 161.3
R22762 XThR.Tn[10].n40 XThR.Tn[10].n39 161.3
R22763 XThR.Tn[10].n35 XThR.Tn[10].n34 161.3
R22764 XThR.Tn[10].n30 XThR.Tn[10].n29 161.3
R22765 XThR.Tn[10].n25 XThR.Tn[10].n24 161.3
R22766 XThR.Tn[10].n20 XThR.Tn[10].n19 161.3
R22767 XThR.Tn[10].n15 XThR.Tn[10].n14 161.3
R22768 XThR.Tn[10].n10 XThR.Tn[10].n9 161.3
R22769 XThR.Tn[10].n78 XThR.Tn[10].t37 161.106
R22770 XThR.Tn[10].n73 XThR.Tn[10].t45 161.106
R22771 XThR.Tn[10].n68 XThR.Tn[10].t27 161.106
R22772 XThR.Tn[10].n63 XThR.Tn[10].t72 161.106
R22773 XThR.Tn[10].n58 XThR.Tn[10].t35 161.106
R22774 XThR.Tn[10].n53 XThR.Tn[10].t61 161.106
R22775 XThR.Tn[10].n48 XThR.Tn[10].t43 161.106
R22776 XThR.Tn[10].n43 XThR.Tn[10].t24 161.106
R22777 XThR.Tn[10].n38 XThR.Tn[10].t69 161.106
R22778 XThR.Tn[10].n33 XThR.Tn[10].t15 161.106
R22779 XThR.Tn[10].n28 XThR.Tn[10].t59 161.106
R22780 XThR.Tn[10].n23 XThR.Tn[10].t26 161.106
R22781 XThR.Tn[10].n18 XThR.Tn[10].t58 161.106
R22782 XThR.Tn[10].n13 XThR.Tn[10].t41 161.106
R22783 XThR.Tn[10].n8 XThR.Tn[10].t63 161.106
R22784 XThR.Tn[10].n6 XThR.Tn[10].t47 161.106
R22785 XThR.Tn[10].n79 XThR.Tn[10].t34 159.978
R22786 XThR.Tn[10].n74 XThR.Tn[10].t39 159.978
R22787 XThR.Tn[10].n69 XThR.Tn[10].t22 159.978
R22788 XThR.Tn[10].n64 XThR.Tn[10].t68 159.978
R22789 XThR.Tn[10].n59 XThR.Tn[10].t32 159.978
R22790 XThR.Tn[10].n54 XThR.Tn[10].t57 159.978
R22791 XThR.Tn[10].n49 XThR.Tn[10].t38 159.978
R22792 XThR.Tn[10].n44 XThR.Tn[10].t20 159.978
R22793 XThR.Tn[10].n39 XThR.Tn[10].t66 159.978
R22794 XThR.Tn[10].n34 XThR.Tn[10].t12 159.978
R22795 XThR.Tn[10].n29 XThR.Tn[10].t56 159.978
R22796 XThR.Tn[10].n24 XThR.Tn[10].t21 159.978
R22797 XThR.Tn[10].n19 XThR.Tn[10].t55 159.978
R22798 XThR.Tn[10].n14 XThR.Tn[10].t36 159.978
R22799 XThR.Tn[10].n9 XThR.Tn[10].t60 159.978
R22800 XThR.Tn[10].n78 XThR.Tn[10].t29 145.038
R22801 XThR.Tn[10].n73 XThR.Tn[10].t49 145.038
R22802 XThR.Tn[10].n68 XThR.Tn[10].t31 145.038
R22803 XThR.Tn[10].n63 XThR.Tn[10].t16 145.038
R22804 XThR.Tn[10].n58 XThR.Tn[10].t46 145.038
R22805 XThR.Tn[10].n53 XThR.Tn[10].t28 145.038
R22806 XThR.Tn[10].n48 XThR.Tn[10].t33 145.038
R22807 XThR.Tn[10].n43 XThR.Tn[10].t17 145.038
R22808 XThR.Tn[10].n38 XThR.Tn[10].t14 145.038
R22809 XThR.Tn[10].n33 XThR.Tn[10].t44 145.038
R22810 XThR.Tn[10].n28 XThR.Tn[10].t67 145.038
R22811 XThR.Tn[10].n23 XThR.Tn[10].t30 145.038
R22812 XThR.Tn[10].n18 XThR.Tn[10].t65 145.038
R22813 XThR.Tn[10].n13 XThR.Tn[10].t48 145.038
R22814 XThR.Tn[10].n8 XThR.Tn[10].t13 145.038
R22815 XThR.Tn[10].n6 XThR.Tn[10].t54 145.038
R22816 XThR.Tn[10].n79 XThR.Tn[10].t64 143.911
R22817 XThR.Tn[10].n74 XThR.Tn[10].t25 143.911
R22818 XThR.Tn[10].n69 XThR.Tn[10].t71 143.911
R22819 XThR.Tn[10].n64 XThR.Tn[10].t52 143.911
R22820 XThR.Tn[10].n59 XThR.Tn[10].t19 143.911
R22821 XThR.Tn[10].n54 XThR.Tn[10].t62 143.911
R22822 XThR.Tn[10].n49 XThR.Tn[10].t73 143.911
R22823 XThR.Tn[10].n44 XThR.Tn[10].t53 143.911
R22824 XThR.Tn[10].n39 XThR.Tn[10].t51 143.911
R22825 XThR.Tn[10].n34 XThR.Tn[10].t18 143.911
R22826 XThR.Tn[10].n29 XThR.Tn[10].t42 143.911
R22827 XThR.Tn[10].n24 XThR.Tn[10].t70 143.911
R22828 XThR.Tn[10].n19 XThR.Tn[10].t40 143.911
R22829 XThR.Tn[10].n14 XThR.Tn[10].t23 143.911
R22830 XThR.Tn[10].n9 XThR.Tn[10].t50 143.911
R22831 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R22832 XThR.Tn[10].n85 XThR.Tn[10].t5 26.5955
R22833 XThR.Tn[10].n85 XThR.Tn[10].t3 26.5955
R22834 XThR.Tn[10].n0 XThR.Tn[10].t10 26.5955
R22835 XThR.Tn[10].n0 XThR.Tn[10].t8 26.5955
R22836 XThR.Tn[10].n1 XThR.Tn[10].t11 26.5955
R22837 XThR.Tn[10].n1 XThR.Tn[10].t9 26.5955
R22838 XThR.Tn[10].n86 XThR.Tn[10].t0 26.5955
R22839 XThR.Tn[10].n86 XThR.Tn[10].t6 26.5955
R22840 XThR.Tn[10].n4 XThR.Tn[10].t2 24.9236
R22841 XThR.Tn[10].n4 XThR.Tn[10].t7 24.9236
R22842 XThR.Tn[10].n3 XThR.Tn[10].t1 24.9236
R22843 XThR.Tn[10].n3 XThR.Tn[10].t4 24.9236
R22844 XThR.Tn[10] XThR.Tn[10].n5 18.8943
R22845 XThR.Tn[10].n88 XThR.Tn[10].n87 13.5534
R22846 XThR.Tn[10].n84 XThR.Tn[10] 7.84567
R22847 XThR.Tn[10].n84 XThR.Tn[10] 6.34069
R22848 XThR.Tn[10] XThR.Tn[10].n7 5.34038
R22849 XThR.Tn[10].n12 XThR.Tn[10].n11 4.5005
R22850 XThR.Tn[10].n17 XThR.Tn[10].n16 4.5005
R22851 XThR.Tn[10].n22 XThR.Tn[10].n21 4.5005
R22852 XThR.Tn[10].n27 XThR.Tn[10].n26 4.5005
R22853 XThR.Tn[10].n32 XThR.Tn[10].n31 4.5005
R22854 XThR.Tn[10].n37 XThR.Tn[10].n36 4.5005
R22855 XThR.Tn[10].n42 XThR.Tn[10].n41 4.5005
R22856 XThR.Tn[10].n47 XThR.Tn[10].n46 4.5005
R22857 XThR.Tn[10].n52 XThR.Tn[10].n51 4.5005
R22858 XThR.Tn[10].n57 XThR.Tn[10].n56 4.5005
R22859 XThR.Tn[10].n62 XThR.Tn[10].n61 4.5005
R22860 XThR.Tn[10].n67 XThR.Tn[10].n66 4.5005
R22861 XThR.Tn[10].n72 XThR.Tn[10].n71 4.5005
R22862 XThR.Tn[10].n77 XThR.Tn[10].n76 4.5005
R22863 XThR.Tn[10].n82 XThR.Tn[10].n81 4.5005
R22864 XThR.Tn[10].n83 XThR.Tn[10] 3.70586
R22865 XThR.Tn[10].n12 XThR.Tn[10] 2.52282
R22866 XThR.Tn[10].n17 XThR.Tn[10] 2.52282
R22867 XThR.Tn[10].n22 XThR.Tn[10] 2.52282
R22868 XThR.Tn[10].n27 XThR.Tn[10] 2.52282
R22869 XThR.Tn[10].n32 XThR.Tn[10] 2.52282
R22870 XThR.Tn[10].n37 XThR.Tn[10] 2.52282
R22871 XThR.Tn[10].n42 XThR.Tn[10] 2.52282
R22872 XThR.Tn[10].n47 XThR.Tn[10] 2.52282
R22873 XThR.Tn[10].n52 XThR.Tn[10] 2.52282
R22874 XThR.Tn[10].n57 XThR.Tn[10] 2.52282
R22875 XThR.Tn[10].n62 XThR.Tn[10] 2.52282
R22876 XThR.Tn[10].n67 XThR.Tn[10] 2.52282
R22877 XThR.Tn[10].n72 XThR.Tn[10] 2.52282
R22878 XThR.Tn[10].n77 XThR.Tn[10] 2.52282
R22879 XThR.Tn[10].n82 XThR.Tn[10] 2.52282
R22880 XThR.Tn[10] XThR.Tn[10].n84 1.79489
R22881 XThR.Tn[10] XThR.Tn[10].n88 1.50638
R22882 XThR.Tn[10].n88 XThR.Tn[10] 1.19676
R22883 XThR.Tn[10].n80 XThR.Tn[10] 1.08677
R22884 XThR.Tn[10].n75 XThR.Tn[10] 1.08677
R22885 XThR.Tn[10].n70 XThR.Tn[10] 1.08677
R22886 XThR.Tn[10].n65 XThR.Tn[10] 1.08677
R22887 XThR.Tn[10].n60 XThR.Tn[10] 1.08677
R22888 XThR.Tn[10].n55 XThR.Tn[10] 1.08677
R22889 XThR.Tn[10].n50 XThR.Tn[10] 1.08677
R22890 XThR.Tn[10].n45 XThR.Tn[10] 1.08677
R22891 XThR.Tn[10].n40 XThR.Tn[10] 1.08677
R22892 XThR.Tn[10].n35 XThR.Tn[10] 1.08677
R22893 XThR.Tn[10].n30 XThR.Tn[10] 1.08677
R22894 XThR.Tn[10].n25 XThR.Tn[10] 1.08677
R22895 XThR.Tn[10].n20 XThR.Tn[10] 1.08677
R22896 XThR.Tn[10].n15 XThR.Tn[10] 1.08677
R22897 XThR.Tn[10].n10 XThR.Tn[10] 1.08677
R22898 XThR.Tn[10] XThR.Tn[10].n12 0.839786
R22899 XThR.Tn[10] XThR.Tn[10].n17 0.839786
R22900 XThR.Tn[10] XThR.Tn[10].n22 0.839786
R22901 XThR.Tn[10] XThR.Tn[10].n27 0.839786
R22902 XThR.Tn[10] XThR.Tn[10].n32 0.839786
R22903 XThR.Tn[10] XThR.Tn[10].n37 0.839786
R22904 XThR.Tn[10] XThR.Tn[10].n42 0.839786
R22905 XThR.Tn[10] XThR.Tn[10].n47 0.839786
R22906 XThR.Tn[10] XThR.Tn[10].n52 0.839786
R22907 XThR.Tn[10] XThR.Tn[10].n57 0.839786
R22908 XThR.Tn[10] XThR.Tn[10].n62 0.839786
R22909 XThR.Tn[10] XThR.Tn[10].n67 0.839786
R22910 XThR.Tn[10] XThR.Tn[10].n72 0.839786
R22911 XThR.Tn[10] XThR.Tn[10].n77 0.839786
R22912 XThR.Tn[10] XThR.Tn[10].n82 0.839786
R22913 XThR.Tn[10].n7 XThR.Tn[10] 0.499542
R22914 XThR.Tn[10].n81 XThR.Tn[10] 0.063
R22915 XThR.Tn[10].n76 XThR.Tn[10] 0.063
R22916 XThR.Tn[10].n71 XThR.Tn[10] 0.063
R22917 XThR.Tn[10].n66 XThR.Tn[10] 0.063
R22918 XThR.Tn[10].n61 XThR.Tn[10] 0.063
R22919 XThR.Tn[10].n56 XThR.Tn[10] 0.063
R22920 XThR.Tn[10].n51 XThR.Tn[10] 0.063
R22921 XThR.Tn[10].n46 XThR.Tn[10] 0.063
R22922 XThR.Tn[10].n41 XThR.Tn[10] 0.063
R22923 XThR.Tn[10].n36 XThR.Tn[10] 0.063
R22924 XThR.Tn[10].n31 XThR.Tn[10] 0.063
R22925 XThR.Tn[10].n26 XThR.Tn[10] 0.063
R22926 XThR.Tn[10].n21 XThR.Tn[10] 0.063
R22927 XThR.Tn[10].n16 XThR.Tn[10] 0.063
R22928 XThR.Tn[10].n11 XThR.Tn[10] 0.063
R22929 XThR.Tn[10].n83 XThR.Tn[10] 0.0540714
R22930 XThR.Tn[10] XThR.Tn[10].n83 0.038
R22931 XThR.Tn[10].n7 XThR.Tn[10] 0.0143889
R22932 XThR.Tn[10].n81 XThR.Tn[10].n80 0.00771154
R22933 XThR.Tn[10].n76 XThR.Tn[10].n75 0.00771154
R22934 XThR.Tn[10].n71 XThR.Tn[10].n70 0.00771154
R22935 XThR.Tn[10].n66 XThR.Tn[10].n65 0.00771154
R22936 XThR.Tn[10].n61 XThR.Tn[10].n60 0.00771154
R22937 XThR.Tn[10].n56 XThR.Tn[10].n55 0.00771154
R22938 XThR.Tn[10].n51 XThR.Tn[10].n50 0.00771154
R22939 XThR.Tn[10].n46 XThR.Tn[10].n45 0.00771154
R22940 XThR.Tn[10].n41 XThR.Tn[10].n40 0.00771154
R22941 XThR.Tn[10].n36 XThR.Tn[10].n35 0.00771154
R22942 XThR.Tn[10].n31 XThR.Tn[10].n30 0.00771154
R22943 XThR.Tn[10].n26 XThR.Tn[10].n25 0.00771154
R22944 XThR.Tn[10].n21 XThR.Tn[10].n20 0.00771154
R22945 XThR.Tn[10].n16 XThR.Tn[10].n15 0.00771154
R22946 XThR.Tn[10].n11 XThR.Tn[10].n10 0.00771154
R22947 XThC.Tn[14].n5 XThC.Tn[14].n4 256.104
R22948 XThC.Tn[14].n8 XThC.Tn[14].n6 243.68
R22949 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22950 XThC.Tn[14].n8 XThC.Tn[14].n7 205.28
R22951 XThC.Tn[14].n5 XThC.Tn[14].n3 202.095
R22952 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22953 XThC.Tn[14].n71 XThC.Tn[14].n69 161.365
R22954 XThC.Tn[14].n67 XThC.Tn[14].n65 161.365
R22955 XThC.Tn[14].n63 XThC.Tn[14].n61 161.365
R22956 XThC.Tn[14].n59 XThC.Tn[14].n57 161.365
R22957 XThC.Tn[14].n55 XThC.Tn[14].n53 161.365
R22958 XThC.Tn[14].n51 XThC.Tn[14].n49 161.365
R22959 XThC.Tn[14].n47 XThC.Tn[14].n45 161.365
R22960 XThC.Tn[14].n43 XThC.Tn[14].n41 161.365
R22961 XThC.Tn[14].n39 XThC.Tn[14].n37 161.365
R22962 XThC.Tn[14].n35 XThC.Tn[14].n33 161.365
R22963 XThC.Tn[14].n31 XThC.Tn[14].n29 161.365
R22964 XThC.Tn[14].n27 XThC.Tn[14].n25 161.365
R22965 XThC.Tn[14].n23 XThC.Tn[14].n21 161.365
R22966 XThC.Tn[14].n19 XThC.Tn[14].n17 161.365
R22967 XThC.Tn[14].n15 XThC.Tn[14].n13 161.365
R22968 XThC.Tn[14].n12 XThC.Tn[14].n10 161.365
R22969 XThC.Tn[14].n69 XThC.Tn[14].t12 161.202
R22970 XThC.Tn[14].n65 XThC.Tn[14].t33 161.202
R22971 XThC.Tn[14].n61 XThC.Tn[14].t21 161.202
R22972 XThC.Tn[14].n57 XThC.Tn[14].t19 161.202
R22973 XThC.Tn[14].n53 XThC.Tn[14].t42 161.202
R22974 XThC.Tn[14].n49 XThC.Tn[14].t30 161.202
R22975 XThC.Tn[14].n45 XThC.Tn[14].t27 161.202
R22976 XThC.Tn[14].n41 XThC.Tn[14].t41 161.202
R22977 XThC.Tn[14].n37 XThC.Tn[14].t39 161.202
R22978 XThC.Tn[14].n33 XThC.Tn[14].t31 161.202
R22979 XThC.Tn[14].n29 XThC.Tn[14].t17 161.202
R22980 XThC.Tn[14].n25 XThC.Tn[14].t14 161.202
R22981 XThC.Tn[14].n21 XThC.Tn[14].t26 161.202
R22982 XThC.Tn[14].n17 XThC.Tn[14].t25 161.202
R22983 XThC.Tn[14].n13 XThC.Tn[14].t22 161.202
R22984 XThC.Tn[14].n10 XThC.Tn[14].t38 161.202
R22985 XThC.Tn[14].n69 XThC.Tn[14].t18 145.137
R22986 XThC.Tn[14].n65 XThC.Tn[14].t40 145.137
R22987 XThC.Tn[14].n61 XThC.Tn[14].t28 145.137
R22988 XThC.Tn[14].n57 XThC.Tn[14].t24 145.137
R22989 XThC.Tn[14].n53 XThC.Tn[14].t16 145.137
R22990 XThC.Tn[14].n49 XThC.Tn[14].t36 145.137
R22991 XThC.Tn[14].n45 XThC.Tn[14].t35 145.137
R22992 XThC.Tn[14].n41 XThC.Tn[14].t15 145.137
R22993 XThC.Tn[14].n37 XThC.Tn[14].t13 145.137
R22994 XThC.Tn[14].n33 XThC.Tn[14].t37 145.137
R22995 XThC.Tn[14].n29 XThC.Tn[14].t23 145.137
R22996 XThC.Tn[14].n25 XThC.Tn[14].t20 145.137
R22997 XThC.Tn[14].n21 XThC.Tn[14].t34 145.137
R22998 XThC.Tn[14].n17 XThC.Tn[14].t32 145.137
R22999 XThC.Tn[14].n13 XThC.Tn[14].t29 145.137
R23000 XThC.Tn[14].n10 XThC.Tn[14].t43 145.137
R23001 XThC.Tn[14].n3 XThC.Tn[14].t4 26.5955
R23002 XThC.Tn[14].n3 XThC.Tn[14].t5 26.5955
R23003 XThC.Tn[14].n4 XThC.Tn[14].t7 26.5955
R23004 XThC.Tn[14].n4 XThC.Tn[14].t6 26.5955
R23005 XThC.Tn[14].n6 XThC.Tn[14].t11 26.5955
R23006 XThC.Tn[14].n6 XThC.Tn[14].t10 26.5955
R23007 XThC.Tn[14].n7 XThC.Tn[14].t9 26.5955
R23008 XThC.Tn[14].n7 XThC.Tn[14].t8 26.5955
R23009 XThC.Tn[14].n0 XThC.Tn[14].t0 24.9236
R23010 XThC.Tn[14].n0 XThC.Tn[14].t2 24.9236
R23011 XThC.Tn[14].n1 XThC.Tn[14].t1 24.9236
R23012 XThC.Tn[14].n1 XThC.Tn[14].t3 24.9236
R23013 XThC.Tn[14] XThC.Tn[14].n8 22.9652
R23014 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R23015 XThC.Tn[14].n9 XThC.Tn[14].n5 13.9299
R23016 XThC.Tn[14].n9 XThC.Tn[14] 13.9299
R23017 XThC.Tn[14] XThC.Tn[14].n12 8.0245
R23018 XThC.Tn[14].n72 XThC.Tn[14].n71 7.9105
R23019 XThC.Tn[14].n68 XThC.Tn[14].n67 7.9105
R23020 XThC.Tn[14].n64 XThC.Tn[14].n63 7.9105
R23021 XThC.Tn[14].n60 XThC.Tn[14].n59 7.9105
R23022 XThC.Tn[14].n56 XThC.Tn[14].n55 7.9105
R23023 XThC.Tn[14].n52 XThC.Tn[14].n51 7.9105
R23024 XThC.Tn[14].n48 XThC.Tn[14].n47 7.9105
R23025 XThC.Tn[14].n44 XThC.Tn[14].n43 7.9105
R23026 XThC.Tn[14].n40 XThC.Tn[14].n39 7.9105
R23027 XThC.Tn[14].n36 XThC.Tn[14].n35 7.9105
R23028 XThC.Tn[14].n32 XThC.Tn[14].n31 7.9105
R23029 XThC.Tn[14].n28 XThC.Tn[14].n27 7.9105
R23030 XThC.Tn[14].n24 XThC.Tn[14].n23 7.9105
R23031 XThC.Tn[14].n20 XThC.Tn[14].n19 7.9105
R23032 XThC.Tn[14].n16 XThC.Tn[14].n15 7.9105
R23033 XThC.Tn[14].n74 XThC.Tn[14].n73 7.51947
R23034 XThC.Tn[14].n73 XThC.Tn[14] 5.85107
R23035 XThC.Tn[14].n74 XThC.Tn[14].n9 2.99115
R23036 XThC.Tn[14].n9 XThC.Tn[14] 2.87153
R23037 XThC.Tn[14] XThC.Tn[14].n74 2.2734
R23038 XThC.Tn[14].n73 XThC.Tn[14] 1.06164
R23039 XThC.Tn[14].n16 XThC.Tn[14] 0.235138
R23040 XThC.Tn[14].n20 XThC.Tn[14] 0.235138
R23041 XThC.Tn[14].n24 XThC.Tn[14] 0.235138
R23042 XThC.Tn[14].n28 XThC.Tn[14] 0.235138
R23043 XThC.Tn[14].n32 XThC.Tn[14] 0.235138
R23044 XThC.Tn[14].n36 XThC.Tn[14] 0.235138
R23045 XThC.Tn[14].n40 XThC.Tn[14] 0.235138
R23046 XThC.Tn[14].n44 XThC.Tn[14] 0.235138
R23047 XThC.Tn[14].n48 XThC.Tn[14] 0.235138
R23048 XThC.Tn[14].n52 XThC.Tn[14] 0.235138
R23049 XThC.Tn[14].n56 XThC.Tn[14] 0.235138
R23050 XThC.Tn[14].n60 XThC.Tn[14] 0.235138
R23051 XThC.Tn[14].n64 XThC.Tn[14] 0.235138
R23052 XThC.Tn[14].n68 XThC.Tn[14] 0.235138
R23053 XThC.Tn[14].n72 XThC.Tn[14] 0.235138
R23054 XThC.Tn[14] XThC.Tn[14].n16 0.114505
R23055 XThC.Tn[14] XThC.Tn[14].n20 0.114505
R23056 XThC.Tn[14] XThC.Tn[14].n24 0.114505
R23057 XThC.Tn[14] XThC.Tn[14].n28 0.114505
R23058 XThC.Tn[14] XThC.Tn[14].n32 0.114505
R23059 XThC.Tn[14] XThC.Tn[14].n36 0.114505
R23060 XThC.Tn[14] XThC.Tn[14].n40 0.114505
R23061 XThC.Tn[14] XThC.Tn[14].n44 0.114505
R23062 XThC.Tn[14] XThC.Tn[14].n48 0.114505
R23063 XThC.Tn[14] XThC.Tn[14].n52 0.114505
R23064 XThC.Tn[14] XThC.Tn[14].n56 0.114505
R23065 XThC.Tn[14] XThC.Tn[14].n60 0.114505
R23066 XThC.Tn[14] XThC.Tn[14].n64 0.114505
R23067 XThC.Tn[14] XThC.Tn[14].n68 0.114505
R23068 XThC.Tn[14] XThC.Tn[14].n72 0.114505
R23069 XThC.Tn[14].n71 XThC.Tn[14].n70 0.0599512
R23070 XThC.Tn[14].n67 XThC.Tn[14].n66 0.0599512
R23071 XThC.Tn[14].n63 XThC.Tn[14].n62 0.0599512
R23072 XThC.Tn[14].n59 XThC.Tn[14].n58 0.0599512
R23073 XThC.Tn[14].n55 XThC.Tn[14].n54 0.0599512
R23074 XThC.Tn[14].n51 XThC.Tn[14].n50 0.0599512
R23075 XThC.Tn[14].n47 XThC.Tn[14].n46 0.0599512
R23076 XThC.Tn[14].n43 XThC.Tn[14].n42 0.0599512
R23077 XThC.Tn[14].n39 XThC.Tn[14].n38 0.0599512
R23078 XThC.Tn[14].n35 XThC.Tn[14].n34 0.0599512
R23079 XThC.Tn[14].n31 XThC.Tn[14].n30 0.0599512
R23080 XThC.Tn[14].n27 XThC.Tn[14].n26 0.0599512
R23081 XThC.Tn[14].n23 XThC.Tn[14].n22 0.0599512
R23082 XThC.Tn[14].n19 XThC.Tn[14].n18 0.0599512
R23083 XThC.Tn[14].n15 XThC.Tn[14].n14 0.0599512
R23084 XThC.Tn[14].n12 XThC.Tn[14].n11 0.0599512
R23085 XThC.Tn[14].n70 XThC.Tn[14] 0.0469286
R23086 XThC.Tn[14].n66 XThC.Tn[14] 0.0469286
R23087 XThC.Tn[14].n62 XThC.Tn[14] 0.0469286
R23088 XThC.Tn[14].n58 XThC.Tn[14] 0.0469286
R23089 XThC.Tn[14].n54 XThC.Tn[14] 0.0469286
R23090 XThC.Tn[14].n50 XThC.Tn[14] 0.0469286
R23091 XThC.Tn[14].n46 XThC.Tn[14] 0.0469286
R23092 XThC.Tn[14].n42 XThC.Tn[14] 0.0469286
R23093 XThC.Tn[14].n38 XThC.Tn[14] 0.0469286
R23094 XThC.Tn[14].n34 XThC.Tn[14] 0.0469286
R23095 XThC.Tn[14].n30 XThC.Tn[14] 0.0469286
R23096 XThC.Tn[14].n26 XThC.Tn[14] 0.0469286
R23097 XThC.Tn[14].n22 XThC.Tn[14] 0.0469286
R23098 XThC.Tn[14].n18 XThC.Tn[14] 0.0469286
R23099 XThC.Tn[14].n14 XThC.Tn[14] 0.0469286
R23100 XThC.Tn[14].n11 XThC.Tn[14] 0.0469286
R23101 XThC.Tn[14].n70 XThC.Tn[14] 0.0401341
R23102 XThC.Tn[14].n66 XThC.Tn[14] 0.0401341
R23103 XThC.Tn[14].n62 XThC.Tn[14] 0.0401341
R23104 XThC.Tn[14].n58 XThC.Tn[14] 0.0401341
R23105 XThC.Tn[14].n54 XThC.Tn[14] 0.0401341
R23106 XThC.Tn[14].n50 XThC.Tn[14] 0.0401341
R23107 XThC.Tn[14].n46 XThC.Tn[14] 0.0401341
R23108 XThC.Tn[14].n42 XThC.Tn[14] 0.0401341
R23109 XThC.Tn[14].n38 XThC.Tn[14] 0.0401341
R23110 XThC.Tn[14].n34 XThC.Tn[14] 0.0401341
R23111 XThC.Tn[14].n30 XThC.Tn[14] 0.0401341
R23112 XThC.Tn[14].n26 XThC.Tn[14] 0.0401341
R23113 XThC.Tn[14].n22 XThC.Tn[14] 0.0401341
R23114 XThC.Tn[14].n18 XThC.Tn[14] 0.0401341
R23115 XThC.Tn[14].n14 XThC.Tn[14] 0.0401341
R23116 XThC.Tn[14].n11 XThC.Tn[14] 0.0401341
R23117 XThC.TB1.n6 XThC.TB1.t11 212.081
R23118 XThC.TB1.n5 XThC.TB1.t8 212.081
R23119 XThC.TB1.n11 XThC.TB1.t6 212.081
R23120 XThC.TB1.n3 XThC.TB1.t17 212.081
R23121 XThC.TB1.n15 XThC.TB1.t10 212.081
R23122 XThC.TB1.n16 XThC.TB1.t14 212.081
R23123 XThC.TB1.n18 XThC.TB1.t7 212.081
R23124 XThC.TB1.n14 XThC.TB1.t18 212.081
R23125 XThC.TB1.n22 XThC.TB1.n2 201.288
R23126 XThC.TB1.n8 XThC.TB1.n7 173.761
R23127 XThC.TB1.n17 XThC.TB1 158.656
R23128 XThC.TB1.n10 XThC.TB1.n9 152
R23129 XThC.TB1.n8 XThC.TB1.n4 152
R23130 XThC.TB1.n13 XThC.TB1.n12 152
R23131 XThC.TB1.n20 XThC.TB1.n19 152
R23132 XThC.TB1.n6 XThC.TB1.t16 139.78
R23133 XThC.TB1.n5 XThC.TB1.t13 139.78
R23134 XThC.TB1.n11 XThC.TB1.t12 139.78
R23135 XThC.TB1.n3 XThC.TB1.t5 139.78
R23136 XThC.TB1.n15 XThC.TB1.t4 139.78
R23137 XThC.TB1.n16 XThC.TB1.t3 139.78
R23138 XThC.TB1.n18 XThC.TB1.t15 139.78
R23139 XThC.TB1.n14 XThC.TB1.t9 139.78
R23140 XThC.TB1.n0 XThC.TB1.t1 132.067
R23141 XThC.TB1.n21 XThC.TB1.n13 61.4091
R23142 XThC.TB1.n16 XThC.TB1.n15 61.346
R23143 XThC.TB1.n10 XThC.TB1.n4 49.6611
R23144 XThC.TB1.n12 XThC.TB1.n11 45.2793
R23145 XThC.TB1.n7 XThC.TB1.n5 42.3581
R23146 XThC.TB1.n19 XThC.TB1.n14 30.6732
R23147 XThC.TB1.n19 XThC.TB1.n18 30.6732
R23148 XThC.TB1.n18 XThC.TB1.n17 30.6732
R23149 XThC.TB1.n17 XThC.TB1.n16 30.6732
R23150 XThC.TB1.n2 XThC.TB1.t0 26.5955
R23151 XThC.TB1.n2 XThC.TB1.t2 26.5955
R23152 XThC.TB1 XThC.TB1.n22 23.489
R23153 XThC.TB1.n9 XThC.TB1.n8 21.7605
R23154 XThC.TB1.n7 XThC.TB1.n6 18.9884
R23155 XThC.TB1.n12 XThC.TB1.n3 16.0672
R23156 XThC.TB1.n20 XThC.TB1 14.8485
R23157 XThC.TB1.n13 XThC.TB1 11.5205
R23158 XThC.TB1.n22 XThC.TB1.n21 10.7939
R23159 XThC.TB1.n9 XThC.TB1 10.2405
R23160 XThC.TB1 XThC.TB1.n20 8.7045
R23161 XThC.TB1.n21 XThC.TB1 8.41671
R23162 XThC.TB1.n5 XThC.TB1.n4 7.30353
R23163 XThC.TB1.n11 XThC.TB1.n10 4.38232
R23164 XThC.TB1.n1 XThC.TB1.n0 4.15748
R23165 XThC.TB1 XThC.TB1.n1 3.76521
R23166 XThC.TB1.n0 XThC.TB1 1.17559
R23167 XThC.TB1.n1 XThC.TB1 0.921363
R23168 XThC.Tn[8].n71 XThC.Tn[8].n70 256.104
R23169 XThC.Tn[8].n75 XThC.Tn[8].n74 243.679
R23170 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R23171 XThC.Tn[8].n75 XThC.Tn[8].n73 205.28
R23172 XThC.Tn[8].n71 XThC.Tn[8].n69 202.095
R23173 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R23174 XThC.Tn[8].n65 XThC.Tn[8].n63 161.365
R23175 XThC.Tn[8].n61 XThC.Tn[8].n59 161.365
R23176 XThC.Tn[8].n57 XThC.Tn[8].n55 161.365
R23177 XThC.Tn[8].n53 XThC.Tn[8].n51 161.365
R23178 XThC.Tn[8].n49 XThC.Tn[8].n47 161.365
R23179 XThC.Tn[8].n45 XThC.Tn[8].n43 161.365
R23180 XThC.Tn[8].n41 XThC.Tn[8].n39 161.365
R23181 XThC.Tn[8].n37 XThC.Tn[8].n35 161.365
R23182 XThC.Tn[8].n33 XThC.Tn[8].n31 161.365
R23183 XThC.Tn[8].n29 XThC.Tn[8].n27 161.365
R23184 XThC.Tn[8].n25 XThC.Tn[8].n23 161.365
R23185 XThC.Tn[8].n21 XThC.Tn[8].n19 161.365
R23186 XThC.Tn[8].n17 XThC.Tn[8].n15 161.365
R23187 XThC.Tn[8].n13 XThC.Tn[8].n11 161.365
R23188 XThC.Tn[8].n9 XThC.Tn[8].n7 161.365
R23189 XThC.Tn[8].n6 XThC.Tn[8].n4 161.365
R23190 XThC.Tn[8].n63 XThC.Tn[8].t15 161.202
R23191 XThC.Tn[8].n59 XThC.Tn[8].t37 161.202
R23192 XThC.Tn[8].n55 XThC.Tn[8].t24 161.202
R23193 XThC.Tn[8].n51 XThC.Tn[8].t21 161.202
R23194 XThC.Tn[8].n47 XThC.Tn[8].t13 161.202
R23195 XThC.Tn[8].n43 XThC.Tn[8].t32 161.202
R23196 XThC.Tn[8].n39 XThC.Tn[8].t31 161.202
R23197 XThC.Tn[8].n35 XThC.Tn[8].t12 161.202
R23198 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R23199 XThC.Tn[8].n27 XThC.Tn[8].t33 161.202
R23200 XThC.Tn[8].n23 XThC.Tn[8].t20 161.202
R23201 XThC.Tn[8].n19 XThC.Tn[8].t19 161.202
R23202 XThC.Tn[8].n15 XThC.Tn[8].t30 161.202
R23203 XThC.Tn[8].n11 XThC.Tn[8].t28 161.202
R23204 XThC.Tn[8].n7 XThC.Tn[8].t26 161.202
R23205 XThC.Tn[8].n4 XThC.Tn[8].t41 161.202
R23206 XThC.Tn[8].n63 XThC.Tn[8].t18 145.137
R23207 XThC.Tn[8].n59 XThC.Tn[8].t40 145.137
R23208 XThC.Tn[8].n55 XThC.Tn[8].t27 145.137
R23209 XThC.Tn[8].n51 XThC.Tn[8].t25 145.137
R23210 XThC.Tn[8].n47 XThC.Tn[8].t17 145.137
R23211 XThC.Tn[8].n43 XThC.Tn[8].t38 145.137
R23212 XThC.Tn[8].n39 XThC.Tn[8].t36 145.137
R23213 XThC.Tn[8].n35 XThC.Tn[8].t16 145.137
R23214 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R23215 XThC.Tn[8].n27 XThC.Tn[8].t39 145.137
R23216 XThC.Tn[8].n23 XThC.Tn[8].t23 145.137
R23217 XThC.Tn[8].n19 XThC.Tn[8].t22 145.137
R23218 XThC.Tn[8].n15 XThC.Tn[8].t35 145.137
R23219 XThC.Tn[8].n11 XThC.Tn[8].t34 145.137
R23220 XThC.Tn[8].n7 XThC.Tn[8].t29 145.137
R23221 XThC.Tn[8].n4 XThC.Tn[8].t43 145.137
R23222 XThC.Tn[8].n69 XThC.Tn[8].t9 26.5955
R23223 XThC.Tn[8].n69 XThC.Tn[8].t10 26.5955
R23224 XThC.Tn[8].n70 XThC.Tn[8].t8 26.5955
R23225 XThC.Tn[8].n70 XThC.Tn[8].t11 26.5955
R23226 XThC.Tn[8].n73 XThC.Tn[8].t2 26.5955
R23227 XThC.Tn[8].n73 XThC.Tn[8].t1 26.5955
R23228 XThC.Tn[8].n74 XThC.Tn[8].t0 26.5955
R23229 XThC.Tn[8].n74 XThC.Tn[8].t3 26.5955
R23230 XThC.Tn[8].n1 XThC.Tn[8].t7 24.9236
R23231 XThC.Tn[8].n1 XThC.Tn[8].t6 24.9236
R23232 XThC.Tn[8].n0 XThC.Tn[8].t5 24.9236
R23233 XThC.Tn[8].n0 XThC.Tn[8].t4 24.9236
R23234 XThC.Tn[8] XThC.Tn[8].n75 22.9652
R23235 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R23236 XThC.Tn[8].n72 XThC.Tn[8].n71 13.9299
R23237 XThC.Tn[8] XThC.Tn[8].n72 13.9299
R23238 XThC.Tn[8] XThC.Tn[8].n6 8.0245
R23239 XThC.Tn[8].n66 XThC.Tn[8].n65 7.9105
R23240 XThC.Tn[8].n62 XThC.Tn[8].n61 7.9105
R23241 XThC.Tn[8].n58 XThC.Tn[8].n57 7.9105
R23242 XThC.Tn[8].n54 XThC.Tn[8].n53 7.9105
R23243 XThC.Tn[8].n50 XThC.Tn[8].n49 7.9105
R23244 XThC.Tn[8].n46 XThC.Tn[8].n45 7.9105
R23245 XThC.Tn[8].n42 XThC.Tn[8].n41 7.9105
R23246 XThC.Tn[8].n38 XThC.Tn[8].n37 7.9105
R23247 XThC.Tn[8].n34 XThC.Tn[8].n33 7.9105
R23248 XThC.Tn[8].n30 XThC.Tn[8].n29 7.9105
R23249 XThC.Tn[8].n26 XThC.Tn[8].n25 7.9105
R23250 XThC.Tn[8].n22 XThC.Tn[8].n21 7.9105
R23251 XThC.Tn[8].n18 XThC.Tn[8].n17 7.9105
R23252 XThC.Tn[8].n14 XThC.Tn[8].n13 7.9105
R23253 XThC.Tn[8].n10 XThC.Tn[8].n9 7.9105
R23254 XThC.Tn[8].n68 XThC.Tn[8].n67 7.42331
R23255 XThC.Tn[8].n67 XThC.Tn[8] 4.24005
R23256 XThC.Tn[8].n72 XThC.Tn[8].n68 2.99115
R23257 XThC.Tn[8].n72 XThC.Tn[8] 2.87153
R23258 XThC.Tn[8].n68 XThC.Tn[8] 2.2734
R23259 XThC.Tn[8].n3 XThC.Tn[8] 0.672375
R23260 XThC.Tn[8].n10 XThC.Tn[8] 0.235138
R23261 XThC.Tn[8].n14 XThC.Tn[8] 0.235138
R23262 XThC.Tn[8].n18 XThC.Tn[8] 0.235138
R23263 XThC.Tn[8].n22 XThC.Tn[8] 0.235138
R23264 XThC.Tn[8].n26 XThC.Tn[8] 0.235138
R23265 XThC.Tn[8].n30 XThC.Tn[8] 0.235138
R23266 XThC.Tn[8].n34 XThC.Tn[8] 0.235138
R23267 XThC.Tn[8].n38 XThC.Tn[8] 0.235138
R23268 XThC.Tn[8].n42 XThC.Tn[8] 0.235138
R23269 XThC.Tn[8].n46 XThC.Tn[8] 0.235138
R23270 XThC.Tn[8].n50 XThC.Tn[8] 0.235138
R23271 XThC.Tn[8].n54 XThC.Tn[8] 0.235138
R23272 XThC.Tn[8].n58 XThC.Tn[8] 0.235138
R23273 XThC.Tn[8].n62 XThC.Tn[8] 0.235138
R23274 XThC.Tn[8].n66 XThC.Tn[8] 0.235138
R23275 XThC.Tn[8].n67 XThC.Tn[8].n3 0.220435
R23276 XThC.Tn[8].n3 XThC.Tn[8] 0.168469
R23277 XThC.Tn[8] XThC.Tn[8].n10 0.114505
R23278 XThC.Tn[8] XThC.Tn[8].n14 0.114505
R23279 XThC.Tn[8] XThC.Tn[8].n18 0.114505
R23280 XThC.Tn[8] XThC.Tn[8].n22 0.114505
R23281 XThC.Tn[8] XThC.Tn[8].n26 0.114505
R23282 XThC.Tn[8] XThC.Tn[8].n30 0.114505
R23283 XThC.Tn[8] XThC.Tn[8].n34 0.114505
R23284 XThC.Tn[8] XThC.Tn[8].n38 0.114505
R23285 XThC.Tn[8] XThC.Tn[8].n42 0.114505
R23286 XThC.Tn[8] XThC.Tn[8].n46 0.114505
R23287 XThC.Tn[8] XThC.Tn[8].n50 0.114505
R23288 XThC.Tn[8] XThC.Tn[8].n54 0.114505
R23289 XThC.Tn[8] XThC.Tn[8].n58 0.114505
R23290 XThC.Tn[8] XThC.Tn[8].n62 0.114505
R23291 XThC.Tn[8] XThC.Tn[8].n66 0.114505
R23292 XThC.Tn[8].n65 XThC.Tn[8].n64 0.0599512
R23293 XThC.Tn[8].n61 XThC.Tn[8].n60 0.0599512
R23294 XThC.Tn[8].n57 XThC.Tn[8].n56 0.0599512
R23295 XThC.Tn[8].n53 XThC.Tn[8].n52 0.0599512
R23296 XThC.Tn[8].n49 XThC.Tn[8].n48 0.0599512
R23297 XThC.Tn[8].n45 XThC.Tn[8].n44 0.0599512
R23298 XThC.Tn[8].n41 XThC.Tn[8].n40 0.0599512
R23299 XThC.Tn[8].n37 XThC.Tn[8].n36 0.0599512
R23300 XThC.Tn[8].n33 XThC.Tn[8].n32 0.0599512
R23301 XThC.Tn[8].n29 XThC.Tn[8].n28 0.0599512
R23302 XThC.Tn[8].n25 XThC.Tn[8].n24 0.0599512
R23303 XThC.Tn[8].n21 XThC.Tn[8].n20 0.0599512
R23304 XThC.Tn[8].n17 XThC.Tn[8].n16 0.0599512
R23305 XThC.Tn[8].n13 XThC.Tn[8].n12 0.0599512
R23306 XThC.Tn[8].n9 XThC.Tn[8].n8 0.0599512
R23307 XThC.Tn[8].n6 XThC.Tn[8].n5 0.0599512
R23308 XThC.Tn[8].n64 XThC.Tn[8] 0.0469286
R23309 XThC.Tn[8].n60 XThC.Tn[8] 0.0469286
R23310 XThC.Tn[8].n56 XThC.Tn[8] 0.0469286
R23311 XThC.Tn[8].n52 XThC.Tn[8] 0.0469286
R23312 XThC.Tn[8].n48 XThC.Tn[8] 0.0469286
R23313 XThC.Tn[8].n44 XThC.Tn[8] 0.0469286
R23314 XThC.Tn[8].n40 XThC.Tn[8] 0.0469286
R23315 XThC.Tn[8].n36 XThC.Tn[8] 0.0469286
R23316 XThC.Tn[8].n32 XThC.Tn[8] 0.0469286
R23317 XThC.Tn[8].n28 XThC.Tn[8] 0.0469286
R23318 XThC.Tn[8].n24 XThC.Tn[8] 0.0469286
R23319 XThC.Tn[8].n20 XThC.Tn[8] 0.0469286
R23320 XThC.Tn[8].n16 XThC.Tn[8] 0.0469286
R23321 XThC.Tn[8].n12 XThC.Tn[8] 0.0469286
R23322 XThC.Tn[8].n8 XThC.Tn[8] 0.0469286
R23323 XThC.Tn[8].n5 XThC.Tn[8] 0.0469286
R23324 XThC.Tn[8].n64 XThC.Tn[8] 0.0401341
R23325 XThC.Tn[8].n60 XThC.Tn[8] 0.0401341
R23326 XThC.Tn[8].n56 XThC.Tn[8] 0.0401341
R23327 XThC.Tn[8].n52 XThC.Tn[8] 0.0401341
R23328 XThC.Tn[8].n48 XThC.Tn[8] 0.0401341
R23329 XThC.Tn[8].n44 XThC.Tn[8] 0.0401341
R23330 XThC.Tn[8].n40 XThC.Tn[8] 0.0401341
R23331 XThC.Tn[8].n36 XThC.Tn[8] 0.0401341
R23332 XThC.Tn[8].n32 XThC.Tn[8] 0.0401341
R23333 XThC.Tn[8].n28 XThC.Tn[8] 0.0401341
R23334 XThC.Tn[8].n24 XThC.Tn[8] 0.0401341
R23335 XThC.Tn[8].n20 XThC.Tn[8] 0.0401341
R23336 XThC.Tn[8].n16 XThC.Tn[8] 0.0401341
R23337 XThC.Tn[8].n12 XThC.Tn[8] 0.0401341
R23338 XThC.Tn[8].n8 XThC.Tn[8] 0.0401341
R23339 XThC.Tn[8].n5 XThC.Tn[8] 0.0401341
R23340 XThR.Tn[1].n88 XThR.Tn[1].n87 332.334
R23341 XThR.Tn[1].n88 XThR.Tn[1].n86 296.493
R23342 XThR.Tn[1] XThR.Tn[1].n79 161.363
R23343 XThR.Tn[1] XThR.Tn[1].n74 161.363
R23344 XThR.Tn[1] XThR.Tn[1].n69 161.363
R23345 XThR.Tn[1] XThR.Tn[1].n64 161.363
R23346 XThR.Tn[1] XThR.Tn[1].n59 161.363
R23347 XThR.Tn[1] XThR.Tn[1].n54 161.363
R23348 XThR.Tn[1] XThR.Tn[1].n49 161.363
R23349 XThR.Tn[1] XThR.Tn[1].n44 161.363
R23350 XThR.Tn[1] XThR.Tn[1].n39 161.363
R23351 XThR.Tn[1] XThR.Tn[1].n34 161.363
R23352 XThR.Tn[1] XThR.Tn[1].n29 161.363
R23353 XThR.Tn[1] XThR.Tn[1].n24 161.363
R23354 XThR.Tn[1] XThR.Tn[1].n19 161.363
R23355 XThR.Tn[1] XThR.Tn[1].n14 161.363
R23356 XThR.Tn[1] XThR.Tn[1].n9 161.363
R23357 XThR.Tn[1] XThR.Tn[1].n7 161.363
R23358 XThR.Tn[1].n81 XThR.Tn[1].n80 161.3
R23359 XThR.Tn[1].n76 XThR.Tn[1].n75 161.3
R23360 XThR.Tn[1].n71 XThR.Tn[1].n70 161.3
R23361 XThR.Tn[1].n66 XThR.Tn[1].n65 161.3
R23362 XThR.Tn[1].n61 XThR.Tn[1].n60 161.3
R23363 XThR.Tn[1].n56 XThR.Tn[1].n55 161.3
R23364 XThR.Tn[1].n51 XThR.Tn[1].n50 161.3
R23365 XThR.Tn[1].n46 XThR.Tn[1].n45 161.3
R23366 XThR.Tn[1].n41 XThR.Tn[1].n40 161.3
R23367 XThR.Tn[1].n36 XThR.Tn[1].n35 161.3
R23368 XThR.Tn[1].n31 XThR.Tn[1].n30 161.3
R23369 XThR.Tn[1].n26 XThR.Tn[1].n25 161.3
R23370 XThR.Tn[1].n21 XThR.Tn[1].n20 161.3
R23371 XThR.Tn[1].n16 XThR.Tn[1].n15 161.3
R23372 XThR.Tn[1].n11 XThR.Tn[1].n10 161.3
R23373 XThR.Tn[1].n79 XThR.Tn[1].t70 161.106
R23374 XThR.Tn[1].n74 XThR.Tn[1].t14 161.106
R23375 XThR.Tn[1].n69 XThR.Tn[1].t56 161.106
R23376 XThR.Tn[1].n64 XThR.Tn[1].t42 161.106
R23377 XThR.Tn[1].n59 XThR.Tn[1].t68 161.106
R23378 XThR.Tn[1].n54 XThR.Tn[1].t31 161.106
R23379 XThR.Tn[1].n49 XThR.Tn[1].t12 161.106
R23380 XThR.Tn[1].n44 XThR.Tn[1].t54 161.106
R23381 XThR.Tn[1].n39 XThR.Tn[1].t41 161.106
R23382 XThR.Tn[1].n34 XThR.Tn[1].t46 161.106
R23383 XThR.Tn[1].n29 XThR.Tn[1].t29 161.106
R23384 XThR.Tn[1].n24 XThR.Tn[1].t55 161.106
R23385 XThR.Tn[1].n19 XThR.Tn[1].t28 161.106
R23386 XThR.Tn[1].n14 XThR.Tn[1].t73 161.106
R23387 XThR.Tn[1].n9 XThR.Tn[1].t34 161.106
R23388 XThR.Tn[1].n7 XThR.Tn[1].t18 161.106
R23389 XThR.Tn[1].n80 XThR.Tn[1].t66 159.978
R23390 XThR.Tn[1].n75 XThR.Tn[1].t72 159.978
R23391 XThR.Tn[1].n70 XThR.Tn[1].t52 159.978
R23392 XThR.Tn[1].n65 XThR.Tn[1].t39 159.978
R23393 XThR.Tn[1].n60 XThR.Tn[1].t63 159.978
R23394 XThR.Tn[1].n55 XThR.Tn[1].t27 159.978
R23395 XThR.Tn[1].n50 XThR.Tn[1].t71 159.978
R23396 XThR.Tn[1].n45 XThR.Tn[1].t49 159.978
R23397 XThR.Tn[1].n40 XThR.Tn[1].t36 159.978
R23398 XThR.Tn[1].n35 XThR.Tn[1].t43 159.978
R23399 XThR.Tn[1].n30 XThR.Tn[1].t26 159.978
R23400 XThR.Tn[1].n25 XThR.Tn[1].t51 159.978
R23401 XThR.Tn[1].n20 XThR.Tn[1].t25 159.978
R23402 XThR.Tn[1].n15 XThR.Tn[1].t69 159.978
R23403 XThR.Tn[1].n10 XThR.Tn[1].t30 159.978
R23404 XThR.Tn[1].n79 XThR.Tn[1].t58 145.038
R23405 XThR.Tn[1].n74 XThR.Tn[1].t20 145.038
R23406 XThR.Tn[1].n69 XThR.Tn[1].t62 145.038
R23407 XThR.Tn[1].n64 XThR.Tn[1].t47 145.038
R23408 XThR.Tn[1].n59 XThR.Tn[1].t15 145.038
R23409 XThR.Tn[1].n54 XThR.Tn[1].t57 145.038
R23410 XThR.Tn[1].n49 XThR.Tn[1].t64 145.038
R23411 XThR.Tn[1].n44 XThR.Tn[1].t48 145.038
R23412 XThR.Tn[1].n39 XThR.Tn[1].t45 145.038
R23413 XThR.Tn[1].n34 XThR.Tn[1].t13 145.038
R23414 XThR.Tn[1].n29 XThR.Tn[1].t37 145.038
R23415 XThR.Tn[1].n24 XThR.Tn[1].t59 145.038
R23416 XThR.Tn[1].n19 XThR.Tn[1].t35 145.038
R23417 XThR.Tn[1].n14 XThR.Tn[1].t19 145.038
R23418 XThR.Tn[1].n9 XThR.Tn[1].t44 145.038
R23419 XThR.Tn[1].n7 XThR.Tn[1].t24 145.038
R23420 XThR.Tn[1].n80 XThR.Tn[1].t17 143.911
R23421 XThR.Tn[1].n75 XThR.Tn[1].t40 143.911
R23422 XThR.Tn[1].n70 XThR.Tn[1].t22 143.911
R23423 XThR.Tn[1].n65 XThR.Tn[1].t65 143.911
R23424 XThR.Tn[1].n60 XThR.Tn[1].t33 143.911
R23425 XThR.Tn[1].n55 XThR.Tn[1].t16 143.911
R23426 XThR.Tn[1].n50 XThR.Tn[1].t23 143.911
R23427 XThR.Tn[1].n45 XThR.Tn[1].t67 143.911
R23428 XThR.Tn[1].n40 XThR.Tn[1].t60 143.911
R23429 XThR.Tn[1].n35 XThR.Tn[1].t32 143.911
R23430 XThR.Tn[1].n30 XThR.Tn[1].t53 143.911
R23431 XThR.Tn[1].n25 XThR.Tn[1].t21 143.911
R23432 XThR.Tn[1].n20 XThR.Tn[1].t50 143.911
R23433 XThR.Tn[1].n15 XThR.Tn[1].t38 143.911
R23434 XThR.Tn[1].n10 XThR.Tn[1].t61 143.911
R23435 XThR.Tn[1].n2 XThR.Tn[1].n0 135.249
R23436 XThR.Tn[1].n2 XThR.Tn[1].n1 98.981
R23437 XThR.Tn[1].n4 XThR.Tn[1].n3 98.981
R23438 XThR.Tn[1].n6 XThR.Tn[1].n5 98.981
R23439 XThR.Tn[1].n4 XThR.Tn[1].n2 36.2672
R23440 XThR.Tn[1].n6 XThR.Tn[1].n4 36.2672
R23441 XThR.Tn[1].n85 XThR.Tn[1].n6 32.6405
R23442 XThR.Tn[1].n86 XThR.Tn[1].t0 26.5955
R23443 XThR.Tn[1].n86 XThR.Tn[1].t1 26.5955
R23444 XThR.Tn[1].n87 XThR.Tn[1].t3 26.5955
R23445 XThR.Tn[1].n87 XThR.Tn[1].t2 26.5955
R23446 XThR.Tn[1].n0 XThR.Tn[1].t11 24.9236
R23447 XThR.Tn[1].n0 XThR.Tn[1].t8 24.9236
R23448 XThR.Tn[1].n1 XThR.Tn[1].t10 24.9236
R23449 XThR.Tn[1].n1 XThR.Tn[1].t9 24.9236
R23450 XThR.Tn[1].n3 XThR.Tn[1].t6 24.9236
R23451 XThR.Tn[1].n3 XThR.Tn[1].t5 24.9236
R23452 XThR.Tn[1].n5 XThR.Tn[1].t7 24.9236
R23453 XThR.Tn[1].n5 XThR.Tn[1].t4 24.9236
R23454 XThR.Tn[1].n89 XThR.Tn[1].n88 18.5605
R23455 XThR.Tn[1].n89 XThR.Tn[1].n85 11.5205
R23456 XThR.Tn[1].n85 XThR.Tn[1] 6.42118
R23457 XThR.Tn[1] XThR.Tn[1].n8 5.34038
R23458 XThR.Tn[1].n13 XThR.Tn[1].n12 4.5005
R23459 XThR.Tn[1].n18 XThR.Tn[1].n17 4.5005
R23460 XThR.Tn[1].n23 XThR.Tn[1].n22 4.5005
R23461 XThR.Tn[1].n28 XThR.Tn[1].n27 4.5005
R23462 XThR.Tn[1].n33 XThR.Tn[1].n32 4.5005
R23463 XThR.Tn[1].n38 XThR.Tn[1].n37 4.5005
R23464 XThR.Tn[1].n43 XThR.Tn[1].n42 4.5005
R23465 XThR.Tn[1].n48 XThR.Tn[1].n47 4.5005
R23466 XThR.Tn[1].n53 XThR.Tn[1].n52 4.5005
R23467 XThR.Tn[1].n58 XThR.Tn[1].n57 4.5005
R23468 XThR.Tn[1].n63 XThR.Tn[1].n62 4.5005
R23469 XThR.Tn[1].n68 XThR.Tn[1].n67 4.5005
R23470 XThR.Tn[1].n73 XThR.Tn[1].n72 4.5005
R23471 XThR.Tn[1].n78 XThR.Tn[1].n77 4.5005
R23472 XThR.Tn[1].n83 XThR.Tn[1].n82 4.5005
R23473 XThR.Tn[1].n84 XThR.Tn[1] 3.70586
R23474 XThR.Tn[1].n13 XThR.Tn[1] 2.52282
R23475 XThR.Tn[1].n18 XThR.Tn[1] 2.52282
R23476 XThR.Tn[1].n23 XThR.Tn[1] 2.52282
R23477 XThR.Tn[1].n28 XThR.Tn[1] 2.52282
R23478 XThR.Tn[1].n33 XThR.Tn[1] 2.52282
R23479 XThR.Tn[1].n38 XThR.Tn[1] 2.52282
R23480 XThR.Tn[1].n43 XThR.Tn[1] 2.52282
R23481 XThR.Tn[1].n48 XThR.Tn[1] 2.52282
R23482 XThR.Tn[1].n53 XThR.Tn[1] 2.52282
R23483 XThR.Tn[1].n58 XThR.Tn[1] 2.52282
R23484 XThR.Tn[1].n63 XThR.Tn[1] 2.52282
R23485 XThR.Tn[1].n68 XThR.Tn[1] 2.52282
R23486 XThR.Tn[1].n73 XThR.Tn[1] 2.52282
R23487 XThR.Tn[1].n78 XThR.Tn[1] 2.52282
R23488 XThR.Tn[1].n83 XThR.Tn[1] 2.52282
R23489 XThR.Tn[1].n81 XThR.Tn[1] 1.08677
R23490 XThR.Tn[1].n76 XThR.Tn[1] 1.08677
R23491 XThR.Tn[1].n71 XThR.Tn[1] 1.08677
R23492 XThR.Tn[1].n66 XThR.Tn[1] 1.08677
R23493 XThR.Tn[1].n61 XThR.Tn[1] 1.08677
R23494 XThR.Tn[1].n56 XThR.Tn[1] 1.08677
R23495 XThR.Tn[1].n51 XThR.Tn[1] 1.08677
R23496 XThR.Tn[1].n46 XThR.Tn[1] 1.08677
R23497 XThR.Tn[1].n41 XThR.Tn[1] 1.08677
R23498 XThR.Tn[1].n36 XThR.Tn[1] 1.08677
R23499 XThR.Tn[1].n31 XThR.Tn[1] 1.08677
R23500 XThR.Tn[1].n26 XThR.Tn[1] 1.08677
R23501 XThR.Tn[1].n21 XThR.Tn[1] 1.08677
R23502 XThR.Tn[1].n16 XThR.Tn[1] 1.08677
R23503 XThR.Tn[1].n11 XThR.Tn[1] 1.08677
R23504 XThR.Tn[1] XThR.Tn[1].n13 0.839786
R23505 XThR.Tn[1] XThR.Tn[1].n18 0.839786
R23506 XThR.Tn[1] XThR.Tn[1].n23 0.839786
R23507 XThR.Tn[1] XThR.Tn[1].n28 0.839786
R23508 XThR.Tn[1] XThR.Tn[1].n33 0.839786
R23509 XThR.Tn[1] XThR.Tn[1].n38 0.839786
R23510 XThR.Tn[1] XThR.Tn[1].n43 0.839786
R23511 XThR.Tn[1] XThR.Tn[1].n48 0.839786
R23512 XThR.Tn[1] XThR.Tn[1].n53 0.839786
R23513 XThR.Tn[1] XThR.Tn[1].n58 0.839786
R23514 XThR.Tn[1] XThR.Tn[1].n63 0.839786
R23515 XThR.Tn[1] XThR.Tn[1].n68 0.839786
R23516 XThR.Tn[1] XThR.Tn[1].n73 0.839786
R23517 XThR.Tn[1] XThR.Tn[1].n78 0.839786
R23518 XThR.Tn[1] XThR.Tn[1].n83 0.839786
R23519 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R23520 XThR.Tn[1].n8 XThR.Tn[1] 0.499542
R23521 XThR.Tn[1].n82 XThR.Tn[1] 0.063
R23522 XThR.Tn[1].n77 XThR.Tn[1] 0.063
R23523 XThR.Tn[1].n72 XThR.Tn[1] 0.063
R23524 XThR.Tn[1].n67 XThR.Tn[1] 0.063
R23525 XThR.Tn[1].n62 XThR.Tn[1] 0.063
R23526 XThR.Tn[1].n57 XThR.Tn[1] 0.063
R23527 XThR.Tn[1].n52 XThR.Tn[1] 0.063
R23528 XThR.Tn[1].n47 XThR.Tn[1] 0.063
R23529 XThR.Tn[1].n42 XThR.Tn[1] 0.063
R23530 XThR.Tn[1].n37 XThR.Tn[1] 0.063
R23531 XThR.Tn[1].n32 XThR.Tn[1] 0.063
R23532 XThR.Tn[1].n27 XThR.Tn[1] 0.063
R23533 XThR.Tn[1].n22 XThR.Tn[1] 0.063
R23534 XThR.Tn[1].n17 XThR.Tn[1] 0.063
R23535 XThR.Tn[1].n12 XThR.Tn[1] 0.063
R23536 XThR.Tn[1].n84 XThR.Tn[1] 0.0540714
R23537 XThR.Tn[1] XThR.Tn[1].n84 0.038
R23538 XThR.Tn[1].n8 XThR.Tn[1] 0.0143889
R23539 XThR.Tn[1].n82 XThR.Tn[1].n81 0.00771154
R23540 XThR.Tn[1].n77 XThR.Tn[1].n76 0.00771154
R23541 XThR.Tn[1].n72 XThR.Tn[1].n71 0.00771154
R23542 XThR.Tn[1].n67 XThR.Tn[1].n66 0.00771154
R23543 XThR.Tn[1].n62 XThR.Tn[1].n61 0.00771154
R23544 XThR.Tn[1].n57 XThR.Tn[1].n56 0.00771154
R23545 XThR.Tn[1].n52 XThR.Tn[1].n51 0.00771154
R23546 XThR.Tn[1].n47 XThR.Tn[1].n46 0.00771154
R23547 XThR.Tn[1].n42 XThR.Tn[1].n41 0.00771154
R23548 XThR.Tn[1].n37 XThR.Tn[1].n36 0.00771154
R23549 XThR.Tn[1].n32 XThR.Tn[1].n31 0.00771154
R23550 XThR.Tn[1].n27 XThR.Tn[1].n26 0.00771154
R23551 XThR.Tn[1].n22 XThR.Tn[1].n21 0.00771154
R23552 XThR.Tn[1].n17 XThR.Tn[1].n16 0.00771154
R23553 XThR.Tn[1].n12 XThR.Tn[1].n11 0.00771154
R23554 XThC.Tn[7].n2 XThC.Tn[7].n1 255.096
R23555 XThC.Tn[7].n69 XThC.Tn[7].n67 236.589
R23556 XThC.Tn[7].n2 XThC.Tn[7].n0 201.845
R23557 XThC.Tn[7].n69 XThC.Tn[7].n68 200.321
R23558 XThC.Tn[7].n64 XThC.Tn[7].n62 161.365
R23559 XThC.Tn[7].n60 XThC.Tn[7].n58 161.365
R23560 XThC.Tn[7].n56 XThC.Tn[7].n54 161.365
R23561 XThC.Tn[7].n52 XThC.Tn[7].n50 161.365
R23562 XThC.Tn[7].n48 XThC.Tn[7].n46 161.365
R23563 XThC.Tn[7].n44 XThC.Tn[7].n42 161.365
R23564 XThC.Tn[7].n40 XThC.Tn[7].n38 161.365
R23565 XThC.Tn[7].n36 XThC.Tn[7].n34 161.365
R23566 XThC.Tn[7].n32 XThC.Tn[7].n30 161.365
R23567 XThC.Tn[7].n28 XThC.Tn[7].n26 161.365
R23568 XThC.Tn[7].n24 XThC.Tn[7].n22 161.365
R23569 XThC.Tn[7].n20 XThC.Tn[7].n18 161.365
R23570 XThC.Tn[7].n16 XThC.Tn[7].n14 161.365
R23571 XThC.Tn[7].n12 XThC.Tn[7].n10 161.365
R23572 XThC.Tn[7].n8 XThC.Tn[7].n6 161.365
R23573 XThC.Tn[7].n5 XThC.Tn[7].n3 161.365
R23574 XThC.Tn[7].n62 XThC.Tn[7].t19 161.202
R23575 XThC.Tn[7].n58 XThC.Tn[7].t9 161.202
R23576 XThC.Tn[7].n54 XThC.Tn[7].t28 161.202
R23577 XThC.Tn[7].n50 XThC.Tn[7].t26 161.202
R23578 XThC.Tn[7].n46 XThC.Tn[7].t17 161.202
R23579 XThC.Tn[7].n42 XThC.Tn[7].t38 161.202
R23580 XThC.Tn[7].n38 XThC.Tn[7].t36 161.202
R23581 XThC.Tn[7].n34 XThC.Tn[7].t16 161.202
R23582 XThC.Tn[7].n30 XThC.Tn[7].t14 161.202
R23583 XThC.Tn[7].n26 XThC.Tn[7].t39 161.202
R23584 XThC.Tn[7].n22 XThC.Tn[7].t23 161.202
R23585 XThC.Tn[7].n18 XThC.Tn[7].t22 161.202
R23586 XThC.Tn[7].n14 XThC.Tn[7].t35 161.202
R23587 XThC.Tn[7].n10 XThC.Tn[7].t34 161.202
R23588 XThC.Tn[7].n6 XThC.Tn[7].t30 161.202
R23589 XThC.Tn[7].n3 XThC.Tn[7].t11 161.202
R23590 XThC.Tn[7].n62 XThC.Tn[7].t15 145.137
R23591 XThC.Tn[7].n58 XThC.Tn[7].t37 145.137
R23592 XThC.Tn[7].n54 XThC.Tn[7].t24 145.137
R23593 XThC.Tn[7].n50 XThC.Tn[7].t21 145.137
R23594 XThC.Tn[7].n46 XThC.Tn[7].t13 145.137
R23595 XThC.Tn[7].n42 XThC.Tn[7].t32 145.137
R23596 XThC.Tn[7].n38 XThC.Tn[7].t31 145.137
R23597 XThC.Tn[7].n34 XThC.Tn[7].t12 145.137
R23598 XThC.Tn[7].n30 XThC.Tn[7].t10 145.137
R23599 XThC.Tn[7].n26 XThC.Tn[7].t33 145.137
R23600 XThC.Tn[7].n22 XThC.Tn[7].t20 145.137
R23601 XThC.Tn[7].n18 XThC.Tn[7].t18 145.137
R23602 XThC.Tn[7].n14 XThC.Tn[7].t29 145.137
R23603 XThC.Tn[7].n10 XThC.Tn[7].t27 145.137
R23604 XThC.Tn[7].n6 XThC.Tn[7].t25 145.137
R23605 XThC.Tn[7].n3 XThC.Tn[7].t8 145.137
R23606 XThC.Tn[7].n0 XThC.Tn[7].t4 26.5955
R23607 XThC.Tn[7].n0 XThC.Tn[7].t7 26.5955
R23608 XThC.Tn[7].n1 XThC.Tn[7].t6 26.5955
R23609 XThC.Tn[7].n1 XThC.Tn[7].t5 26.5955
R23610 XThC.Tn[7] XThC.Tn[7].n2 26.5002
R23611 XThC.Tn[7].n67 XThC.Tn[7].t2 24.9236
R23612 XThC.Tn[7].n67 XThC.Tn[7].t1 24.9236
R23613 XThC.Tn[7].n68 XThC.Tn[7].t0 24.9236
R23614 XThC.Tn[7].n68 XThC.Tn[7].t3 24.9236
R23615 XThC.Tn[7].n70 XThC.Tn[7].n69 12.0894
R23616 XThC.Tn[7].n70 XThC.Tn[7] 9.64206
R23617 XThC.Tn[7].n66 XThC.Tn[7] 8.14595
R23618 XThC.Tn[7] XThC.Tn[7].n5 8.0245
R23619 XThC.Tn[7].n65 XThC.Tn[7].n64 7.9105
R23620 XThC.Tn[7].n61 XThC.Tn[7].n60 7.9105
R23621 XThC.Tn[7].n57 XThC.Tn[7].n56 7.9105
R23622 XThC.Tn[7].n53 XThC.Tn[7].n52 7.9105
R23623 XThC.Tn[7].n49 XThC.Tn[7].n48 7.9105
R23624 XThC.Tn[7].n45 XThC.Tn[7].n44 7.9105
R23625 XThC.Tn[7].n41 XThC.Tn[7].n40 7.9105
R23626 XThC.Tn[7].n37 XThC.Tn[7].n36 7.9105
R23627 XThC.Tn[7].n33 XThC.Tn[7].n32 7.9105
R23628 XThC.Tn[7].n29 XThC.Tn[7].n28 7.9105
R23629 XThC.Tn[7].n25 XThC.Tn[7].n24 7.9105
R23630 XThC.Tn[7].n21 XThC.Tn[7].n20 7.9105
R23631 XThC.Tn[7].n17 XThC.Tn[7].n16 7.9105
R23632 XThC.Tn[7].n13 XThC.Tn[7].n12 7.9105
R23633 XThC.Tn[7].n9 XThC.Tn[7].n8 7.9105
R23634 XThC.Tn[7].n66 XThC.Tn[7] 5.30358
R23635 XThC.Tn[7] XThC.Tn[7].n66 3.15894
R23636 XThC.Tn[7] XThC.Tn[7].n70 1.66284
R23637 XThC.Tn[7].n9 XThC.Tn[7] 0.235138
R23638 XThC.Tn[7].n13 XThC.Tn[7] 0.235138
R23639 XThC.Tn[7].n17 XThC.Tn[7] 0.235138
R23640 XThC.Tn[7].n21 XThC.Tn[7] 0.235138
R23641 XThC.Tn[7].n25 XThC.Tn[7] 0.235138
R23642 XThC.Tn[7].n29 XThC.Tn[7] 0.235138
R23643 XThC.Tn[7].n33 XThC.Tn[7] 0.235138
R23644 XThC.Tn[7].n37 XThC.Tn[7] 0.235138
R23645 XThC.Tn[7].n41 XThC.Tn[7] 0.235138
R23646 XThC.Tn[7].n45 XThC.Tn[7] 0.235138
R23647 XThC.Tn[7].n49 XThC.Tn[7] 0.235138
R23648 XThC.Tn[7].n53 XThC.Tn[7] 0.235138
R23649 XThC.Tn[7].n57 XThC.Tn[7] 0.235138
R23650 XThC.Tn[7].n61 XThC.Tn[7] 0.235138
R23651 XThC.Tn[7].n65 XThC.Tn[7] 0.235138
R23652 XThC.Tn[7] XThC.Tn[7].n9 0.114505
R23653 XThC.Tn[7] XThC.Tn[7].n13 0.114505
R23654 XThC.Tn[7] XThC.Tn[7].n17 0.114505
R23655 XThC.Tn[7] XThC.Tn[7].n21 0.114505
R23656 XThC.Tn[7] XThC.Tn[7].n25 0.114505
R23657 XThC.Tn[7] XThC.Tn[7].n29 0.114505
R23658 XThC.Tn[7] XThC.Tn[7].n33 0.114505
R23659 XThC.Tn[7] XThC.Tn[7].n37 0.114505
R23660 XThC.Tn[7] XThC.Tn[7].n41 0.114505
R23661 XThC.Tn[7] XThC.Tn[7].n45 0.114505
R23662 XThC.Tn[7] XThC.Tn[7].n49 0.114505
R23663 XThC.Tn[7] XThC.Tn[7].n53 0.114505
R23664 XThC.Tn[7] XThC.Tn[7].n57 0.114505
R23665 XThC.Tn[7] XThC.Tn[7].n61 0.114505
R23666 XThC.Tn[7] XThC.Tn[7].n65 0.114505
R23667 XThC.Tn[7].n64 XThC.Tn[7].n63 0.0599512
R23668 XThC.Tn[7].n60 XThC.Tn[7].n59 0.0599512
R23669 XThC.Tn[7].n56 XThC.Tn[7].n55 0.0599512
R23670 XThC.Tn[7].n52 XThC.Tn[7].n51 0.0599512
R23671 XThC.Tn[7].n48 XThC.Tn[7].n47 0.0599512
R23672 XThC.Tn[7].n44 XThC.Tn[7].n43 0.0599512
R23673 XThC.Tn[7].n40 XThC.Tn[7].n39 0.0599512
R23674 XThC.Tn[7].n36 XThC.Tn[7].n35 0.0599512
R23675 XThC.Tn[7].n32 XThC.Tn[7].n31 0.0599512
R23676 XThC.Tn[7].n28 XThC.Tn[7].n27 0.0599512
R23677 XThC.Tn[7].n24 XThC.Tn[7].n23 0.0599512
R23678 XThC.Tn[7].n20 XThC.Tn[7].n19 0.0599512
R23679 XThC.Tn[7].n16 XThC.Tn[7].n15 0.0599512
R23680 XThC.Tn[7].n12 XThC.Tn[7].n11 0.0599512
R23681 XThC.Tn[7].n8 XThC.Tn[7].n7 0.0599512
R23682 XThC.Tn[7].n5 XThC.Tn[7].n4 0.0599512
R23683 XThC.Tn[7].n63 XThC.Tn[7] 0.0469286
R23684 XThC.Tn[7].n59 XThC.Tn[7] 0.0469286
R23685 XThC.Tn[7].n55 XThC.Tn[7] 0.0469286
R23686 XThC.Tn[7].n51 XThC.Tn[7] 0.0469286
R23687 XThC.Tn[7].n47 XThC.Tn[7] 0.0469286
R23688 XThC.Tn[7].n43 XThC.Tn[7] 0.0469286
R23689 XThC.Tn[7].n39 XThC.Tn[7] 0.0469286
R23690 XThC.Tn[7].n35 XThC.Tn[7] 0.0469286
R23691 XThC.Tn[7].n31 XThC.Tn[7] 0.0469286
R23692 XThC.Tn[7].n27 XThC.Tn[7] 0.0469286
R23693 XThC.Tn[7].n23 XThC.Tn[7] 0.0469286
R23694 XThC.Tn[7].n19 XThC.Tn[7] 0.0469286
R23695 XThC.Tn[7].n15 XThC.Tn[7] 0.0469286
R23696 XThC.Tn[7].n11 XThC.Tn[7] 0.0469286
R23697 XThC.Tn[7].n7 XThC.Tn[7] 0.0469286
R23698 XThC.Tn[7].n4 XThC.Tn[7] 0.0469286
R23699 XThC.Tn[7].n63 XThC.Tn[7] 0.0401341
R23700 XThC.Tn[7].n59 XThC.Tn[7] 0.0401341
R23701 XThC.Tn[7].n55 XThC.Tn[7] 0.0401341
R23702 XThC.Tn[7].n51 XThC.Tn[7] 0.0401341
R23703 XThC.Tn[7].n47 XThC.Tn[7] 0.0401341
R23704 XThC.Tn[7].n43 XThC.Tn[7] 0.0401341
R23705 XThC.Tn[7].n39 XThC.Tn[7] 0.0401341
R23706 XThC.Tn[7].n35 XThC.Tn[7] 0.0401341
R23707 XThC.Tn[7].n31 XThC.Tn[7] 0.0401341
R23708 XThC.Tn[7].n27 XThC.Tn[7] 0.0401341
R23709 XThC.Tn[7].n23 XThC.Tn[7] 0.0401341
R23710 XThC.Tn[7].n19 XThC.Tn[7] 0.0401341
R23711 XThC.Tn[7].n15 XThC.Tn[7] 0.0401341
R23712 XThC.Tn[7].n11 XThC.Tn[7] 0.0401341
R23713 XThC.Tn[7].n7 XThC.Tn[7] 0.0401341
R23714 XThC.Tn[7].n4 XThC.Tn[7] 0.0401341
R23715 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R23716 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R23717 XThR.Tn[4] XThR.Tn[4].n82 161.363
R23718 XThR.Tn[4] XThR.Tn[4].n77 161.363
R23719 XThR.Tn[4] XThR.Tn[4].n72 161.363
R23720 XThR.Tn[4] XThR.Tn[4].n67 161.363
R23721 XThR.Tn[4] XThR.Tn[4].n62 161.363
R23722 XThR.Tn[4] XThR.Tn[4].n57 161.363
R23723 XThR.Tn[4] XThR.Tn[4].n52 161.363
R23724 XThR.Tn[4] XThR.Tn[4].n47 161.363
R23725 XThR.Tn[4] XThR.Tn[4].n42 161.363
R23726 XThR.Tn[4] XThR.Tn[4].n37 161.363
R23727 XThR.Tn[4] XThR.Tn[4].n32 161.363
R23728 XThR.Tn[4] XThR.Tn[4].n27 161.363
R23729 XThR.Tn[4] XThR.Tn[4].n22 161.363
R23730 XThR.Tn[4] XThR.Tn[4].n17 161.363
R23731 XThR.Tn[4] XThR.Tn[4].n12 161.363
R23732 XThR.Tn[4] XThR.Tn[4].n10 161.363
R23733 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R23734 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R23735 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R23736 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R23737 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R23738 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R23739 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R23740 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R23741 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R23742 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R23743 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R23744 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R23745 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R23746 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R23747 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R23748 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R23749 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R23750 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R23751 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R23752 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R23753 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R23754 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R23755 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R23756 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R23757 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R23758 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R23759 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R23760 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R23761 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R23762 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R23763 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R23764 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R23765 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R23766 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R23767 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R23768 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R23769 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R23770 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R23771 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R23772 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R23773 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R23774 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R23775 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R23776 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R23777 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R23778 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R23779 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R23780 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R23781 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R23782 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R23783 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R23784 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R23785 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R23786 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R23787 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R23788 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R23789 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R23790 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R23791 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R23792 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R23793 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R23794 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R23795 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R23796 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R23797 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R23798 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R23799 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R23800 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R23801 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R23802 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R23803 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R23804 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R23805 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R23806 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R23807 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R23808 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R23809 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R23810 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R23811 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R23812 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R23813 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R23814 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R23815 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R23816 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R23817 XThR.Tn[4].n1 XThR.Tn[4].t4 26.5955
R23818 XThR.Tn[4].n1 XThR.Tn[4].t7 26.5955
R23819 XThR.Tn[4].n0 XThR.Tn[4].t5 26.5955
R23820 XThR.Tn[4].n0 XThR.Tn[4].t6 26.5955
R23821 XThR.Tn[4].n3 XThR.Tn[4].t11 24.9236
R23822 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R23823 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R23824 XThR.Tn[4].n4 XThR.Tn[4].t9 24.9236
R23825 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R23826 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R23827 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R23828 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R23829 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R23830 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R23831 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R23832 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R23833 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R23834 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R23835 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R23836 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R23837 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R23838 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R23839 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R23840 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R23841 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R23842 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R23843 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R23844 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R23845 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R23846 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R23847 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R23848 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R23849 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R23850 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R23851 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R23852 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R23853 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R23854 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R23855 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R23856 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R23857 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R23858 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R23859 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R23860 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R23861 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R23862 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R23863 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R23864 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R23865 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R23866 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R23867 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R23868 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R23869 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R23870 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R23871 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R23872 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R23873 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R23874 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R23875 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R23876 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R23877 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R23878 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R23879 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R23880 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R23881 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R23882 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R23883 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R23884 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R23885 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R23886 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R23887 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R23888 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R23889 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R23890 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R23891 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R23892 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R23893 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R23894 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R23895 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R23896 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R23897 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R23898 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R23899 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R23900 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R23901 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R23902 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R23903 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R23904 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R23905 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R23906 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R23907 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R23908 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R23909 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R23910 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R23911 XThR.Tn[4] XThR.Tn[4].n87 0.038
R23912 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R23913 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R23914 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R23915 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R23916 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R23917 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R23918 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R23919 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R23920 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R23921 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R23922 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R23923 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R23924 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R23925 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R23926 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R23927 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R23928 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R23929 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R23930 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R23931 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R23932 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R23933 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R23934 XThR.Tn[11] XThR.Tn[11].n82 161.363
R23935 XThR.Tn[11] XThR.Tn[11].n77 161.363
R23936 XThR.Tn[11] XThR.Tn[11].n72 161.363
R23937 XThR.Tn[11] XThR.Tn[11].n67 161.363
R23938 XThR.Tn[11] XThR.Tn[11].n62 161.363
R23939 XThR.Tn[11] XThR.Tn[11].n57 161.363
R23940 XThR.Tn[11] XThR.Tn[11].n52 161.363
R23941 XThR.Tn[11] XThR.Tn[11].n47 161.363
R23942 XThR.Tn[11] XThR.Tn[11].n42 161.363
R23943 XThR.Tn[11] XThR.Tn[11].n37 161.363
R23944 XThR.Tn[11] XThR.Tn[11].n32 161.363
R23945 XThR.Tn[11] XThR.Tn[11].n27 161.363
R23946 XThR.Tn[11] XThR.Tn[11].n22 161.363
R23947 XThR.Tn[11] XThR.Tn[11].n17 161.363
R23948 XThR.Tn[11] XThR.Tn[11].n12 161.363
R23949 XThR.Tn[11] XThR.Tn[11].n10 161.363
R23950 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R23951 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R23952 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R23953 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R23954 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R23955 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R23956 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R23957 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R23958 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R23959 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R23960 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R23961 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R23962 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R23963 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R23964 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R23965 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R23966 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R23967 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R23968 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R23969 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R23970 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R23971 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R23972 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R23973 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R23974 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R23975 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R23976 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R23977 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R23978 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R23979 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R23980 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R23981 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R23982 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R23983 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R23984 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R23985 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R23986 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R23987 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R23988 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R23989 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R23990 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R23991 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R23992 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R23993 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R23994 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R23995 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R23996 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R23997 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R23998 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R23999 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R24000 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R24001 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R24002 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R24003 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R24004 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R24005 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R24006 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R24007 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R24008 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R24009 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R24010 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R24011 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R24012 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R24013 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R24014 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R24015 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R24016 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R24017 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R24018 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R24019 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R24020 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R24021 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R24022 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R24023 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R24024 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R24025 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R24026 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R24027 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R24028 XThR.Tn[11].n6 XThR.Tn[11].t4 26.5955
R24029 XThR.Tn[11].n6 XThR.Tn[11].t6 26.5955
R24030 XThR.Tn[11].n7 XThR.Tn[11].t5 26.5955
R24031 XThR.Tn[11].n7 XThR.Tn[11].t7 26.5955
R24032 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R24033 XThR.Tn[11].n3 XThR.Tn[11].t10 26.5955
R24034 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R24035 XThR.Tn[11].n4 XThR.Tn[11].t11 26.5955
R24036 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R24037 XThR.Tn[11].n0 XThR.Tn[11].t0 24.9236
R24038 XThR.Tn[11].n1 XThR.Tn[11].t3 24.9236
R24039 XThR.Tn[11].n1 XThR.Tn[11].t1 24.9236
R24040 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R24041 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R24042 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R24043 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R24044 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R24045 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R24046 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R24047 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R24048 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R24049 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R24050 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R24051 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R24052 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R24053 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R24054 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R24055 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R24056 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R24057 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R24058 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R24059 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R24060 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R24061 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R24062 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R24063 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R24064 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R24065 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R24066 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R24067 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R24068 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R24069 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R24070 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R24071 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R24072 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R24073 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R24074 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R24075 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R24076 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R24077 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R24078 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R24079 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R24080 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R24081 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R24082 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R24083 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R24084 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R24085 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R24086 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R24087 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R24088 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R24089 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R24090 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R24091 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R24092 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R24093 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R24094 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R24095 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R24096 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R24097 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R24098 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R24099 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R24100 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R24101 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R24102 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R24103 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R24104 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R24105 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R24106 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R24107 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R24108 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R24109 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R24110 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R24111 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R24112 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R24113 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R24114 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R24115 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R24116 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R24117 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R24118 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R24119 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R24120 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R24121 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R24122 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R24123 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R24124 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R24125 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R24126 XThR.Tn[11] XThR.Tn[11].n87 0.038
R24127 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R24128 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R24129 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R24130 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R24131 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R24132 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R24133 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R24134 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R24135 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R24136 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R24137 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R24138 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R24139 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R24140 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R24141 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R24142 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R24143 XThR.Tn[7].n5 XThR.Tn[7].n3 244.069
R24144 XThR.Tn[7].n2 XThR.Tn[7].n1 236.589
R24145 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R24146 XThR.Tn[7].n2 XThR.Tn[7].n0 200.321
R24147 XThR.Tn[7] XThR.Tn[7].n79 161.363
R24148 XThR.Tn[7] XThR.Tn[7].n74 161.363
R24149 XThR.Tn[7] XThR.Tn[7].n69 161.363
R24150 XThR.Tn[7] XThR.Tn[7].n64 161.363
R24151 XThR.Tn[7] XThR.Tn[7].n59 161.363
R24152 XThR.Tn[7] XThR.Tn[7].n54 161.363
R24153 XThR.Tn[7] XThR.Tn[7].n49 161.363
R24154 XThR.Tn[7] XThR.Tn[7].n44 161.363
R24155 XThR.Tn[7] XThR.Tn[7].n39 161.363
R24156 XThR.Tn[7] XThR.Tn[7].n34 161.363
R24157 XThR.Tn[7] XThR.Tn[7].n29 161.363
R24158 XThR.Tn[7] XThR.Tn[7].n24 161.363
R24159 XThR.Tn[7] XThR.Tn[7].n19 161.363
R24160 XThR.Tn[7] XThR.Tn[7].n14 161.363
R24161 XThR.Tn[7] XThR.Tn[7].n9 161.363
R24162 XThR.Tn[7] XThR.Tn[7].n7 161.363
R24163 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R24164 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R24165 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R24166 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R24167 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R24168 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R24169 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R24170 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R24171 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R24172 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R24173 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R24174 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R24175 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R24176 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R24177 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R24178 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R24179 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R24180 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R24181 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R24182 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R24183 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R24184 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R24185 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R24186 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R24187 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R24188 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R24189 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R24190 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R24191 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R24192 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R24193 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R24194 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R24195 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R24196 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R24197 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R24198 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R24199 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R24200 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R24201 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R24202 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R24203 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R24204 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R24205 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R24206 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R24207 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R24208 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R24209 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R24210 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R24211 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R24212 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R24213 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R24214 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R24215 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R24216 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R24217 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R24218 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R24219 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R24220 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R24221 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R24222 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R24223 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R24224 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R24225 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R24226 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R24227 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R24228 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R24229 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R24230 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R24231 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R24232 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R24233 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R24234 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R24235 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R24236 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R24237 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R24238 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R24239 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R24240 XThR.Tn[7].n4 XThR.Tn[7].t5 26.5955
R24241 XThR.Tn[7].n4 XThR.Tn[7].t4 26.5955
R24242 XThR.Tn[7].n3 XThR.Tn[7].t6 26.5955
R24243 XThR.Tn[7].n3 XThR.Tn[7].t7 26.5955
R24244 XThR.Tn[7].n0 XThR.Tn[7].t2 24.9236
R24245 XThR.Tn[7].n0 XThR.Tn[7].t1 24.9236
R24246 XThR.Tn[7].n1 XThR.Tn[7].t3 24.9236
R24247 XThR.Tn[7].n1 XThR.Tn[7].t0 24.9236
R24248 XThR.Tn[7] XThR.Tn[7].n2 16.079
R24249 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R24250 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R24251 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R24252 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R24253 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R24254 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R24255 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R24256 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R24257 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R24258 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R24259 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R24260 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R24261 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R24262 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R24263 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R24264 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R24265 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R24266 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R24267 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R24268 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R24269 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R24270 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R24271 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R24272 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R24273 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R24274 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R24275 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R24276 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R24277 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R24278 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R24279 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R24280 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R24281 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R24282 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R24283 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R24284 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R24285 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R24286 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R24287 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R24288 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R24289 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R24290 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R24291 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R24292 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R24293 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R24294 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R24295 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R24296 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R24297 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R24298 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R24299 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R24300 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R24301 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R24302 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R24303 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R24304 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R24305 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R24306 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R24307 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R24308 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R24309 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R24310 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R24311 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R24312 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R24313 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R24314 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R24315 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R24316 XThR.Tn[7].n6 XThR.Tn[7] 0.829611
R24317 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R24318 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R24319 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R24320 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R24321 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R24322 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R24323 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R24324 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R24325 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R24326 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R24327 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R24328 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R24329 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R24330 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R24331 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R24332 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R24333 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R24334 XThR.Tn[7] XThR.Tn[7].n84 0.038
R24335 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R24336 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R24337 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R24338 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R24339 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R24340 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R24341 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R24342 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R24343 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R24344 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R24345 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R24346 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R24347 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R24348 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R24349 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R24350 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R24351 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R24352 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R24353 XThR.Tn[0] XThR.Tn[0].n82 161.363
R24354 XThR.Tn[0] XThR.Tn[0].n77 161.363
R24355 XThR.Tn[0] XThR.Tn[0].n72 161.363
R24356 XThR.Tn[0] XThR.Tn[0].n67 161.363
R24357 XThR.Tn[0] XThR.Tn[0].n62 161.363
R24358 XThR.Tn[0] XThR.Tn[0].n57 161.363
R24359 XThR.Tn[0] XThR.Tn[0].n52 161.363
R24360 XThR.Tn[0] XThR.Tn[0].n47 161.363
R24361 XThR.Tn[0] XThR.Tn[0].n42 161.363
R24362 XThR.Tn[0] XThR.Tn[0].n37 161.363
R24363 XThR.Tn[0] XThR.Tn[0].n32 161.363
R24364 XThR.Tn[0] XThR.Tn[0].n27 161.363
R24365 XThR.Tn[0] XThR.Tn[0].n22 161.363
R24366 XThR.Tn[0] XThR.Tn[0].n17 161.363
R24367 XThR.Tn[0] XThR.Tn[0].n12 161.363
R24368 XThR.Tn[0] XThR.Tn[0].n10 161.363
R24369 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R24370 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R24371 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R24372 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R24373 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R24374 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R24375 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R24376 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R24377 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R24378 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R24379 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R24380 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R24381 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R24382 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R24383 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R24384 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R24385 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R24386 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R24387 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R24388 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R24389 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R24390 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R24391 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R24392 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R24393 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R24394 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R24395 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R24396 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R24397 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R24398 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R24399 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R24400 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R24401 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R24402 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R24403 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R24404 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R24405 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R24406 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R24407 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R24408 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R24409 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R24410 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R24411 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R24412 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R24413 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R24414 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R24415 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R24416 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R24417 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R24418 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R24419 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R24420 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R24421 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R24422 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R24423 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R24424 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R24425 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R24426 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R24427 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R24428 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R24429 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R24430 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R24431 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R24432 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R24433 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R24434 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R24435 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R24436 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R24437 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R24438 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R24439 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R24440 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R24441 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R24442 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R24443 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R24444 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R24445 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R24446 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R24447 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R24448 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R24449 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R24450 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R24451 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R24452 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R24453 XThR.Tn[0].n1 XThR.Tn[0].t5 26.5955
R24454 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R24455 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R24456 XThR.Tn[0].n0 XThR.Tn[0].t7 26.5955
R24457 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R24458 XThR.Tn[0].n3 XThR.Tn[0].t10 24.9236
R24459 XThR.Tn[0].n4 XThR.Tn[0].t8 24.9236
R24460 XThR.Tn[0].n4 XThR.Tn[0].t11 24.9236
R24461 XThR.Tn[0].n5 XThR.Tn[0].t3 24.9236
R24462 XThR.Tn[0].n5 XThR.Tn[0].t2 24.9236
R24463 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R24464 XThR.Tn[0].n6 XThR.Tn[0].t1 24.9236
R24465 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R24466 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R24467 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R24468 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R24469 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R24470 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R24471 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R24472 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R24473 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R24474 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R24475 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R24476 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R24477 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R24478 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R24479 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R24480 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R24481 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R24482 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R24483 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R24484 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R24485 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R24486 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R24487 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R24488 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R24489 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R24490 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R24491 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R24492 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R24493 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R24494 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R24495 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R24496 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R24497 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R24498 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R24499 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R24500 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R24501 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R24502 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R24503 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R24504 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R24505 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R24506 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R24507 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R24508 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R24509 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R24510 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R24511 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R24512 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R24513 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R24514 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R24515 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R24516 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R24517 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R24518 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R24519 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R24520 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R24521 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R24522 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R24523 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R24524 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R24525 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R24526 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R24527 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R24528 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R24529 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R24530 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R24531 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R24532 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R24533 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R24534 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R24535 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R24536 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R24537 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R24538 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R24539 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R24540 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R24541 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R24542 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R24543 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R24544 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R24545 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R24546 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R24547 XThR.Tn[0] XThR.Tn[0].n87 0.038
R24548 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R24549 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R24550 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R24551 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R24552 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R24553 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R24554 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R24555 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R24556 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R24557 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R24558 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R24559 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R24560 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R24561 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R24562 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R24563 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R24564 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R24565 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R24566 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R24567 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R24568 XThR.Tn[8].n87 XThR.Tn[8].n85 202.094
R24569 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R24570 XThR.Tn[8] XThR.Tn[8].n78 161.363
R24571 XThR.Tn[8] XThR.Tn[8].n73 161.363
R24572 XThR.Tn[8] XThR.Tn[8].n68 161.363
R24573 XThR.Tn[8] XThR.Tn[8].n63 161.363
R24574 XThR.Tn[8] XThR.Tn[8].n58 161.363
R24575 XThR.Tn[8] XThR.Tn[8].n53 161.363
R24576 XThR.Tn[8] XThR.Tn[8].n48 161.363
R24577 XThR.Tn[8] XThR.Tn[8].n43 161.363
R24578 XThR.Tn[8] XThR.Tn[8].n38 161.363
R24579 XThR.Tn[8] XThR.Tn[8].n33 161.363
R24580 XThR.Tn[8] XThR.Tn[8].n28 161.363
R24581 XThR.Tn[8] XThR.Tn[8].n23 161.363
R24582 XThR.Tn[8] XThR.Tn[8].n18 161.363
R24583 XThR.Tn[8] XThR.Tn[8].n13 161.363
R24584 XThR.Tn[8] XThR.Tn[8].n8 161.363
R24585 XThR.Tn[8] XThR.Tn[8].n6 161.363
R24586 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R24587 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R24588 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R24589 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R24590 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R24591 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R24592 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R24593 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R24594 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R24595 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R24596 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R24597 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R24598 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R24599 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R24600 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R24601 XThR.Tn[8].n78 XThR.Tn[8].t23 161.106
R24602 XThR.Tn[8].n73 XThR.Tn[8].t29 161.106
R24603 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R24604 XThR.Tn[8].n63 XThR.Tn[8].t57 161.106
R24605 XThR.Tn[8].n58 XThR.Tn[8].t21 161.106
R24606 XThR.Tn[8].n53 XThR.Tn[8].t46 161.106
R24607 XThR.Tn[8].n48 XThR.Tn[8].t27 161.106
R24608 XThR.Tn[8].n43 XThR.Tn[8].t69 161.106
R24609 XThR.Tn[8].n38 XThR.Tn[8].t56 161.106
R24610 XThR.Tn[8].n33 XThR.Tn[8].t61 161.106
R24611 XThR.Tn[8].n28 XThR.Tn[8].t44 161.106
R24612 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R24613 XThR.Tn[8].n18 XThR.Tn[8].t43 161.106
R24614 XThR.Tn[8].n13 XThR.Tn[8].t26 161.106
R24615 XThR.Tn[8].n8 XThR.Tn[8].t49 161.106
R24616 XThR.Tn[8].n6 XThR.Tn[8].t33 161.106
R24617 XThR.Tn[8].n79 XThR.Tn[8].t19 159.978
R24618 XThR.Tn[8].n74 XThR.Tn[8].t25 159.978
R24619 XThR.Tn[8].n69 XThR.Tn[8].t67 159.978
R24620 XThR.Tn[8].n64 XThR.Tn[8].t54 159.978
R24621 XThR.Tn[8].n59 XThR.Tn[8].t16 159.978
R24622 XThR.Tn[8].n54 XThR.Tn[8].t42 159.978
R24623 XThR.Tn[8].n49 XThR.Tn[8].t24 159.978
R24624 XThR.Tn[8].n44 XThR.Tn[8].t64 159.978
R24625 XThR.Tn[8].n39 XThR.Tn[8].t51 159.978
R24626 XThR.Tn[8].n34 XThR.Tn[8].t58 159.978
R24627 XThR.Tn[8].n29 XThR.Tn[8].t41 159.978
R24628 XThR.Tn[8].n24 XThR.Tn[8].t66 159.978
R24629 XThR.Tn[8].n19 XThR.Tn[8].t40 159.978
R24630 XThR.Tn[8].n14 XThR.Tn[8].t22 159.978
R24631 XThR.Tn[8].n9 XThR.Tn[8].t45 159.978
R24632 XThR.Tn[8].n78 XThR.Tn[8].t73 145.038
R24633 XThR.Tn[8].n73 XThR.Tn[8].t35 145.038
R24634 XThR.Tn[8].n68 XThR.Tn[8].t15 145.038
R24635 XThR.Tn[8].n63 XThR.Tn[8].t62 145.038
R24636 XThR.Tn[8].n58 XThR.Tn[8].t30 145.038
R24637 XThR.Tn[8].n53 XThR.Tn[8].t72 145.038
R24638 XThR.Tn[8].n48 XThR.Tn[8].t17 145.038
R24639 XThR.Tn[8].n43 XThR.Tn[8].t63 145.038
R24640 XThR.Tn[8].n38 XThR.Tn[8].t60 145.038
R24641 XThR.Tn[8].n33 XThR.Tn[8].t28 145.038
R24642 XThR.Tn[8].n28 XThR.Tn[8].t52 145.038
R24643 XThR.Tn[8].n23 XThR.Tn[8].t12 145.038
R24644 XThR.Tn[8].n18 XThR.Tn[8].t50 145.038
R24645 XThR.Tn[8].n13 XThR.Tn[8].t34 145.038
R24646 XThR.Tn[8].n8 XThR.Tn[8].t59 145.038
R24647 XThR.Tn[8].n6 XThR.Tn[8].t39 145.038
R24648 XThR.Tn[8].n79 XThR.Tn[8].t32 143.911
R24649 XThR.Tn[8].n74 XThR.Tn[8].t55 143.911
R24650 XThR.Tn[8].n69 XThR.Tn[8].t37 143.911
R24651 XThR.Tn[8].n64 XThR.Tn[8].t18 143.911
R24652 XThR.Tn[8].n59 XThR.Tn[8].t48 143.911
R24653 XThR.Tn[8].n54 XThR.Tn[8].t31 143.911
R24654 XThR.Tn[8].n49 XThR.Tn[8].t38 143.911
R24655 XThR.Tn[8].n44 XThR.Tn[8].t20 143.911
R24656 XThR.Tn[8].n39 XThR.Tn[8].t14 143.911
R24657 XThR.Tn[8].n34 XThR.Tn[8].t47 143.911
R24658 XThR.Tn[8].n29 XThR.Tn[8].t68 143.911
R24659 XThR.Tn[8].n24 XThR.Tn[8].t36 143.911
R24660 XThR.Tn[8].n19 XThR.Tn[8].t65 143.911
R24661 XThR.Tn[8].n14 XThR.Tn[8].t53 143.911
R24662 XThR.Tn[8].n9 XThR.Tn[8].t13 143.911
R24663 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R24664 XThR.Tn[8].n86 XThR.Tn[8].t5 26.5955
R24665 XThR.Tn[8].n86 XThR.Tn[8].t7 26.5955
R24666 XThR.Tn[8].n0 XThR.Tn[8].t10 26.5955
R24667 XThR.Tn[8].n0 XThR.Tn[8].t8 26.5955
R24668 XThR.Tn[8].n1 XThR.Tn[8].t11 26.5955
R24669 XThR.Tn[8].n1 XThR.Tn[8].t9 26.5955
R24670 XThR.Tn[8].n85 XThR.Tn[8].t6 26.5955
R24671 XThR.Tn[8].n85 XThR.Tn[8].t0 26.5955
R24672 XThR.Tn[8].n4 XThR.Tn[8].t2 24.9236
R24673 XThR.Tn[8].n4 XThR.Tn[8].t4 24.9236
R24674 XThR.Tn[8].n3 XThR.Tn[8].t1 24.9236
R24675 XThR.Tn[8].n3 XThR.Tn[8].t3 24.9236
R24676 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R24677 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R24678 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R24679 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R24680 XThR.Tn[8] XThR.Tn[8].n7 5.34038
R24681 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R24682 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R24683 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R24684 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R24685 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R24686 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R24687 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R24688 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R24689 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R24690 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R24691 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R24692 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R24693 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R24694 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R24695 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R24696 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R24697 XThR.Tn[8].n12 XThR.Tn[8] 2.52282
R24698 XThR.Tn[8].n17 XThR.Tn[8] 2.52282
R24699 XThR.Tn[8].n22 XThR.Tn[8] 2.52282
R24700 XThR.Tn[8].n27 XThR.Tn[8] 2.52282
R24701 XThR.Tn[8].n32 XThR.Tn[8] 2.52282
R24702 XThR.Tn[8].n37 XThR.Tn[8] 2.52282
R24703 XThR.Tn[8].n42 XThR.Tn[8] 2.52282
R24704 XThR.Tn[8].n47 XThR.Tn[8] 2.52282
R24705 XThR.Tn[8].n52 XThR.Tn[8] 2.52282
R24706 XThR.Tn[8].n57 XThR.Tn[8] 2.52282
R24707 XThR.Tn[8].n62 XThR.Tn[8] 2.52282
R24708 XThR.Tn[8].n67 XThR.Tn[8] 2.52282
R24709 XThR.Tn[8].n72 XThR.Tn[8] 2.52282
R24710 XThR.Tn[8].n77 XThR.Tn[8] 2.52282
R24711 XThR.Tn[8].n82 XThR.Tn[8] 2.52282
R24712 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R24713 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R24714 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R24715 XThR.Tn[8].n80 XThR.Tn[8] 1.08677
R24716 XThR.Tn[8].n75 XThR.Tn[8] 1.08677
R24717 XThR.Tn[8].n70 XThR.Tn[8] 1.08677
R24718 XThR.Tn[8].n65 XThR.Tn[8] 1.08677
R24719 XThR.Tn[8].n60 XThR.Tn[8] 1.08677
R24720 XThR.Tn[8].n55 XThR.Tn[8] 1.08677
R24721 XThR.Tn[8].n50 XThR.Tn[8] 1.08677
R24722 XThR.Tn[8].n45 XThR.Tn[8] 1.08677
R24723 XThR.Tn[8].n40 XThR.Tn[8] 1.08677
R24724 XThR.Tn[8].n35 XThR.Tn[8] 1.08677
R24725 XThR.Tn[8].n30 XThR.Tn[8] 1.08677
R24726 XThR.Tn[8].n25 XThR.Tn[8] 1.08677
R24727 XThR.Tn[8].n20 XThR.Tn[8] 1.08677
R24728 XThR.Tn[8].n15 XThR.Tn[8] 1.08677
R24729 XThR.Tn[8].n10 XThR.Tn[8] 1.08677
R24730 XThR.Tn[8] XThR.Tn[8].n12 0.839786
R24731 XThR.Tn[8] XThR.Tn[8].n17 0.839786
R24732 XThR.Tn[8] XThR.Tn[8].n22 0.839786
R24733 XThR.Tn[8] XThR.Tn[8].n27 0.839786
R24734 XThR.Tn[8] XThR.Tn[8].n32 0.839786
R24735 XThR.Tn[8] XThR.Tn[8].n37 0.839786
R24736 XThR.Tn[8] XThR.Tn[8].n42 0.839786
R24737 XThR.Tn[8] XThR.Tn[8].n47 0.839786
R24738 XThR.Tn[8] XThR.Tn[8].n52 0.839786
R24739 XThR.Tn[8] XThR.Tn[8].n57 0.839786
R24740 XThR.Tn[8] XThR.Tn[8].n62 0.839786
R24741 XThR.Tn[8] XThR.Tn[8].n67 0.839786
R24742 XThR.Tn[8] XThR.Tn[8].n72 0.839786
R24743 XThR.Tn[8] XThR.Tn[8].n77 0.839786
R24744 XThR.Tn[8] XThR.Tn[8].n82 0.839786
R24745 XThR.Tn[8].n7 XThR.Tn[8] 0.499542
R24746 XThR.Tn[8].n81 XThR.Tn[8] 0.063
R24747 XThR.Tn[8].n76 XThR.Tn[8] 0.063
R24748 XThR.Tn[8].n71 XThR.Tn[8] 0.063
R24749 XThR.Tn[8].n66 XThR.Tn[8] 0.063
R24750 XThR.Tn[8].n61 XThR.Tn[8] 0.063
R24751 XThR.Tn[8].n56 XThR.Tn[8] 0.063
R24752 XThR.Tn[8].n51 XThR.Tn[8] 0.063
R24753 XThR.Tn[8].n46 XThR.Tn[8] 0.063
R24754 XThR.Tn[8].n41 XThR.Tn[8] 0.063
R24755 XThR.Tn[8].n36 XThR.Tn[8] 0.063
R24756 XThR.Tn[8].n31 XThR.Tn[8] 0.063
R24757 XThR.Tn[8].n26 XThR.Tn[8] 0.063
R24758 XThR.Tn[8].n21 XThR.Tn[8] 0.063
R24759 XThR.Tn[8].n16 XThR.Tn[8] 0.063
R24760 XThR.Tn[8].n11 XThR.Tn[8] 0.063
R24761 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R24762 XThR.Tn[8] XThR.Tn[8].n83 0.038
R24763 XThR.Tn[8].n7 XThR.Tn[8] 0.0143889
R24764 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00771154
R24765 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00771154
R24766 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00771154
R24767 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00771154
R24768 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00771154
R24769 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00771154
R24770 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00771154
R24771 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00771154
R24772 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00771154
R24773 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00771154
R24774 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00771154
R24775 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00771154
R24776 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00771154
R24777 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00771154
R24778 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00771154
R24779 XThC.TB3.n6 XThC.TB3.t3 212.081
R24780 XThC.TB3.n5 XThC.TB3.t15 212.081
R24781 XThC.TB3.n11 XThC.TB3.t14 212.081
R24782 XThC.TB3.n3 XThC.TB3.t10 212.081
R24783 XThC.TB3.n15 XThC.TB3.t11 212.081
R24784 XThC.TB3.n16 XThC.TB3.t12 212.081
R24785 XThC.TB3.n18 XThC.TB3.t4 212.081
R24786 XThC.TB3.n14 XThC.TB3.t16 212.081
R24787 XThC.TB3.n22 XThC.TB3.n2 201.288
R24788 XThC.TB3.n8 XThC.TB3.n7 173.761
R24789 XThC.TB3.n17 XThC.TB3 158.656
R24790 XThC.TB3.n10 XThC.TB3.n9 152
R24791 XThC.TB3.n8 XThC.TB3.n4 152
R24792 XThC.TB3.n13 XThC.TB3.n12 152
R24793 XThC.TB3.n20 XThC.TB3.n19 152
R24794 XThC.TB3.n6 XThC.TB3.t9 139.78
R24795 XThC.TB3.n5 XThC.TB3.t6 139.78
R24796 XThC.TB3.n11 XThC.TB3.t5 139.78
R24797 XThC.TB3.n3 XThC.TB3.t17 139.78
R24798 XThC.TB3.n15 XThC.TB3.t8 139.78
R24799 XThC.TB3.n16 XThC.TB3.t18 139.78
R24800 XThC.TB3.n18 XThC.TB3.t13 139.78
R24801 XThC.TB3.n14 XThC.TB3.t7 139.78
R24802 XThC.TB3.n0 XThC.TB3.t1 132.067
R24803 XThC.TB3.n21 XThC.TB3.n13 61.4096
R24804 XThC.TB3.n16 XThC.TB3.n15 61.346
R24805 XThC.TB3.n10 XThC.TB3.n4 49.6611
R24806 XThC.TB3.n12 XThC.TB3.n11 45.2793
R24807 XThC.TB3.n7 XThC.TB3.n5 42.3581
R24808 XThC.TB3.n19 XThC.TB3.n14 30.6732
R24809 XThC.TB3.n19 XThC.TB3.n18 30.6732
R24810 XThC.TB3.n18 XThC.TB3.n17 30.6732
R24811 XThC.TB3.n17 XThC.TB3.n16 30.6732
R24812 XThC.TB3.n2 XThC.TB3.t2 26.5955
R24813 XThC.TB3.n2 XThC.TB3.t0 26.5955
R24814 XThC.TB3 XThC.TB3.n22 23.489
R24815 XThC.TB3.n9 XThC.TB3.n8 21.7605
R24816 XThC.TB3.n7 XThC.TB3.n6 18.9884
R24817 XThC.TB3.n12 XThC.TB3.n3 16.0672
R24818 XThC.TB3.n20 XThC.TB3 14.8485
R24819 XThC.TB3.n13 XThC.TB3 11.5205
R24820 XThC.TB3.n22 XThC.TB3.n21 10.8207
R24821 XThC.TB3.n9 XThC.TB3 10.2405
R24822 XThC.TB3 XThC.TB3.n20 8.7045
R24823 XThC.TB3.n5 XThC.TB3.n4 7.30353
R24824 XThC.TB3.n21 XThC.TB3 5.33013
R24825 XThC.TB3.n11 XThC.TB3.n10 4.38232
R24826 XThC.TB3.n1 XThC.TB3.n0 4.15748
R24827 XThC.TB3 XThC.TB3.n1 3.76521
R24828 XThC.TB3.n0 XThC.TB3 1.17559
R24829 XThC.TB3.n1 XThC.TB3 0.921363
R24830 data[4].n3 data[4].t0 231.835
R24831 data[4].n0 data[4].t3 230.155
R24832 data[4].n0 data[4].t1 157.856
R24833 data[4].n3 data[4].t2 157.07
R24834 data[4].n1 data[4].n0 152
R24835 data[4].n4 data[4].n3 152
R24836 data[4].n2 data[4].n1 25.6681
R24837 data[4].n4 data[4].n2 10.7642
R24838 data[4].n2 data[4] 2.763
R24839 data[4].n1 data[4] 2.10199
R24840 data[4] data[4].n4 2.01193
R24841 XThR.Tn[13].n87 XThR.Tn[13].n86 256.103
R24842 XThR.Tn[13].n2 XThR.Tn[13].n0 243.68
R24843 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R24844 XThR.Tn[13].n2 XThR.Tn[13].n1 205.28
R24845 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R24846 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R24847 XThR.Tn[13] XThR.Tn[13].n78 161.363
R24848 XThR.Tn[13] XThR.Tn[13].n73 161.363
R24849 XThR.Tn[13] XThR.Tn[13].n68 161.363
R24850 XThR.Tn[13] XThR.Tn[13].n63 161.363
R24851 XThR.Tn[13] XThR.Tn[13].n58 161.363
R24852 XThR.Tn[13] XThR.Tn[13].n53 161.363
R24853 XThR.Tn[13] XThR.Tn[13].n48 161.363
R24854 XThR.Tn[13] XThR.Tn[13].n43 161.363
R24855 XThR.Tn[13] XThR.Tn[13].n38 161.363
R24856 XThR.Tn[13] XThR.Tn[13].n33 161.363
R24857 XThR.Tn[13] XThR.Tn[13].n28 161.363
R24858 XThR.Tn[13] XThR.Tn[13].n23 161.363
R24859 XThR.Tn[13] XThR.Tn[13].n18 161.363
R24860 XThR.Tn[13] XThR.Tn[13].n13 161.363
R24861 XThR.Tn[13] XThR.Tn[13].n8 161.363
R24862 XThR.Tn[13] XThR.Tn[13].n6 161.363
R24863 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R24864 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R24865 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R24866 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R24867 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R24868 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R24869 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R24870 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R24871 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R24872 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R24873 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R24874 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R24875 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R24876 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R24877 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R24878 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R24879 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R24880 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R24881 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R24882 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R24883 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R24884 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R24885 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R24886 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R24887 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R24888 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R24889 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R24890 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R24891 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R24892 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R24893 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R24894 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R24895 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R24896 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R24897 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R24898 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R24899 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R24900 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R24901 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R24902 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R24903 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R24904 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R24905 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R24906 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R24907 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R24908 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R24909 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R24910 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R24911 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R24912 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R24913 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R24914 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R24915 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R24916 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R24917 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R24918 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R24919 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R24920 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R24921 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R24922 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R24923 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R24924 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R24925 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R24926 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R24927 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R24928 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R24929 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R24930 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R24931 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R24932 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R24933 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R24934 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R24935 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R24936 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R24937 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R24938 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R24939 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R24940 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R24941 XThR.Tn[13].n85 XThR.Tn[13].t2 26.5955
R24942 XThR.Tn[13].n85 XThR.Tn[13].t0 26.5955
R24943 XThR.Tn[13].n0 XThR.Tn[13].t9 26.5955
R24944 XThR.Tn[13].n0 XThR.Tn[13].t11 26.5955
R24945 XThR.Tn[13].n1 XThR.Tn[13].t10 26.5955
R24946 XThR.Tn[13].n1 XThR.Tn[13].t8 26.5955
R24947 XThR.Tn[13].n86 XThR.Tn[13].t3 26.5955
R24948 XThR.Tn[13].n86 XThR.Tn[13].t1 26.5955
R24949 XThR.Tn[13].n4 XThR.Tn[13].t6 24.9236
R24950 XThR.Tn[13].n4 XThR.Tn[13].t4 24.9236
R24951 XThR.Tn[13].n3 XThR.Tn[13].t7 24.9236
R24952 XThR.Tn[13].n3 XThR.Tn[13].t5 24.9236
R24953 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R24954 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R24955 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R24956 XThR.Tn[13] XThR.Tn[13].n7 5.34038
R24957 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R24958 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R24959 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R24960 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R24961 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R24962 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R24963 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R24964 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R24965 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R24966 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R24967 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R24968 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R24969 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R24970 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R24971 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R24972 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R24973 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R24974 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R24975 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R24976 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R24977 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R24978 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R24979 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R24980 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R24981 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R24982 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R24983 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R24984 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R24985 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R24986 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R24987 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R24988 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R24989 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R24990 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R24991 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R24992 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R24993 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R24994 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R24995 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R24996 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R24997 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R24998 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R24999 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R25000 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R25001 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R25002 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R25003 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R25004 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R25005 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R25006 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R25007 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R25008 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R25009 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R25010 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R25011 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R25012 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R25013 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R25014 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R25015 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R25016 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R25017 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R25018 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R25019 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R25020 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R25021 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R25022 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R25023 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R25024 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R25025 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R25026 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R25027 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R25028 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R25029 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R25030 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R25031 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R25032 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R25033 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R25034 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R25035 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R25036 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R25037 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R25038 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R25039 XThR.Tn[13] XThR.Tn[13].n83 0.038
R25040 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R25041 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R25042 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R25043 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R25044 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R25045 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R25046 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R25047 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R25048 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R25049 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R25050 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R25051 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R25052 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R25053 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R25054 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R25055 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R25056 data[0].n1 data[0].t0 230.155
R25057 data[0].n0 data[0].t2 228.463
R25058 data[0].n1 data[0].t1 157.856
R25059 data[0].n0 data[0].t3 157.07
R25060 data[0].n2 data[0].n1 152.768
R25061 data[0].n4 data[0].n0 152.256
R25062 data[0].n3 data[0].n2 24.1398
R25063 data[0].n4 data[0].n3 9.48418
R25064 data[0] data[0].n4 6.1445
R25065 data[0].n2 data[0] 5.6325
R25066 data[0].n3 data[0] 2.638
R25067 XThR.TB1.n9 XThR.TB1.t12 212.081
R25068 XThR.TB1.n10 XThR.TB1.t17 212.081
R25069 XThR.TB1.n15 XThR.TB1.t6 212.081
R25070 XThR.TB1.n16 XThR.TB1.t3 212.081
R25071 XThR.TB1.n1 XThR.TB1.t10 212.081
R25072 XThR.TB1.n2 XThR.TB1.t14 212.081
R25073 XThR.TB1.n4 XThR.TB1.t8 212.081
R25074 XThR.TB1.n5 XThR.TB1.t13 212.081
R25075 XThR.TB1.n21 XThR.TB1.n20 201.288
R25076 XThR.TB1.n12 XThR.TB1.n11 173.761
R25077 XThR.TB1.n3 XThR.TB1 167.361
R25078 XThR.TB1.n18 XThR.TB1.n17 152
R25079 XThR.TB1.n14 XThR.TB1.n13 152
R25080 XThR.TB1.n12 XThR.TB1.n8 152
R25081 XThR.TB1.n7 XThR.TB1.n6 152
R25082 XThR.TB1.n9 XThR.TB1.t16 139.78
R25083 XThR.TB1.n10 XThR.TB1.t5 139.78
R25084 XThR.TB1.n15 XThR.TB1.t11 139.78
R25085 XThR.TB1.n16 XThR.TB1.t9 139.78
R25086 XThR.TB1.n1 XThR.TB1.t18 139.78
R25087 XThR.TB1.n2 XThR.TB1.t7 139.78
R25088 XThR.TB1.n4 XThR.TB1.t15 139.78
R25089 XThR.TB1.n5 XThR.TB1.t4 139.78
R25090 XThR.TB1.n0 XThR.TB1.t1 130.548
R25091 XThR.TB1.n19 XThR.TB1.n18 61.4072
R25092 XThR.TB1.n2 XThR.TB1.n1 61.346
R25093 XThR.TB1.n14 XThR.TB1.n8 49.6611
R25094 XThR.TB1.n17 XThR.TB1.n15 45.2793
R25095 XThR.TB1.n11 XThR.TB1.n10 42.3581
R25096 XThR.TB1 XThR.TB1.n21 36.289
R25097 XThR.TB1.n3 XThR.TB1.n2 30.6732
R25098 XThR.TB1.n4 XThR.TB1.n3 30.6732
R25099 XThR.TB1.n6 XThR.TB1.n4 30.6732
R25100 XThR.TB1.n6 XThR.TB1.n5 30.6732
R25101 XThR.TB1.n20 XThR.TB1.t2 26.5955
R25102 XThR.TB1.n20 XThR.TB1.t0 26.5955
R25103 XThR.TB1.n13 XThR.TB1.n12 21.7605
R25104 XThR.TB1.n13 XThR.TB1 21.1205
R25105 XThR.TB1.n11 XThR.TB1.n9 18.9884
R25106 XThR.TB1 XThR.TB1.n7 17.4085
R25107 XThR.TB1.n22 XThR.TB1 16.5652
R25108 XThR.TB1.n17 XThR.TB1.n16 16.0672
R25109 XThR.TB1.n21 XThR.TB1.n19 10.8571
R25110 XThR.TB1 XThR.TB1.n22 9.03579
R25111 XThR.TB1.n19 XThR.TB1 8.65973
R25112 XThR.TB1.n10 XThR.TB1.n8 7.30353
R25113 XThR.TB1.n7 XThR.TB1 6.1445
R25114 XThR.TB1.n15 XThR.TB1.n14 4.38232
R25115 XThR.TB1 XThR.TB1.n0 3.46739
R25116 XThR.TB1.n0 XThR.TB1 2.74112
R25117 XThR.TB1.n22 XThR.TB1 2.21057
R25118 XThR.TB1.n18 XThR.TB1 0.6405
R25119 XThR.TB3.n9 XThR.TB3.t7 212.081
R25120 XThR.TB3.n10 XThR.TB3.t11 212.081
R25121 XThR.TB3.n15 XThR.TB3.t18 212.081
R25122 XThR.TB3.n16 XThR.TB3.t14 212.081
R25123 XThR.TB3.n1 XThR.TB3.t9 212.081
R25124 XThR.TB3.n2 XThR.TB3.t13 212.081
R25125 XThR.TB3.n4 XThR.TB3.t8 212.081
R25126 XThR.TB3.n5 XThR.TB3.t12 212.081
R25127 XThR.TB3.n21 XThR.TB3.n20 201.288
R25128 XThR.TB3.n12 XThR.TB3.n11 173.761
R25129 XThR.TB3.n3 XThR.TB3 167.361
R25130 XThR.TB3.n18 XThR.TB3.n17 152
R25131 XThR.TB3.n14 XThR.TB3.n13 152
R25132 XThR.TB3.n12 XThR.TB3.n8 152
R25133 XThR.TB3.n7 XThR.TB3.n6 152
R25134 XThR.TB3.n9 XThR.TB3.t10 139.78
R25135 XThR.TB3.n10 XThR.TB3.t16 139.78
R25136 XThR.TB3.n15 XThR.TB3.t5 139.78
R25137 XThR.TB3.n16 XThR.TB3.t3 139.78
R25138 XThR.TB3.n1 XThR.TB3.t17 139.78
R25139 XThR.TB3.n2 XThR.TB3.t6 139.78
R25140 XThR.TB3.n4 XThR.TB3.t15 139.78
R25141 XThR.TB3.n5 XThR.TB3.t4 139.78
R25142 XThR.TB3.n0 XThR.TB3.t2 130.548
R25143 XThR.TB3.n19 XThR.TB3.n18 61.4096
R25144 XThR.TB3.n2 XThR.TB3.n1 61.346
R25145 XThR.TB3.n14 XThR.TB3.n8 49.6611
R25146 XThR.TB3.n17 XThR.TB3.n15 45.2793
R25147 XThR.TB3.n11 XThR.TB3.n10 42.3581
R25148 XThR.TB3 XThR.TB3.n21 36.289
R25149 XThR.TB3.n3 XThR.TB3.n2 30.6732
R25150 XThR.TB3.n4 XThR.TB3.n3 30.6732
R25151 XThR.TB3.n6 XThR.TB3.n4 30.6732
R25152 XThR.TB3.n6 XThR.TB3.n5 30.6732
R25153 XThR.TB3.n20 XThR.TB3.t0 26.5955
R25154 XThR.TB3.n20 XThR.TB3.t1 26.5955
R25155 XThR.TB3.n13 XThR.TB3.n12 21.7605
R25156 XThR.TB3.n13 XThR.TB3 21.1205
R25157 XThR.TB3.n11 XThR.TB3.n9 18.9884
R25158 XThR.TB3 XThR.TB3.n7 17.4085
R25159 XThR.TB3.n22 XThR.TB3 16.5652
R25160 XThR.TB3.n17 XThR.TB3.n16 16.0672
R25161 XThR.TB3.n21 XThR.TB3.n19 10.8207
R25162 XThR.TB3 XThR.TB3.n22 9.03579
R25163 XThR.TB3.n10 XThR.TB3.n8 7.30353
R25164 XThR.TB3.n7 XThR.TB3 6.1445
R25165 XThR.TB3.n19 XThR.TB3 5.58292
R25166 XThR.TB3.n15 XThR.TB3.n14 4.38232
R25167 XThR.TB3 XThR.TB3.n0 3.46739
R25168 XThR.TB3.n0 XThR.TB3 2.74112
R25169 XThR.TB3.n22 XThR.TB3 2.21057
R25170 XThR.TB3.n18 XThR.TB3 0.6405
R25171 data[6].n0 data[6].t0 230.576
R25172 data[6].n0 data[6].t1 158.275
R25173 data[6].n1 data[6].n0 152
R25174 data[6].n1 data[6] 11.9995
R25175 data[6] data[6].n1 6.66717
R25176 data[1].n4 data[1].t2 230.576
R25177 data[1].n1 data[1].t0 230.363
R25178 data[1].n0 data[1].t4 229.369
R25179 data[1].n4 data[1].t5 158.275
R25180 data[1].n1 data[1].t3 158.064
R25181 data[1].n0 data[1].t1 157.07
R25182 data[1].n2 data[1].n1 153.28
R25183 data[1].n7 data[1].n0 153.147
R25184 data[1].n5 data[1].n4 152
R25185 data[1].n7 data[1].n6 16.3874
R25186 data[1].n6 data[1].n5 14.9641
R25187 data[1].n3 data[1].n2 9.3005
R25188 data[1].n6 data[1].n3 6.49639
R25189 data[1] data[1].n7 3.24826
R25190 data[1].n2 data[1] 2.92621
R25191 data[1].n3 data[1] 2.15819
R25192 data[1].n5 data[1] 2.13383
R25193 data[2].n0 data[2].t0 230.576
R25194 data[2].n0 data[2].t1 158.275
R25195 data[2].n1 data[2].n0 152
R25196 data[2].n1 data[2] 12.7714
R25197 data[2] data[2].n1 2.13383
R25198 data[5].n4 data[5].t2 230.576
R25199 data[5].n1 data[5].t0 230.363
R25200 data[5].n0 data[5].t1 229.369
R25201 data[5].n4 data[5].t5 158.275
R25202 data[5].n1 data[5].t3 158.064
R25203 data[5].n0 data[5].t4 157.07
R25204 data[5].n2 data[5].n1 152.256
R25205 data[5].n7 data[5].n0 152.238
R25206 data[5].n5 data[5].n4 152
R25207 data[5].n7 data[5].n6 16.3874
R25208 data[5].n6 data[5].n5 14.6005
R25209 data[5].n3 data[5].n2 9.3005
R25210 data[5].n5 data[5] 6.66717
R25211 data[5].n6 data[5].n3 6.49639
R25212 data[5].n2 data[5] 6.1445
R25213 data[5] data[5].n7 5.68939
R25214 data[5].n3 data[5] 2.28319
R25215 data[3].n0 data[3].t1 230.576
R25216 data[3].n0 data[3].t0 158.275
R25217 data[3].n1 data[3].n0 153.553
R25218 data[3].n1 data[3] 11.6078
R25219 data[3] data[3].n1 2.90959
R25220 data[7].n0 data[7].t0 230.576
R25221 data[7].n0 data[7].t1 158.275
R25222 data[7].n1 data[7].n0 152
R25223 data[7].n1 data[7] 11.9995
R25224 data[7] data[7].n1 6.66717
R25225 bias[1] bias[1].t0 23.8076
R25226 bias[2] bias[2].t0 57.7456
R25227 bias[0] bias[0].t0 12.1467
C0 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02762f
C1 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C2 XA.XIR[6].XIC[9].icell.SM VPWR 0.00158f
C3 XA.XIR[7].XIC[10].icell.SM Vbias 0.00701f
C4 XA.XIR[4].XIC[6].icell.PDM VPWR 0.00799f
C5 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C6 XThR.TA2 XThR.TB6 0.10153f
C7 XA.XIR[6].XIC[5].icell.SM Iout 0.00388f
C8 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02762f
C9 XA.XIR[1].XIC[5].icell.PUM VPWR 0.00937f
C10 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7] 0.00341f
C11 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.15202f
C12 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.03425f
C13 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C14 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.SM 0.0039f
C15 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.SM 0.0039f
C16 XA.XIR[13].XIC[11].icell.Ien VPWR 0.1903f
C17 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.SM 0.00168f
C18 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04031f
C19 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.03431f
C20 XThR.Tn[3] VPWR 6.64542f
C21 XThR.Tn[13] XA.XIR[14].XIC[5].icell.Ien 0.00338f
C22 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00214f
C23 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.SM 0.00168f
C24 XThC.TB7 a_7651_9569# 0.00477f
C25 XA.XIR[15].XIC[0].icell.SM VPWR 0.00158f
C26 XA.XIR[2].XIC[14].icell.PDM Iout 0.00117f
C27 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.03023f
C28 XA.XIR[0].XIC[10].icell.Ien Vbias 0.2113f
C29 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.15202f
C30 XThC.Tn[12] XThC.Tn[13] 0.23689f
C31 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.SM 0.00168f
C32 XA.XIR[7].XIC[13].icell.Ien Iout 0.06417f
C33 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.04036f
C34 XA.XIR[5].XIC[0].icell.Ien Iout 0.06411f
C35 XThR.Tn[6] XA.XIR[7].XIC[7].icell.Ien 0.00338f
C36 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C37 XA.XIR[11].XIC[0].icell.SM Vbias 0.00675f
C38 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00584f
C39 XA.XIR[11].XIC[1].icell.PDM VPWR 0.00799f
C40 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C41 XThR.Tn[4] XA.XIR[5].XIC[9].icell.SM 0.00121f
C42 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00584f
C43 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00214f
C44 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Iout 0.00347f
C45 XA.XIR[7].XIC_dummy_right.icell.Ien Vbias 0.00288f
C46 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.03425f
C47 XA.XIR[12].XIC[12].icell.PUM Vbias 0.0031f
C48 XA.XIR[3].XIC_dummy_right.icell.PUM Vbias 0.00223f
C49 XA.XIR[5].XIC[2].icell.Ien Vbias 0.21098f
C50 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Ien 0.00584f
C51 XThR.TB7 a_n997_3979# 0.00477f
C52 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.03425f
C53 XThR.Tn[7] XA.XIR[8].XIC[14].icell.Ien 0.00338f
C54 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00214f
C55 XThR.Tn[3] XA.XIR[4].XIC[11].icell.SM 0.00121f
C56 XA.XIR[10].XIC[5].icell.PDM VPWR 0.00799f
C57 XThR.Tn[13] a_n997_1803# 0.0021f
C58 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04031f
C59 XA.XIR[13].XIC[0].icell.Ien Iout 0.06411f
C60 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5] 0.00341f
C61 XA.XIR[15].XIC[4].icell.PDM Vbias 0.04261f
C62 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.SM 0.00168f
C63 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.SM 0.0039f
C64 XA.XIR[1].XIC[13].icell.PUM Vbias 0.0031f
C65 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.SM 0.00168f
C66 a_7651_9569# VPWR 0.00385f
C67 XA.XIR[14].XIC[10].icell.PDM Vbias 0.04261f
C68 XA.XIR[15].XIC[5].icell.SM VPWR 0.00158f
C69 XA.XIR[5].XIC[9].icell.PUM VPWR 0.00937f
C70 XA.XIR[15].XIC[13].icell.SM Vbias 0.00701f
C71 XA.XIR[3].XIC[3].icell.PDM VPWR 0.00799f
C72 XA.XIR[12].XIC[11].icell.PDM VPWR 0.00799f
C73 XThC.TB6 XThC.Tn[13] 0.32552f
C74 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PUM 0.00465f
C75 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.SM 0.0039f
C76 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38993f
C77 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00584f
C78 XA.XIR[15].XIC[1].icell.SM Iout 0.00388f
C79 XA.XIR[9].XIC[2].icell.PDM Vbias 0.04261f
C80 XThC.TB5 a_8739_9569# 0.00424f
C81 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C82 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00584f
C83 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.15202f
C84 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C85 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6] 0.00341f
C86 XA.XIR[15].XIC[12].icell.PDM VPWR 0.0114f
C87 XThR.TB3 XThR.Tn[5] 0.00381f
C88 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00214f
C89 XA.XIR[9].XIC[6].icell.PUM Vbias 0.0031f
C90 XA.XIR[12].XIC[13].icell.Ien Vbias 0.21098f
C91 XA.XIR[1].XIC[14].icell.SM Iout 0.00388f
C92 XA.XIR[8].XIC[2].icell.SM VPWR 0.00158f
C93 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02823f
C94 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C95 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00584f
C96 XThR.Tn[13] XA.XIR[14].XIC[0].icell.Ien 0.0037f
C97 XThC.TAN XThC.Tn[6] 0.05039f
C98 XThR.TA2 XThR.Tn[1] 0.00411f
C99 XA.XIR[11].XIC[3].icell.Ien VPWR 0.1903f
C100 XA.XIR[9].XIC[9].icell.PDM Iout 0.00117f
C101 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.SM 0.0039f
C102 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.SM 0.00168f
C103 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9] 0.00341f
C104 XA.XIR[2].XIC[4].icell.SM Vbias 0.00701f
C105 XA.XIR[9].XIC[11].icell.SM VPWR 0.00158f
C106 XA.XIR[10].XIC[5].icell.Ien VPWR 0.1903f
C107 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02762f
C108 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11] 0.00341f
C109 XThR.TB7 XThR.Tn[7] 0.0835f
C110 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.15202f
C111 XThR.TB7 a_n997_2891# 0.00474f
C112 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C113 XThR.Tn[2] XA.XIR[2].XIC[7].icell.PDM 0.00341f
C114 XA.XIR[5].XIC_15.icell.PDM Vbias 0.04401f
C115 XThR.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.00338f
C116 XA.XIR[9].XIC[7].icell.SM Iout 0.00388f
C117 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02762f
C118 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.SM 0.0039f
C119 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04031f
C120 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02762f
C121 XA.XIR[0].XIC[7].icell.PDM Vbias 0.04278f
C122 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Ien 0.00232f
C123 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00214f
C124 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04031f
C125 XA.XIR[7].XIC[14].icell.PDM VPWR 0.00809f
C126 XThR.Tn[0] XA.XIR[1].XIC[12].icell.SM 0.00121f
C127 XThR.Tn[0] XThR.Tn[1] 0.22353f
C128 XA.XIR[4].XIC[7].icell.Ien VPWR 0.1903f
C129 XA.XIR[14].XIC[6].icell.Ien Vbias 0.21098f
C130 XThC.TB4 XThC.TAN 0.33064f
C131 XA.XIR[2].XIC[11].icell.Ien VPWR 0.1903f
C132 XA.XIR[7].XIC[2].icell.PDM Iout 0.00117f
C133 XThC.TA3 XThC.TB5 0.11935f
C134 XA.XIR[12].XIC[14].icell.SM Vbias 0.00701f
C135 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.SM 0.00168f
C136 XA.XIR[13].XIC[8].icell.Ien Vbias 0.21098f
C137 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C138 XThC.TB1 XThC.TB5 0.05054f
C139 XA.XIR[4].XIC[3].icell.Ien Iout 0.06417f
C140 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.SM 0.00168f
C141 XA.XIR[10].XIC[14].icell.PDM Iout 0.00117f
C142 XA.XIR[8].XIC[10].icell.SM Vbias 0.00701f
C143 XA.XIR[7].XIC[7].icell.SM VPWR 0.00158f
C144 XA.XIR[10].XIC_15.icell.SM VPWR 0.00275f
C145 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.SM 0.0039f
C146 XA.XIR[2].XIC[7].icell.Ien Iout 0.06417f
C147 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04052f
C148 XThC.TB5 XThC.Tn[11] 0.02206f
C149 XA.XIR[12].XIC[10].icell.PUM Vbias 0.0031f
C150 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00214f
C151 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.SM 0.0039f
C152 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C153 XA.XIR[7].XIC[3].icell.SM Iout 0.00388f
C154 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.SM 0.00168f
C155 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.15202f
C156 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C157 XThC.Tn[9] XThR.Tn[5] 0.28739f
C158 XA.XIR[1].XIC[14].icell.PDM Vbias 0.04261f
C159 XThC.Tn[0] XA.XIR[7].XIC_dummy_left.icell.Iout 0.00109f
C160 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.03425f
C161 XA.XIR[3].XIC[0].icell.SM VPWR 0.00158f
C162 XA.XIR[13].XIC_15.icell.PDM Iout 0.00133f
C163 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02762f
C164 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.03425f
C165 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.SM 0.00168f
C166 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.SM 0.0039f
C167 XA.XIR[3].XIC[6].icell.Ien Vbias 0.21098f
C168 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02762f
C169 XThR.Tn[7] XA.XIR[8].XIC[4].icell.SM 0.00121f
C170 XA.XIR[9].XIC[1].icell.PUM Vbias 0.0031f
C171 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.SM 0.0039f
C172 XA.XIR[6].XIC[9].icell.PUM Vbias 0.0031f
C173 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02762f
C174 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18965f
C175 a_n1049_6699# XThR.TB5 0.0021f
C176 XA.XIR[8].XIC[13].icell.Ien Iout 0.06417f
C177 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PUM 0.00465f
C178 a_10915_9569# XThC.Tn[13] 0.01061f
C179 XThC.TA3 a_4067_9615# 0.0127f
C180 XThR.Tn[8] XA.XIR[9].XIC[13].icell.Ien 0.00338f
C181 XThR.Tn[11] XA.XIR[12].XIC[2].icell.Ien 0.00338f
C182 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.15202f
C183 XA.XIR[15].XIC[11].icell.SM Vbias 0.00701f
C184 XA.XIR[4].XIC[2].icell.PDM Vbias 0.04261f
C185 XA.XIR[7].XIC[0].icell.PUM VPWR 0.00937f
C186 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.SM 0.00168f
C187 XA.XIR[0].XIC[3].icell.Ien Iout 0.06389f
C188 XA.XIR[1].XIC[3].icell.Ien Vbias 0.21104f
C189 XA.XIR[8].XIC_dummy_right.icell.Ien Vbias 0.00288f
C190 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.PDM 0.00591f
C191 XA.XIR[3].XIC[13].icell.PUM VPWR 0.00937f
C192 XA.XIR[4].XIC_15.icell.Ien Vbias 0.21234f
C193 a_n1049_5317# VPWR 0.72036f
C194 XThR.Tn[1] a_n1049_7493# 0.00444f
C195 XThR.Tn[10] XA.XIR[11].XIC[5].icell.SM 0.00121f
C196 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00214f
C197 XThR.Tn[0] XA.XIR[0].XIC[8].icell.PDM 0.00341f
C198 XA.XIR[6].XIC[10].icell.PDM VPWR 0.00799f
C199 XA.XIR[6].XIC[14].icell.SM VPWR 0.00207f
C200 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.03547f
C201 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C202 XA.XIR[12].XIC[11].icell.Ien Vbias 0.21098f
C203 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.SM 0.0039f
C204 XA.XIR[6].XIC[10].icell.SM Iout 0.00388f
C205 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00584f
C206 XThR.TB4 a_n1049_6405# 0.01546f
C207 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PUM 0.00465f
C208 XA.XIR[1].XIC[10].icell.PUM VPWR 0.00937f
C209 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.15202f
C210 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C211 XThR.TA2 a_n997_3755# 0.00149f
C212 XA.XIR[4].XIC[9].icell.PDM Iout 0.00117f
C213 XThC.Tn[11] XThR.Tn[11] 0.28739f
C214 XA.XIR[14].XIC[1].icell.PDM VPWR 0.00799f
C215 XA.XIR[14].XIC[0].icell.SM Vbias 0.00675f
C216 XThR.TB5 XThR.Tn[9] 0.01732f
C217 XThR.TBN XThR.Tn[4] 0.60351f
C218 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00584f
C219 XA.XIR[13].XIC[5].icell.PDM VPWR 0.00799f
C220 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.03425f
C221 XThC.Tn[1] XThR.Tn[7] 0.28739f
C222 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C223 XThC.Tn[9] Vbias 2.3038f
C224 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00584f
C225 XA.XIR[10].XIC[1].icell.PDM Vbias 0.04261f
C226 XA.XIR[0].XIC_15.icell.Ien Vbias 0.21286f
C227 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.SM 0.0039f
C228 XA.XIR[15].XIC[14].icell.PUM Vbias 0.0031f
C229 XA.XIR[12].XIC[10].icell.PDM VPWR 0.00799f
C230 XThC.TBN Vbias 0.16617f
C231 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PDM 0.00172f
C232 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C233 XThR.Tn[6] XA.XIR[7].XIC[12].icell.Ien 0.00338f
C234 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00214f
C235 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.SM 0.00168f
C236 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.0353f
C237 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04031f
C238 XThC.Tn[10] XThR.Tn[6] 0.28739f
C239 XA.XIR[9].XIC[3].icell.PUM VPWR 0.00937f
C240 XThR.Tn[4] XA.XIR[5].XIC[14].icell.SM 0.00121f
C241 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PUM 0.00465f
C242 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04031f
C243 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PUM 0.00465f
C244 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C245 XA.XIR[15].XIC[11].icell.PDM VPWR 0.0114f
C246 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[9].icell.SM 0.0039f
C247 XA.XIR[5].XIC[7].icell.Ien Vbias 0.21098f
C248 XA.XIR[15].XIC[5].icell.PUM Vbias 0.0031f
C249 XA.XIR[11].XIC[4].icell.PDM Iout 0.00117f
C250 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.SM 0.0039f
C251 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04031f
C252 a_n1049_7787# XThR.Tn[2] 0.00158f
C253 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PUM 0.00465f
C254 XThC.TA3 XThC.Tn[3] 0.03065f
C255 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00584f
C256 XThR.TBN XThR.TB6 0.1894f
C257 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.SM 0.00168f
C258 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.03425f
C259 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.03425f
C260 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.SM 0.00168f
C261 XA.XIR[10].XIC[8].icell.PDM Iout 0.00117f
C262 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04031f
C263 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.03425f
C264 XA.XIR[2].XIC[1].icell.SM VPWR 0.00158f
C265 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02762f
C266 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.SM 0.0039f
C267 XThC.TBN XThC.Tn[5] 0.60785f
C268 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.SM 0.00168f
C269 XA.XIR[5].XIC[14].icell.PUM VPWR 0.00937f
C270 a_4861_9615# XThC.Tn[4] 0.00198f
C271 XA.XIR[5].XIC[6].icell.PDM VPWR 0.00799f
C272 XThC.Tn[14] XThR.Tn[12] 0.28745f
C273 XA.XIR[4].XIC[0].icell.SM Vbias 0.00675f
C274 XThR.TB4 data[6] 0.0086f
C275 XThR.Tn[10] a_n997_2891# 0.1927f
C276 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00584f
C277 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00584f
C278 XA.XIR[15].XIC[6].icell.SM Iout 0.00388f
C279 XA.XIR[6].XIC[1].icell.PUM VPWR 0.00937f
C280 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.SM 0.00168f
C281 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00214f
C282 XA.XIR[8].XIC[8].icell.PDM VPWR 0.00799f
C283 XA.XIR[3].XIC[6].icell.PDM Iout 0.00117f
C284 XA.XIR[14].XIC[3].icell.Ien VPWR 0.19084f
C285 XThC.TB3 a_5949_9615# 0.009f
C286 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PUM 0.00465f
C287 XThR.TB3 XThR.Tn[2] 0.18254f
C288 XA.XIR[7].XIC[2].icell.PUM Vbias 0.0031f
C289 XThC.TA2 XThC.Tn[9] 0.00838f
C290 XA.XIR[11].XIC[1].icell.SM Vbias 0.00701f
C291 XA.XIR[15].XIC[9].icell.SM Vbias 0.00701f
C292 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C293 XA.XIR[13].XIC[5].icell.Ien VPWR 0.1903f
C294 XThC.TA2 XThC.TBN 0.03867f
C295 XA.XIR[9].XIC[11].icell.PUM Vbias 0.0031f
C296 XThC.TB4 XThC.Tn[8] 0.01306f
C297 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04031f
C298 XThR.TB7 a_n997_1579# 0.013f
C299 XA.XIR[10].XIC[3].icell.SM Vbias 0.00701f
C300 XA.XIR[8].XIC[7].icell.SM VPWR 0.00158f
C301 XThR.Tn[2] XA.XIR[3].XIC[6].icell.Ien 0.00338f
C302 XThC.TA1 XThC.TBN 0.00282f
C303 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PUM 0.00465f
C304 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PUM 0.00465f
C305 XA.XIR[12].XIC[7].icell.PUM VPWR 0.00937f
C306 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00584f
C307 XA.XIR[8].XIC[3].icell.SM Iout 0.00388f
C308 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12] 0.00341f
C309 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PUM 0.00465f
C310 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00584f
C311 XThR.Tn[8] XA.XIR[9].XIC[3].icell.SM 0.00121f
C312 XA.XIR[10].XIC[13].icell.PDM Iout 0.00117f
C313 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C314 XThC.Tn[0] XA.XIR[8].XIC_dummy_left.icell.Iout 0.00109f
C315 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.04036f
C316 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C317 XThR.Tn[3] XA.XIR[3].XIC[4].icell.PDM 0.00341f
C318 XThR.TAN XThR.TB5 0.30227f
C319 XA.XIR[7].XIC[10].icell.PDM Vbias 0.04261f
C320 XA.XIR[11].XIC[8].icell.Ien VPWR 0.1903f
C321 XThC.Tn[13] XThR.Tn[10] 0.2874f
C322 XThR.TBN XThR.Tn[8] 0.47811f
C323 XA.XIR[1].XIC[5].icell.PDM VPWR 0.00799f
C324 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PUM 0.00465f
C325 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.SM 0.00168f
C326 XA.XIR[0].XIC[0].icell.SM Vbias 0.00691f
C327 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.SM 0.0039f
C328 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04031f
C329 XA.XIR[3].XIC[3].icell.Ien VPWR 0.1903f
C330 XA.XIR[4].XIC[5].icell.SM Vbias 0.00701f
C331 XA.XIR[11].XIC[4].icell.Ien Iout 0.06417f
C332 XA.XIR[2].XIC[9].icell.SM Vbias 0.00701f
C333 XThC.Tn[2] XA.XIR[0].XIC[4].icell.Ien 0.00191f
C334 XA.XIR[13].XIC[14].icell.PDM Iout 0.00117f
C335 XA.XIR[6].XIC[6].icell.PUM VPWR 0.00937f
C336 XA.XIR[13].XIC_15.icell.SM VPWR 0.00275f
C337 XA.XIR[9].XIC[12].icell.SM Iout 0.00388f
C338 XThC.TB7 a_5949_9615# 0.00153f
C339 XA.XIR[7].XIC[7].icell.PUM Vbias 0.0031f
C340 XA.XIR[10].XIC[6].icell.Ien Iout 0.06417f
C341 XThR.Tn[9] XA.XIR[10].XIC[6].icell.Ien 0.00338f
C342 XThC.TBN a_10051_9569# 0.23006f
C343 XA.XIR[9].XIC_15.icell.SM Vbias 0.00701f
C344 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00584f
C345 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02762f
C346 XA.XIR[4].XIC[12].icell.Ien VPWR 0.1903f
C347 XA.XIR[15].XIC[12].icell.PUM Vbias 0.0031f
C348 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.389f
C349 XA.XIR[2].XIC[13].icell.PDM VPWR 0.00799f
C350 XA.XIR[4].XIC[8].icell.Ien Iout 0.06417f
C351 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8] 0.00341f
C352 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C353 XThR.TBN XThR.Tn[1] 0.61094f
C354 XA.XIR[7].XIC[12].icell.SM VPWR 0.00158f
C355 XThC.Tn[9] XThR.Tn[2] 0.28739f
C356 XA.XIR[2].XIC[1].icell.PDM Iout 0.00117f
C357 XA.XIR[2].XIC[12].icell.Ien Iout 0.06417f
C358 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00214f
C359 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PUM 0.00465f
C360 XThR.TB6 a_n1049_5611# 0.26831f
C361 XA.XIR[0].XIC[5].icell.SM Vbias 0.00716f
C362 XA.XIR[10].XIC[0].icell.PUM VPWR 0.00937f
C363 XA.XIR[7].XIC[8].icell.SM Iout 0.00388f
C364 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C365 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.SM 0.00168f
C366 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04052f
C367 XThR.Tn[6] XA.XIR[7].XIC[2].icell.SM 0.00121f
C368 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.15202f
C369 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.SM 0.0039f
C370 XThR.Tn[12] XA.XIR[13].XIC[4].icell.Ien 0.00338f
C371 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02762f
C372 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.03425f
C373 a_5949_9615# VPWR 0.7053f
C374 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.03425f
C375 XA.XIR[3].XIC[11].icell.Ien Vbias 0.21098f
C376 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00584f
C377 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C378 XA.XIR[1].XIC_dummy_left.icell.Ien Vbias 0.00329f
C379 XThR.Tn[1] XA.XIR[2].XIC[3].icell.Ien 0.00338f
C380 XThR.Tn[7] XA.XIR[8].XIC[9].icell.SM 0.00121f
C381 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.0353f
C382 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C383 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PUM 0.00465f
C384 XA.XIR[6].XIC[14].icell.PUM Vbias 0.0031f
C385 XA.XIR[0].XIC[12].icell.Ien VPWR 0.19211f
C386 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C387 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00214f
C388 XA.XIR[12].XIC[1].icell.Ien VPWR 0.1903f
C389 XA.XIR[6].XIC[6].icell.PDM Vbias 0.04261f
C390 XThR.Tn[11] XA.XIR[12].XIC[7].icell.Ien 0.00338f
C391 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C392 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.15202f
C393 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.15202f
C394 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5] 0.00341f
C395 XA.XIR[0].XIC[8].icell.Ien Iout 0.06389f
C396 XThC.TAN2 XThC.Tn[9] 0.12399f
C397 XA.XIR[1].XIC[8].icell.Ien Vbias 0.21104f
C398 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C399 XThC.Tn[11] XThR.Tn[14] 0.28739f
C400 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PUM 0.00465f
C401 XA.XIR[15].XIC[13].icell.Ien Vbias 0.17899f
C402 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00214f
C403 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PUM 0.00465f
C404 XThC.TA3 data[0] 0.86893f
C405 XThC.TAN2 XThC.TBN 0.77125f
C406 XA.XIR[5].XIC[4].icell.Ien VPWR 0.1903f
C407 XThC.TB1 data[0] 0.06453f
C408 XThC.Tn[7] XThR.Tn[5] 0.28739f
C409 XA.XIR[13].XIC[1].icell.PDM Vbias 0.04261f
C410 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.15202f
C411 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C412 XA.XIR[15].XIC[10].icell.PDM VPWR 0.0114f
C413 XA.XIR[10].XIC[0].icell.SM Iout 0.00388f
C414 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.SM 0.00168f
C415 XThR.Tn[9] XA.XIR[10].XIC[0].icell.SM 0.00127f
C416 XA.XIR[12].XIC[6].icell.PDM Vbias 0.04261f
C417 XA.XIR[6].XIC[13].icell.PDM Iout 0.00117f
C418 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01577f
C419 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C420 XThR.Tn[1] XA.XIR[1].XIC[9].icell.PDM 0.00341f
C421 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02762f
C422 XThC.Tn[12] XThR.Tn[4] 0.28739f
C423 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.SM 0.0039f
C424 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C425 XA.XIR[14].XIC[4].icell.PDM Iout 0.00117f
C426 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.15202f
C427 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.1106f
C428 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.SM 0.00168f
C429 XA.XIR[9].XIC[8].icell.PDM VPWR 0.00799f
C430 XThR.TB3 XThR.TB4 2.13136f
C431 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C432 XA.XIR[13].XIC[8].icell.PDM Iout 0.00117f
C433 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Iout 0.00347f
C434 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C435 XA.XIR[8].XIC[2].icell.PUM Vbias 0.0031f
C436 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.SM 0.0039f
C437 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.03425f
C438 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.03425f
C439 XThR.Tn[5] XA.XIR[6].XIC[4].icell.Ien 0.00338f
C440 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.15202f
C441 XA.XIR[15].XIC[14].icell.SM Vbias 0.00701f
C442 XA.XIR[2].XIC[0].icell.Ien Iout 0.06411f
C443 XA.XIR[9].XIC[8].icell.PUM VPWR 0.00937f
C444 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00256f
C445 XThC.Tn[0] XThR.Tn[11] 0.28744f
C446 XA.XIR[5].XIC[12].icell.Ien Vbias 0.21098f
C447 XA.XIR[5].XIC[2].icell.PDM Vbias 0.04261f
C448 XThC.Tn[4] XThR.Tn[3] 0.28739f
C449 XA.XIR[15].XIC[10].icell.PUM Vbias 0.0031f
C450 XA.XIR[3].XIC[14].icell.PDM Vbias 0.04261f
C451 XThC.Tn[14] XThR.Tn[0] 0.28766f
C452 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.15202f
C453 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PUM 0.00465f
C454 XThR.TBN a_n997_3755# 0.229f
C455 XA.XIR[7].XIC[1].icell.PDM VPWR 0.00799f
C456 XA.XIR[11].XIC[12].icell.SM Iout 0.00388f
C457 XThR.Tn[11] XThR.Tn[12] 0.11452f
C458 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.SM 0.0039f
C459 XA.XIR[8].XIC[4].icell.PDM Vbias 0.04261f
C460 XA.XIR[14].XIC[1].icell.SM Vbias 0.00701f
C461 XA.XIR[1].XIC_15.icell.SM Iout 0.0047f
C462 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10] 0.00341f
C463 XThC.Tn[7] Vbias 2.28836f
C464 XA.XIR[4].XIC[2].icell.SM VPWR 0.00158f
C465 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.SM 0.00168f
C466 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.SM 0.00168f
C467 XThR.TA2 data[4] 0.48493f
C468 XA.XIR[10].XIC[12].icell.PDM Iout 0.00117f
C469 XA.XIR[2].XIC[6].icell.SM VPWR 0.00158f
C470 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04031f
C471 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14] 0.00341f
C472 XA.XIR[13].XIC[3].icell.SM Vbias 0.00701f
C473 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.03425f
C474 XA.XIR[8].XIC[7].icell.PUM Vbias 0.0031f
C475 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C476 XA.XIR[2].XIC[2].icell.SM Iout 0.00388f
C477 XA.XIR[7].XIC[4].icell.PUM VPWR 0.00937f
C478 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C479 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04031f
C480 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.SM 0.0039f
C481 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PUM 0.00465f
C482 XA.XIR[0].XIC[13].icell.PDM VPWR 0.00774f
C483 XA.XIR[12].XIC[5].icell.Ien Vbias 0.21098f
C484 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00584f
C485 XA.XIR[13].XIC[13].icell.PDM Iout 0.00117f
C486 XA.XIR[5].XIC[9].icell.PDM Iout 0.00117f
C487 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C488 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01451f
C489 XThC.Tn[13] XThR.Tn[13] 0.2874f
C490 XA.XIR[14].XIC[8].icell.Ien VPWR 0.19084f
C491 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C492 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00584f
C493 XA.XIR[11].XIC[6].icell.SM Vbias 0.00701f
C494 XA.XIR[1].XIC[1].icell.PDM Vbias 0.04261f
C495 XThC.Tn[0] XThC.Tn[3] 0.12427f
C496 XThC.Tn[1] XThC.Tn[2] 0.72045f
C497 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PUM 0.00465f
C498 XA.XIR[8].XIC[11].icell.PDM Iout 0.00117f
C499 XA.XIR[3].XIC[1].icell.SM Vbias 0.00701f
C500 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04031f
C501 XA.XIR[14].XIC[4].icell.Ien Iout 0.06417f
C502 XA.XIR[9].XIC_dummy_right.icell.PUM Vbias 0.00223f
C503 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C504 XA.XIR[10].XIC[8].icell.SM Vbias 0.00701f
C505 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.SM 0.0039f
C506 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PUM 0.00429f
C507 XThR.Tn[2] XA.XIR[3].XIC[11].icell.Ien 0.00338f
C508 XA.XIR[8].XIC[12].icell.SM VPWR 0.00158f
C509 XA.XIR[15].XIC[11].icell.Ien Vbias 0.17899f
C510 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00256f
C511 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.SM 0.00168f
C512 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C513 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C514 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C515 XA.XIR[13].XIC[6].icell.Ien Iout 0.06417f
C516 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C517 XA.XIR[6].XIC[4].icell.Ien Vbias 0.21098f
C518 XA.XIR[0].XIC[2].icell.SM VPWR 0.00158f
C519 XThR.Tn[12] XA.XIR[13].XIC[12].icell.SM 0.00121f
C520 XA.XIR[8].XIC[8].icell.SM Iout 0.00388f
C521 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C522 XThC.Tn[3] XThR.Tn[12] 0.28739f
C523 XThR.Tn[4] XA.XIR[4].XIC[12].icell.PDM 0.00341f
C524 XThR.Tn[8] XA.XIR[9].XIC[8].icell.SM 0.00121f
C525 XThC.Tn[12] XThR.Tn[8] 0.28739f
C526 XThC.TB3 a_8739_9569# 0.07285f
C527 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PUM 0.00465f
C528 XA.XIR[5].XIC[0].icell.PUM VPWR 0.00937f
C529 XA.XIR[12].XIC_15.icell.SM Vbias 0.00701f
C530 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PUM 0.00465f
C531 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.03425f
C532 XA.XIR[4].XIC[10].icell.SM Vbias 0.00701f
C533 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39003f
C534 XThR.TB2 a_n1049_5317# 0.00844f
C535 XA.XIR[3].XIC[8].icell.Ien VPWR 0.1903f
C536 XA.XIR[1].XIC[8].icell.PDM Iout 0.00117f
C537 XA.XIR[11].XIC[9].icell.Ien Iout 0.06417f
C538 XA.XIR[2].XIC[14].icell.SM Vbias 0.00701f
C539 XA.XIR[2].XIC[9].icell.PDM Vbias 0.04261f
C540 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.SM 0.0039f
C541 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C542 XA.XIR[6].XIC[11].icell.PUM VPWR 0.00937f
C543 XA.XIR[3].XIC[4].icell.Ien Iout 0.06417f
C544 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PUM 0.00465f
C545 XA.XIR[7].XIC[12].icell.PUM Vbias 0.0031f
C546 XA.XIR[13].XIC[0].icell.PUM VPWR 0.00937f
C547 XA.XIR[4].XIC[8].icell.PDM VPWR 0.00799f
C548 XThC.TB4 XThC.Tn[6] 0.00608f
C549 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.SM 0.00168f
C550 XA.XIR[1].XIC[5].icell.Ien VPWR 0.1903f
C551 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7] 0.00341f
C552 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C553 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C554 XThC.Tn[2] XThR.Tn[10] 0.28739f
C555 a_3773_9615# Vbias 0.00846f
C556 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04052f
C557 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C558 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C559 XThR.Tn[13] XA.XIR[14].XIC[5].icell.SM 0.00121f
C560 XThC.Tn[12] XThR.Tn[1] 0.28739f
C561 XA.XIR[4].XIC[13].icell.Ien Iout 0.06417f
C562 XThC.TB7 a_8739_9569# 0.00474f
C563 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.SM 0.00168f
C564 XA.XIR[15].XIC[2].icell.PUM VPWR 0.00937f
C565 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PUM 0.00186f
C566 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C567 XA.XIR[0].XIC[10].icell.SM Vbias 0.00716f
C568 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.SM 0.0039f
C569 XA.XIR[4].XIC_dummy_right.icell.Ien Vbias 0.00288f
C570 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04031f
C571 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C572 XA.XIR[7].XIC[13].icell.SM Iout 0.00388f
C573 XThR.Tn[6] XA.XIR[7].XIC[7].icell.SM 0.00121f
C574 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.SM 0.0039f
C575 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.15202f
C576 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C577 XThR.Tn[12] XA.XIR[13].XIC[9].icell.Ien 0.00338f
C578 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.SM 0.00168f
C579 XA.XIR[6].XIC_15.icell.SM VPWR 0.00275f
C580 XA.XIR[11].XIC[3].icell.PDM VPWR 0.00799f
C581 XA.XIR[11].XIC[2].icell.PUM Vbias 0.0031f
C582 XA.XIR[11].XIC[10].icell.SM Iout 0.00388f
C583 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Ien 0.00232f
C584 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.SM 0.0039f
C585 XThC.TA3 XThC.TB3 0.57441f
C586 XThR.Tn[1] XA.XIR[2].XIC[8].icell.Ien 0.00338f
C587 XThR.TB6 XThR.TB7 2.05133f
C588 XA.XIR[5].XIC[2].icell.SM Vbias 0.00701f
C589 XThR.Tn[7] XA.XIR[8].XIC[14].icell.SM 0.00121f
C590 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C591 XThC.TB1 XThC.TB3 0.04033f
C592 XA.XIR[10].XIC[7].icell.PDM VPWR 0.00799f
C593 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C594 XA.XIR[9].XIC[1].icell.Ien Vbias 0.21098f
C595 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04052f
C596 XA.XIR[1].XIC[1].icell.PUM Vbias 0.0031f
C597 XA.XIR[13].XIC[0].icell.SM Iout 0.00388f
C598 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02762f
C599 XA.XIR[15].XIC[6].icell.PDM Vbias 0.04261f
C600 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C601 XA.XIR[0].XIC[13].icell.Ien Iout 0.06389f
C602 XThR.TB1 XThR.TB4 0.05121f
C603 XA.XIR[1].XIC[13].icell.Ien Vbias 0.21104f
C604 XThC.Tn[7] XThR.Tn[2] 0.28746f
C605 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C606 a_8739_9569# VPWR 0.00583f
C607 XA.XIR[5].XIC[9].icell.Ien VPWR 0.1903f
C608 XA.XIR[15].XIC[7].icell.PUM VPWR 0.00937f
C609 XA.XIR[0].XIC_dummy_right.icell.Ien Vbias 0.00307f
C610 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C611 XA.XIR[3].XIC[5].icell.PDM VPWR 0.00799f
C612 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.03425f
C613 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00214f
C614 XA.XIR[5].XIC[5].icell.Ien Iout 0.06417f
C615 a_n1049_5317# XThR.Tn[6] 0.26047f
C616 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.SM 0.00168f
C617 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C618 XA.XIR[9].XIC[4].icell.PDM Vbias 0.04261f
C619 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.SM 0.0039f
C620 XThC.TB5 a_9827_9569# 0.06458f
C621 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00584f
C622 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C623 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6] 0.00341f
C624 XThC.TA3 XThC.TB7 0.37429f
C625 XThR.TBN a_n997_715# 0.21503f
C626 XThR.Tn[12] XA.XIR[13].XIC[10].icell.SM 0.00121f
C627 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00584f
C628 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00214f
C629 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.03425f
C630 XThC.TB2 XThC.TB6 0.04959f
C631 XThC.TB1 XThC.TB7 0.05222f
C632 XThC.Tn[0] XThR.Tn[14] 0.28742f
C633 XA.XIR[9].XIC[6].icell.Ien Vbias 0.21098f
C634 XA.XIR[8].XIC[4].icell.PUM VPWR 0.00937f
C635 XThR.TA2 XThR.TA3 0.44014f
C636 XThC.Tn[2] XA.XIR[0].XIC[4].icell.PDM 0.00353f
C637 XThC.TB7 XThC.Tn[11] 0.07471f
C638 XThR.Tn[2] XA.XIR[3].XIC[1].icell.SM 0.00121f
C639 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02762f
C640 XThC.TAN2 XThC.Tn[7] 0.01439f
C641 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.SM 0.00168f
C642 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02762f
C643 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00214f
C644 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.15202f
C645 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00584f
C646 XThR.Tn[13] a_n997_1579# 0.19413f
C647 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C648 XA.XIR[10].XIC[11].icell.PDM Iout 0.00117f
C649 XA.XIR[12].XIC[2].icell.Ien VPWR 0.1903f
C650 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04031f
C651 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02762f
C652 XThR.Tn[5] Iout 1.16233f
C653 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C654 XA.XIR[14].XIC[12].icell.SM Iout 0.00388f
C655 XThR.TB7 XThR.Tn[8] 0.07806f
C656 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C657 XA.XIR[11].XIC[3].icell.SM VPWR 0.00158f
C658 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00214f
C659 XThR.Tn[5] XA.XIR[6].XIC[9].icell.Ien 0.00338f
C660 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.15202f
C661 XA.XIR[9].XIC[11].icell.PDM Iout 0.00117f
C662 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9] 0.00341f
C663 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PUM 0.00465f
C664 XA.XIR[13].XIC[12].icell.PDM Iout 0.00117f
C665 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PUM 0.00465f
C666 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C667 XA.XIR[9].XIC[13].icell.PUM VPWR 0.00937f
C668 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.SM 0.0039f
C669 XA.XIR[2].XIC[6].icell.PUM Vbias 0.0031f
C670 XThC.Tn[1] XThR.Tn[4] 0.28739f
C671 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11] 0.00341f
C672 XA.XIR[10].XIC[5].icell.SM VPWR 0.00158f
C673 XA.XIR[10].XIC[13].icell.SM Vbias 0.00701f
C674 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC[14].icell.SM 0.0039f
C675 XThR.Tn[14] XA.XIR[15].XIC[2].icell.Ien 0.00338f
C676 XThR.Tn[2] XA.XIR[2].XIC[9].icell.PDM 0.00341f
C677 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C678 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C679 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.SM 0.0039f
C680 XThC.TA3 VPWR 0.87301f
C681 XA.XIR[10].XIC[1].icell.SM Iout 0.00388f
C682 XA.XIR[7].XIC[2].icell.Ien Vbias 0.21098f
C683 XThC.TB1 VPWR 1.1176f
C684 XThR.Tn[9] XA.XIR[10].XIC[1].icell.SM 0.00121f
C685 XA.XIR[0].XIC[9].icell.PDM Vbias 0.04282f
C686 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C687 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.03023f
C688 XThC.Tn[11] VPWR 6.86576f
C689 XA.XIR[14].XIC[6].icell.SM Vbias 0.00701f
C690 XA.XIR[4].XIC[7].icell.SM VPWR 0.00158f
C691 XA.XIR[11].XIC[14].icell.Ien Iout 0.06417f
C692 XA.XIR[2].XIC[11].icell.SM VPWR 0.00158f
C693 XA.XIR[12].XIC_15.icell.PDM Vbias 0.04401f
C694 XA.XIR[7].XIC[4].icell.PDM Iout 0.00117f
C695 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38936f
C696 XA.XIR[2].XIC[0].icell.PDM VPWR 0.00799f
C697 XA.XIR[12].XIC_dummy_right.icell.PUM Vbias 0.00223f
C698 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C699 XA.XIR[13].XIC[8].icell.SM Vbias 0.00701f
C700 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C701 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.SM 0.00168f
C702 XA.XIR[4].XIC[3].icell.SM Iout 0.00388f
C703 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C704 XA.XIR[2].XIC[7].icell.SM Iout 0.00388f
C705 XA.XIR[7].XIC[9].icell.PUM VPWR 0.00937f
C706 XA.XIR[8].XIC[12].icell.PUM Vbias 0.0031f
C707 XThC.Tn[0] XA.XIR[4].XIC_dummy_left.icell.Iout 0.00109f
C708 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.03433f
C709 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.SM 0.0039f
C710 XThC.Tn[3] XThR.Tn[0] 0.28743f
C711 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00214f
C712 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C713 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.SM 0.00168f
C714 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04031f
C715 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PUM 0.00465f
C716 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39f
C717 XA.XIR[3].XIC[2].icell.PUM VPWR 0.00937f
C718 XA.XIR[14].XIC[9].icell.Ien Iout 0.06417f
C719 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C720 XA.XIR[3].XIC[6].icell.SM Vbias 0.00701f
C721 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[3].icell.Ien 0.00214f
C722 Vbias Iout 83.1596f
C723 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.SM 0.0039f
C724 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00214f
C725 XThR.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.00338f
C726 XThR.Tn[9] Vbias 3.74874f
C727 XThC.TAN XThC.Tn[9] 0.09571f
C728 XA.XIR[1].XIC[1].icell.Ien Iout 0.06417f
C729 XA.XIR[6].XIC[9].icell.Ien Vbias 0.21098f
C730 XA.XIR[0].XIC[7].icell.SM VPWR 0.00158f
C731 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Iout 0.00347f
C732 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.03425f
C733 XThR.Tn[11] XA.XIR[12].XIC[2].icell.SM 0.00121f
C734 XThR.TA3 a_n1049_7493# 0.0127f
C735 XA.XIR[8].XIC[13].icell.SM Iout 0.00388f
C736 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C737 XThC.TA3 a_5155_9615# 0.02287f
C738 XThR.Tn[8] XA.XIR[9].XIC[13].icell.SM 0.00121f
C739 XThC.TAN XThC.TBN 0.38751f
C740 XA.XIR[4].XIC[4].icell.PDM Vbias 0.04261f
C741 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C742 XA.XIR[0].XIC[3].icell.SM Iout 0.00367f
C743 XThR.Tn[12] XA.XIR[13].XIC[14].icell.Ien 0.00338f
C744 XA.XIR[1].XIC[3].icell.SM Vbias 0.00704f
C745 XThC.Tn[2] XThR.Tn[13] 0.28739f
C746 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.SM 0.0039f
C747 XThC.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00109f
C748 XA.XIR[3].XIC[13].icell.Ien VPWR 0.1903f
C749 XA.XIR[10].XIC[1].icell.PUM VPWR 0.00937f
C750 XA.XIR[3].XIC[9].icell.Ien Iout 0.06417f
C751 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Ien 0.00584f
C752 XThR.Tn[0] XA.XIR[0].XIC[10].icell.PDM 0.00341f
C753 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C754 XThR.TAN XThR.Tn[5] 0.00705f
C755 XThR.TB6 XThR.Tn[10] 0.02461f
C756 XA.XIR[6].XIC[12].icell.PDM VPWR 0.00799f
C757 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PUM 0.00465f
C758 XThC.Tn[5] Iout 0.83957f
C759 XA.XIR[15].XIC[0].icell.Ien Vbias 0.17752f
C760 XThC.Tn[5] XThR.Tn[9] 0.28739f
C761 XA.XIR[6].XIC[0].icell.PDM Iout 0.00117f
C762 XA.XIR[1].XIC[10].icell.Ien VPWR 0.1903f
C763 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.SM 0.00168f
C764 XThC.Tn[1] XThR.Tn[8] 0.28739f
C765 XA.XIR[4].XIC[11].icell.PDM Iout 0.00117f
C766 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00256f
C767 XA.XIR[14].XIC[3].icell.PDM VPWR 0.00799f
C768 XA.XIR[14].XIC[2].icell.PUM Vbias 0.0031f
C769 XA.XIR[14].XIC[10].icell.SM Iout 0.00388f
C770 XA.XIR[1].XIC[6].icell.Ien Iout 0.06417f
C771 XA.XIR[13].XIC[7].icell.PDM VPWR 0.00799f
C772 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.SM 0.00168f
C773 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C774 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Ien 0.00232f
C775 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.03425f
C776 XA.XIR[10].XIC[3].icell.PDM Vbias 0.04261f
C777 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C778 XA.XIR[10].XIC[11].icell.SM Vbias 0.00701f
C779 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00214f
C780 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C781 XThR.Tn[6] XA.XIR[7].XIC[12].icell.SM 0.00121f
C782 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.SM 0.00168f
C783 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PUM 0.00465f
C784 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C785 XA.XIR[12].XIC[0].icell.PDM Iout 0.00117f
C786 XA.XIR[9].XIC[3].icell.Ien VPWR 0.1903f
C787 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04031f
C788 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00584f
C789 XA.XIR[5].XIC[7].icell.SM Vbias 0.00701f
C790 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.03425f
C791 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00584f
C792 XThR.Tn[1] XA.XIR[2].XIC[13].icell.Ien 0.00338f
C793 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04031f
C794 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04031f
C795 XA.XIR[15].XIC[5].icell.Ien Vbias 0.17899f
C796 XA.XIR[11].XIC[6].icell.PDM Iout 0.00117f
C797 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.03425f
C798 XThC.Tn[1] XThR.Tn[1] 0.28739f
C799 XA.XIR[11].XIC[12].icell.Ien Iout 0.06417f
C800 XA.XIR[3].XIC[1].icell.PDM Vbias 0.04261f
C801 XThR.TB7 a_n997_3755# 0.00476f
C802 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00214f
C803 XThR.Tn[0] XA.XIR[1].XIC[4].icell.Ien 0.00338f
C804 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C805 XA.XIR[10].XIC[10].icell.PDM Iout 0.00117f
C806 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04031f
C807 XThR.Tn[8] XThR.Tn[10] 0.00255f
C808 XA.XIR[2].XIC[3].icell.PUM VPWR 0.00937f
C809 XThR.TBN a_n997_2667# 0.22784f
C810 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C811 XA.XIR[5].XIC[14].icell.Ien VPWR 0.19036f
C812 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02762f
C813 XA.XIR[5].XIC[8].icell.PDM VPWR 0.00799f
C814 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C815 XA.XIR[4].XIC[2].icell.PUM Vbias 0.0031f
C816 XA.XIR[13].XIC[11].icell.PDM Iout 0.00117f
C817 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PUM 0.00442f
C818 XA.XIR[8].XIC[2].icell.Ien Vbias 0.21098f
C819 XThR.Tn[10] XA.XIR[11].XIC[1].icell.Ien 0.00338f
C820 XThC.TB2 XThC.Tn[1] 0.17879f
C821 XA.XIR[15].XIC_15.icell.SM Vbias 0.00701f
C822 XA.XIR[10].XIC[14].icell.PUM Vbias 0.0031f
C823 XA.XIR[5].XIC[10].icell.Ien Iout 0.06417f
C824 XThC.TAN data[2] 0.07481f
C825 XA.XIR[0].XIC[0].icell.PDM VPWR 0.00774f
C826 XA.XIR[8].XIC[10].icell.PDM VPWR 0.00799f
C827 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.03023f
C828 XA.XIR[6].XIC[1].icell.Ien VPWR 0.1903f
C829 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C830 XA.XIR[3].XIC[8].icell.PDM Iout 0.00117f
C831 XA.XIR[14].XIC[3].icell.SM VPWR 0.00158f
C832 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.0353f
C833 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13] 0.00341f
C834 XA.XIR[11].XIC[3].icell.PUM Vbias 0.0031f
C835 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00584f
C836 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C837 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.SM 0.00168f
C838 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C839 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00214f
C840 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04031f
C841 XA.XIR[13].XIC[5].icell.SM VPWR 0.00158f
C842 XA.XIR[13].XIC[13].icell.SM Vbias 0.00701f
C843 XA.XIR[8].XIC[9].icell.PUM VPWR 0.00937f
C844 XA.XIR[9].XIC[11].icell.Ien Vbias 0.21098f
C845 XThR.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.00338f
C846 XThR.Tn[2] Iout 1.16236f
C847 XA.XIR[10].XIC[5].icell.PUM Vbias 0.0031f
C848 XThR.Tn[2] XA.XIR[3].XIC[6].icell.SM 0.00121f
C849 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.03425f
C850 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.03425f
C851 XA.XIR[13].XIC[1].icell.SM Iout 0.00388f
C852 XThC.Tn[13] XThR.Tn[7] 0.2874f
C853 XA.XIR[12].XIC[14].icell.PDM Vbias 0.04261f
C854 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C855 XA.XIR[12].XIC[7].icell.Ien VPWR 0.1903f
C856 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C857 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12] 0.00341f
C858 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.03425f
C859 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Iout 0.00347f
C860 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C861 XThR.Tn[3] XA.XIR[3].XIC[6].icell.PDM 0.00341f
C862 XA.XIR[12].XIC[3].icell.Ien Iout 0.06417f
C863 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C864 XA.XIR[11].XIC[8].icell.SM VPWR 0.00158f
C865 XA.XIR[1].XIC[7].icell.PDM VPWR 0.00799f
C866 XA.XIR[7].XIC[12].icell.PDM Vbias 0.04261f
C867 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.15202f
C868 XThR.Tn[5] XA.XIR[6].XIC[14].icell.Ien 0.00338f
C869 XA.XIR[0].XIC[2].icell.PUM Vbias 0.0031f
C870 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C871 XA.XIR[15].XIC_15.icell.PDM Vbias 0.04401f
C872 XA.XIR[14].XIC[14].icell.Ien Iout 0.06417f
C873 XA.XIR[4].XIC[7].icell.PUM Vbias 0.0031f
C874 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04031f
C875 XThR.TB6 a_n997_1803# 0.00871f
C876 XA.XIR[3].XIC[3].icell.SM VPWR 0.00158f
C877 XA.XIR[2].XIC[11].icell.PUM Vbias 0.0031f
C878 XA.XIR[11].XIC[4].icell.SM Iout 0.00388f
C879 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C880 XA.XIR[6].XIC[6].icell.Ien VPWR 0.1903f
C881 XThR.Tn[14] XA.XIR[15].XIC[7].icell.Ien 0.00338f
C882 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PUM 0.00465f
C883 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Iout 0.00347f
C884 XThR.TBN XThR.Tn[11] 0.52266f
C885 XThR.Tn[4] XA.XIR[5].XIC[1].icell.Ien 0.00338f
C886 XA.XIR[7].XIC[7].icell.Ien Vbias 0.21098f
C887 XA.XIR[10].XIC[6].icell.SM Iout 0.00388f
C888 XThC.Tn[8] XThC.Tn[9] 0.05322f
C889 XThR.Tn[9] XA.XIR[10].XIC[6].icell.SM 0.00121f
C890 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.15202f
C891 XThC.TB5 data[3] 0.00931f
C892 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PUM 0.00465f
C893 XA.XIR[6].XIC[2].icell.Ien Iout 0.06417f
C894 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.SM 0.00168f
C895 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.03425f
C896 XThC.Tn[12] XThC.Tn[14] 0.03994f
C897 XThC.TBN XThC.Tn[8] 0.50311f
C898 XA.XIR[10].XIC[9].icell.SM Vbias 0.00701f
C899 XThR.TBN XThR.TA3 0.59539f
C900 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00214f
C901 XA.XIR[4].XIC[12].icell.SM VPWR 0.00158f
C902 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04031f
C903 XA.XIR[3].XIC[0].icell.Ien Vbias 0.20951f
C904 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07214f
C905 XA.XIR[4].XIC[8].icell.SM Iout 0.00388f
C906 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8] 0.00341f
C907 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00214f
C908 XA.XIR[7].XIC[14].icell.PUM VPWR 0.00937f
C909 XA.XIR[12].XIC_dummy_left.icell.Ien Vbias 0.00329f
C910 XA.XIR[2].XIC[12].icell.SM Iout 0.00388f
C911 XA.XIR[2].XIC[3].icell.PDM Iout 0.00117f
C912 XA.XIR[5].XIC[1].icell.PUM VPWR 0.00937f
C913 XA.XIR[0].XIC[7].icell.PUM Vbias 0.0031f
C914 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.SM 0.00168f
C915 XA.XIR[11].XIC[10].icell.Ien Iout 0.06417f
C916 XA.XIR[2].XIC_15.icell.SM Vbias 0.00701f
C917 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C918 XThR.Tn[12] XA.XIR[13].XIC[4].icell.SM 0.00121f
C919 XThC.Tn[0] VPWR 5.95931f
C920 XThR.Tn[4] XA.XIR[5].XIC[6].icell.Ien 0.00338f
C921 XA.XIR[3].XIC[11].icell.SM Vbias 0.00701f
C922 XThR.Tn[1] XA.XIR[2].XIC[3].icell.SM 0.00121f
C923 XA.XIR[13].XIC[1].icell.PUM VPWR 0.00937f
C924 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.15202f
C925 XThR.Tn[3] XA.XIR[4].XIC[8].icell.Ien 0.00338f
C926 XThR.TB6 XThR.Tn[13] 0.32265f
C927 XA.XIR[6].XIC[14].icell.Ien Vbias 0.21098f
C928 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04031f
C929 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C930 XA.XIR[0].XIC[12].icell.SM VPWR 0.00158f
C931 XA.XIR[6].XIC[8].icell.PDM Vbias 0.04261f
C932 XThR.Tn[11] XA.XIR[12].XIC[7].icell.SM 0.00121f
C933 XThC.TB6 XThC.Tn[14] 0.00128f
C934 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PUM 0.00465f
C935 XThR.Tn[12] VPWR 7.57625f
C936 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C937 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C938 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.04494f
C939 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5] 0.00341f
C940 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C941 XA.XIR[0].XIC[8].icell.SM Iout 0.00367f
C942 Vbias data[1] 0.00255f
C943 XA.XIR[1].XIC[8].icell.SM Vbias 0.00704f
C944 XA.XIR[10].XIC[12].icell.PUM Vbias 0.0031f
C945 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.SM 0.00168f
C946 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.03425f
C947 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C948 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.03425f
C949 XA.XIR[2].XIC[0].icell.PUM VPWR 0.00937f
C950 XA.XIR[5].XIC[4].icell.SM VPWR 0.00158f
C951 XA.XIR[15].XIC[2].icell.Ien VPWR 0.32895f
C952 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C953 XA.XIR[11].XIC[0].icell.Ien Iout 0.06411f
C954 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C955 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.03425f
C956 XA.XIR[13].XIC[3].icell.PDM Vbias 0.04261f
C957 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.04498f
C958 XA.XIR[3].XIC[14].icell.Ien Iout 0.06417f
C959 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.SM 0.0039f
C960 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00214f
C961 XA.XIR[13].XIC[11].icell.SM Vbias 0.00701f
C962 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C963 XThR.Tn[12] XA.XIR[13].XIC[10].icell.Ien 0.00338f
C964 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C965 XThR.TB4 a_n1049_6699# 0.23756f
C966 XA.XIR[12].XIC[8].icell.PDM Vbias 0.04261f
C967 XThR.TB7 a_n997_715# 0.06874f
C968 XA.XIR[6].XIC_15.icell.PDM Iout 0.00133f
C969 XA.XIR[1].XIC_15.icell.Ien VPWR 0.25566f
C970 XThC.TAN XThC.Tn[7] 0.08407f
C971 XA.XIR[15].XIC[0].icell.PDM Iout 0.00117f
C972 XThR.TA2 a_n1319_5317# 0.00295f
C973 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C974 XThR.Tn[1] XA.XIR[1].XIC[11].icell.PDM 0.00341f
C975 XThR.TB5 a_n1049_5317# 0.00907f
C976 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.SM 0.00168f
C977 XA.XIR[1].XIC[11].icell.Ien Iout 0.06417f
C978 XA.XIR[9].XIC[1].icell.SM Vbias 0.00701f
C979 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.SM 0.0039f
C980 XA.XIR[14].XIC[6].icell.PDM Iout 0.00117f
C981 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02762f
C982 XA.XIR[14].XIC[12].icell.Ien Iout 0.06417f
C983 XA.XIR[9].XIC[10].icell.PDM VPWR 0.00799f
C984 XA.XIR[13].XIC[10].icell.PDM Iout 0.00117f
C985 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00214f
C986 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.SM 0.00168f
C987 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PUM 0.00465f
C988 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00214f
C989 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.SM 0.0039f
C990 XThR.Tn[5] XA.XIR[6].XIC[4].icell.SM 0.00121f
C991 XA.XIR[15].XIC_dummy_right.icell.PUM Vbias 0.00223f
C992 XA.XIR[10].XIC[13].icell.Ien Vbias 0.21098f
C993 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08441f
C994 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.15202f
C995 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.15202f
C996 XA.XIR[9].XIC[8].icell.Ien VPWR 0.1903f
C997 XThR.TA3 a_n1049_5611# 0.01824f
C998 XThR.TB4 XThR.Tn[9] 0.01318f
C999 XA.XIR[5].XIC[12].icell.SM Vbias 0.00701f
C1000 XThC.TA2 data[1] 0.37233f
C1001 XA.XIR[5].XIC[4].icell.PDM Vbias 0.04261f
C1002 XA.XIR[9].XIC[4].icell.Ien Iout 0.06417f
C1003 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C1004 XA.XIR[13].XIC[14].icell.PUM Vbias 0.0031f
C1005 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.15202f
C1006 XThC.TA1 data[1] 0.11102f
C1007 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00214f
C1008 XThR.Tn[0] XA.XIR[1].XIC[9].icell.Ien 0.00338f
C1009 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.SM 0.0039f
C1010 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.03425f
C1011 XA.XIR[7].XIC[3].icell.PDM VPWR 0.00799f
C1012 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C1013 XA.XIR[12].XIC[13].icell.PDM Vbias 0.04261f
C1014 XThC.TB5 XThC.Tn[12] 0.32495f
C1015 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.0353f
C1016 XA.XIR[11].XIC[13].icell.SM VPWR 0.00158f
C1017 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1018 XA.XIR[8].XIC[6].icell.PDM Vbias 0.04261f
C1019 XA.XIR[14].XIC[3].icell.PUM Vbias 0.0031f
C1020 XA.XIR[4].XIC[4].icell.PUM VPWR 0.00937f
C1021 XThR.TB1 bias[2] 0.00266f
C1022 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10] 0.00341f
C1023 XThC.Tn[10] XThR.Tn[5] 0.28739f
C1024 XA.XIR[2].XIC[8].icell.PUM VPWR 0.00937f
C1025 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14] 0.00341f
C1026 XThR.Tn[2] XA.XIR[3].XIC[0].icell.Ien 0.00338f
C1027 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00584f
C1028 XA.XIR[13].XIC[5].icell.PUM Vbias 0.0031f
C1029 XA.XIR[8].XIC[7].icell.Ien Vbias 0.21098f
C1030 XA.XIR[15].XIC[14].icell.PDM Vbias 0.04261f
C1031 XA.XIR[7].XIC[4].icell.Ien VPWR 0.1903f
C1032 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00584f
C1033 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C1034 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07079f
C1035 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.03425f
C1036 XA.XIR[5].XIC_15.icell.Ien Iout 0.0642f
C1037 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C1038 XA.XIR[5].XIC[11].icell.PDM Iout 0.00117f
C1039 XA.XIR[12].XIC[5].icell.SM Vbias 0.00701f
C1040 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C1041 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1042 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.SM 0.0039f
C1043 XA.XIR[14].XIC[8].icell.SM VPWR 0.00158f
C1044 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00584f
C1045 a_10915_9569# XThC.Tn[14] 0.20278f
C1046 XA.XIR[10].XIC[14].icell.SM Vbias 0.00701f
C1047 XA.XIR[11].XIC[8].icell.PUM Vbias 0.0031f
C1048 XA.XIR[1].XIC[3].icell.PDM Vbias 0.04261f
C1049 XA.XIR[8].XIC[13].icell.PDM Iout 0.00117f
C1050 XA.XIR[14].XIC[4].icell.SM Iout 0.00388f
C1051 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.03425f
C1052 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00214f
C1053 XA.XIR[1].XIC[0].icell.SM VPWR 0.00158f
C1054 XA.XIR[3].XIC[3].icell.PUM Vbias 0.0031f
C1055 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04052f
C1056 XThR.Tn[2] XA.XIR[3].XIC[11].icell.SM 0.00121f
C1057 XA.XIR[8].XIC[14].icell.PUM VPWR 0.00937f
C1058 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.SM 0.00168f
C1059 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.03589f
C1060 XA.XIR[10].XIC[10].icell.PUM Vbias 0.0031f
C1061 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C1062 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.SM 0.00168f
C1063 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00214f
C1064 XThR.TBN XThR.Tn[14] 0.47807f
C1065 XA.XIR[6].XIC[4].icell.SM Vbias 0.00701f
C1066 XA.XIR[13].XIC[6].icell.SM Iout 0.00388f
C1067 XThC.TB5 XThC.TB6 2.12831f
C1068 XA.XIR[0].XIC[4].icell.PUM VPWR 0.00882f
C1069 XThR.Tn[4] XA.XIR[4].XIC[14].icell.PDM 0.00341f
C1070 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PUM 0.00465f
C1071 XA.XIR[11].XIC_15.icell.PDM Iout 0.00133f
C1072 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.SM 0.00168f
C1073 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.15202f
C1074 XA.XIR[11].XIC_15.icell.Ien Iout 0.0642f
C1075 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.03425f
C1076 XA.XIR[12].XIC[8].icell.Ien Iout 0.06417f
C1077 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02762f
C1078 XA.XIR[13].XIC[9].icell.SM Vbias 0.00701f
C1079 VPWR data[7] 0.212f
C1080 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00214f
C1081 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PUM 0.00465f
C1082 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.SM 0.00168f
C1083 XA.XIR[4].XIC[12].icell.PUM Vbias 0.0031f
C1084 XA.XIR[3].XIC[8].icell.SM VPWR 0.00158f
C1085 XA.XIR[1].XIC[10].icell.PDM Iout 0.00117f
C1086 XA.XIR[2].XIC_dummy_right.icell.PUM Vbias 0.00223f
C1087 XThC.Tn[12] XThR.Tn[11] 0.28739f
C1088 XA.XIR[2].XIC[11].icell.PDM Vbias 0.04261f
C1089 XThR.Tn[10] XA.XIR[11].XIC[2].icell.Ien 0.00338f
C1090 XA.XIR[3].XIC[4].icell.SM Iout 0.00388f
C1091 XA.XIR[6].XIC[11].icell.Ien VPWR 0.1903f
C1092 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PUM 0.00465f
C1093 XThR.TA2 VPWR 0.68638f
C1094 XA.XIR[7].XIC[12].icell.Ien Vbias 0.21098f
C1095 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C1096 XThC.Tn[2] XThR.Tn[7] 0.28739f
C1097 XA.XIR[4].XIC[10].icell.PDM VPWR 0.00799f
C1098 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C1099 XThC.Tn[10] Vbias 2.36503f
C1100 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.15202f
C1101 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7] 0.00341f
C1102 XA.XIR[6].XIC[7].icell.Ien Iout 0.06417f
C1103 XA.XIR[14].XIC[10].icell.Ien Iout 0.06417f
C1104 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Iout 0.00347f
C1105 XA.XIR[1].XIC[5].icell.SM VPWR 0.00158f
C1106 XThR.TAN XThR.TB4 0.33064f
C1107 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C1108 a_4861_9615# Vbias 0.00548f
C1109 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.SM 0.00168f
C1110 XA.XIR[1].XIC[1].icell.SM Iout 0.00388f
C1111 XThC.Tn[11] XThR.Tn[6] 0.28739f
C1112 XA.XIR[10].XIC[11].icell.Ien Vbias 0.21098f
C1113 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.SM 0.00168f
C1114 XThC.TAN2 data[1] 0.01444f
C1115 XA.XIR[4].XIC[13].icell.SM Iout 0.00388f
C1116 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.15202f
C1117 XThR.Tn[12] XA.XIR[13].XIC_15.icell.Ien 0.00117f
C1118 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.15202f
C1119 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.389f
C1120 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02762f
C1121 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C1122 XThC.TB7 a_9827_9569# 0.00571f
C1123 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00584f
C1124 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.01438f
C1125 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.SM 0.0039f
C1126 XA.XIR[0].XIC[12].icell.PUM Vbias 0.0031f
C1127 XThR.Tn[0] VPWR 6.66912f
C1128 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.SM 0.00168f
C1129 XThC.TA3 XThC.Tn[4] 0.0274f
C1130 XA.XIR[12].XIC[1].icell.PUM Vbias 0.0031f
C1131 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C1132 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04031f
C1133 XA.XIR[5].XIC[0].icell.SM Iout 0.00388f
C1134 XA.XIR[13].XIC[12].icell.PUM Vbias 0.0031f
C1135 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.SM 0.0039f
C1136 XA.XIR[11].XIC[5].icell.PDM VPWR 0.00799f
C1137 XThC.TB3 a_4387_10575# 0.00941f
C1138 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C1139 XThC.Tn[7] XThC.Tn[8] 0.07597f
C1140 XThR.Tn[4] XA.XIR[5].XIC[11].icell.Ien 0.00338f
C1141 XA.XIR[11].XIC[11].icell.SM VPWR 0.00158f
C1142 XThR.Tn[1] XA.XIR[2].XIC[8].icell.SM 0.00121f
C1143 XA.XIR[5].XIC[4].icell.PUM Vbias 0.0031f
C1144 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[8].icell.Ien 0.00214f
C1145 XThC.TBN XThC.Tn[6] 0.61358f
C1146 XThR.Tn[3] XA.XIR[4].XIC[13].icell.Ien 0.00338f
C1147 XA.XIR[10].XIC[9].icell.PDM VPWR 0.00799f
C1148 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00214f
C1149 a_4861_9615# XThC.Tn[5] 0.00208f
C1150 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C1151 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.SM 0.0039f
C1152 XA.XIR[15].XIC[8].icell.PDM Vbias 0.04261f
C1153 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C1154 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01432f
C1155 XA.XIR[0].XIC[13].icell.SM Iout 0.00367f
C1156 XA.XIR[1].XIC[13].icell.SM Vbias 0.00704f
C1157 a_9827_9569# VPWR 0.0017f
C1158 XThR.TB7 a_n997_2667# 0.00474f
C1159 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00584f
C1160 XA.XIR[5].XIC[9].icell.SM VPWR 0.00158f
C1161 XA.XIR[15].XIC[7].icell.Ien VPWR 0.32895f
C1162 XThR.TBN XA.XIR[0].XIC_dummy_left.icell.Iout 0.00137f
C1163 XA.XIR[3].XIC[7].icell.PDM VPWR 0.00799f
C1164 XThC.TB4 XThC.Tn[9] 0.01318f
C1165 XA.XIR[2].XIC[1].icell.Ien Vbias 0.21098f
C1166 XA.XIR[5].XIC[5].icell.SM Iout 0.00388f
C1167 XA.XIR[15].XIC[3].icell.Ien Iout 0.06807f
C1168 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00584f
C1169 XThC.TB4 XThC.TBN 0.15636f
C1170 XA.XIR[9].XIC[6].icell.PDM Vbias 0.04261f
C1171 XA.XIR[13].XIC[13].icell.Ien Vbias 0.21098f
C1172 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6] 0.00341f
C1173 a_n1049_7493# VPWR 0.72084f
C1174 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00214f
C1175 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Iout 0.00347f
C1176 XThC.Tn[14] XThR.Tn[10] 0.28745f
C1177 XA.XIR[12].XIC[12].icell.PDM Vbias 0.04261f
C1178 XA.XIR[11].XIC[14].icell.PUM VPWR 0.00937f
C1179 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.SM 0.0039f
C1180 XA.XIR[1].XIC_dummy_right.icell.SM VPWR 0.00123f
C1181 XA.XIR[9].XIC[6].icell.SM Vbias 0.00701f
C1182 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C1183 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02762f
C1184 XA.XIR[8].XIC[4].icell.Ien VPWR 0.1903f
C1185 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C1186 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.SM 0.00168f
C1187 XThR.Tn[13] XA.XIR[14].XIC[1].icell.Ien 0.00338f
C1188 XA.XIR[12].XIC[2].icell.SM VPWR 0.00158f
C1189 XA.XIR[14].XIC[13].icell.SM VPWR 0.00158f
C1190 XA.XIR[15].XIC[13].icell.PDM Vbias 0.04261f
C1191 XA.XIR[11].XIC[5].icell.PUM VPWR 0.00937f
C1192 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04031f
C1193 XA.XIR[9].XIC[13].icell.PDM Iout 0.00117f
C1194 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00214f
C1195 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.03425f
C1196 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.03425f
C1197 XThR.Tn[5] XA.XIR[6].XIC[9].icell.SM 0.00121f
C1198 XThR.TB6 a_n997_3979# 0.0046f
C1199 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9] 0.00341f
C1200 XA.XIR[4].XIC[2].icell.Ien Vbias 0.21098f
C1201 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.15202f
C1202 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00214f
C1203 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.SM 0.0039f
C1204 XA.XIR[9].XIC[13].icell.Ien VPWR 0.1903f
C1205 XA.XIR[7].XIC[0].icell.Ien Iout 0.06411f
C1206 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.SM 0.00168f
C1207 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00214f
C1208 XA.XIR[10].XIC[7].icell.PUM VPWR 0.00937f
C1209 XA.XIR[2].XIC[6].icell.Ien Vbias 0.21098f
C1210 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11] 0.00341f
C1211 XThC.TAN Iout 0.00967f
C1212 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00584f
C1213 XThR.Tn[2] XA.XIR[2].XIC[11].icell.PDM 0.00341f
C1214 XA.XIR[6].XIC[1].icell.SM VPWR 0.00158f
C1215 XThR.Tn[14] XA.XIR[15].XIC[2].icell.SM 0.00121f
C1216 XThR.TB7 XThR.Tn[11] 0.07412f
C1217 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00584f
C1218 XA.XIR[9].XIC[9].icell.Ien Iout 0.06417f
C1219 XA.XIR[7].XIC[2].icell.SM Vbias 0.00701f
C1220 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.15202f
C1221 XThR.Tn[7] XA.XIR[8].XIC[1].icell.Ien 0.00338f
C1222 XA.XIR[0].XIC[11].icell.PDM Vbias 0.04282f
C1223 XThC.Tn[10] XThR.Tn[2] 0.28739f
C1224 XThR.Tn[0] XA.XIR[1].XIC[14].icell.Ien 0.00338f
C1225 XA.XIR[13].XIC[14].icell.SM Vbias 0.00701f
C1226 XThR.TA3 XThR.TB7 0.37429f
C1227 XA.XIR[14].XIC[8].icell.PUM Vbias 0.0031f
C1228 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.SM 0.0039f
C1229 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00584f
C1230 XA.XIR[4].XIC[9].icell.PUM VPWR 0.00937f
C1231 XA.XIR[11].XIC[14].icell.PDM Iout 0.00117f
C1232 XA.XIR[7].XIC[6].icell.PDM Iout 0.00117f
C1233 XA.XIR[2].XIC[13].icell.PUM VPWR 0.00937f
C1234 XA.XIR[2].XIC[2].icell.PDM VPWR 0.00799f
C1235 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.SM 0.00168f
C1236 XA.XIR[13].XIC[10].icell.PUM Vbias 0.0031f
C1237 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8] 0.00341f
C1238 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C1239 XA.XIR[8].XIC[12].icell.Ien Vbias 0.21098f
C1240 XA.XIR[7].XIC[9].icell.Ien VPWR 0.1903f
C1241 XA.XIR[11].XIC[9].icell.SM VPWR 0.00158f
C1242 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.15202f
C1243 XA.XIR[14].XIC_15.icell.PDM Iout 0.00133f
C1244 XA.XIR[0].XIC[2].icell.Ien Vbias 0.2113f
C1245 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.SM 0.00168f
C1246 XA.XIR[14].XIC_15.icell.Ien Iout 0.0642f
C1247 XA.XIR[7].XIC[5].icell.Ien Iout 0.06417f
C1248 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04031f
C1249 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.SM 0.00168f
C1250 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00584f
C1251 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.SM 0.0039f
C1252 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00584f
C1253 XThC.TAN2 XThC.Tn[10] 0.12148f
C1254 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C1255 XThR.Tn[4] XA.XIR[5].XIC[1].icell.SM 0.00121f
C1256 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.SM 0.00168f
C1257 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C1258 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.15202f
C1259 XThC.Tn[12] XThR.Tn[14] 0.28739f
C1260 XA.XIR[3].XIC[8].icell.PUM Vbias 0.0031f
C1261 XThR.Tn[7] XA.XIR[8].XIC[6].icell.Ien 0.00338f
C1262 XThR.Tn[3] XA.XIR[4].XIC[3].icell.SM 0.00121f
C1263 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C1264 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C1265 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.0353f
C1266 XThR.Tn[8] a_n997_3979# 0.1927f
C1267 XA.XIR[6].XIC[9].icell.SM Vbias 0.00701f
C1268 XA.XIR[0].XIC[9].icell.PUM VPWR 0.00877f
C1269 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02762f
C1270 XThC.TB4 data[2] 0.0086f
C1271 XThC.TA3 a_6243_9615# 0.02018f
C1272 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PUM 0.00186f
C1273 XA.XIR[4].XIC[6].icell.PDM Vbias 0.04261f
C1274 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00584f
C1275 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.03425f
C1276 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.SM 0.00168f
C1277 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00214f
C1278 XA.XIR[1].XIC[5].icell.PUM Vbias 0.0031f
C1279 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02762f
C1280 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Ien 0.00232f
C1281 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01734f
C1282 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.15202f
C1283 XThR.TB6 XThR.Tn[7] 0.01462f
C1284 XThR.TB6 a_n997_2891# 0.00466f
C1285 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PUM 0.00465f
C1286 XA.XIR[3].XIC[13].icell.SM VPWR 0.00158f
C1287 XA.XIR[13].XIC[11].icell.Ien Vbias 0.21098f
C1288 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02762f
C1289 XA.XIR[10].XIC[1].icell.Ien VPWR 0.1903f
C1290 XThR.Tn[3] Vbias 3.74868f
C1291 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.03425f
C1292 XThC.Tn[13] XThR.Tn[4] 0.2874f
C1293 XThR.Tn[10] XA.XIR[11].XIC[7].icell.Ien 0.00338f
C1294 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00214f
C1295 XThR.Tn[0] XA.XIR[0].XIC[12].icell.PDM 0.00341f
C1296 XA.XIR[3].XIC[9].icell.SM Iout 0.00388f
C1297 a_4067_9615# XThC.Tn[1] 0.00584f
C1298 XA.XIR[11].XIC[12].icell.PUM VPWR 0.00937f
C1299 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.15202f
C1300 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00584f
C1301 XA.XIR[6].XIC[14].icell.PDM VPWR 0.00809f
C1302 XThR.TA1 XThR.TA2 1.80461f
C1303 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.03425f
C1304 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C1305 XA.XIR[15].XIC[0].icell.SM Vbias 0.00675f
C1306 XA.XIR[6].XIC[12].icell.Ien Iout 0.06417f
C1307 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.SM 0.0039f
C1308 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.15202f
C1309 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.15202f
C1310 XA.XIR[6].XIC[2].icell.PDM Iout 0.00117f
C1311 XA.XIR[1].XIC[10].icell.SM VPWR 0.00158f
C1312 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C1313 XA.XIR[4].XIC[13].icell.PDM Iout 0.00117f
C1314 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00214f
C1315 XA.XIR[14].XIC[5].icell.PDM VPWR 0.00799f
C1316 XA.XIR[14].XIC[11].icell.SM VPWR 0.00158f
C1317 XA.XIR[1].XIC[6].icell.SM Iout 0.00388f
C1318 XA.XIR[11].XIC[1].icell.PDM Vbias 0.04261f
C1319 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PUM 0.00465f
C1320 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00584f
C1321 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C1322 XA.XIR[13].XIC[9].icell.PDM VPWR 0.00799f
C1323 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00214f
C1324 XThC.Tn[1] XThR.Tn[11] 0.28739f
C1325 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.15202f
C1326 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02762f
C1327 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.15202f
C1328 XA.XIR[10].XIC[5].icell.PDM Vbias 0.04261f
C1329 XThC.Tn[5] XThR.Tn[3] 0.28739f
C1330 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.03425f
C1331 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C1332 XA.XIR[2].XIC[1].icell.PUM VPWR 0.00937f
C1333 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.SM 0.00168f
C1334 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04031f
C1335 XA.XIR[9].XIC[3].icell.SM VPWR 0.00158f
C1336 XA.XIR[12].XIC[2].icell.PDM Iout 0.00117f
C1337 a_7651_9569# Vbias 0.00376f
C1338 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.SM 0.00168f
C1339 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C1340 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.15202f
C1341 XA.XIR[5].XIC[9].icell.PUM Vbias 0.0031f
C1342 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04052f
C1343 XThR.Tn[1] XA.XIR[2].XIC[13].icell.SM 0.00121f
C1344 XThR.TBN VPWR 4.54127f
C1345 XA.XIR[15].XIC[5].icell.SM Vbias 0.00701f
C1346 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PUM 0.00465f
C1347 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04031f
C1348 XThC.Tn[0] XThR.Tn[6] 0.28741f
C1349 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C1350 XThR.Tn[7] XThR.Tn[8] 0.07425f
C1351 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PUM 0.00465f
C1352 XA.XIR[11].XIC[13].icell.Ien VPWR 0.1903f
C1353 XA.XIR[11].XIC[8].icell.PDM Iout 0.00117f
C1354 XA.XIR[3].XIC[3].icell.PDM Vbias 0.04261f
C1355 XA.XIR[12].XIC[11].icell.PDM Vbias 0.04261f
C1356 XA.XIR[6].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1357 XThR.TAN2 XThR.Tn[12] 0.22096f
C1358 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.SM 0.0039f
C1359 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.03425f
C1360 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1361 XThR.Tn[0] XA.XIR[1].XIC[4].icell.SM 0.00121f
C1362 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00214f
C1363 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02762f
C1364 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.15202f
C1365 XA.XIR[2].XIC[3].icell.Ien VPWR 0.1903f
C1366 XThC.Tn[14] XThR.Tn[13] 0.28745f
C1367 XA.XIR[15].XIC[12].icell.PDM Vbias 0.04261f
C1368 XA.XIR[14].XIC[14].icell.PUM VPWR 0.00937f
C1369 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.SM 0.00168f
C1370 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02762f
C1371 XA.XIR[5].XIC[14].icell.SM VPWR 0.00207f
C1372 XThC.Tn[1] XThC.Tn[3] 0.10977f
C1373 XA.XIR[5].XIC[10].icell.PDM VPWR 0.00799f
C1374 XA.XIR[8].XIC[2].icell.SM Vbias 0.00701f
C1375 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.0355f
C1376 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00214f
C1377 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.SM 0.0039f
C1378 XThC.Tn[8] Iout 0.8379f
C1379 XThR.Tn[10] XThR.Tn[11] 0.05908f
C1380 XA.XIR[5].XIC[10].icell.SM Iout 0.00388f
C1381 XA.XIR[0].XIC[2].icell.PDM VPWR 0.00774f
C1382 XThR.TB3 a_n1049_6405# 0.00913f
C1383 XThC.Tn[8] XThR.Tn[9] 0.28739f
C1384 XThC.Tn[6] XThC.Tn[7] 0.1602f
C1385 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C1386 XA.XIR[15].XIC[8].icell.Ien Iout 0.06807f
C1387 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.SM 0.00168f
C1388 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.SM 0.00168f
C1389 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PUM 0.00465f
C1390 XA.XIR[8].XIC[12].icell.PDM VPWR 0.00799f
C1391 XA.XIR[3].XIC[10].icell.PDM Iout 0.00117f
C1392 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11115f
C1393 XA.XIR[14].XIC[5].icell.PUM VPWR 0.00937f
C1394 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13] 0.00341f
C1395 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[0].icell.SM 0.0039f
C1396 XThC.Tn[4] XThR.Tn[12] 0.28739f
C1397 XA.XIR[11].XIC[3].icell.Ien Vbias 0.21098f
C1398 XThC.Tn[13] XThR.Tn[8] 0.2874f
C1399 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C1400 XA.XIR[8].XIC[0].icell.PDM Iout 0.00117f
C1401 XThR.TA3 XThR.Tn[10] 0.00404f
C1402 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.SM 0.0039f
C1403 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04031f
C1404 XA.XIR[9].XIC[11].icell.SM Vbias 0.00701f
C1405 XA.XIR[13].XIC[7].icell.PUM VPWR 0.00937f
C1406 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04031f
C1407 XA.XIR[8].XIC[9].icell.Ien VPWR 0.1903f
C1408 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.SM 0.0039f
C1409 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C1410 XThR.TB7 XThR.Tn[14] 0.4222f
C1411 XA.XIR[10].XIC[5].icell.Ien Vbias 0.21098f
C1412 XA.XIR[11].XIC[14].icell.SM VPWR 0.00207f
C1413 XA.XIR[11].XIC[13].icell.PDM Iout 0.00117f
C1414 XA.XIR[12].XIC[7].icell.SM VPWR 0.00158f
C1415 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C1416 XThR.Tn[4] XA.XIR[4].XIC[1].icell.PDM 0.00341f
C1417 XThR.Tn[8] XA.XIR[9].XIC[5].icell.Ien 0.00338f
C1418 XA.XIR[8].XIC[5].icell.Ien Iout 0.06417f
C1419 XThR.Tn[5] a_n1049_5317# 0.00158f
C1420 XThR.Tn[3] XA.XIR[3].XIC[8].icell.PDM 0.00341f
C1421 XA.XIR[12].XIC[3].icell.SM Iout 0.00388f
C1422 XA.XIR[11].XIC[10].icell.PUM VPWR 0.00937f
C1423 XA.XIR[7].XIC[14].icell.PDM Vbias 0.04261f
C1424 XA.XIR[1].XIC[9].icell.PDM VPWR 0.00799f
C1425 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.SM 0.0039f
C1426 XThC.TB4 XThC.Tn[7] 0.01797f
C1427 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00214f
C1428 VPWR data[3] 0.20846f
C1429 XA.XIR[14].XIC[14].icell.PDM Iout 0.00117f
C1430 XThR.Tn[5] XA.XIR[6].XIC[14].icell.SM 0.00121f
C1431 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.15202f
C1432 XA.XIR[4].XIC[7].icell.Ien Vbias 0.21098f
C1433 XThC.Tn[0] XA.XIR[12].XIC_dummy_left.icell.Iout 0.00109f
C1434 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04031f
C1435 XA.XIR[3].XIC[5].icell.PUM VPWR 0.00937f
C1436 XA.XIR[2].XIC[11].icell.Ien Vbias 0.21098f
C1437 XThR.TA2 XThR.TB2 0.18237f
C1438 XThC.Tn[3] XThR.Tn[10] 0.28739f
C1439 XThR.Tn[2] XThR.Tn[3] 0.10553f
C1440 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00214f
C1441 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02762f
C1442 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.03425f
C1443 XThR.Tn[14] XA.XIR[15].XIC[7].icell.SM 0.00121f
C1444 XA.XIR[6].XIC[6].icell.SM VPWR 0.00158f
C1445 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.SM 0.0039f
C1446 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C1447 XA.XIR[9].XIC[14].icell.Ien Iout 0.06417f
C1448 XA.XIR[14].XIC[9].icell.SM VPWR 0.00158f
C1449 XA.XIR[7].XIC[7].icell.SM Vbias 0.00701f
C1450 XThC.Tn[13] XThR.Tn[1] 0.2874f
C1451 XA.XIR[10].XIC_15.icell.SM Vbias 0.00701f
C1452 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.15202f
C1453 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.0404f
C1454 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.03425f
C1455 XA.XIR[6].XIC[2].icell.SM Iout 0.00388f
C1456 XThC.TAN data[1] 0.00593f
C1457 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.SM 0.00168f
C1458 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00214f
C1459 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C1460 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PUM 0.00465f
C1461 XA.XIR[4].XIC[14].icell.PUM VPWR 0.00937f
C1462 XA.XIR[3].XIC[0].icell.SM Vbias 0.00675f
C1463 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04031f
C1464 XThR.Tn[13] XA.XIR[14].XIC[2].icell.Ien 0.00338f
C1465 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.SM 0.0039f
C1466 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00584f
C1467 XA.XIR[11].XIC[0].icell.PUM VPWR 0.00937f
C1468 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00584f
C1469 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C1470 XA.XIR[7].XIC[14].icell.Ien VPWR 0.19036f
C1471 XThR.Tn[0] XThR.TB2 0.00125f
C1472 a_n1049_5611# VPWR 0.71817f
C1473 XA.XIR[2].XIC[5].icell.PDM Iout 0.00117f
C1474 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.15202f
C1475 XA.XIR[0].XIC[7].icell.Ien Vbias 0.21134f
C1476 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02762f
C1477 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.15202f
C1478 XA.XIR[7].XIC[10].icell.Ien Iout 0.06417f
C1479 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00214f
C1480 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.03425f
C1481 XA.XIR[11].XIC[11].icell.Ien VPWR 0.1903f
C1482 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C1483 XThR.Tn[6] XA.XIR[7].XIC[4].icell.Ien 0.00338f
C1484 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.SM 0.00168f
C1485 XThR.TB6 a_n997_1579# 0.07626f
C1486 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PUM 0.00465f
C1487 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C1488 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00214f
C1489 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PUM 0.00465f
C1490 XThR.Tn[4] XA.XIR[5].XIC[6].icell.SM 0.00121f
C1491 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.03425f
C1492 XA.XIR[3].XIC[13].icell.PUM Vbias 0.0031f
C1493 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[5].icell.SM 0.0039f
C1494 XA.XIR[13].XIC[1].icell.Ien VPWR 0.1903f
C1495 XThR.Tn[7] XA.XIR[8].XIC[11].icell.Ien 0.00338f
C1496 XThR.Tn[3] XA.XIR[4].XIC[8].icell.SM 0.00121f
C1497 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.SM 0.0039f
C1498 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00584f
C1499 XA.XIR[14].XIC[12].icell.PUM VPWR 0.00937f
C1500 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00584f
C1501 XA.XIR[0].XIC[14].icell.PUM VPWR 0.00877f
C1502 XA.XIR[6].XIC[14].icell.SM Vbias 0.00701f
C1503 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04031f
C1504 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.03425f
C1505 XA.XIR[6].XIC[10].icell.PDM Vbias 0.04261f
C1506 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C1507 XA.XIR[8].XIC[0].icell.Ien Iout 0.06411f
C1508 XThR.Tn[8] XA.XIR[9].XIC[0].icell.Ien 0.00338f
C1509 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.SM 0.0039f
C1510 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5] 0.00341f
C1511 XThR.TAN2 data[7] 0.07741f
C1512 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.SM 0.0039f
C1513 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C1514 XA.XIR[1].XIC[10].icell.PUM Vbias 0.0031f
C1515 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C1516 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PUM 0.00465f
C1517 XA.XIR[14].XIC[1].icell.PDM Vbias 0.04261f
C1518 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.SM 0.00168f
C1519 XA.XIR[5].XIC[6].icell.PUM VPWR 0.00937f
C1520 XA.XIR[15].XIC[2].icell.SM VPWR 0.00158f
C1521 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C1522 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02762f
C1523 XThR.TA2 XThR.TAN2 0.0512f
C1524 XThC.Tn[1] XThR.Tn[14] 0.28739f
C1525 XA.XIR[13].XIC[5].icell.PDM Vbias 0.04261f
C1526 XThC.TB7 XThC.Tn[12] 0.07222f
C1527 XA.XIR[3].XIC[14].icell.SM Iout 0.00388f
C1528 XThC.TAN2 a_7651_9569# 0.02087f
C1529 XThC.TB3 XThC.TB6 0.04428f
C1530 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00214f
C1531 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.SM 0.0039f
C1532 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.03425f
C1533 XThR.TB2 a_n1049_7493# 0.02133f
C1534 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PUM 0.00429f
C1535 XA.XIR[12].XIC[10].icell.PDM Vbias 0.04261f
C1536 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.SM 0.0039f
C1537 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.15202f
C1538 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Iout 0.00347f
C1539 XA.XIR[15].XIC[2].icell.PDM Iout 0.00117f
C1540 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C1541 XThR.Tn[1] XA.XIR[1].XIC[13].icell.PDM 0.00341f
C1542 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C1543 a_8963_9569# XThC.Tn[11] 0.19413f
C1544 XA.XIR[9].XIC[3].icell.PUM Vbias 0.0031f
C1545 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00584f
C1546 XA.XIR[1].XIC[11].icell.SM Iout 0.00388f
C1547 XA.XIR[14].XIC[8].icell.PDM Iout 0.00117f
C1548 XA.XIR[15].XIC[11].icell.PDM Vbias 0.04261f
C1549 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02762f
C1550 XA.XIR[14].XIC[13].icell.Ien VPWR 0.19084f
C1551 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.15202f
C1552 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00584f
C1553 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.03425f
C1554 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00584f
C1555 XThC.Tn[2] XThR.Tn[4] 0.28739f
C1556 XA.XIR[9].XIC[12].icell.PDM VPWR 0.00799f
C1557 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.03425f
C1558 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C1559 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02762f
C1560 XA.XIR[9].XIC[0].icell.PDM Iout 0.00117f
C1561 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9] 0.00341f
C1562 XThR.Tn[12] XA.XIR[13].XIC[0].icell.Ien 0.00368f
C1563 XThC.Tn[12] VPWR 6.85795f
C1564 XA.XIR[9].XIC[8].icell.SM VPWR 0.00158f
C1565 XA.XIR[2].XIC[1].icell.SM Vbias 0.00701f
C1566 XA.XIR[10].XIC[2].icell.Ien VPWR 0.1903f
C1567 XThC.TB6 XThC.TB7 2.05133f
C1568 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.15202f
C1569 XA.XIR[5].XIC[14].icell.PUM Vbias 0.0031f
C1570 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[13].icell.Ien 0.00214f
C1571 XThR.TA1 XThR.TBN 0.00282f
C1572 XA.XIR[5].XIC[6].icell.PDM Vbias 0.04261f
C1573 XThR.Tn[11] XThR.Tn[13] 0.00153f
C1574 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.SM 0.00168f
C1575 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00214f
C1576 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C1577 XA.XIR[9].XIC[4].icell.SM Iout 0.00388f
C1578 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C1579 XThR.TB7 a_n1319_5317# 0.01283f
C1580 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04031f
C1581 XA.XIR[11].XIC[12].icell.PDM Iout 0.00117f
C1582 XThR.Tn[0] XA.XIR[1].XIC[9].icell.SM 0.00121f
C1583 XA.XIR[7].XIC[5].icell.PDM VPWR 0.00799f
C1584 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04031f
C1585 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00584f
C1586 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PUM 0.00465f
C1587 XA.XIR[8].XIC[8].icell.PDM Vbias 0.04261f
C1588 XA.XIR[6].XIC[1].icell.PUM Vbias 0.0031f
C1589 XA.XIR[14].XIC[3].icell.Ien Vbias 0.21098f
C1590 XThC.Tn[4] XThR.Tn[0] 0.28741f
C1591 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10] 0.00341f
C1592 XA.XIR[4].XIC[4].icell.Ien VPWR 0.1903f
C1593 a_n1049_7787# XThR.TB3 0.00124f
C1594 XA.XIR[2].XIC[8].icell.Ien VPWR 0.1903f
C1595 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.15202f
C1596 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14] 0.00341f
C1597 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00584f
C1598 XThR.TB4 XThR.Tn[3] 0.1895f
C1599 XThR.Tn[2] XA.XIR[3].XIC[0].icell.SM 0.00121f
C1600 XA.XIR[13].XIC[5].icell.Ien Vbias 0.21098f
C1601 XA.XIR[8].XIC[7].icell.SM Vbias 0.00701f
C1602 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C1603 XA.XIR[14].XIC[13].icell.PDM Iout 0.00117f
C1604 XA.XIR[14].XIC[14].icell.SM VPWR 0.00207f
C1605 XA.XIR[7].XIC[4].icell.SM VPWR 0.00158f
C1606 XA.XIR[2].XIC[4].icell.Ien Iout 0.06417f
C1607 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02762f
C1608 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00214f
C1609 XThC.TAN XThC.Tn[10] 0.14845f
C1610 XA.XIR[5].XIC[13].icell.PDM Iout 0.00117f
C1611 XA.XIR[12].XIC[7].icell.PUM Vbias 0.0031f
C1612 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02762f
C1613 XA.XIR[10].XIC_dummy_right.icell.PUM Vbias 0.00223f
C1614 XThC.TB6 VPWR 1.03148f
C1615 XA.XIR[14].XIC[10].icell.PUM VPWR 0.00937f
C1616 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C1617 XA.XIR[1].XIC[5].icell.PDM Vbias 0.04261f
C1618 XA.XIR[11].XIC[8].icell.Ien Vbias 0.21098f
C1619 XThC.TAN a_4861_9615# 0.0036f
C1620 XA.XIR[8].XIC_15.icell.PDM Iout 0.00133f
C1621 XA.XIR[1].XIC[2].icell.PUM VPWR 0.00937f
C1622 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C1623 XA.XIR[3].XIC[3].icell.Ien Vbias 0.21098f
C1624 XThC.Tn[3] XThR.Tn[13] 0.28739f
C1625 XA.XIR[8].XIC[14].icell.Ien VPWR 0.19036f
C1626 XThR.Tn[7] XA.XIR[8].XIC[1].icell.SM 0.00121f
C1627 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.SM 0.00168f
C1628 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C1629 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C1630 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18982f
C1631 XA.XIR[13].XIC_15.icell.SM Vbias 0.00701f
C1632 XA.XIR[6].XIC[6].icell.PUM Vbias 0.0031f
C1633 XA.XIR[8].XIC[10].icell.Ien Iout 0.06417f
C1634 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C1635 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38912f
C1636 XThR.Tn[8] XA.XIR[9].XIC[10].icell.Ien 0.00338f
C1637 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.03425f
C1638 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Iout 0.00347f
C1639 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.15202f
C1640 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04675f
C1641 XThC.Tn[6] Iout 0.83892f
C1642 XA.XIR[12].XIC[8].icell.SM Iout 0.00388f
C1643 XThC.Tn[6] XThR.Tn[9] 0.28739f
C1644 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02762f
C1645 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00214f
C1646 XA.XIR[4].XIC[12].icell.Ien Vbias 0.21098f
C1647 XThC.Tn[2] XThR.Tn[8] 0.28739f
C1648 XA.XIR[7].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1649 XA.XIR[3].XIC[10].icell.PUM VPWR 0.00937f
C1650 XA.XIR[1].XIC[12].icell.PDM Iout 0.00117f
C1651 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C1652 XA.XIR[2].XIC[13].icell.PDM Vbias 0.04261f
C1653 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02762f
C1654 XThR.Tn[10] XA.XIR[11].XIC[2].icell.SM 0.00121f
C1655 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.03425f
C1656 XA.XIR[6].XIC[11].icell.SM VPWR 0.00158f
C1657 XA.XIR[7].XIC[12].icell.SM Vbias 0.00701f
C1658 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PUM 0.00465f
C1659 XA.XIR[6].XIC[1].icell.PDM VPWR 0.00799f
C1660 XA.XIR[4].XIC[12].icell.PDM VPWR 0.00799f
C1661 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.SM 0.00168f
C1662 XA.XIR[6].XIC[7].icell.SM Iout 0.00388f
C1663 XA.XIR[14].XIC[11].icell.Ien VPWR 0.19084f
C1664 XA.XIR[1].XIC[7].icell.PUM VPWR 0.00937f
C1665 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7] 0.00341f
C1666 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C1667 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.15202f
C1668 XA.XIR[4].XIC[0].icell.PDM Iout 0.00117f
C1669 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.SM 0.0039f
C1670 a_5949_9615# Vbias 0.00634f
C1671 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C1672 XThR.Tn[13] XA.XIR[14].XIC[7].icell.Ien 0.00338f
C1673 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C1674 XThC.TB7 a_10915_9569# 0.06874f
C1675 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PDM 0.00172f
C1676 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.15202f
C1677 XThC.Tn[2] XThR.Tn[1] 0.28742f
C1678 XA.XIR[12].XIC[1].icell.PDM VPWR 0.00799f
C1679 XA.XIR[0].XIC[12].icell.Ien Vbias 0.2113f
C1680 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C1681 XA.XIR[7].XIC_15.icell.Ien Iout 0.0642f
C1682 XA.XIR[12].XIC[1].icell.Ien Vbias 0.21098f
C1683 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C1684 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04031f
C1685 XThR.Tn[6] XA.XIR[7].XIC[9].icell.Ien 0.00338f
C1686 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PUM 0.00471f
C1687 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C1688 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00584f
C1689 XThR.Tn[13] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00107f
C1690 XA.XIR[11].XIC[7].icell.PDM VPWR 0.00799f
C1691 XThR.TBN XThR.TB2 0.2075f
C1692 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00584f
C1693 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.SM 0.00168f
C1694 XThR.TB7 VPWR 1.14768f
C1695 XThR.Tn[4] XA.XIR[5].XIC[11].icell.SM 0.00121f
C1696 XA.XIR[5].XIC[4].icell.Ien Vbias 0.21098f
C1697 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04031f
C1698 XThR.Tn[3] XA.XIR[4].XIC[13].icell.SM 0.00121f
C1699 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.15202f
C1700 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C1701 a_5949_9615# XThC.Tn[5] 0.27124f
C1702 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PUM 0.00429f
C1703 XThC.TB2 XThC.Tn[2] 0.01113f
C1704 XA.XIR[15].XIC[10].icell.PDM Vbias 0.04261f
C1705 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PUM 0.00465f
C1706 XA.XIR[1].XIC_15.icell.PUM Vbias 0.0031f
C1707 a_10915_9569# VPWR 0.00307f
C1708 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PUM 0.00465f
C1709 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C1710 XA.XIR[5].XIC[11].icell.PUM VPWR 0.00937f
C1711 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.SM 0.0039f
C1712 XA.XIR[15].XIC[7].icell.SM VPWR 0.00158f
C1713 XA.XIR[3].XIC[9].icell.PDM VPWR 0.00799f
C1714 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.SM 0.0039f
C1715 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C1716 XThR.TB5 XThR.Tn[12] 0.32095f
C1717 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00584f
C1718 XA.XIR[15].XIC[3].icell.SM Iout 0.00388f
C1719 XA.XIR[9].XIC[8].icell.PDM Vbias 0.04261f
C1720 XThC.Tn[14] XThR.Tn[7] 0.28745f
C1721 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C1722 XThC.Tn[0] XA.XIR[15].XIC_dummy_left.icell.Iout 0.00109f
C1723 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00584f
C1724 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C1725 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.02762f
C1726 XThR.Tn[4] XThR.TB6 0.00264f
C1727 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00214f
C1728 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6] 0.00341f
C1729 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PDM 0.00555f
C1730 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.15202f
C1731 XA.XIR[13].XIC[2].icell.Ien VPWR 0.1903f
C1732 XA.XIR[11].XIC[11].icell.PDM Iout 0.00117f
C1733 XA.XIR[9].XIC[8].icell.PUM Vbias 0.0031f
C1734 XA.XIR[8].XIC[4].icell.SM VPWR 0.00158f
C1735 XThR.Tn[2] XA.XIR[3].XIC[3].icell.Ien 0.00338f
C1736 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.SM 0.00168f
C1737 XThR.Tn[13] XThR.Tn[14] 0.1554f
C1738 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C1739 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00584f
C1740 XA.XIR[12].XIC[4].icell.PUM VPWR 0.00937f
C1741 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C1742 XA.XIR[4].XIC[0].icell.Ien Iout 0.06411f
C1743 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C1744 XA.XIR[14].XIC[12].icell.PDM Iout 0.00117f
C1745 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00214f
C1746 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02762f
C1747 XThC.Tn[8] XThC.Tn[10] 0.00465f
C1748 XA.XIR[7].XIC[1].icell.PDM Vbias 0.04261f
C1749 XA.XIR[11].XIC[5].icell.Ien VPWR 0.1903f
C1750 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.SM 0.0039f
C1751 XA.XIR[9].XIC_15.icell.PDM Iout 0.00133f
C1752 XA.XIR[5].XIC_15.icell.SM VPWR 0.00275f
C1753 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04031f
C1754 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9] 0.00341f
C1755 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C1756 XA.XIR[4].XIC[2].icell.SM Vbias 0.00701f
C1757 XA.XIR[7].XIC[0].icell.SM Iout 0.00388f
C1758 XThC.TBN XThC.Tn[9] 0.49745f
C1759 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.15202f
C1760 XA.XIR[9].XIC[13].icell.SM VPWR 0.00158f
C1761 XA.XIR[10].XIC[7].icell.Ien VPWR 0.1903f
C1762 XThR.TBN XThR.TAN2 0.77119f
C1763 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02762f
C1764 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.SM 0.00168f
C1765 XThR.TB4 a_n1049_5317# 0.00463f
C1766 XA.XIR[2].XIC[6].icell.SM Vbias 0.00701f
C1767 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02762f
C1768 XThC.Tn[13] XThC.Tn[14] 0.38789f
C1769 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11] 0.00341f
C1770 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.SM 0.0039f
C1771 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C1772 XThR.Tn[2] XA.XIR[2].XIC[13].icell.PDM 0.00341f
C1773 XA.XIR[6].XIC[3].icell.PUM VPWR 0.00937f
C1774 XA.XIR[9].XIC[9].icell.SM Iout 0.00388f
C1775 XA.XIR[7].XIC[4].icell.PUM Vbias 0.0031f
C1776 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02762f
C1777 XA.XIR[10].XIC[3].icell.Ien Iout 0.06417f
C1778 XThR.Tn[9] XA.XIR[10].XIC[3].icell.Ien 0.00338f
C1779 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C1780 XA.XIR[0].XIC[13].icell.PDM Vbias 0.04282f
C1781 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.SM 0.0039f
C1782 XThR.TB1 XThR.TB3 0.04033f
C1783 XThR.TBN XThR.Tn[6] 0.59882f
C1784 XA.XIR[12].XIC[13].icell.SM Iout 0.00388f
C1785 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00214f
C1786 XThR.Tn[0] XA.XIR[1].XIC[14].icell.SM 0.00121f
C1787 XA.XIR[13].XIC_dummy_right.icell.PUM Vbias 0.00223f
C1788 XA.XIR[14].XIC[8].icell.Ien Vbias 0.21098f
C1789 XA.XIR[4].XIC[9].icell.Ien VPWR 0.1903f
C1790 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1791 XA.XIR[11].XIC_15.icell.SM VPWR 0.00275f
C1792 XA.XIR[7].XIC[8].icell.PDM Iout 0.00117f
C1793 XA.XIR[2].XIC[13].icell.Ien VPWR 0.1903f
C1794 XA.XIR[2].XIC[4].icell.PDM VPWR 0.00799f
C1795 XA.XIR[0].XIC[0].icell.Ien Iout 0.06382f
C1796 XA.XIR[4].XIC[5].icell.Ien Iout 0.06417f
C1797 XThC.Tn[1] VPWR 5.91915f
C1798 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C1799 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8] 0.00341f
C1800 XThR.TB2 a_n1049_5611# 0.00844f
C1801 XA.XIR[8].XIC[12].icell.SM Vbias 0.00701f
C1802 XA.XIR[2].XIC[9].icell.Ien Iout 0.06417f
C1803 XA.XIR[7].XIC[9].icell.SM VPWR 0.00158f
C1804 XA.XIR[0].XIC[2].icell.SM Vbias 0.00716f
C1805 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C1806 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.SM 0.0039f
C1807 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02762f
C1808 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C1809 XA.XIR[7].XIC[5].icell.SM Iout 0.00388f
C1810 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.15202f
C1811 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04031f
C1812 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02762f
C1813 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02762f
C1814 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.SM 0.0039f
C1815 XA.XIR[10].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1816 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C1817 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.04432f
C1818 XA.XIR[3].XIC[8].icell.Ien Vbias 0.21098f
C1819 XThR.Tn[7] XA.XIR[8].XIC[6].icell.SM 0.00121f
C1820 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.SM 0.0039f
C1821 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C1822 XA.XIR[0].XIC[9].icell.Ien VPWR 0.19115f
C1823 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.15202f
C1824 XA.XIR[6].XIC[11].icell.PUM Vbias 0.0031f
C1825 XThR.TB6 XThR.Tn[8] 0.02461f
C1826 XA.XIR[8].XIC_15.icell.Ien Iout 0.0642f
C1827 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C1828 XThR.Tn[8] XA.XIR[9].XIC_15.icell.Ien 0.00117f
C1829 XThR.Tn[11] XA.XIR[12].XIC[4].icell.Ien 0.00338f
C1830 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PUM 0.00465f
C1831 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PUM 0.00465f
C1832 XA.XIR[4].XIC[8].icell.PDM Vbias 0.04261f
C1833 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.15202f
C1834 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C1835 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C1836 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04052f
C1837 XA.XIR[0].XIC[5].icell.Ien Iout 0.06389f
C1838 XA.XIR[11].XIC[1].icell.PUM VPWR 0.00937f
C1839 XA.XIR[1].XIC[5].icell.Ien Vbias 0.21104f
C1840 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01577f
C1841 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02762f
C1842 XThC.TAN a_7651_9569# 0.01152f
C1843 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.03425f
C1844 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C1845 XThR.Tn[10] VPWR 7.53208f
C1846 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00214f
C1847 XThR.Tn[10] XA.XIR[11].XIC[7].icell.SM 0.00121f
C1848 XThR.Tn[0] XA.XIR[0].XIC[14].icell.PDM 0.00341f
C1849 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.04497f
C1850 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C1851 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1852 XA.XIR[15].XIC[1].icell.PDM VPWR 0.0114f
C1853 XA.XIR[15].XIC[2].icell.PUM Vbias 0.0031f
C1854 XThR.TB5 data[7] 0.00931f
C1855 XA.XIR[6].XIC[12].icell.SM Iout 0.00388f
C1856 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00584f
C1857 XA.XIR[1].XIC[12].icell.PUM VPWR 0.00937f
C1858 XA.XIR[6].XIC[4].icell.PDM Iout 0.00117f
C1859 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.SM 0.00168f
C1860 XA.XIR[4].XIC_15.icell.PDM Iout 0.00133f
C1861 XA.XIR[14].XIC[7].icell.PDM VPWR 0.00799f
C1862 XThR.Tn[1] XA.XIR[1].XIC[0].icell.PDM 0.00347f
C1863 XA.XIR[11].XIC[3].icell.PDM Vbias 0.04261f
C1864 XA.XIR[6].XIC_15.icell.SM Vbias 0.00701f
C1865 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00584f
C1866 XThC.Tn[0] XA.XIR[3].XIC_dummy_left.icell.Iout 0.00109f
C1867 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00214f
C1868 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.03425f
C1869 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PUM 0.0044f
C1870 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00256f
C1871 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.SM 0.00168f
C1872 XThR.TA2 XThR.TB5 0.01866f
C1873 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.15202f
C1874 XA.XIR[10].XIC[7].icell.PDM Vbias 0.04261f
C1875 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.SM 0.0039f
C1876 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C1877 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C1878 XThR.Tn[6] XA.XIR[7].XIC[14].icell.Ien 0.00338f
C1879 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00214f
C1880 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C1881 a_n1049_5611# XThR.Tn[6] 0.00158f
C1882 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.04036f
C1883 XThC.TB5 XThC.Tn[13] 0.00145f
C1884 XA.XIR[12].XIC[4].icell.PDM Iout 0.00117f
C1885 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PUM 0.00465f
C1886 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02762f
C1887 XThC.TB6 a_7875_9569# 0.0046f
C1888 XA.XIR[9].XIC[5].icell.PUM VPWR 0.00937f
C1889 XA.XIR[12].XIC[11].icell.SM Iout 0.00388f
C1890 a_8739_9569# Vbias 0.00278f
C1891 XA.XIR[3].XIC_15.icell.SM Iout 0.0047f
C1892 data[5] data[6] 0.01513f
C1893 XThR.TA1 XThR.TB7 0.00179f
C1894 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[10].icell.SM 0.0039f
C1895 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C1896 XA.XIR[5].XIC[9].icell.Ien Vbias 0.21098f
C1897 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PUM 0.00186f
C1898 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.03425f
C1899 XA.XIR[15].XIC[7].icell.PUM Vbias 0.0031f
C1900 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.03425f
C1901 XThC.Tn[11] XThR.Tn[5] 0.28739f
C1902 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.SM 0.0039f
C1903 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04031f
C1904 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00584f
C1905 XA.XIR[11].XIC[10].icell.PDM Iout 0.00117f
C1906 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.03425f
C1907 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02893f
C1908 XA.XIR[3].XIC[5].icell.PDM Vbias 0.04261f
C1909 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02762f
C1910 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01721f
C1911 XA.XIR[8].XIC[0].icell.SM Iout 0.00388f
C1912 XThR.Tn[8] XA.XIR[9].XIC[0].icell.SM 0.00121f
C1913 XA.XIR[2].XIC[3].icell.SM VPWR 0.00158f
C1914 XA.XIR[14].XIC[11].icell.PDM Iout 0.00117f
C1915 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C1916 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C1917 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1918 XA.XIR[5].XIC[12].icell.PDM VPWR 0.00799f
C1919 XA.XIR[8].XIC[4].icell.PUM Vbias 0.0031f
C1920 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PUM 0.00465f
C1921 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PUM 0.00465f
C1922 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02762f
C1923 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00584f
C1924 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04037f
C1925 XA.XIR[0].XIC[4].icell.PDM VPWR 0.00777f
C1926 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.SM 0.0039f
C1927 XThR.TA3 XThR.Tn[7] 0.00182f
C1928 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C1929 XA.XIR[12].XIC[2].icell.Ien Vbias 0.21098f
C1930 XA.XIR[15].XIC[8].icell.SM Iout 0.00388f
C1931 XA.XIR[5].XIC[0].icell.PDM Iout 0.00117f
C1932 a_n1049_8581# XThR.Tn[0] 0.2685f
C1933 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C1934 XThR.TA3 a_n997_2891# 0.00342f
C1935 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C1936 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00214f
C1937 XA.XIR[3].XIC[12].icell.PDM Iout 0.00117f
C1938 XA.XIR[8].XIC[14].icell.PDM VPWR 0.00809f
C1939 XA.XIR[14].XIC[5].icell.Ien VPWR 0.19084f
C1940 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13] 0.00341f
C1941 XA.XIR[11].XIC[3].icell.SM Vbias 0.00701f
C1942 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.15202f
C1943 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02762f
C1944 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C1945 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.03425f
C1946 XA.XIR[8].XIC[2].icell.PDM Iout 0.00117f
C1947 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04031f
C1948 XA.XIR[13].XIC[7].icell.Ien VPWR 0.1903f
C1949 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04031f
C1950 XA.XIR[9].XIC[13].icell.PUM Vbias 0.0031f
C1951 XA.XIR[10].XIC[5].icell.SM Vbias 0.00701f
C1952 XA.XIR[8].XIC[9].icell.SM VPWR 0.00158f
C1953 XThR.Tn[2] XA.XIR[3].XIC[8].icell.Ien 0.00338f
C1954 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1955 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1956 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Iout 0.00347f
C1957 XThC.Tn[8] XThR.Tn[3] 0.28739f
C1958 XA.XIR[13].XIC[3].icell.Ien Iout 0.06417f
C1959 XA.XIR[12].XIC[9].icell.PUM VPWR 0.00937f
C1960 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00584f
C1961 XA.XIR[8].XIC[5].icell.SM Iout 0.00388f
C1962 XThR.Tn[4] XA.XIR[4].XIC[3].icell.PDM 0.00341f
C1963 XThC.Tn[13] XThR.Tn[11] 0.2874f
C1964 XThC.TA3 Vbias 0.0149f
C1965 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00584f
C1966 XThR.Tn[8] XA.XIR[9].XIC[5].icell.SM 0.00121f
C1967 XThC.TB1 Vbias 0.01234f
C1968 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.15235f
C1969 XThR.Tn[3] XA.XIR[3].XIC[10].icell.PDM 0.00341f
C1970 XA.XIR[1].XIC[11].icell.PDM VPWR 0.00799f
C1971 XThC.Tn[3] XThR.Tn[7] 0.28739f
C1972 XThC.Tn[11] Vbias 2.46509f
C1973 a_n997_1803# VPWR 0.01991f
C1974 XA.XIR[14].XIC_15.icell.SM VPWR 0.00275f
C1975 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.SM 0.0039f
C1976 XA.XIR[3].XIC[5].icell.Ien VPWR 0.1903f
C1977 XA.XIR[4].XIC[7].icell.SM Vbias 0.00701f
C1978 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04031f
C1979 XA.XIR[2].XIC[11].icell.SM Vbias 0.00701f
C1980 XA.XIR[2].XIC[0].icell.PDM Vbias 0.04207f
C1981 XA.XIR[11].XIC[6].icell.Ien Iout 0.06417f
C1982 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01432f
C1983 XA.XIR[5].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1984 XThR.Tn[11] XA.XIR[12].XIC[12].icell.SM 0.00121f
C1985 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C1986 XThR.TB6 a_n997_3755# 0.0046f
C1987 XA.XIR[9].XIC[14].icell.SM Iout 0.00388f
C1988 XA.XIR[6].XIC[8].icell.PUM VPWR 0.00937f
C1989 XA.XIR[7].XIC[9].icell.PUM Vbias 0.0031f
C1990 XA.XIR[10].XIC[8].icell.Ien Iout 0.06417f
C1991 XThC.Tn[12] XThR.Tn[6] 0.28739f
C1992 XThR.Tn[9] XA.XIR[10].XIC[8].icell.Ien 0.00338f
C1993 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02762f
C1994 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PUM 0.00465f
C1995 XA.XIR[8].XIC[0].icell.PUM VPWR 0.00937f
C1996 XA.XIR[1].XIC[2].icell.Ien VPWR 0.1903f
C1997 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00584f
C1998 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.SM 0.00168f
C1999 XThC.TA3 XThC.Tn[5] 0.02758f
C2000 XA.XIR[4].XIC[14].icell.Ien VPWR 0.19036f
C2001 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.SM 0.0039f
C2002 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.03425f
C2003 XA.XIR[13].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2004 XA.XIR[3].XIC[2].icell.PUM Vbias 0.0031f
C2005 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04031f
C2006 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.04036f
C2007 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PUM 0.00465f
C2008 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.03425f
C2009 XThR.Tn[13] XA.XIR[14].XIC[2].icell.SM 0.00121f
C2010 a_7651_9569# XThC.Tn[8] 0.1927f
C2011 XA.XIR[4].XIC[10].icell.Ien Iout 0.06417f
C2012 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.SM 0.00168f
C2013 XA.XIR[2].XIC[14].icell.Ien Iout 0.06417f
C2014 XA.XIR[7].XIC[14].icell.SM VPWR 0.00207f
C2015 XA.XIR[5].XIC[1].icell.Ien VPWR 0.1903f
C2016 XA.XIR[2].XIC[7].icell.PDM Iout 0.00117f
C2017 XA.XIR[12].XIC[9].icell.SM Iout 0.00388f
C2018 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.SM 0.0039f
C2019 XThC.TBN XThC.Tn[7] 0.91493f
C2020 XA.XIR[0].XIC[7].icell.SM Vbias 0.00716f
C2021 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00214f
C2022 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02762f
C2023 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.SM 0.00168f
C2024 XA.XIR[7].XIC[10].icell.SM Iout 0.00388f
C2025 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C2026 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.15202f
C2027 XThR.Tn[6] XA.XIR[7].XIC[4].icell.SM 0.00121f
C2028 XA.XIR[14].XIC[0].icell.Ien VPWR 0.19084f
C2029 XThR.Tn[12] XA.XIR[13].XIC[6].icell.Ien 0.00338f
C2030 XThR.TB2 XThR.TB7 0.0437f
C2031 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.SM 0.0039f
C2032 XThC.TA2 XThC.TA3 0.44014f
C2033 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02762f
C2034 XThC.TB1 XThC.TA2 0.01609f
C2035 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.03425f
C2036 XThC.TA1 XThC.TA3 0.07824f
C2037 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00584f
C2038 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.03425f
C2039 XA.XIR[3].XIC[13].icell.Ien Vbias 0.21098f
C2040 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PUM 0.00186f
C2041 XThR.Tn[1] XA.XIR[2].XIC[5].icell.Ien 0.00338f
C2042 XThR.Tn[13] VPWR 7.61336f
C2043 XThR.Tn[7] XA.XIR[8].XIC[11].icell.SM 0.00121f
C2044 XThC.TA1 XThC.TB1 0.1098f
C2045 XA.XIR[10].XIC[1].icell.PUM Vbias 0.0031f
C2046 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04031f
C2047 XA.XIR[6].XIC_dummy_right.icell.PUM Vbias 0.00223f
C2048 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18971f
C2049 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Iout 0.00347f
C2050 XA.XIR[6].XIC[12].icell.PDM Vbias 0.04261f
C2051 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C2052 XThC.TB4 XThC.Tn[10] 0.01391f
C2053 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Iout 0.00347f
C2054 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C2055 XThR.Tn[11] XA.XIR[12].XIC[9].icell.Ien 0.00338f
C2056 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.15202f
C2057 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5] 0.00341f
C2058 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.SM 0.00168f
C2059 XA.XIR[0].XIC[10].icell.Ien Iout 0.06389f
C2060 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Ien 0.00584f
C2061 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C2062 XA.XIR[1].XIC[10].icell.Ien Vbias 0.21104f
C2063 XThR.TAN a_n1049_6405# 0.00268f
C2064 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.SM 0.00168f
C2065 XThC.TB6 XThC.Tn[4] 0.00264f
C2066 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00214f
C2067 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.03023f
C2068 XThC.TB4 a_4861_9615# 0.23756f
C2069 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C2070 XA.XIR[5].XIC[6].icell.Ien VPWR 0.1903f
C2071 XA.XIR[14].XIC[3].icell.PDM Vbias 0.04261f
C2072 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.15202f
C2073 XA.XIR[15].XIC[4].icell.PUM VPWR 0.00937f
C2074 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.15202f
C2075 XA.XIR[11].XIC[0].icell.SM Iout 0.00388f
C2076 XThR.Tn[5] XA.XIR[6].XIC[1].icell.Ien 0.00338f
C2077 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00214f
C2078 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C2079 XA.XIR[13].XIC[7].icell.PDM Vbias 0.04261f
C2080 XA.XIR[5].XIC[2].icell.Ien Iout 0.06417f
C2081 XThC.TAN2 a_8739_9569# 0.01719f
C2082 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02762f
C2083 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01746f
C2084 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.03529f
C2085 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00214f
C2086 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6] 0.00341f
C2087 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C2088 XA.XIR[15].XIC[4].icell.PDM Iout 0.00117f
C2089 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.SM 0.0039f
C2090 XThR.Tn[1] XA.XIR[1].XIC_15.icell.PDM 0.00341f
C2091 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02762f
C2092 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.SM 0.00168f
C2093 XA.XIR[9].XIC[3].icell.Ien Vbias 0.21098f
C2094 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00214f
C2095 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.SM 0.00168f
C2096 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02762f
C2097 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C2098 XA.XIR[14].XIC[10].icell.PDM Iout 0.00117f
C2099 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.15202f
C2100 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.03425f
C2101 XA.XIR[15].XIC[13].icell.SM Iout 0.00388f
C2102 XA.XIR[9].XIC[14].icell.PDM VPWR 0.00809f
C2103 a_7331_10587# data[0] 0.00451f
C2104 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C2105 XThR.Tn[11] XA.XIR[12].XIC[10].icell.SM 0.00121f
C2106 XA.XIR[7].XIC[1].icell.PUM VPWR 0.00937f
C2107 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00214f
C2108 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PDM 0.0059f
C2109 XThC.TBN a_3773_9615# 0.08456f
C2110 XA.XIR[9].XIC[2].icell.PDM Iout 0.00117f
C2111 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.15202f
C2112 XThC.Tn[11] XThR.Tn[2] 0.28739f
C2113 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9] 0.00341f
C2114 XThR.Tn[5] XA.XIR[6].XIC[6].icell.Ien 0.00338f
C2115 XA.XIR[9].XIC[10].icell.PUM VPWR 0.00937f
C2116 XThR.Tn[12] XA.XIR[13].XIC[0].icell.SM 0.00127f
C2117 XThR.TB7 XThR.TAN2 1.11559f
C2118 XA.XIR[2].XIC[3].icell.PUM Vbias 0.0031f
C2119 XA.XIR[10].XIC[2].icell.SM VPWR 0.00158f
C2120 XA.XIR[5].XIC[14].icell.Ien Vbias 0.21098f
C2121 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.SM 0.0039f
C2122 XThR.Tn[2] XA.XIR[2].XIC[0].icell.PDM 0.00347f
C2123 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C2124 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PUM 0.00465f
C2125 XA.XIR[5].XIC[8].icell.PDM Vbias 0.04261f
C2126 XA.XIR[12].XIC[13].icell.Ien Iout 0.06417f
C2127 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04031f
C2128 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02787f
C2129 XThR.TAN data[6] 0.07481f
C2130 XThR.TB7 XThR.Tn[6] 0.21438f
C2131 XA.XIR[0].XIC[0].icell.PDM Vbias 0.04227f
C2132 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04031f
C2133 XA.XIR[7].XIC[7].icell.PDM VPWR 0.00799f
C2134 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C2135 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.SM 0.0039f
C2136 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.03425f
C2137 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.03425f
C2138 XA.XIR[6].XIC[1].icell.Ien Vbias 0.21098f
C2139 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.SM 0.00168f
C2140 XA.XIR[8].XIC[10].icell.PDM Vbias 0.04261f
C2141 XA.XIR[4].XIC[4].icell.SM VPWR 0.00158f
C2142 XA.XIR[14].XIC[3].icell.SM Vbias 0.00701f
C2143 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10] 0.00341f
C2144 XThC.TA3 XThC.TAN2 0.197f
C2145 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C2146 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00214f
C2147 XA.XIR[2].XIC[8].icell.SM VPWR 0.00158f
C2148 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C2149 XThC.TB1 XThC.TAN2 0.12307f
C2150 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14] 0.00341f
C2151 XThR.TBN XThR.TB5 0.16186f
C2152 XA.XIR[13].XIC[5].icell.SM Vbias 0.00701f
C2153 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2154 XThC.TAN2 XThC.Tn[11] 0.12129f
C2155 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2156 XA.XIR[8].XIC[9].icell.PUM Vbias 0.0031f
C2157 XA.XIR[7].XIC[6].icell.PUM VPWR 0.00937f
C2158 XA.XIR[2].XIC[4].icell.SM Iout 0.00388f
C2159 XThR.TB3 a_n1049_6699# 0.0093f
C2160 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.SM 0.0039f
C2161 XThC.Tn[13] XThR.Tn[14] 0.2874f
C2162 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00214f
C2163 XA.XIR[12].XIC[7].icell.Ien Vbias 0.21098f
C2164 XThC.Tn[0] XThR.Tn[5] 0.28743f
C2165 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00584f
C2166 XA.XIR[5].XIC_15.icell.PDM Iout 0.00133f
C2167 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.SM 0.00168f
C2168 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00584f
C2169 XA.XIR[1].XIC[7].icell.PDM Vbias 0.04261f
C2170 XA.XIR[11].XIC[8].icell.SM Vbias 0.00701f
C2171 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Ien 0.00214f
C2172 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38997f
C2173 XThC.TAN a_5949_9615# 0.00927f
C2174 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00214f
C2175 XThR.TBN a_n1049_8581# 0.0607f
C2176 XA.XIR[14].XIC[6].icell.Ien Iout 0.06417f
C2177 XA.XIR[3].XIC[3].icell.SM Vbias 0.00701f
C2178 XThR.Tn[2] XA.XIR[3].XIC[13].icell.Ien 0.00338f
C2179 XA.XIR[8].XIC[14].icell.SM VPWR 0.00207f
C2180 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C2181 XA.XIR[12].XIC[14].icell.SM Iout 0.00388f
C2182 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.SM 0.00168f
C2183 XA.XIR[0].XIC[4].icell.SM VPWR 0.00158f
C2184 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04031f
C2185 XA.XIR[13].XIC[8].icell.Ien Iout 0.06417f
C2186 XA.XIR[6].XIC[6].icell.Ien Vbias 0.21098f
C2187 XThC.Tn[14] XThR.Tn[4] 0.28745f
C2188 XA.XIR[8].XIC[10].icell.SM Iout 0.00388f
C2189 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PUM 0.00465f
C2190 XThR.Tn[8] XA.XIR[9].XIC[10].icell.SM 0.00121f
C2191 a_4067_9615# XThC.Tn[2] 0.27699f
C2192 XThR.TB3 XThR.Tn[9] 0.00285f
C2193 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00214f
C2194 XThR.TB2 XThR.Tn[10] 0.00106f
C2195 XA.XIR[4].XIC[12].icell.SM Vbias 0.00701f
C2196 XA.XIR[3].XIC[10].icell.Ien VPWR 0.1903f
C2197 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C2198 XA.XIR[1].XIC[14].icell.PDM Iout 0.00117f
C2199 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PUM 0.00465f
C2200 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.SM 0.00168f
C2201 XA.XIR[2].XIC_15.icell.PDM Vbias 0.04401f
C2202 XA.XIR[14].XIC_dummy_left.icell.SM VPWR 0.00269f
C2203 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C2204 XThR.Tn[0] XA.XIR[0].XIC[1].icell.PDM 0.00341f
C2205 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02762f
C2206 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C2207 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.SM 0.0039f
C2208 XA.XIR[3].XIC[6].icell.Ien Iout 0.06417f
C2209 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.03425f
C2210 XA.XIR[6].XIC[3].icell.PDM VPWR 0.00799f
C2211 XA.XIR[6].XIC[13].icell.PUM VPWR 0.00937f
C2212 XA.XIR[7].XIC[14].icell.PUM Vbias 0.0031f
C2213 XThR.Tn[11] XA.XIR[12].XIC[14].icell.Ien 0.00338f
C2214 XA.XIR[4].XIC[14].icell.PDM VPWR 0.00809f
C2215 XA.XIR[5].XIC[1].icell.PUM Vbias 0.0031f
C2216 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PUM 0.00465f
C2217 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C2218 XThC.Tn[2] XThR.Tn[11] 0.28739f
C2219 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7] 0.00341f
C2220 XA.XIR[1].XIC[7].icell.Ien VPWR 0.1903f
C2221 XThC.Tn[6] XThR.Tn[3] 0.28739f
C2222 XA.XIR[15].XIC[11].icell.SM Iout 0.00388f
C2223 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C2224 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C2225 XA.XIR[4].XIC[2].icell.PDM Iout 0.00117f
C2226 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C2227 XThC.TB6 a_6243_9615# 0.01199f
C2228 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02834f
C2229 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C2230 XA.XIR[1].XIC[3].icell.Ien Iout 0.06417f
C2231 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PUM 0.00465f
C2232 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.SM 0.00168f
C2233 XThC.Tn[0] Vbias 1.91132f
C2234 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C2235 XThR.Tn[13] XA.XIR[14].XIC[7].icell.SM 0.00121f
C2236 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.SM 0.00168f
C2237 XA.XIR[4].XIC_15.icell.Ien Iout 0.0642f
C2238 XA.XIR[13].XIC[1].icell.PUM Vbias 0.0031f
C2239 XA.XIR[0].XIC[12].icell.SM Vbias 0.00716f
C2240 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.SM 0.00168f
C2241 XA.XIR[12].XIC[3].icell.PDM VPWR 0.00799f
C2242 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04031f
C2243 XThR.Tn[12] Vbias 3.74784f
C2244 XThC.Tn[1] XThR.Tn[6] 0.28739f
C2245 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.03431f
C2246 XThR.Tn[6] XA.XIR[7].XIC[9].icell.SM 0.00121f
C2247 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.SM 0.0039f
C2248 XA.XIR[12].XIC[11].icell.Ien Iout 0.06417f
C2249 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02762f
C2250 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.04036f
C2251 XA.XIR[11].XIC[9].icell.PDM VPWR 0.00799f
C2252 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C2253 XThR.TA2 a_n1319_5611# 0.00467f
C2254 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04031f
C2255 XA.XIR[5].XIC[4].icell.SM Vbias 0.00701f
C2256 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02762f
C2257 XThR.Tn[1] XA.XIR[2].XIC[10].icell.Ien 0.00338f
C2258 XA.XIR[14].XIC[0].icell.SM Iout 0.00388f
C2259 XA.XIR[15].XIC[2].icell.Ien Vbias 0.17899f
C2260 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PUM 0.00186f
C2261 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02762f
C2262 XThR.TB5 a_n1049_5611# 0.0093f
C2263 XThC.Tn[2] XThC.Tn[3] 0.33669f
C2264 XA.XIR[4].XIC[0].icell.PUM VPWR 0.00937f
C2265 XThC.Tn[9] Iout 0.83793f
C2266 XThC.Tn[9] XThR.Tn[9] 0.28739f
C2267 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02762f
C2268 XA.XIR[10].XIC[1].icell.PDM Iout 0.00117f
C2269 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.SM 0.00168f
C2270 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04031f
C2271 XA.XIR[0].XIC_15.icell.Ien Iout 0.06388f
C2272 XA.XIR[1].XIC_15.icell.Ien Vbias 0.2124f
C2273 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.03425f
C2274 XThC.TBN Iout 0.00167f
C2275 XThC.Tn[5] XThR.Tn[12] 0.28739f
C2276 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.03425f
C2277 XThC.Tn[14] XThR.Tn[8] 0.28745f
C2278 XA.XIR[5].XIC[11].icell.Ien VPWR 0.1903f
C2279 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PUM 0.00465f
C2280 XThR.TAN2 XThR.Tn[10] 0.12147f
C2281 XA.XIR[15].XIC[9].icell.PUM VPWR 0.00937f
C2282 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C2283 XA.XIR[3].XIC[11].icell.PDM VPWR 0.00799f
C2284 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00214f
C2285 XA.XIR[5].XIC[7].icell.Ien Iout 0.06417f
C2286 XA.XIR[9].XIC[10].icell.PDM Vbias 0.04261f
C2287 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.SM 0.0039f
C2288 XThR.TAN XThR.TB3 0.23315f
C2289 a_n1319_6405# VPWR 0.00676f
C2290 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C2291 XA.XIR[8].XIC[1].icell.PDM VPWR 0.00799f
C2292 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00584f
C2293 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.15202f
C2294 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02762f
C2295 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02762f
C2296 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00214f
C2297 XA.XIR[13].XIC[2].icell.SM VPWR 0.00158f
C2298 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.SM 0.0039f
C2299 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C2300 XThC.TB4 a_7651_9569# 0.00497f
C2301 XA.XIR[9].XIC[8].icell.Ien Vbias 0.21098f
C2302 XA.XIR[8].XIC[6].icell.PUM VPWR 0.00937f
C2303 XThR.Tn[2] XA.XIR[3].XIC[3].icell.SM 0.00121f
C2304 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00214f
C2305 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C2306 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00214f
C2307 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02762f
C2308 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.SM 0.0039f
C2309 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.SM 0.00168f
C2310 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.15202f
C2311 XA.XIR[12].XIC[4].icell.Ien VPWR 0.1903f
C2312 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12] 0.00341f
C2313 XThC.Tn[4] XThR.Tn[10] 0.28739f
C2314 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.SM 0.00168f
C2315 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C2316 XA.XIR[4].XIC[0].icell.SM Iout 0.00388f
C2317 XThC.Tn[14] XThR.Tn[1] 0.28745f
C2318 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C2319 XA.XIR[7].XIC[3].icell.PDM Vbias 0.04261f
C2320 XA.XIR[11].XIC[13].icell.SM Vbias 0.00701f
C2321 XThR.Tn[8] data[4] 0.01643f
C2322 XA.XIR[11].XIC[5].icell.SM VPWR 0.00158f
C2323 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.SM 0.0039f
C2324 XThR.Tn[5] XA.XIR[6].XIC[11].icell.Ien 0.00338f
C2325 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.15202f
C2326 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04031f
C2327 a_n997_3979# VPWR 0.01662f
C2328 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00214f
C2329 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.03023f
C2330 XThR.Tn[11] XA.XIR[12].XIC[12].icell.Ien 0.00338f
C2331 XA.XIR[4].XIC[4].icell.PUM Vbias 0.0031f
C2332 XThR.TA2 XThR.Tn[5] 0.00361f
C2333 XA.XIR[2].XIC[8].icell.PUM Vbias 0.0031f
C2334 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.04617f
C2335 XA.XIR[11].XIC[1].icell.SM Iout 0.00388f
C2336 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01577f
C2337 XA.XIR[10].XIC[7].icell.SM VPWR 0.00158f
C2338 XA.XIR[15].XIC[9].icell.SM Iout 0.00388f
C2339 XThR.Tn[2] XA.XIR[2].XIC_15.icell.PDM 0.00341f
C2340 XThR.Tn[14] XA.XIR[15].XIC[4].icell.Ien 0.00338f
C2341 XA.XIR[6].XIC[3].icell.Ien VPWR 0.1903f
C2342 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2343 XA.XIR[10].XIC[3].icell.SM Iout 0.00388f
C2344 XA.XIR[7].XIC[4].icell.Ien Vbias 0.21098f
C2345 XThR.Tn[9] XA.XIR[10].XIC[3].icell.SM 0.00121f
C2346 XThR.Tn[3] XA.XIR[4].XIC[0].icell.Ien 0.00338f
C2347 XA.XIR[0].XIC_15.icell.PDM Vbias 0.04438f
C2348 XThC.Tn[0] XA.XIR[10].XIC_dummy_left.icell.Iout 0.00109f
C2349 XThR.TB6 a_n997_2667# 0.00468f
C2350 XA.XIR[14].XIC[8].icell.SM Vbias 0.00701f
C2351 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04031f
C2352 XA.XIR[4].XIC[9].icell.SM VPWR 0.00158f
C2353 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C2354 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C2355 XA.XIR[2].XIC[13].icell.SM VPWR 0.00158f
C2356 XA.XIR[7].XIC[10].icell.PDM Iout 0.00117f
C2357 XThC.Tn[0] XThR.Tn[2] 0.28748f
C2358 XA.XIR[0].XIC[0].icell.SM Iout 0.00367f
C2359 XA.XIR[2].XIC[6].icell.PDM VPWR 0.00799f
C2360 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.SM 0.00168f
C2361 XA.XIR[1].XIC[0].icell.SM Vbias 0.00679f
C2362 XA.XIR[4].XIC[5].icell.SM Iout 0.00388f
C2363 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8] 0.00341f
C2364 XA.XIR[8].XIC[14].icell.PUM Vbias 0.0031f
C2365 XA.XIR[2].XIC[9].icell.SM Iout 0.00388f
C2366 XA.XIR[7].XIC[11].icell.PUM VPWR 0.00937f
C2367 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.SM 0.0039f
C2368 XA.XIR[0].XIC[4].icell.PUM Vbias 0.0031f
C2369 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.SM 0.0039f
C2370 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.SM 0.00168f
C2371 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00214f
C2372 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04031f
C2373 XThR.Tn[12] XA.XIR[13].XIC[1].icell.SM 0.00121f
C2374 a_7331_10587# VPWR 0.0063f
C2375 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.SM 0.00168f
C2376 XA.XIR[9].XIC_15.icell.SM Iout 0.0047f
C2377 XThR.Tn[4] XA.XIR[5].XIC[3].icell.Ien 0.00338f
C2378 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00214f
C2379 XA.XIR[3].XIC[8].icell.SM Vbias 0.00701f
C2380 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[4].icell.Ien 0.00214f
C2381 XThC.Tn[6] XA.XIR[0].XIC[7].icell.Ien 0.002f
C2382 XThR.Tn[3] XA.XIR[4].XIC[5].icell.Ien 0.00338f
C2383 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.15202f
C2384 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.SM 0.0039f
C2385 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00214f
C2386 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.SM 0.0039f
C2387 XA.XIR[8].XIC[1].icell.PUM VPWR 0.00937f
C2388 XThR.TA3 XThR.Tn[4] 0.02736f
C2389 XA.XIR[6].XIC[11].icell.Ien Vbias 0.21098f
C2390 XA.XIR[0].XIC[9].icell.SM VPWR 0.00158f
C2391 XThC.Tn[2] XThR.Tn[14] 0.28739f
C2392 XA.XIR[4].XIC[10].icell.PDM Vbias 0.04261f
C2393 XThR.Tn[11] XA.XIR[12].XIC[4].icell.SM 0.00121f
C2394 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.03425f
C2395 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.SM 0.00168f
C2396 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02809f
C2397 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.03425f
C2398 XThC.TB7 XThC.Tn[13] 0.11626f
C2399 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02762f
C2400 XThR.Tn[7] VPWR 6.97893f
C2401 XThR.TAN2 a_n997_1803# 0.09118f
C2402 XA.XIR[0].XIC[5].icell.SM Iout 0.00367f
C2403 XA.XIR[1].XIC[5].icell.SM Vbias 0.00704f
C2404 a_n997_2891# VPWR 0.01347f
C2405 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.SM 0.0039f
C2406 XA.XIR[5].XIC[1].icell.SM VPWR 0.00158f
C2407 XThR.TB6 XThR.Tn[11] 0.02465f
C2408 XA.XIR[7].XIC_15.icell.SM VPWR 0.00275f
C2409 XA.XIR[3].XIC_15.icell.Ien VPWR 0.25566f
C2410 XThC.TAN a_8739_9569# 0.0168f
C2411 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10] 0.00341f
C2412 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PUM 0.00465f
C2413 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.PDM 0.00591f
C2414 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C2415 XA.XIR[3].XIC[11].icell.Ien Iout 0.06417f
C2416 XA.XIR[2].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2417 XThR.TA3 XThR.TB6 0.19112f
C2418 XA.XIR[15].XIC[3].icell.PDM VPWR 0.0114f
C2419 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Iout 0.00347f
C2420 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02762f
C2421 XThC.Tn[3] XThR.Tn[4] 0.28739f
C2422 XThR.Tn[0] Vbias 3.75791f
C2423 XA.XIR[1].XIC[12].icell.Ien VPWR 0.1903f
C2424 XA.XIR[6].XIC[6].icell.PDM Iout 0.00117f
C2425 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.3891f
C2426 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C2427 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C2428 XThR.Tn[1] XA.XIR[1].XIC[2].icell.PDM 0.00341f
C2429 XA.XIR[14].XIC[9].icell.PDM VPWR 0.00799f
C2430 XThR.Tn[0] XA.XIR[1].XIC[1].icell.Ien 0.00338f
C2431 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02762f
C2432 XA.XIR[11].XIC[5].icell.PDM Vbias 0.04261f
C2433 XA.XIR[1].XIC[8].icell.Ien Iout 0.06417f
C2434 XA.XIR[15].XIC[13].icell.Ien Iout 0.06807f
C2435 XA.XIR[11].XIC[11].icell.SM Vbias 0.00701f
C2436 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.03554f
C2437 XThC.Tn[13] VPWR 6.87751f
C2438 XThR.Tn[11] XA.XIR[12].XIC[10].icell.Ien 0.00338f
C2439 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C2440 XA.XIR[10].XIC[9].icell.PDM Vbias 0.04261f
C2441 XA.XIR[9].XIC[1].icell.PDM VPWR 0.00799f
C2442 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00214f
C2443 XA.XIR[13].XIC[1].icell.PDM Iout 0.00117f
C2444 XThR.Tn[5] XA.XIR[6].XIC[1].icell.SM 0.00121f
C2445 XThR.Tn[6] XA.XIR[7].XIC[14].icell.SM 0.00121f
C2446 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.SM 0.00168f
C2447 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PDM 0.00172f
C2448 XThR.TAN XThR.TB1 1.61695f
C2449 XA.XIR[12].XIC[6].icell.PDM Iout 0.00117f
C2450 XThC.TB6 a_8963_9569# 0.00468f
C2451 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2452 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.03425f
C2453 XA.XIR[9].XIC[5].icell.Ien VPWR 0.1903f
C2454 XA.XIR[12].XIC[12].icell.SM VPWR 0.00158f
C2455 XThR.TAN2 XThR.Tn[13] 0.00106f
C2456 a_9827_9569# Vbias 0.00491f
C2457 XThC.Tn[5] XThR.Tn[0] 0.28744f
C2458 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.03425f
C2459 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00584f
C2460 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C2461 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00584f
C2462 XThR.Tn[1] XA.XIR[2].XIC_15.icell.Ien 0.00117f
C2463 XA.XIR[15].XIC[7].icell.Ien Vbias 0.17899f
C2464 XA.XIR[5].XIC[9].icell.SM Vbias 0.00701f
C2465 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04031f
C2466 XA.XIR[3].XIC[7].icell.PDM Vbias 0.04261f
C2467 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02762f
C2468 XThC.TA3 XThC.TAN 0.35844f
C2469 XThR.Tn[0] XA.XIR[1].XIC[6].icell.Ien 0.00338f
C2470 XThC.TB1 XThC.TAN 1.61695f
C2471 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00584f
C2472 XThC.TB2 XThC.TB5 0.0451f
C2473 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02762f
C2474 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02762f
C2475 XThC.TAN XThC.Tn[11] 0.03903f
C2476 XThR.Tn[14] XA.XIR[15].XIC[12].icell.SM 0.00121f
C2477 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PUM 0.00465f
C2478 XThR.TB5 XThR.TB7 0.036f
C2479 XA.XIR[2].XIC[5].icell.PUM VPWR 0.00937f
C2480 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02762f
C2481 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.15202f
C2482 XA.XIR[15].XIC[14].icell.SM Iout 0.00388f
C2483 XA.XIR[11].XIC[14].icell.PUM Vbias 0.0031f
C2484 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.SM 0.00168f
C2485 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2486 XA.XIR[5].XIC[14].icell.PDM VPWR 0.00809f
C2487 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.03425f
C2488 XA.XIR[8].XIC[4].icell.Ien Vbias 0.21098f
C2489 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.03425f
C2490 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C2491 XThC.Tn[4] XThR.Tn[13] 0.28739f
C2492 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04031f
C2493 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.0353f
C2494 XA.XIR[0].XIC[6].icell.PDM VPWR 0.0078f
C2495 XA.XIR[12].XIC[2].icell.SM Vbias 0.00701f
C2496 XA.XIR[5].XIC[12].icell.Ien Iout 0.06417f
C2497 XA.XIR[5].XIC[2].icell.PDM Iout 0.00117f
C2498 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.SM 0.00168f
C2499 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2500 XA.XIR[3].XIC[14].icell.PDM Iout 0.00117f
C2501 XA.XIR[14].XIC[13].icell.SM Vbias 0.00701f
C2502 XA.XIR[14].XIC[5].icell.SM VPWR 0.00158f
C2503 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13] 0.00341f
C2504 XA.XIR[11].XIC[5].icell.PUM Vbias 0.0031f
C2505 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02762f
C2506 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C2507 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00584f
C2508 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C2509 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01577f
C2510 XA.XIR[8].XIC[4].icell.PDM Iout 0.00117f
C2511 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.SM 0.00168f
C2512 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00584f
C2513 XA.XIR[14].XIC[1].icell.SM Iout 0.00388f
C2514 XThC.Tn[7] Iout 0.84037f
C2515 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04031f
C2516 XA.XIR[13].XIC[7].icell.SM VPWR 0.00158f
C2517 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00584f
C2518 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04031f
C2519 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00214f
C2520 XThC.TB2 a_4067_9615# 0.02133f
C2521 XThC.Tn[7] XThR.Tn[9] 0.28739f
C2522 XA.XIR[9].XIC[13].icell.Ien Vbias 0.21098f
C2523 XA.XIR[10].XIC[7].icell.PUM Vbias 0.0031f
C2524 XThR.Tn[2] XA.XIR[3].XIC[8].icell.SM 0.00121f
C2525 XA.XIR[8].XIC[11].icell.PUM VPWR 0.00937f
C2526 XThC.Tn[3] XThR.Tn[8] 0.28739f
C2527 XA.XIR[13].XIC[3].icell.SM Iout 0.00388f
C2528 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PUM 0.00465f
C2529 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.SM 0.00168f
C2530 XA.XIR[6].XIC[1].icell.SM Vbias 0.00701f
C2531 XA.XIR[12].XIC[9].icell.Ien VPWR 0.1903f
C2532 XThR.Tn[4] XA.XIR[4].XIC[5].icell.PDM 0.00341f
C2533 XThR.TB4 XThR.Tn[12] 0.00209f
C2534 XThC.Tn[0] XA.XIR[13].XIC_dummy_left.icell.Iout 0.00109f
C2535 XThR.Tn[3] XA.XIR[3].XIC[12].icell.PDM 0.00341f
C2536 XA.XIR[12].XIC[5].icell.Ien Iout 0.06417f
C2537 XA.XIR[1].XIC[13].icell.PDM VPWR 0.00799f
C2538 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PUM 0.00186f
C2539 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.SM 0.00168f
C2540 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04052f
C2541 XA.XIR[4].XIC[9].icell.PUM Vbias 0.0031f
C2542 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00214f
C2543 XA.XIR[3].XIC[5].icell.SM VPWR 0.00158f
C2544 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PUM 0.00465f
C2545 XA.XIR[11].XIC[6].icell.SM Iout 0.00388f
C2546 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PUM 0.00465f
C2547 XThR.Tn[3] a_n1049_6405# 0.00542f
C2548 XA.XIR[1].XIC[1].icell.PDM Iout 0.00117f
C2549 XA.XIR[2].XIC[13].icell.PUM Vbias 0.0031f
C2550 XA.XIR[2].XIC[2].icell.PDM Vbias 0.04261f
C2551 XA.XIR[9].XIC[0].icell.Ien VPWR 0.1903f
C2552 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PUM 0.00465f
C2553 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C2554 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.SM 0.00168f
C2555 XA.XIR[3].XIC[1].icell.SM Iout 0.00388f
C2556 XThR.Tn[14] XA.XIR[15].XIC[9].icell.Ien 0.00338f
C2557 XA.XIR[6].XIC[8].icell.Ien VPWR 0.1903f
C2558 XA.XIR[10].XIC[8].icell.SM Iout 0.00388f
C2559 XA.XIR[7].XIC[9].icell.Ien Vbias 0.21098f
C2560 XA.XIR[11].XIC[9].icell.SM Vbias 0.00701f
C2561 XThR.Tn[9] XA.XIR[10].XIC[8].icell.SM 0.00121f
C2562 XThR.Tn[1] XA.XIR[2].XIC[0].icell.SM 0.00121f
C2563 XA.XIR[15].XIC[11].icell.Ien Iout 0.06807f
C2564 XA.XIR[4].XIC[1].icell.PDM VPWR 0.00799f
C2565 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.SM 0.0039f
C2566 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01757f
C2567 XA.XIR[6].XIC[4].icell.Ien Iout 0.06417f
C2568 XThR.Tn[0] XThR.Tn[2] 0.00536f
C2569 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7] 0.00341f
C2570 XA.XIR[1].XIC[2].icell.SM VPWR 0.00158f
C2571 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C2572 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00214f
C2573 XA.XIR[4].XIC[14].icell.SM VPWR 0.00207f
C2574 XThC.Tn[3] XThR.Tn[1] 0.28739f
C2575 XA.XIR[8].XIC_15.icell.SM VPWR 0.00275f
C2576 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00214f
C2577 XThC.TB7 a_6243_10571# 0.01283f
C2578 XA.XIR[12].XIC_15.icell.SM Iout 0.0047f
C2579 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04031f
C2580 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00584f
C2581 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PUM 0.00465f
C2582 XA.XIR[4].XIC[10].icell.SM Iout 0.00388f
C2583 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C2584 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C2585 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2586 XA.XIR[2].XIC[14].icell.SM Iout 0.00388f
C2587 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.15202f
C2588 XA.XIR[2].XIC[9].icell.PDM Iout 0.00117f
C2589 XA.XIR[12].XIC[10].icell.SM VPWR 0.00158f
C2590 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11117f
C2591 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02762f
C2592 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10] 0.00341f
C2593 XA.XIR[0].XIC[9].icell.PUM Vbias 0.0031f
C2594 a_5949_9615# XThC.Tn[6] 0.0018f
C2595 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C2596 XThR.TBN XThR.Tn[5] 0.59912f
C2597 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.SM 0.00168f
C2598 a_n997_1579# VPWR 0.02417f
C2599 XThR.Tn[12] XA.XIR[13].XIC[6].icell.SM 0.00121f
C2600 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.SM 0.00168f
C2601 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C2602 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00584f
C2603 XThR.TB6 XThR.Tn[14] 0.00128f
C2604 XThR.Tn[4] XA.XIR[5].XIC[8].icell.Ien 0.00338f
C2605 XA.XIR[3].XIC[13].icell.SM Vbias 0.00701f
C2606 XThR.Tn[11] XA.XIR[12].XIC_15.icell.Ien 0.00117f
C2607 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C2608 XThR.Tn[1] XA.XIR[2].XIC[5].icell.SM 0.00121f
C2609 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2610 XThC.TB3 XThC.Tn[2] 0.1864f
C2611 XThR.Tn[14] XA.XIR[15].XIC[10].icell.SM 0.00121f
C2612 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.15202f
C2613 XThR.Tn[3] XA.XIR[4].XIC[10].icell.Ien 0.00338f
C2614 data[1] data[2] 0.01393f
C2615 XA.XIR[10].XIC[0].icell.PDM VPWR 0.00799f
C2616 XA.XIR[10].XIC[1].icell.Ien Vbias 0.21098f
C2617 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C2618 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04031f
C2619 XA.XIR[11].XIC[12].icell.PUM Vbias 0.0031f
C2620 XA.XIR[0].XIC[14].icell.SM VPWR 0.00207f
C2621 a_6243_10571# VPWR 0.00653f
C2622 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C2623 XA.XIR[6].XIC[14].icell.PDM Vbias 0.04261f
C2624 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.03425f
C2625 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5] 0.00341f
C2626 XA.XIR[0].XIC[10].icell.SM Iout 0.00367f
C2627 XA.XIR[1].XIC[10].icell.SM Vbias 0.00704f
C2628 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C2629 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02762f
C2630 XA.XIR[14].XIC[5].icell.PDM Vbias 0.04261f
C2631 a_n1049_7493# XThR.Tn[2] 0.26564f
C2632 XThC.TB4 a_5949_9615# 0.00465f
C2633 XA.XIR[5].XIC[6].icell.SM VPWR 0.00158f
C2634 XA.XIR[14].XIC[11].icell.SM Vbias 0.00701f
C2635 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00214f
C2636 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.SM 0.00168f
C2637 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C2638 XA.XIR[15].XIC[4].icell.Ien VPWR 0.32895f
C2639 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.04563f
C2640 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00214f
C2641 XA.XIR[13].XIC[9].icell.PDM Vbias 0.04261f
C2642 XA.XIR[3].XIC_dummy_right.icell.SM VPWR 0.00123f
C2643 XA.XIR[12].XIC[13].icell.PUM VPWR 0.00937f
C2644 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.SM 0.0039f
C2645 XA.XIR[5].XIC[2].icell.SM Iout 0.00388f
C2646 XThC.TAN2 a_9827_9569# 0.09118f
C2647 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.SM 0.00168f
C2648 XA.XIR[9].XIC[1].icell.Ien Iout 0.06417f
C2649 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.15202f
C2650 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PUM 0.00465f
C2651 XThC.TB1 XThC.Tn[8] 0.29191f
C2652 XA.XIR[2].XIC[1].icell.PUM Vbias 0.0031f
C2653 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6] 0.00341f
C2654 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C2655 XA.XIR[15].XIC[6].icell.PDM Iout 0.00117f
C2656 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C2657 XThC.Tn[9] XThC.Tn[10] 0.07959f
C2658 XA.XIR[1].XIC[13].icell.Ien Iout 0.06417f
C2659 XA.XIR[9].XIC[3].icell.SM Vbias 0.00701f
C2660 XThR.TB5 XThR.Tn[10] 0.01742f
C2661 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C2662 XA.XIR[4].XIC[1].icell.PUM VPWR 0.00937f
C2663 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.SM 0.0039f
C2664 XThC.TBN XThC.Tn[10] 0.51405f
C2665 XThR.TBN Vbias 0.00722f
C2666 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00584f
C2667 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02762f
C2668 XA.XIR[11].XIC[13].icell.Ien Vbias 0.21098f
C2669 XA.XIR[1].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2670 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2671 XA.XIR[7].XIC[1].icell.Ien VPWR 0.1903f
C2672 XThR.TB2 a_n997_3979# 0.00191f
C2673 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00584f
C2674 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.15202f
C2675 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00214f
C2676 XThC.TBN a_4861_9615# 0.07601f
C2677 XA.XIR[9].XIC[4].icell.PDM Iout 0.00117f
C2678 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PUM 0.00465f
C2679 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.SM 0.0039f
C2680 XThR.Tn[5] XA.XIR[6].XIC[6].icell.SM 0.00121f
C2681 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.15202f
C2682 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9] 0.00341f
C2683 XA.XIR[9].XIC[10].icell.Ien VPWR 0.1903f
C2684 XA.XIR[14].XIC[14].icell.PUM Vbias 0.0031f
C2685 XA.XIR[2].XIC[3].icell.Ien Vbias 0.21098f
C2686 XA.XIR[10].XIC[4].icell.PUM VPWR 0.00937f
C2687 XA.XIR[5].XIC[14].icell.SM Vbias 0.00701f
C2688 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.SM 0.0039f
C2689 XA.XIR[5].XIC[10].icell.PDM Vbias 0.04261f
C2690 XThR.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.00341f
C2691 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.03425f
C2692 XA.XIR[9].XIC[6].icell.Ien Iout 0.06417f
C2693 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.0353f
C2694 XA.XIR[12].XIC[14].icell.Ien VPWR 0.19036f
C2695 XThR.TA2 XThR.TB4 0.04137f
C2696 XThC.Tn[2] VPWR 5.93664f
C2697 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.15202f
C2698 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02762f
C2699 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00214f
C2700 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04031f
C2701 XA.XIR[0].XIC[2].icell.PDM Vbias 0.04282f
C2702 XA.XIR[7].XIC[9].icell.PDM VPWR 0.00799f
C2703 XThR.Tn[0] XA.XIR[1].XIC[11].icell.Ien 0.00338f
C2704 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04031f
C2705 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C2706 XA.XIR[8].XIC[12].icell.PDM Vbias 0.04261f
C2707 XA.XIR[14].XIC[5].icell.PUM Vbias 0.0031f
C2708 XA.XIR[0].XIC[1].icell.PUM VPWR 0.00877f
C2709 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10] 0.00341f
C2710 XA.XIR[4].XIC[6].icell.PUM VPWR 0.00937f
C2711 XThR.Tn[5] a_n1049_5611# 0.27042f
C2712 XA.XIR[2].XIC[10].icell.PUM VPWR 0.00937f
C2713 XA.XIR[13].XIC[7].icell.PUM Vbias 0.0031f
C2714 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00584f
C2715 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C2716 XThR.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.00338f
C2717 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00584f
C2718 XA.XIR[8].XIC[9].icell.Ien Vbias 0.21098f
C2719 XA.XIR[7].XIC[6].icell.Ien VPWR 0.1903f
C2720 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00584f
C2721 XA.XIR[10].XIC[13].icell.SM Iout 0.00388f
C2722 XA.XIR[9].XIC_dummy_left.icell.SM VPWR 0.00269f
C2723 XThR.Tn[9] XA.XIR[10].XIC[13].icell.SM 0.00121f
C2724 XA.XIR[11].XIC[14].icell.SM Vbias 0.00701f
C2725 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PUM 0.00429f
C2726 XA.XIR[12].XIC[7].icell.SM Vbias 0.00701f
C2727 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00214f
C2728 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C2729 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.SM 0.0039f
C2730 XA.XIR[7].XIC[2].icell.Ien Iout 0.06417f
C2731 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00584f
C2732 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C2733 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C2734 XA.XIR[11].XIC[10].icell.PUM Vbias 0.0031f
C2735 XA.XIR[1].XIC[9].icell.PDM Vbias 0.04261f
C2736 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.03425f
C2737 XA.XIR[14].XIC[6].icell.SM Iout 0.00388f
C2738 XThC.TAN XThC.Tn[0] 0.00139f
C2739 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00214f
C2740 XA.XIR[3].XIC[5].icell.PUM Vbias 0.0031f
C2741 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2742 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PUM 0.00465f
C2743 XThR.Tn[2] XA.XIR[3].XIC[13].icell.SM 0.00121f
C2744 XThR.Tn[7] XA.XIR[8].XIC[3].icell.Ien 0.00338f
C2745 XA.XIR[12].XIC_15.icell.PDM Iout 0.00133f
C2746 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.SM 0.00168f
C2747 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00214f
C2748 XA.XIR[13].XIC[8].icell.SM Iout 0.00388f
C2749 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C2750 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.SM 0.0039f
C2751 XA.XIR[0].XIC[6].icell.PUM VPWR 0.00877f
C2752 XA.XIR[14].XIC[9].icell.SM Vbias 0.00701f
C2753 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C2754 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02762f
C2755 XA.XIR[6].XIC[6].icell.SM Vbias 0.00701f
C2756 XThC.TB2 data[0] 0.00267f
C2757 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02762f
C2758 XThR.TAN data[5] 0.00593f
C2759 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00214f
C2760 XThR.TAN2 a_n997_3979# 0.02087f
C2761 XA.XIR[12].XIC[11].icell.PUM VPWR 0.00937f
C2762 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10] 0.00341f
C2763 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.15202f
C2764 XA.XIR[4].XIC[14].icell.PUM Vbias 0.0031f
C2765 XA.XIR[3].XIC[10].icell.SM VPWR 0.00158f
C2766 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.SM 0.0039f
C2767 XThR.Tn[10] XA.XIR[11].XIC[4].icell.Ien 0.00338f
C2768 XA.XIR[6].XIC[13].icell.Ien VPWR 0.1903f
C2769 XA.XIR[3].XIC[6].icell.SM Iout 0.00388f
C2770 XThR.Tn[0] XA.XIR[0].XIC[3].icell.PDM 0.00341f
C2771 XA.XIR[6].XIC[5].icell.PDM VPWR 0.00799f
C2772 XA.XIR[7].XIC[14].icell.Ien Vbias 0.21098f
C2773 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PUM 0.00465f
C2774 XThR.Tn[9] Iout 1.16233f
C2775 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2776 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.15202f
C2777 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.SM 0.00168f
C2778 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.03425f
C2779 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Ien 0.00584f
C2780 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2781 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7] 0.00341f
C2782 XA.XIR[6].XIC[9].icell.Ien Iout 0.06417f
C2783 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.15202f
C2784 XA.XIR[1].XIC[7].icell.SM VPWR 0.00158f
C2785 XA.XIR[15].XIC[12].icell.SM VPWR 0.00158f
C2786 XThR.TB5 a_n997_1803# 0.06458f
C2787 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C2788 XA.XIR[4].XIC[4].icell.PDM Iout 0.00117f
C2789 XThR.TB3 XThR.Tn[3] 0.01287f
C2790 XA.XIR[11].XIC[11].icell.Ien Vbias 0.21098f
C2791 XThR.TBN XA.XIR[10].XIC_dummy_left.icell.Iout 0.00376f
C2792 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.SM 0.00168f
C2793 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C2794 XA.XIR[1].XIC[3].icell.SM Iout 0.00388f
C2795 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13] 0.00341f
C2796 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C2797 XA.XIR[13].XIC[0].icell.PDM VPWR 0.00799f
C2798 XThC.TBN XA.XIR[0].XIC[11].icell.PDM 0.00104f
C2799 XA.XIR[13].XIC[1].icell.Ien Vbias 0.21098f
C2800 XThC.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.00109f
C2801 XThR.TBN XThR.Tn[2] 0.6189f
C2802 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.15202f
C2803 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.15202f
C2804 XA.XIR[14].XIC[12].icell.PUM Vbias 0.0031f
C2805 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02762f
C2806 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00584f
C2807 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.SM 0.0039f
C2808 XA.XIR[0].XIC[14].icell.PUM Vbias 0.0031f
C2809 XThC.Tn[12] XThR.Tn[5] 0.28739f
C2810 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C2811 XA.XIR[12].XIC[5].icell.PDM VPWR 0.00799f
C2812 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04031f
C2813 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C2814 XA.XIR[12].XIC[12].icell.Ien VPWR 0.1903f
C2815 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2816 XA.XIR[15].XIC[0].icell.Ien Iout 0.06801f
C2817 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02762f
C2818 XThR.Tn[1] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00122f
C2819 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04031f
C2820 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.SM 0.00168f
C2821 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PUM 0.00465f
C2822 XThR.Tn[4] XA.XIR[5].XIC[13].icell.Ien 0.00338f
C2823 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.15202f
C2824 XThR.Tn[1] XA.XIR[2].XIC[10].icell.SM 0.00121f
C2825 XA.XIR[5].XIC[6].icell.PUM Vbias 0.0031f
C2826 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04031f
C2827 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[9].icell.Ien 0.00214f
C2828 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.SM 0.00168f
C2829 XA.XIR[15].XIC[2].icell.SM Vbias 0.00701f
C2830 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00214f
C2831 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.SM 0.0039f
C2832 XThR.Tn[3] XA.XIR[4].XIC_15.icell.Ien 0.00117f
C2833 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PUM 0.00465f
C2834 XA.XIR[8].XIC[1].icell.Ien VPWR 0.1903f
C2835 XThR.Tn[14] XA.XIR[15].XIC[12].icell.Ien 0.00338f
C2836 XThR.Tn[0] XA.XIR[1].XIC[1].icell.SM 0.00121f
C2837 XThR.TAN2 XThR.Tn[7] 0.01439f
C2838 XA.XIR[10].XIC[3].icell.PDM Iout 0.00117f
C2839 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04031f
C2840 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00584f
C2841 XA.XIR[10].XIC[11].icell.SM Iout 0.00388f
C2842 XThR.TAN a_n1049_6699# 0.0036f
C2843 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01577f
C2844 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00584f
C2845 XThR.TAN2 a_n997_2891# 0.01719f
C2846 XThR.Tn[9] XA.XIR[10].XIC[11].icell.SM 0.00121f
C2847 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00584f
C2848 XA.XIR[5].XIC[11].icell.SM VPWR 0.00158f
C2849 XThR.TB5 XThR.Tn[13] 0.00145f
C2850 XA.XIR[5].XIC[1].icell.PDM VPWR 0.00799f
C2851 XA.XIR[15].XIC[9].icell.Ien VPWR 0.32895f
C2852 XThR.Tn[6] XThR.Tn[7] 0.06617f
C2853 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.03425f
C2854 XA.XIR[3].XIC[13].icell.PDM VPWR 0.00799f
C2855 XA.XIR[14].XIC[13].icell.Ien Vbias 0.21098f
C2856 XA.XIR[15].XIC[5].icell.Ien Iout 0.06807f
C2857 XA.XIR[5].XIC[7].icell.SM Iout 0.00388f
C2858 XA.XIR[9].XIC[12].icell.PDM Vbias 0.04261f
C2859 XA.XIR[8].XIC[3].icell.PDM VPWR 0.00799f
C2860 XThC.Tn[9] XThR.Tn[3] 0.28739f
C2861 XA.XIR[3].XIC[1].icell.PDM Iout 0.00117f
C2862 XThC.Tn[14] XThR.Tn[11] 0.28745f
C2863 XThR.Tn[4] VPWR 6.61651f
C2864 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C2865 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.15202f
C2866 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.SM 0.0039f
C2867 XThC.Tn[4] XThR.Tn[7] 0.28739f
C2868 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00214f
C2869 XA.XIR[13].XIC[4].icell.PUM VPWR 0.00937f
C2870 XThC.Tn[12] Vbias 2.48611f
C2871 XThC.TB4 a_8739_9569# 0.00813f
C2872 XA.XIR[9].XIC[8].icell.SM Vbias 0.00701f
C2873 XA.XIR[8].XIC[6].icell.Ien VPWR 0.1903f
C2874 XA.XIR[10].XIC[2].icell.Ien Vbias 0.21098f
C2875 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.SM 0.00168f
C2876 XThR.TAN XThR.Tn[9] 0.0565f
C2877 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C2878 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C2879 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12] 0.00341f
C2880 XA.XIR[12].XIC[4].icell.SM VPWR 0.00158f
C2881 XA.XIR[8].XIC[2].icell.Ien Iout 0.06417f
C2882 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PUM 0.00471f
C2883 XThR.Tn[8] XA.XIR[9].XIC[2].icell.Ien 0.00338f
C2884 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C2885 XA.XIR[15].XIC_15.icell.SM Iout 0.0047f
C2886 XA.XIR[7].XIC[5].icell.PDM Vbias 0.04261f
C2887 XThC.Tn[13] XThR.Tn[6] 0.2874f
C2888 XA.XIR[1].XIC[0].icell.PDM VPWR 0.00799f
C2889 XA.XIR[11].XIC[7].icell.PUM VPWR 0.00937f
C2890 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04031f
C2891 XThR.Tn[5] XA.XIR[6].XIC[11].icell.SM 0.00121f
C2892 XThR.TB6 VPWR 1.05512f
C2893 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00214f
C2894 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PUM 0.00465f
C2895 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.15202f
C2896 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02812f
C2897 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C2898 XA.XIR[4].XIC[4].icell.Ien Vbias 0.21098f
C2899 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04031f
C2900 XA.XIR[9].XIC_15.icell.Ien VPWR 0.25566f
C2901 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00256f
C2902 XA.XIR[2].XIC[8].icell.Ien Vbias 0.21098f
C2903 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00584f
C2904 XThC.TA3 XThC.Tn[6] 0.10589f
C2905 XA.XIR[10].XIC[9].icell.PUM VPWR 0.00937f
C2906 XA.XIR[15].XIC[10].icell.SM VPWR 0.00158f
C2907 XA.XIR[6].XIC[3].icell.SM VPWR 0.00158f
C2908 XThR.Tn[14] XA.XIR[15].XIC[4].icell.SM 0.00121f
C2909 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C2910 XA.XIR[13].XIC[13].icell.SM Iout 0.00388f
C2911 XA.XIR[14].XIC[14].icell.SM Vbias 0.00701f
C2912 XA.XIR[9].XIC[11].icell.Ien Iout 0.06417f
C2913 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.15202f
C2914 XThC.TAN2 data[3] 0.07741f
C2915 XA.XIR[7].XIC[4].icell.SM Vbias 0.00701f
C2916 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[1].icell.SM 0.0039f
C2917 XThR.Tn[3] XA.XIR[4].XIC[0].icell.SM 0.00121f
C2918 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PUM 0.00465f
C2919 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.SM 0.0039f
C2920 XA.XIR[12].XIC[14].icell.PDM Iout 0.00117f
C2921 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PUM 0.00465f
C2922 XA.XIR[14].XIC[10].icell.PUM Vbias 0.0031f
C2923 XThC.TBN a_7651_9569# 0.23021f
C2924 XThC.Tn[8] XThR.Tn[12] 0.28739f
C2925 XA.XIR[4].XIC[11].icell.PUM VPWR 0.00937f
C2926 XThR.Tn[10] XA.XIR[11].XIC[12].icell.SM 0.00121f
C2927 XThR.TA3 data[4] 0.8689f
C2928 XThC.TB6 Vbias 0.01776f
C2929 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.SM 0.0039f
C2930 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02762f
C2931 XA.XIR[7].XIC[12].icell.PDM Iout 0.00117f
C2932 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01577f
C2933 XA.XIR[12].XIC[10].icell.Ien VPWR 0.1903f
C2934 XA.XIR[2].XIC[8].icell.PDM VPWR 0.00799f
C2935 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C2936 XA.XIR[15].XIC_15.icell.PDM Iout 0.00133f
C2937 XA.XIR[1].XIC[2].icell.PUM Vbias 0.0031f
C2938 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10] 0.00341f
C2939 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02762f
C2940 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8] 0.00341f
C2941 XA.XIR[7].XIC[11].icell.Ien VPWR 0.1903f
C2942 XA.XIR[8].XIC[14].icell.Ien Vbias 0.21098f
C2943 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.SM 0.00168f
C2944 XThC.TA3 XThC.TB4 0.14536f
C2945 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.SM 0.0039f
C2946 XA.XIR[0].XIC[4].icell.Ien Vbias 0.21127f
C2947 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C2948 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C2949 XThC.TB1 XThC.TB4 0.05121f
C2950 XThC.TB2 XThC.TB3 2.04808f
C2951 XA.XIR[11].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2952 XA.XIR[7].XIC[7].icell.Ien Iout 0.06417f
C2953 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04031f
C2954 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.03425f
C2955 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00584f
C2956 XThC.TB4 XThC.Tn[11] 0.30582f
C2957 a_2979_9615# VPWR 0.70527f
C2958 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.SM 0.00168f
C2959 XThR.Tn[14] XA.XIR[15].XIC[10].icell.Ien 0.00338f
C2960 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00584f
C2961 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2962 XThR.Tn[4] XA.XIR[5].XIC[3].icell.SM 0.00121f
C2963 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C2964 XA.XIR[10].XIC[9].icell.SM Iout 0.00388f
C2965 XA.XIR[3].XIC[10].icell.PUM Vbias 0.0031f
C2966 XA.XIR[15].XIC[13].icell.PUM VPWR 0.00937f
C2967 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00584f
C2968 XThR.Tn[9] XA.XIR[10].XIC[9].icell.SM 0.00121f
C2969 XThR.TBN XThR.TB4 0.15627f
C2970 XThC.TB6 XThC.Tn[5] 0.20189f
C2971 XThR.Tn[3] XA.XIR[4].XIC[5].icell.SM 0.00121f
C2972 XThR.Tn[7] XA.XIR[8].XIC[8].icell.Ien 0.00338f
C2973 XThR.Tn[8] VPWR 7.51456f
C2974 XA.XIR[3].XIC[0].icell.Ien Iout 0.06411f
C2975 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.03425f
C2976 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C2977 XA.XIR[6].XIC[11].icell.SM Vbias 0.00701f
C2978 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13] 0.00341f
C2979 XA.XIR[0].XIC[11].icell.PUM VPWR 0.00878f
C2980 XA.XIR[6].XIC[1].icell.PDM Vbias 0.04261f
C2981 XA.XIR[4].XIC_15.icell.SM VPWR 0.00275f
C2982 XA.XIR[4].XIC[12].icell.PDM Vbias 0.04261f
C2983 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2984 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C2985 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C2986 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02762f
C2987 XA.XIR[14].XIC[11].icell.Ien Vbias 0.21098f
C2988 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C2989 XA.XIR[1].XIC[7].icell.PUM Vbias 0.0031f
C2990 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PUM 0.00186f
C2991 XThR.TBN XA.XIR[13].XIC_dummy_left.icell.Iout 0.00446f
C2992 XA.XIR[11].XIC[1].icell.Ien VPWR 0.1903f
C2993 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.15202f
C2994 XThR.TB3 a_n1049_5317# 0.00899f
C2995 XA.XIR[2].XIC_15.icell.SM Iout 0.0047f
C2996 XA.XIR[5].XIC[3].icell.PUM VPWR 0.00937f
C2997 XThC.TAN a_9827_9569# 0.00228f
C2998 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02762f
C2999 XThC.TB2 XThC.TB7 0.0437f
C3000 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.03425f
C3001 XA.XIR[9].XIC[0].icell.SM VPWR 0.00158f
C3002 a_10051_9569# XThC.Tn[12] 0.00623f
C3003 XThR.Tn[10] XA.XIR[11].XIC[9].icell.Ien 0.00338f
C3004 XThC.TA2 XThC.TB6 0.10153f
C3005 XA.XIR[3].XIC[11].icell.SM Iout 0.00388f
C3006 XThC.TA1 XThC.TB6 0.00193f
C3007 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00214f
C3008 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00584f
C3009 XA.XIR[1].XIC[0].icell.Ien VPWR 0.1903f
C3010 XThR.Tn[14] a_n997_715# 0.1927f
C3011 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C3012 XA.XIR[15].XIC[5].icell.PDM VPWR 0.0114f
C3013 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00584f
C3014 XA.XIR[12].XIC[1].icell.PDM Vbias 0.04261f
C3015 XThR.Tn[11] a_n997_2667# 0.19413f
C3016 XA.XIR[6].XIC[14].icell.Ien Iout 0.06417f
C3017 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.15202f
C3018 XA.XIR[1].XIC[12].icell.SM VPWR 0.00158f
C3019 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.SM 0.00168f
C3020 XA.XIR[6].XIC[8].icell.PDM Iout 0.00117f
C3021 XThR.Tn[1] VPWR 6.67344f
C3022 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00214f
C3023 XThR.Tn[1] XA.XIR[1].XIC[4].icell.PDM 0.00341f
C3024 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C3025 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C3026 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.SM 0.0039f
C3027 XA.XIR[11].XIC[7].icell.PDM Vbias 0.04261f
C3028 XA.XIR[15].XIC[14].icell.Ien VPWR 0.329f
C3029 XA.XIR[1].XIC[8].icell.SM Iout 0.00388f
C3030 XA.XIR[0].XIC_15.icell.SM VPWR 0.00257f
C3031 XThC.Tn[12] XThR.Tn[2] 0.28739f
C3032 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PUM 0.00465f
C3033 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00214f
C3034 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00584f
C3035 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C3036 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.15202f
C3037 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.15202f
C3038 XA.XIR[9].XIC[3].icell.PDM VPWR 0.00799f
C3039 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.03425f
C3040 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C3041 XA.XIR[13].XIC[3].icell.PDM Iout 0.00117f
C3042 XA.XIR[13].XIC[11].icell.SM Iout 0.00388f
C3043 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02762f
C3044 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.SM 0.0039f
C3045 XThR.TAN2 a_n997_1579# 0.00199f
C3046 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C3047 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.SM 0.00168f
C3048 XThC.TB2 VPWR 0.97668f
C3049 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PUM 0.00102f
C3050 XA.XIR[12].XIC[8].icell.PDM Iout 0.00117f
C3051 XA.XIR[9].XIC[5].icell.SM VPWR 0.00158f
C3052 XThC.TB6 a_10051_9569# 0.07626f
C3053 a_10915_9569# Vbias 0.01295f
C3054 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.15202f
C3055 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C3056 XA.XIR[5].XIC[11].icell.PUM Vbias 0.0031f
C3057 XThR.Tn[10] XA.XIR[11].XIC[10].icell.SM 0.00121f
C3058 XA.XIR[15].XIC[7].icell.SM Vbias 0.00701f
C3059 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04031f
C3060 XA.XIR[9].XIC[1].icell.SM Iout 0.00388f
C3061 XA.XIR[3].XIC[9].icell.PDM Vbias 0.04261f
C3062 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PUM 0.00465f
C3063 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.SM 0.0039f
C3064 XThC.TAN2 XThC.Tn[12] 0.22686f
C3065 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.SM 0.00168f
C3066 XThC.Tn[14] XThR.Tn[14] 0.28745f
C3067 XThR.Tn[0] XA.XIR[1].XIC[6].icell.SM 0.00121f
C3068 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00214f
C3069 XThC.Tn[1] XThR.Tn[5] 0.28739f
C3070 XThR.Tn[11] XA.XIR[12].XIC[0].icell.Ien 0.0037f
C3071 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C3072 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.03425f
C3073 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.SM 0.00168f
C3074 XA.XIR[2].XIC[5].icell.Ien VPWR 0.1903f
C3075 XA.XIR[10].XIC[13].icell.Ien Iout 0.06417f
C3076 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Iout 0.00347f
C3077 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3078 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C3079 XThR.Tn[9] XA.XIR[10].XIC[13].icell.Ien 0.00338f
C3080 XA.XIR[13].XIC[2].icell.Ien Vbias 0.21098f
C3081 a_n1049_7493# XA.XIR[1].XIC_dummy_left.icell.Iout 0.0013f
C3082 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3083 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.SM 0.0039f
C3084 XA.XIR[7].XIC[1].icell.SM VPWR 0.00158f
C3085 XA.XIR[8].XIC[4].icell.SM Vbias 0.00701f
C3086 XA.XIR[5].XIC[12].icell.SM Iout 0.00388f
C3087 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04031f
C3088 XThR.TB4 a_n1049_5611# 0.00465f
C3089 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01093f
C3090 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00214f
C3091 XA.XIR[12].XIC[4].icell.PUM Vbias 0.0031f
C3092 XA.XIR[15].XIC[11].icell.PUM VPWR 0.00937f
C3093 XA.XIR[5].XIC[4].icell.PDM Iout 0.00117f
C3094 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C3095 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13] 0.00341f
C3096 XA.XIR[14].XIC[7].icell.PUM VPWR 0.00937f
C3097 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02762f
C3098 XA.XIR[11].XIC[5].icell.Ien Vbias 0.21098f
C3099 XA.XIR[5].XIC_15.icell.SM Vbias 0.00701f
C3100 XA.XIR[12].XIC[13].icell.PDM Iout 0.00117f
C3101 XA.XIR[12].XIC_15.icell.Ien VPWR 0.25566f
C3102 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C3103 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PUM 0.00441f
C3104 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.SM 0.0039f
C3105 XA.XIR[8].XIC[6].icell.PDM Iout 0.00117f
C3106 XThC.TB2 a_5155_9615# 0.00847f
C3107 XA.XIR[13].XIC[9].icell.PUM VPWR 0.00937f
C3108 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04031f
C3109 XA.XIR[8].XIC[11].icell.Ien VPWR 0.1903f
C3110 XA.XIR[9].XIC[13].icell.SM Vbias 0.00701f
C3111 XThC.TAN2 XThC.TB6 0.06405f
C3112 XA.XIR[10].XIC[7].icell.Ien Vbias 0.21098f
C3113 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.SM 0.0039f
C3114 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.03023f
C3115 XA.XIR[6].XIC[3].icell.PUM Vbias 0.0031f
C3116 XA.XIR[8].XIC[7].icell.Ien Iout 0.06417f
C3117 XThR.Tn[4] XA.XIR[4].XIC[7].icell.PDM 0.00341f
C3118 XA.XIR[15].XIC[14].icell.PDM Iout 0.00117f
C3119 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10] 0.00341f
C3120 XThR.Tn[8] XA.XIR[9].XIC[7].icell.Ien 0.00338f
C3121 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C3122 XThR.TB5 a_n1319_6405# 0.01188f
C3123 XThR.Tn[3] XA.XIR[3].XIC[14].icell.PDM 0.00341f
C3124 XA.XIR[12].XIC[5].icell.SM Iout 0.00388f
C3125 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.SM 0.0039f
C3126 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C3127 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07214f
C3128 XThR.TA1 XThR.TB6 0.00193f
C3129 XThC.Tn[3] XThR.Tn[11] 0.28739f
C3130 XThR.Tn[14] XA.XIR[15].XIC_15.icell.Ien 0.00117f
C3131 XThC.Tn[8] XThR.Tn[0] 0.28773f
C3132 XA.XIR[4].XIC[9].icell.Ien Vbias 0.21098f
C3133 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.15202f
C3134 XThR.Tn[6] XA.XIR[7].XIC[1].icell.Ien 0.00338f
C3135 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.03425f
C3136 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.03425f
C3137 XA.XIR[3].XIC[7].icell.PUM VPWR 0.00937f
C3138 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Ien 0.00584f
C3139 XA.XIR[10].XIC[14].icell.SM Iout 0.00388f
C3140 XThR.Tn[9] XA.XIR[10].XIC[14].icell.SM 0.00121f
C3141 XThC.Tn[7] XThR.Tn[3] 0.28739f
C3142 XA.XIR[1].XIC[3].icell.PDM Iout 0.00117f
C3143 a_n997_3755# VPWR 0.0133f
C3144 XA.XIR[2].XIC[13].icell.Ien Vbias 0.21098f
C3145 XA.XIR[11].XIC_15.icell.SM Vbias 0.00701f
C3146 XA.XIR[2].XIC[4].icell.PDM Vbias 0.04261f
C3147 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.03425f
C3148 XThC.Tn[1] Vbias 2.40656f
C3149 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00214f
C3150 XA.XIR[6].XIC[8].icell.SM VPWR 0.00158f
C3151 XA.XIR[9].XIC_dummy_right.icell.SM VPWR 0.00123f
C3152 XA.XIR[7].XIC[9].icell.SM Vbias 0.00701f
C3153 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.SM 0.0039f
C3154 XA.XIR[15].XIC[12].icell.Ien VPWR 0.32895f
C3155 XA.XIR[4].XIC[3].icell.PDM VPWR 0.00799f
C3156 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.03425f
C3157 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00214f
C3158 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7] 0.00341f
C3159 XThR.TB5 a_n997_3979# 0.00418f
C3160 XA.XIR[6].XIC[4].icell.SM Iout 0.00388f
C3161 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13] 0.00341f
C3162 XA.XIR[1].XIC[4].icell.PUM VPWR 0.00937f
C3163 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.SM 0.00168f
C3164 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.03425f
C3165 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.15202f
C3166 XThC.Tn[2] XThR.Tn[6] 0.28739f
C3167 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3168 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3169 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04031f
C3170 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PUM 0.00465f
C3171 XA.XIR[13].XIC[9].icell.SM Iout 0.00388f
C3172 XThR.Tn[10] XA.XIR[11].XIC[14].icell.Ien 0.00338f
C3173 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00584f
C3174 XThR.Tn[13] XA.XIR[14].XIC[4].icell.Ien 0.00338f
C3175 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.SM 0.00168f
C3176 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.03425f
C3177 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00584f
C3178 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PUM 0.00465f
C3179 XA.XIR[2].XIC[11].icell.PDM Iout 0.00117f
C3180 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.15202f
C3181 XA.XIR[0].XIC[9].icell.Ien Vbias 0.2113f
C3182 XThC.Tn[2] XThC.Tn[4] 0.02725f
C3183 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02762f
C3184 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00214f
C3185 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.SM 0.00168f
C3186 XA.XIR[7].XIC[12].icell.Ien Iout 0.06417f
C3187 XThR.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.00338f
C3188 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C3189 XA.XIR[1].XIC_dummy_left.icell.SM VPWR 0.00269f
C3190 XThC.Tn[10] Iout 0.83837f
C3191 XA.XIR[14].XIC[1].icell.Ien VPWR 0.19084f
C3192 XThC.Tn[10] XThR.Tn[9] 0.28739f
C3193 XA.XIR[11].XIC[1].icell.PUM Vbias 0.0031f
C3194 XThR.Tn[4] XA.XIR[5].XIC[8].icell.SM 0.00121f
C3195 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00214f
C3196 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[6].icell.SM 0.0039f
C3197 XA.XIR[3].XIC_15.icell.PUM Vbias 0.0031f
C3198 XThR.Tn[7] XA.XIR[8].XIC[13].icell.Ien 0.00338f
C3199 XA.XIR[10].XIC[2].icell.PDM VPWR 0.00799f
C3200 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.SM 0.0039f
C3201 XThR.Tn[3] XA.XIR[4].XIC[10].icell.SM 0.00121f
C3202 XThC.Tn[6] XThR.Tn[12] 0.28739f
C3203 XThR.TA1 XThR.Tn[8] 0.00204f
C3204 XThR.Tn[10] Vbias 3.7463f
C3205 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00584f
C3206 XA.XIR[10].XIC[11].icell.Ien Iout 0.06417f
C3207 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C3208 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00214f
C3209 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04031f
C3210 XThR.Tn[9] XA.XIR[10].XIC[11].icell.Ien 0.00338f
C3211 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C3212 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.SM 0.00168f
C3213 XA.XIR[15].XIC[1].icell.PDM Vbias 0.04261f
C3214 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5] 0.00341f
C3215 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02762f
C3216 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00214f
C3217 XThC.TA2 XThC.Tn[1] 0.00411f
C3218 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C3219 XA.XIR[1].XIC[12].icell.PUM Vbias 0.0031f
C3220 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.SM 0.00168f
C3221 XA.XIR[14].XIC[7].icell.PDM Vbias 0.04261f
C3222 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C3223 XA.XIR[5].XIC[8].icell.PUM VPWR 0.00937f
C3224 XA.XIR[15].XIC[4].icell.SM VPWR 0.00158f
C3225 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PUM 0.00465f
C3226 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Ien 0.00618f
C3227 XA.XIR[3].XIC[0].icell.PDM VPWR 0.00799f
C3228 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C3229 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02762f
C3230 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00214f
C3231 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.03425f
C3232 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.0353f
C3233 XThR.TB5 XThR.Tn[7] 0.00912f
C3234 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.15202f
C3235 XThC.Tn[5] XThR.Tn[10] 0.28739f
C3236 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.03425f
C3237 XThR.TB5 a_n997_2891# 0.00424f
C3238 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.04041f
C3239 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6] 0.00341f
C3240 XA.XIR[15].XIC[8].icell.PDM Iout 0.00117f
C3241 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C3242 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.SM 0.00168f
C3243 XA.XIR[9].XIC[5].icell.PUM Vbias 0.0031f
C3244 XA.XIR[1].XIC[13].icell.SM Iout 0.00388f
C3245 XA.XIR[8].XIC[1].icell.SM VPWR 0.00158f
C3246 XA.XIR[4].XIC[1].icell.Ien VPWR 0.1903f
C3247 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C3248 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00584f
C3249 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C3250 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00584f
C3251 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Iout 0.00347f
C3252 XThR.TB2 XThR.TB6 0.04959f
C3253 XA.XIR[2].XIC[1].icell.Ien Iout 0.06417f
C3254 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.1106f
C3255 XThC.TBN a_5949_9615# 0.0768f
C3256 XA.XIR[11].XIC[2].icell.Ien VPWR 0.1903f
C3257 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.SM 0.0039f
C3258 XA.XIR[15].XIC[10].icell.Ien VPWR 0.32895f
C3259 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.SM 0.0039f
C3260 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.03425f
C3261 XA.XIR[9].XIC[6].icell.PDM Iout 0.00117f
C3262 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9] 0.00341f
C3263 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00214f
C3264 XA.XIR[9].XIC[10].icell.SM VPWR 0.00158f
C3265 XA.XIR[13].XIC[13].icell.Ien Iout 0.06417f
C3266 XA.XIR[10].XIC[4].icell.Ien VPWR 0.1903f
C3267 XA.XIR[2].XIC[3].icell.SM Vbias 0.00701f
C3268 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.15202f
C3269 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11] 0.00341f
C3270 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[14].icell.Ien 0.00214f
C3271 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.SM 0.00168f
C3272 XThR.Tn[2] XA.XIR[2].XIC[4].icell.PDM 0.00341f
C3273 XA.XIR[5].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3274 XA.XIR[5].XIC[12].icell.PDM Vbias 0.04261f
C3275 XA.XIR[12].XIC[12].icell.PDM Iout 0.00117f
C3276 XA.XIR[9].XIC[6].icell.SM Iout 0.00388f
C3277 XThC.Tn[1] XThR.Tn[2] 0.28739f
C3278 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00214f
C3279 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PUM 0.00465f
C3280 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04031f
C3281 XThR.Tn[10] XA.XIR[11].XIC[12].icell.Ien 0.00338f
C3282 XA.XIR[0].XIC[4].icell.PDM Vbias 0.04271f
C3283 XThR.Tn[0] XA.XIR[1].XIC[11].icell.SM 0.00121f
C3284 XA.XIR[7].XIC[11].icell.PDM VPWR 0.00799f
C3285 XA.XIR[8].XIC[14].icell.PDM Vbias 0.04261f
C3286 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04031f
C3287 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00584f
C3288 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18966f
C3289 XA.XIR[14].XIC[5].icell.Ien Vbias 0.21098f
C3290 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10] 0.00341f
C3291 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00256f
C3292 XA.XIR[4].XIC[6].icell.Ien VPWR 0.1903f
C3293 XA.XIR[15].XIC[13].icell.PDM Iout 0.00117f
C3294 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.15202f
C3295 XA.XIR[2].XIC[10].icell.Ien VPWR 0.1903f
C3296 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00584f
C3297 XA.XIR[4].XIC[2].icell.Ien Iout 0.06417f
C3298 XA.XIR[13].XIC[7].icell.Ien Vbias 0.21098f
C3299 XA.XIR[8].XIC[9].icell.SM Vbias 0.00701f
C3300 XA.XIR[7].XIC[6].icell.SM VPWR 0.00158f
C3301 XA.XIR[2].XIC[6].icell.Ien Iout 0.06417f
C3302 a_n997_715# VPWR 0.02818f
C3303 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.03425f
C3304 XA.XIR[11].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3305 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.03504f
C3306 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00214f
C3307 XA.XIR[12].XIC[9].icell.PUM Vbias 0.0031f
C3308 XA.XIR[7].XIC[2].icell.SM Iout 0.00388f
C3309 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3310 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.15202f
C3311 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.SM 0.00168f
C3312 XThR.Tn[13] XA.XIR[14].XIC[12].icell.SM 0.00121f
C3313 XThC.Tn[3] XThR.Tn[14] 0.28739f
C3314 XA.XIR[1].XIC[11].icell.PDM Vbias 0.04261f
C3315 XA.XIR[13].XIC[14].icell.SM Iout 0.00388f
C3316 XThC.TB7 XThC.Tn[14] 0.4237f
C3317 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.0404f
C3318 XA.XIR[14].XIC_15.icell.SM Vbias 0.00701f
C3319 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13] 0.00341f
C3320 XA.XIR[3].XIC[5].icell.Ien Vbias 0.21098f
C3321 XThR.TB2 XThR.Tn[8] 0.00167f
C3322 XThR.TB4 XThR.TB7 0.03475f
C3323 XThR.Tn[7] XA.XIR[8].XIC[3].icell.SM 0.00121f
C3324 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00214f
C3325 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PUM 0.00186f
C3326 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.03425f
C3327 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C3328 XA.XIR[12].XIC_dummy_right.icell.SM VPWR 0.00123f
C3329 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.SM 0.00168f
C3330 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00584f
C3331 XA.XIR[0].XIC[6].icell.Ien VPWR 0.18973f
C3332 XA.XIR[6].XIC[8].icell.PUM Vbias 0.0031f
C3333 XThC.TA3 a_8739_10571# 0.00995f
C3334 XA.XIR[8].XIC[12].icell.Ien Iout 0.06417f
C3335 XThR.Tn[8] XA.XIR[9].XIC[12].icell.Ien 0.00338f
C3336 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.15202f
C3337 XThR.TB6 XThR.TAN2 0.06405f
C3338 XA.XIR[0].XIC[2].icell.Ien Iout 0.06389f
C3339 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C3340 XA.XIR[1].XIC[2].icell.Ien Vbias 0.21104f
C3341 XA.XIR[15].XIC[0].icell.PUM VPWR 0.00937f
C3342 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.SM 0.00168f
C3343 XThC.Tn[4] XThR.Tn[4] 0.28739f
C3344 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00214f
C3345 XA.XIR[4].XIC[14].icell.Ien Vbias 0.21098f
C3346 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.03589f
C3347 XThR.Tn[3] a_n1049_6699# 0.27008f
C3348 XA.XIR[3].XIC[12].icell.PUM VPWR 0.00937f
C3349 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00214f
C3350 XThC.TB2 a_7875_9569# 0.06476f
C3351 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C3352 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PUM 0.00465f
C3353 XThR.TB6 XThR.Tn[6] 0.00639f
C3354 XThR.Tn[10] XA.XIR[11].XIC[4].icell.SM 0.00121f
C3355 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PUM 0.00465f
C3356 XA.XIR[6].XIC[13].icell.SM VPWR 0.00158f
C3357 XThR.Tn[0] XA.XIR[0].XIC[5].icell.PDM 0.00341f
C3358 XA.XIR[6].XIC[7].icell.PDM VPWR 0.00799f
C3359 XA.XIR[7].XIC[14].icell.SM Vbias 0.00701f
C3360 XA.XIR[5].XIC[1].icell.Ien Vbias 0.21098f
C3361 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.03425f
C3362 XThC.Tn[14] VPWR 6.85545f
C3363 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C3364 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PUM 0.00465f
C3365 XA.XIR[6].XIC[9].icell.SM Iout 0.00388f
C3366 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PUM 0.00186f
C3367 XA.XIR[1].XIC[9].icell.PUM VPWR 0.00937f
C3368 XThR.TB2 XThR.Tn[1] 0.17876f
C3369 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C3370 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02762f
C3371 XA.XIR[4].XIC[6].icell.PDM Iout 0.00117f
C3372 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.15202f
C3373 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C3374 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C3375 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00214f
C3376 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.SM 0.0039f
C3377 XA.XIR[14].XIC[0].icell.Ien Vbias 0.20951f
C3378 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.SM 0.00168f
C3379 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PUM 0.00465f
C3380 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.SM 0.0039f
C3381 XThR.Tn[13] XA.XIR[14].XIC[9].icell.Ien 0.00338f
C3382 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.SM 0.0039f
C3383 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.SM 0.00168f
C3384 XA.XIR[13].XIC[2].icell.PDM VPWR 0.00799f
C3385 XThR.Tn[13] Vbias 3.74874f
C3386 XA.XIR[13].XIC[11].icell.Ien Iout 0.06417f
C3387 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00214f
C3388 XThC.Tn[6] XThR.Tn[0] 0.28748f
C3389 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Iout 0.00347f
C3390 XThR.Tn[3] Iout 1.16236f
C3391 XA.XIR[12].XIC[7].icell.PDM VPWR 0.00799f
C3392 XA.XIR[0].XIC[14].icell.Ien Vbias 0.2113f
C3393 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C3394 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.SM 0.00168f
C3395 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04031f
C3396 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3397 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00189f
C3398 XThR.Tn[6] XA.XIR[7].XIC[11].icell.Ien 0.00338f
C3399 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C3400 XA.XIR[15].XIC[0].icell.SM Iout 0.00388f
C3401 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04031f
C3402 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.SM 0.0039f
C3403 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00584f
C3404 XThR.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.00338f
C3405 XThC.TAN XThC.Tn[12] 0.00772f
C3406 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00584f
C3407 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C3408 XThC.TB3 XThC.TB5 0.04438f
C3409 XThR.Tn[4] XA.XIR[5].XIC[13].icell.SM 0.00121f
C3410 XThR.TAN2 XThR.Tn[8] 0.1369f
C3411 VPWR data[4] 0.5303f
C3412 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04031f
C3413 XA.XIR[5].XIC[6].icell.Ien Vbias 0.21098f
C3414 XA.XIR[15].XIC[4].icell.PUM Vbias 0.0031f
C3415 XA.XIR[11].XIC[1].icell.PDM Iout 0.00117f
C3416 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11107f
C3417 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.SM 0.00168f
C3418 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C3419 XThC.Tn[5] XThR.Tn[13] 0.28739f
C3420 XA.XIR[10].XIC[12].icell.SM VPWR 0.00158f
C3421 XThR.TB5 a_n997_1579# 0.00133f
C3422 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.SM 0.0039f
C3423 XA.XIR[10].XIC[5].icell.PDM Iout 0.00117f
C3424 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04031f
C3425 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.SM 0.0039f
C3426 XA.XIR[15].XIC_15.icell.Ien VPWR 0.36724f
C3427 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.SM 0.00168f
C3428 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C3429 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C3430 XA.XIR[5].XIC[13].icell.PUM VPWR 0.00937f
C3431 XThR.Tn[13] XA.XIR[14].XIC[10].icell.SM 0.00121f
C3432 XA.XIR[5].XIC[3].icell.PDM VPWR 0.00799f
C3433 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.SM 0.0039f
C3434 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.SM 0.0039f
C3435 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.SM 0.0039f
C3436 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02762f
C3437 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07214f
C3438 XThR.Tn[10] XA.XIR[11].XIC[0].icell.Ien 0.00338f
C3439 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PUM 0.00465f
C3440 XThC.Tn[4] XThR.Tn[8] 0.28739f
C3441 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00584f
C3442 XA.XIR[15].XIC[5].icell.SM Iout 0.00388f
C3443 XA.XIR[9].XIC[14].icell.PDM Vbias 0.04261f
C3444 XA.XIR[3].XIC[3].icell.PDM Iout 0.00117f
C3445 XA.XIR[12].XIC[11].icell.PDM Iout 0.00117f
C3446 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00584f
C3447 XA.XIR[8].XIC[5].icell.PDM VPWR 0.00799f
C3448 XThC.TB3 a_4067_9615# 0.23056f
C3449 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00584f
C3450 XA.XIR[7].XIC[1].icell.PUM Vbias 0.0031f
C3451 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C3452 XA.XIR[14].XIC[2].icell.Ien VPWR 0.19084f
C3453 XThC.TB5 XThC.TB7 0.036f
C3454 XThC.TAN XThC.TB6 0.30244f
C3455 XThR.TA3 a_n1319_5317# 0.0017f
C3456 XA.XIR[9].XIC[10].icell.PUM Vbias 0.0031f
C3457 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C3458 XA.XIR[13].XIC[4].icell.Ien VPWR 0.1903f
C3459 XA.XIR[8].XIC[6].icell.SM VPWR 0.00158f
C3460 XThR.Tn[2] XA.XIR[3].XIC[5].icell.Ien 0.00338f
C3461 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.SM 0.00168f
C3462 XA.XIR[10].XIC[2].icell.SM Vbias 0.00701f
C3463 XA.XIR[15].XIC[12].icell.PDM Iout 0.00117f
C3464 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C3465 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00584f
C3466 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.SM 0.00168f
C3467 XA.XIR[12].XIC[6].icell.PUM VPWR 0.00937f
C3468 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12] 0.00341f
C3469 XThR.Tn[8] XA.XIR[9].XIC[2].icell.SM 0.00121f
C3470 XA.XIR[8].XIC[2].icell.SM Iout 0.00388f
C3471 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.0343f
C3472 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01577f
C3473 XThR.Tn[3] XA.XIR[3].XIC[1].icell.PDM 0.00341f
C3474 XA.XIR[7].XIC[7].icell.PDM Vbias 0.04261f
C3475 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C3476 XA.XIR[11].XIC[7].icell.Ien VPWR 0.1903f
C3477 XA.XIR[1].XIC[2].icell.PDM VPWR 0.00799f
C3478 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.SM 0.0039f
C3479 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04031f
C3480 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04031f
C3481 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02762f
C3482 XThR.TB2 a_n997_3755# 0.06476f
C3483 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C3484 XA.XIR[4].XIC[4].icell.SM Vbias 0.00701f
C3485 XA.XIR[3].XIC[2].icell.Ien VPWR 0.1903f
C3486 XA.XIR[10].XIC[9].icell.Ien VPWR 0.1903f
C3487 XA.XIR[2].XIC[8].icell.SM Vbias 0.00701f
C3488 XA.XIR[11].XIC[3].icell.Ien Iout 0.06417f
C3489 XThC.Tn[4] XThR.Tn[1] 0.2874f
C3490 XThR.TB4 XThR.Tn[10] 0.01391f
C3491 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.SM 0.0039f
C3492 XThR.TAN XThR.Tn[3] 0.00532f
C3493 XA.XIR[3].XIC[0].icell.PUM VPWR 0.00937f
C3494 XA.XIR[6].XIC[5].icell.PUM VPWR 0.00937f
C3495 XA.XIR[7].XIC[6].icell.PUM Vbias 0.0031f
C3496 XA.XIR[14].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3497 XA.XIR[9].XIC[11].icell.SM Iout 0.00388f
C3498 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02762f
C3499 XThC.TB5 VPWR 1.01191f
C3500 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13] 0.00341f
C3501 XThR.Tn[4] XA.XIR[5].XIC[0].icell.Ien 0.00338f
C3502 XA.XIR[10].XIC[5].icell.Ien Iout 0.06417f
C3503 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.SM 0.00168f
C3504 a_n997_2667# VPWR 0.01642f
C3505 XThR.Tn[9] XA.XIR[10].XIC[5].icell.Ien 0.00338f
C3506 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.03425f
C3507 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3508 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.SM 0.0039f
C3509 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.03425f
C3510 XThC.TBN a_8739_9569# 0.22804f
C3511 XA.XIR[4].XIC[11].icell.Ien VPWR 0.1903f
C3512 XA.XIR[7].XIC[14].icell.PDM Iout 0.00117f
C3513 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.SM 0.00168f
C3514 XA.XIR[2].XIC_15.icell.Ien VPWR 0.25566f
C3515 XA.XIR[2].XIC[10].icell.PDM VPWR 0.00799f
C3516 XA.XIR[8].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3517 XA.XIR[4].XIC[7].icell.Ien Iout 0.06417f
C3518 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8] 0.00341f
C3519 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.SM 0.00168f
C3520 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38708f
C3521 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.SM 0.0039f
C3522 XA.XIR[8].XIC[14].icell.SM Vbias 0.00701f
C3523 XA.XIR[2].XIC[11].icell.Ien Iout 0.06417f
C3524 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.PUM 0.00121f
C3525 XA.XIR[7].XIC[11].icell.SM VPWR 0.00158f
C3526 XThC.TB3 XThC.Tn[3] 0.01287f
C3527 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.SM 0.00168f
C3528 XA.XIR[0].XIC[4].icell.SM Vbias 0.00716f
C3529 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.SM 0.0039f
C3530 XA.XIR[7].XIC[7].icell.SM Iout 0.00388f
C3531 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04031f
C3532 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.15202f
C3533 XThR.Tn[6] XA.XIR[7].XIC[1].icell.SM 0.00121f
C3534 XA.XIR[10].XIC_15.icell.SM Iout 0.0047f
C3535 XThR.Tn[12] XA.XIR[13].XIC[3].icell.Ien 0.00338f
C3536 a_4067_9615# VPWR 0.70648f
C3537 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PUM 0.00465f
C3538 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C3539 XA.XIR[10].XIC[10].icell.SM VPWR 0.00158f
C3540 XThR.Tn[13] XA.XIR[14].XIC[14].icell.Ien 0.00338f
C3541 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.SM 0.0039f
C3542 XA.XIR[3].XIC[10].icell.Ien Vbias 0.21098f
C3543 XThR.Tn[1] XA.XIR[2].XIC[2].icell.Ien 0.00338f
C3544 XThR.Tn[7] XA.XIR[8].XIC[8].icell.SM 0.00121f
C3545 XA.XIR[3].XIC[0].icell.SM Iout 0.00388f
C3546 XA.XIR[6].XIC[13].icell.PUM Vbias 0.0031f
C3547 XA.XIR[0].XIC[11].icell.Ien VPWR 0.19072f
C3548 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.03425f
C3549 XA.XIR[6].XIC[3].icell.PDM Vbias 0.04261f
C3550 XA.XIR[12].XIC[0].icell.Ien VPWR 0.1903f
C3551 XThR.Tn[11] XA.XIR[12].XIC[6].icell.Ien 0.00338f
C3552 XThC.TB5 a_5155_9615# 0.24821f
C3553 XA.XIR[4].XIC[14].icell.PDM Vbias 0.04261f
C3554 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.15235f
C3555 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.15202f
C3556 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.SM 0.00168f
C3557 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PDM 0.00172f
C3558 XA.XIR[0].XIC[7].icell.Ien Iout 0.06389f
C3559 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02762f
C3560 XThR.Tn[10] XA.XIR[11].XIC_15.icell.Ien 0.00117f
C3561 XA.XIR[1].XIC[7].icell.Ien Vbias 0.21104f
C3562 XThR.Tn[11] VPWR 7.58404f
C3563 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3564 XThR.TAN2 a_n997_3755# 0.01939f
C3565 XA.XIR[5].XIC[3].icell.Ien VPWR 0.1903f
C3566 XThC.TA3 XThC.TBN 0.59539f
C3567 XA.XIR[9].XIC[2].icell.PUM VPWR 0.00937f
C3568 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00214f
C3569 XThC.TB1 XThC.TBN 0.1979f
C3570 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.15235f
C3571 XThC.Tn[9] XThC.Tn[11] 0.00252f
C3572 XThR.TA3 VPWR 0.88595f
C3573 XThC.TBN XThC.Tn[11] 0.53369f
C3574 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.SM 0.0039f
C3575 XA.XIR[15].XIC[7].icell.PDM VPWR 0.0114f
C3576 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00584f
C3577 XA.XIR[6].XIC[14].icell.SM Iout 0.00388f
C3578 XA.XIR[1].XIC[14].icell.PUM VPWR 0.00937f
C3579 XA.XIR[6].XIC[10].icell.PDM Iout 0.00117f
C3580 XA.XIR[12].XIC[3].icell.PDM Vbias 0.04261f
C3581 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PUM 0.00465f
C3582 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C3583 XThR.Tn[1] XA.XIR[1].XIC[6].icell.PDM 0.00341f
C3584 XA.XIR[10].XIC[13].icell.PUM VPWR 0.00937f
C3585 XA.XIR[11].XIC[9].icell.PDM Vbias 0.04261f
C3586 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00214f
C3587 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.SM 0.00168f
C3588 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00584f
C3589 XA.XIR[14].XIC[1].icell.PDM Iout 0.00117f
C3590 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.03425f
C3591 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.SM 0.0039f
C3592 XA.XIR[2].XIC[0].icell.SM VPWR 0.00158f
C3593 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.15202f
C3594 XA.XIR[9].XIC[5].icell.PDM VPWR 0.00799f
C3595 XA.XIR[13].XIC[5].icell.PDM Iout 0.00117f
C3596 XA.XIR[13].XIC[12].icell.SM VPWR 0.00158f
C3597 XThC.Tn[3] VPWR 5.90764f
C3598 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00214f
C3599 XThR.Tn[5] XA.XIR[6].XIC[3].icell.Ien 0.00338f
C3600 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.15202f
C3601 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.SM 0.00168f
C3602 XA.XIR[9].XIC[7].icell.PUM VPWR 0.00937f
C3603 XA.XIR[12].XIC[10].icell.PDM Iout 0.00117f
C3604 XThC.TB6 XThC.Tn[8] 0.02461f
C3605 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PUM 0.00465f
C3606 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C3607 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[11].icell.SM 0.0039f
C3608 XA.XIR[5].XIC[11].icell.Ien Vbias 0.21098f
C3609 XA.XIR[15].XIC[9].icell.PUM Vbias 0.0031f
C3610 XThR.TA1 data[4] 0.14415f
C3611 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04052f
C3612 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.SM 0.0039f
C3613 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.SM 0.0039f
C3614 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00584f
C3615 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.03425f
C3616 XA.XIR[3].XIC[11].icell.PDM Vbias 0.04261f
C3617 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C3618 XA.XIR[15].XIC[11].icell.PDM Iout 0.00117f
C3619 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C3620 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.SM 0.0039f
C3621 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C3622 XA.XIR[8].XIC[1].icell.PDM Vbias 0.04261f
C3623 XThR.Tn[11] XA.XIR[12].XIC[0].icell.SM 0.00127f
C3624 XA.XIR[4].XIC[1].icell.SM VPWR 0.00158f
C3625 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.SM 0.00168f
C3626 XA.XIR[2].XIC[5].icell.SM VPWR 0.00158f
C3627 XA.XIR[10].XIC[14].icell.Ien VPWR 0.19036f
C3628 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00214f
C3629 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14] 0.00341f
C3630 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PUM 0.00465f
C3631 XA.XIR[15].XIC_dummy_right.icell.SM VPWR 0.00123f
C3632 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.SM 0.00168f
C3633 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.SM 0.00168f
C3634 XA.XIR[13].XIC[2].icell.SM Vbias 0.00701f
C3635 XA.XIR[8].XIC[6].icell.PUM Vbias 0.0031f
C3636 XThC.TAN XThC.Tn[1] 0.0014f
C3637 XA.XIR[2].XIC[1].icell.SM Iout 0.00388f
C3638 XA.XIR[7].XIC[3].icell.PUM VPWR 0.00937f
C3639 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00584f
C3640 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04031f
C3641 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.SM 0.0039f
C3642 XThR.Tn[13] XA.XIR[14].XIC[12].icell.Ien 0.00338f
C3643 XA.XIR[0].XIC[10].icell.PDM VPWR 0.00774f
C3644 XA.XIR[12].XIC[4].icell.Ien Vbias 0.21098f
C3645 XA.XIR[5].XIC[6].icell.PDM Iout 0.00117f
C3646 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.SM 0.00168f
C3647 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01577f
C3648 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00214f
C3649 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38996f
C3650 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13] 0.00341f
C3651 XA.XIR[14].XIC[7].icell.Ien VPWR 0.19084f
C3652 XA.XIR[11].XIC[5].icell.SM Vbias 0.00701f
C3653 a_5155_9615# XThC.Tn[3] 0.00508f
C3654 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3655 XA.XIR[8].XIC[8].icell.PDM Iout 0.00117f
C3656 XA.XIR[14].XIC[3].icell.Ien Iout 0.06417f
C3657 XThC.TB3 data[0] 0.03253f
C3658 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.SM 0.00168f
C3659 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04031f
C3660 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.03549f
C3661 XThC.TA3 data[2] 0.00198f
C3662 XA.XIR[13].XIC[9].icell.Ien VPWR 0.1903f
C3663 XThC.TB2 a_6243_9615# 0.00844f
C3664 XA.XIR[9].XIC_15.icell.PUM Vbias 0.0031f
C3665 XThR.Tn[2] XA.XIR[3].XIC[10].icell.Ien 0.00338f
C3666 XA.XIR[10].XIC[7].icell.SM Vbias 0.00701f
C3667 XA.XIR[8].XIC[11].icell.SM VPWR 0.00158f
C3668 XThR.TAN a_n1049_5317# 0.01743f
C3669 XA.XIR[0].XIC[1].icell.SM VPWR 0.00158f
C3670 XA.XIR[13].XIC[5].icell.Ien Iout 0.06417f
C3671 XA.XIR[6].XIC[3].icell.Ien Vbias 0.21098f
C3672 XA.XIR[8].XIC[7].icell.SM Iout 0.00388f
C3673 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00584f
C3674 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00584f
C3675 XThR.Tn[4] XA.XIR[4].XIC[9].icell.PDM 0.00341f
C3676 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3677 XThR.TB5 XThR.Tn[4] 0.19957f
C3678 XThR.Tn[8] XA.XIR[9].XIC[7].icell.SM 0.00121f
C3679 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.15202f
C3680 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.0404f
C3681 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.SM 0.0039f
C3682 XA.XIR[4].XIC[9].icell.SM Vbias 0.00701f
C3683 XA.XIR[3].XIC[7].icell.Ien VPWR 0.1903f
C3684 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00214f
C3685 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C3686 XA.XIR[2].XIC[13].icell.SM Vbias 0.00701f
C3687 XA.XIR[1].XIC[5].icell.PDM Iout 0.00117f
C3688 XA.XIR[11].XIC[8].icell.Ien Iout 0.06417f
C3689 XA.XIR[2].XIC[6].icell.PDM Vbias 0.04261f
C3690 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PUM 0.00465f
C3691 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00584f
C3692 XA.XIR[6].XIC[10].icell.PUM VPWR 0.00937f
C3693 XA.XIR[3].XIC[3].icell.Ien Iout 0.06417f
C3694 XA.XIR[10].XIC[11].icell.PUM VPWR 0.00937f
C3695 XA.XIR[7].XIC[11].icell.PUM Vbias 0.0031f
C3696 XA.XIR[4].XIC[5].icell.PDM VPWR 0.00799f
C3697 XA.XIR[13].XIC_15.icell.SM Iout 0.0047f
C3698 XThR.TB5 XThR.TB6 2.12831f
C3699 XA.XIR[1].XIC[4].icell.Ien VPWR 0.1903f
C3700 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7] 0.00341f
C3701 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00584f
C3702 XThC.Tn[13] XThR.Tn[5] 0.2874f
C3703 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C3704 XA.XIR[12].XIC_dummy_left.icell.SM VPWR 0.00269f
C3705 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PUM 0.00465f
C3706 XA.XIR[13].XIC[10].icell.SM VPWR 0.00158f
C3707 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.03425f
C3708 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04031f
C3709 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04052f
C3710 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.SM 0.0039f
C3711 XThR.Tn[13] XA.XIR[14].XIC[4].icell.SM 0.00121f
C3712 XA.XIR[4].XIC[12].icell.Ien Iout 0.06417f
C3713 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02762f
C3714 XA.XIR[2].XIC_dummy_right.icell.SM VPWR 0.00123f
C3715 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C3716 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C3717 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.03425f
C3718 data[6] data[7] 0.04128f
C3719 XA.XIR[8].XIC[1].icell.PUM Vbias 0.0031f
C3720 XA.XIR[2].XIC[13].icell.PDM Iout 0.00117f
C3721 XA.XIR[15].XIC[1].icell.PUM VPWR 0.00937f
C3722 XA.XIR[0].XIC[9].icell.SM Vbias 0.00716f
C3723 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00214f
C3724 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PUM 0.00465f
C3725 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C3726 XA.XIR[7].XIC[12].icell.SM Iout 0.00388f
C3727 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.SM 0.00168f
C3728 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.15202f
C3729 XThR.Tn[6] XA.XIR[7].XIC[6].icell.SM 0.00121f
C3730 XThR.Tn[14] VPWR 7.78627f
C3731 XThR.Tn[7] Vbias 3.74624f
C3732 XThR.Tn[12] XA.XIR[13].XIC[8].icell.Ien 0.00338f
C3733 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PUM 0.00102f
C3734 XA.XIR[11].XIC[0].icell.PDM VPWR 0.00799f
C3735 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.SM 0.0039f
C3736 XThR.TB2 data[4] 0.00267f
C3737 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00584f
C3738 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C3739 XA.XIR[7].XIC_15.icell.SM Vbias 0.00701f
C3740 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PUM 0.00465f
C3741 XA.XIR[5].XIC[1].icell.SM Vbias 0.00701f
C3742 XA.XIR[3].XIC_15.icell.Ien Vbias 0.21234f
C3743 XThR.Tn[1] XA.XIR[2].XIC[7].icell.Ien 0.00338f
C3744 XThR.Tn[7] XA.XIR[8].XIC[13].icell.SM 0.00121f
C3745 XA.XIR[10].XIC[4].icell.PDM VPWR 0.00799f
C3746 VPWR data[0] 0.52929f
C3747 XA.XIR[10].XIC[12].icell.Ien VPWR 0.1903f
C3748 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C3749 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04031f
C3750 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C3751 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02762f
C3752 XA.XIR[15].XIC[3].icell.PDM Vbias 0.04261f
C3753 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5] 0.00341f
C3754 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PUM 0.00465f
C3755 XThR.Tn[13] XA.XIR[14].XIC[10].icell.Ien 0.00338f
C3756 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PUM 0.00465f
C3757 XA.XIR[0].XIC[12].icell.Ien Iout 0.06389f
C3758 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C3759 VPWR bias[1] 1.23968f
C3760 XA.XIR[12].XIC[1].icell.Ien Iout 0.06417f
C3761 XA.XIR[1].XIC[12].icell.Ien Vbias 0.21104f
C3762 XThC.Tn[10] XThR.Tn[3] 0.28739f
C3763 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00214f
C3764 XA.XIR[13].XIC[13].icell.PUM VPWR 0.00937f
C3765 XA.XIR[4].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3766 XThR.TA2 a_n1335_4229# 0.00304f
C3767 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.SM 0.00168f
C3768 XA.XIR[14].XIC[9].icell.PDM Vbias 0.04261f
C3769 XA.XIR[5].XIC[8].icell.Ien VPWR 0.1903f
C3770 XA.XIR[15].XIC[6].icell.PUM VPWR 0.00937f
C3771 XThR.TB5 XThR.Tn[8] 0.01728f
C3772 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.03425f
C3773 XA.XIR[3].XIC[2].icell.PDM VPWR 0.00799f
C3774 XThC.Tn[5] XThR.Tn[7] 0.28739f
C3775 XThC.Tn[13] Vbias 2.40505f
C3776 XA.XIR[5].XIC[4].icell.Ien Iout 0.06417f
C3777 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.SM 0.00168f
C3778 XThC.TA2 a_7331_10587# 0.00304f
C3779 XThR.TA1 XThR.TA3 0.07862f
C3780 XA.XIR[9].XIC[1].icell.PDM Vbias 0.04261f
C3781 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.SM 0.00168f
C3782 XThC.TB5 a_7875_9569# 0.00418f
C3783 XThC.TA1 a_7331_10587# 0.01243f
C3784 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C3785 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6] 0.00341f
C3786 XA.XIR[15].XIC[10].icell.PDM Iout 0.00117f
C3787 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PUM 0.00465f
C3788 XThC.Tn[14] XThR.Tn[6] 0.28745f
C3789 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.SM 0.0039f
C3790 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00214f
C3791 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C3792 XA.XIR[9].XIC[5].icell.Ien Vbias 0.21098f
C3793 XA.XIR[8].XIC[3].icell.PUM VPWR 0.00937f
C3794 XA.XIR[12].XIC[12].icell.SM Vbias 0.00701f
C3795 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.1106f
C3796 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.15202f
C3797 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PUM 0.00429f
C3798 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.15202f
C3799 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PUM 0.00465f
C3800 XThC.TA3 XThC.Tn[7] 0.00184f
C3801 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C3802 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.SM 0.00168f
C3803 XThC.TB1 XThC.Tn[7] 0.0045f
C3804 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.0353f
C3805 XA.XIR[11].XIC[2].icell.SM VPWR 0.00158f
C3806 XThC.TBN XThC.Tn[0] 0.53577f
C3807 XA.XIR[9].XIC[8].icell.PDM Iout 0.00117f
C3808 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.15202f
C3809 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9] 0.00341f
C3810 XThR.Tn[5] XA.XIR[6].XIC[8].icell.Ien 0.00338f
C3811 XA.XIR[13].XIC[14].icell.Ien VPWR 0.19036f
C3812 XA.XIR[9].XIC[12].icell.PUM VPWR 0.00937f
C3813 XA.XIR[10].XIC[4].icell.SM VPWR 0.00158f
C3814 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02762f
C3815 XThC.Tn[9] XThR.Tn[12] 0.28739f
C3816 XA.XIR[2].XIC[5].icell.PUM Vbias 0.0031f
C3817 XThR.TAN2 data[4] 0.02581f
C3818 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11] 0.00341f
C3819 XThR.Tn[2] XA.XIR[2].XIC[6].icell.PDM 0.00341f
C3820 XA.XIR[5].XIC[14].icell.PDM Vbias 0.04261f
C3821 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.03425f
C3822 XA.XIR[0].XIC[6].icell.PDM Vbias 0.04282f
C3823 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04031f
C3824 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C3825 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04031f
C3826 XA.XIR[7].XIC[13].icell.PDM VPWR 0.00799f
C3827 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.SM 0.0039f
C3828 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.11857f
C3829 XA.XIR[14].XIC[5].icell.SM Vbias 0.00701f
C3830 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C3831 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C3832 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00214f
C3833 XA.XIR[4].XIC[6].icell.SM VPWR 0.00158f
C3834 XA.XIR[2].XIC[10].icell.SM VPWR 0.00158f
C3835 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.04591f
C3836 XA.XIR[7].XIC[1].icell.PDM Iout 0.00117f
C3837 XThC.TB4 XThC.Tn[12] 0.00209f
C3838 XA.XIR[12].XIC_15.icell.PUM Vbias 0.0031f
C3839 XA.XIR[4].XIC[2].icell.SM Iout 0.00388f
C3840 XA.XIR[13].XIC[7].icell.SM Vbias 0.00701f
C3841 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.03023f
C3842 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C3843 XA.XIR[8].XIC[11].icell.PUM Vbias 0.0031f
C3844 XA.XIR[7].XIC[8].icell.PUM VPWR 0.00937f
C3845 XA.XIR[2].XIC[6].icell.SM Iout 0.00388f
C3846 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.SM 0.00168f
C3847 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.SM 0.0039f
C3848 XThC.Tn[8] XThR.Tn[10] 0.28739f
C3849 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PUM 0.00465f
C3850 XThC.TB6 XThC.Tn[6] 0.00689f
C3851 XA.XIR[12].XIC[9].icell.Ien Vbias 0.21098f
C3852 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00256f
C3853 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C3854 XA.XIR[10].XIC[10].icell.Ien VPWR 0.1903f
C3855 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.SM 0.00168f
C3856 XA.XIR[1].XIC[13].icell.PDM Vbias 0.04261f
C3857 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C3858 XA.XIR[3].XIC[1].icell.PUM VPWR 0.00937f
C3859 XThC.Tn[5] XA.XIR[0].XIC[6].icell.PDM 0.00343f
C3860 XA.XIR[14].XIC[8].icell.Ien Iout 0.06417f
C3861 XA.XIR[3].XIC[5].icell.SM Vbias 0.00701f
C3862 XThR.Tn[3] XA.XIR[4].XIC[2].icell.Ien 0.00338f
C3863 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.SM 0.00168f
C3864 XThR.Tn[2] XA.XIR[3].XIC_15.icell.Ien 0.00117f
C3865 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00214f
C3866 XA.XIR[9].XIC[0].icell.Ien Vbias 0.20951f
C3867 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PUM 0.00465f
C3868 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.SM 0.00168f
C3869 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C3870 XA.XIR[13].XIC[11].icell.PUM VPWR 0.00937f
C3871 XA.XIR[6].XIC[8].icell.Ien Vbias 0.21098f
C3872 XA.XIR[0].XIC[6].icell.SM VPWR 0.00158f
C3873 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C3874 XA.XIR[8].XIC[12].icell.SM Iout 0.00388f
C3875 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.04036f
C3876 a_10051_9569# XThC.Tn[13] 0.19413f
C3877 XThR.Tn[8] XA.XIR[9].XIC[12].icell.SM 0.00121f
C3878 XThR.Tn[11] XA.XIR[12].XIC[1].icell.SM 0.00121f
C3879 XA.XIR[4].XIC[1].icell.PDM Vbias 0.04261f
C3880 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3881 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C3882 XA.XIR[0].XIC[2].icell.SM Iout 0.00367f
C3883 XA.XIR[1].XIC[2].icell.SM Vbias 0.00704f
C3884 XThC.TB3 XThC.TB7 0.03772f
C3885 XThC.TB4 XThC.TB6 0.04273f
C3886 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C3887 XA.XIR[8].XIC_15.icell.SM Vbias 0.00701f
C3888 XA.XIR[3].XIC[12].icell.Ien VPWR 0.1903f
C3889 XA.XIR[4].XIC[14].icell.SM Vbias 0.00701f
C3890 a_n1319_5317# VPWR 0.00672f
C3891 XThR.TA2 XThR.TB3 0.03869f
C3892 XThR.TB2 XThR.TA3 0.2319f
C3893 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.03425f
C3894 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3895 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.SM 0.0039f
C3896 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Ien 0.00728f
C3897 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02762f
C3898 XA.XIR[3].XIC[8].icell.Ien Iout 0.06417f
C3899 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01577f
C3900 XThR.Tn[0] XA.XIR[0].XIC[7].icell.PDM 0.00341f
C3901 XThR.TAN2 a_n997_2667# 0.01679f
C3902 XA.XIR[7].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3903 XThC.Tn[13] XThR.Tn[2] 0.2874f
C3904 XA.XIR[6].XIC[9].icell.PDM VPWR 0.00799f
C3905 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C3906 XA.XIR[12].XIC[10].icell.SM Vbias 0.00701f
C3907 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.SM 0.00168f
C3908 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PDM 0.00172f
C3909 XA.XIR[1].XIC[9].icell.Ien VPWR 0.1903f
C3910 XThR.Tn[13] XA.XIR[14].XIC_15.icell.Ien 0.00117f
C3911 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C3912 XA.XIR[14].XIC[0].icell.PDM VPWR 0.00799f
C3913 XA.XIR[4].XIC[8].icell.PDM Iout 0.00117f
C3914 XThR.TB5 a_n997_3755# 0.00418f
C3915 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C3916 XA.XIR[1].XIC[5].icell.Ien Iout 0.06417f
C3917 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.03425f
C3918 XThR.TBN a_n1049_6405# 0.07602f
C3919 XA.XIR[13].XIC[4].icell.PDM VPWR 0.00799f
C3920 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C3921 XA.XIR[13].XIC[12].icell.Ien VPWR 0.1903f
C3922 XA.XIR[10].XIC[0].icell.PDM Vbias 0.04207f
C3923 XThC.TB3 VPWR 1.07065f
C3924 XA.XIR[0].XIC[14].icell.SM Vbias 0.00716f
C3925 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02762f
C3926 XThC.TB6 a_5949_10571# 0.01283f
C3927 XThC.TB5 XThC.Tn[4] 0.19958f
C3928 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C3929 XA.XIR[12].XIC[9].icell.PDM VPWR 0.00799f
C3930 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C3931 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04052f
C3932 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.SM 0.0039f
C3933 XThR.Tn[6] XA.XIR[7].XIC[11].icell.SM 0.00121f
C3934 XThR.TB4 a_n997_3979# 0.00497f
C3935 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02762f
C3936 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04031f
C3937 XA.XIR[9].XIC[2].icell.Ien VPWR 0.1903f
C3938 XThC.Tn[2] XThR.Tn[5] 0.28739f
C3939 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PUM 0.00186f
C3940 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04031f
C3941 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02762f
C3942 XThR.Tn[1] XA.XIR[2].XIC[12].icell.Ien 0.00338f
C3943 XA.XIR[5].XIC[6].icell.SM Vbias 0.00701f
C3944 XA.XIR[15].XIC[4].icell.Ien Vbias 0.17899f
C3945 XThR.TBN XA.XIR[9].XIC_dummy_left.icell.Ien 0.00246f
C3946 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04031f
C3947 XA.XIR[6].XIC_15.icell.SM Iout 0.0047f
C3948 XA.XIR[11].XIC[3].icell.PDM Iout 0.00117f
C3949 XA.XIR[12].XIC[13].icell.PUM Vbias 0.0031f
C3950 XThC.TB2 a_3523_10575# 0.01006f
C3951 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00214f
C3952 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C3953 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PUM 0.0047f
C3954 XA.XIR[10].XIC[7].icell.PDM Iout 0.00117f
C3955 XThR.Tn[0] XA.XIR[1].XIC[3].icell.Ien 0.00338f
C3956 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PUM 0.00102f
C3957 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04031f
C3958 XThR.TAN2 XThR.Tn[11] 0.11968f
C3959 XA.XIR[5].XIC[13].icell.Ien VPWR 0.1903f
C3960 XThC.TB7 VPWR 1.07717f
C3961 XA.XIR[5].XIC[5].icell.PDM VPWR 0.00799f
C3962 a_4067_9615# XThC.Tn[4] 0.00141f
C3963 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00584f
C3964 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00584f
C3965 XA.XIR[4].XIC[1].icell.PUM Vbias 0.0031f
C3966 XThR.TA3 XThR.TAN2 0.19736f
C3967 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00214f
C3968 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.03425f
C3969 XA.XIR[5].XIC[9].icell.Ien Iout 0.06417f
C3970 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02762f
C3971 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.SM 0.0039f
C3972 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PUM 0.00465f
C3973 XThR.Tn[14] XA.XIR[15].XIC[1].icell.Ien 0.00338f
C3974 XThR.TB3 a_n1049_7493# 0.23056f
C3975 XA.XIR[6].XIC[0].icell.Ien VPWR 0.1903f
C3976 XA.XIR[8].XIC[7].icell.PDM VPWR 0.00799f
C3977 XThC.TB3 a_5155_9615# 0.00913f
C3978 XA.XIR[14].XIC[2].icell.SM VPWR 0.00158f
C3979 XA.XIR[3].XIC[5].icell.PDM Iout 0.00117f
C3980 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02762f
C3981 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.SM 0.00168f
C3982 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00584f
C3983 XA.XIR[7].XIC[1].icell.Ien Vbias 0.21098f
C3984 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C3985 XThR.TA3 XThR.Tn[6] 0.1056f
C3986 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00214f
C3987 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00214f
C3988 XA.XIR[13].XIC[4].icell.SM VPWR 0.00158f
C3989 XA.XIR[9].XIC[10].icell.Ien Vbias 0.21098f
C3990 XThC.Tn[9] XThR.Tn[0] 0.28777f
C3991 XThC.Tn[4] XThR.Tn[11] 0.28739f
C3992 XThC.TA2 a_6243_10571# 0.00295f
C3993 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04031f
C3994 XA.XIR[8].XIC[8].icell.PUM VPWR 0.00937f
C3995 XThR.Tn[2] XA.XIR[3].XIC[5].icell.SM 0.00121f
C3996 XA.XIR[10].XIC[4].icell.PUM Vbias 0.0031f
C3997 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.SM 0.00168f
C3998 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00214f
C3999 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C4000 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C4001 XA.XIR[12].XIC[6].icell.Ien VPWR 0.1903f
C4002 XA.XIR[12].XIC[14].icell.Ien Vbias 0.21098f
C4003 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C4004 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12] 0.00341f
C4005 XThC.Tn[2] Vbias 2.61718f
C4006 XThR.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.00341f
C4007 XA.XIR[10].XIC_15.icell.Ien VPWR 0.25566f
C4008 XA.XIR[11].XIC[7].icell.SM VPWR 0.00158f
C4009 XA.XIR[1].XIC[4].icell.PDM VPWR 0.00799f
C4010 XA.XIR[12].XIC[2].icell.Ien Iout 0.06417f
C4011 XA.XIR[7].XIC[9].icell.PDM Vbias 0.04261f
C4012 XThR.TB4 XThR.Tn[7] 0.01797f
C4013 XA.XIR[0].XIC[1].icell.PUM Vbias 0.0031f
C4014 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00214f
C4015 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.15202f
C4016 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02762f
C4017 XThR.TB4 a_n997_2891# 0.00813f
C4018 XThR.Tn[5] XA.XIR[6].XIC[13].icell.Ien 0.00338f
C4019 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04031f
C4020 XA.XIR[4].XIC[6].icell.PUM Vbias 0.0031f
C4021 XA.XIR[3].XIC[2].icell.SM VPWR 0.00158f
C4022 XA.XIR[2].XIC[10].icell.PUM Vbias 0.0031f
C4023 XThC.Tn[3] XThR.Tn[6] 0.28739f
C4024 XA.XIR[11].XIC[3].icell.SM Iout 0.00388f
C4025 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C4026 XThC.Tn[0] XA.XIR[11].XIC_dummy_left.icell.Iout 0.00109f
C4027 XThR.Tn[14] XA.XIR[15].XIC[6].icell.Ien 0.00338f
C4028 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C4029 XA.XIR[6].XIC[5].icell.Ien VPWR 0.1903f
C4030 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00584f
C4031 XA.XIR[7].XIC[6].icell.Ien Vbias 0.21098f
C4032 XA.XIR[10].XIC[5].icell.SM Iout 0.00388f
C4033 XThR.Tn[9] XA.XIR[10].XIC[5].icell.SM 0.00121f
C4034 XThC.Tn[8] XThR.Tn[13] 0.28739f
C4035 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C4036 XA.XIR[13].XIC[10].icell.Ien VPWR 0.1903f
C4037 XThC.TBN a_9827_9569# 0.22873f
C4038 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04031f
C4039 XA.XIR[4].XIC[11].icell.SM VPWR 0.00158f
C4040 XThC.Tn[3] XThC.Tn[4] 0.49877f
C4041 XThR.Tn[1] XA.XIR[2].XIC[0].icell.Ien 0.00338f
C4042 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C4043 XA.XIR[2].XIC[12].icell.PDM VPWR 0.00799f
C4044 XThC.Tn[11] Iout 0.84142f
C4045 XThC.Tn[11] XThR.Tn[9] 0.28739f
C4046 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8] 0.00341f
C4047 XA.XIR[4].XIC[7].icell.SM Iout 0.00388f
C4048 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00584f
C4049 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C4050 XA.XIR[8].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4051 XA.XIR[7].XIC[13].icell.PUM VPWR 0.00937f
C4052 XA.XIR[2].XIC[11].icell.SM Iout 0.00388f
C4053 XA.XIR[2].XIC[0].icell.PDM Iout 0.00117f
C4054 XThR.TB6 a_n1319_5611# 0.01283f
C4055 XThC.Tn[7] XThR.Tn[12] 0.28739f
C4056 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C4057 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.SM 0.0039f
C4058 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C4059 XA.XIR[0].XIC[6].icell.PUM Vbias 0.0031f
C4060 XThR.TB1 XThR.TA2 0.01609f
C4061 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C4062 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PUM 0.00179f
C4063 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C4064 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00214f
C4065 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02762f
C4066 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.04036f
C4067 XA.XIR[12].XIC[11].icell.PUM Vbias 0.0031f
C4068 XThR.Tn[12] XA.XIR[13].XIC[3].icell.SM 0.00121f
C4069 a_5155_9615# VPWR 0.7051f
C4070 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.SM 0.00168f
C4071 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04052f
C4072 XThC.TA2 XThC.Tn[2] 0.00108f
C4073 XThR.Tn[4] XA.XIR[5].XIC[5].icell.Ien 0.00338f
C4074 XA.XIR[3].XIC[10].icell.SM Vbias 0.00701f
C4075 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[5].icell.Ien 0.00214f
C4076 XThR.Tn[1] XA.XIR[2].XIC[2].icell.SM 0.00121f
C4077 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00214f
C4078 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C4079 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.15202f
C4080 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02762f
C4081 XThR.Tn[3] XA.XIR[4].XIC[7].icell.Ien 0.00338f
C4082 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C4083 XA.XIR[6].XIC[13].icell.Ien Vbias 0.21098f
C4084 XA.XIR[0].XIC[11].icell.SM VPWR 0.00158f
C4085 XA.XIR[6].XIC[5].icell.PDM Vbias 0.04261f
C4086 XA.XIR[12].XIC[0].icell.SM VPWR 0.00158f
C4087 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.SM 0.0039f
C4088 XThR.Tn[11] XA.XIR[12].XIC[6].icell.SM 0.00121f
C4089 XThC.TB5 a_6243_9615# 0.00907f
C4090 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C4091 XThR.TB1 XThR.Tn[0] 0.1837f
C4092 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00584f
C4093 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00584f
C4094 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5] 0.00341f
C4095 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C4096 XA.XIR[0].XIC[7].icell.SM Iout 0.00367f
C4097 XA.XIR[1].XIC[7].icell.SM Vbias 0.00704f
C4098 XA.XIR[15].XIC[12].icell.SM Vbias 0.00701f
C4099 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.SM 0.0039f
C4100 XThC.Tn[6] XThR.Tn[10] 0.28739f
C4101 XA.XIR[5].XIC[3].icell.SM VPWR 0.00158f
C4102 XThR.Tn[4] XThR.Tn[5] 0.07388f
C4103 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02762f
C4104 XA.XIR[13].XIC[0].icell.PDM Vbias 0.04207f
C4105 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PUM 0.00465f
C4106 XA.XIR[3].XIC[13].icell.Ien Iout 0.06417f
C4107 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PUM 0.00465f
C4108 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PUM 0.00465f
C4109 XA.XIR[15].XIC[9].icell.PDM VPWR 0.0114f
C4110 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00214f
C4111 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02762f
C4112 XThR.TBN a_n1049_7787# 0.08456f
C4113 XA.XIR[12].XIC[5].icell.PDM Vbias 0.04261f
C4114 XA.XIR[6].XIC[12].icell.PDM Iout 0.00117f
C4115 XA.XIR[12].XIC[12].icell.Ien Vbias 0.21098f
C4116 XA.XIR[1].XIC[14].icell.Ien VPWR 0.19036f
C4117 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.03425f
C4118 XA.XIR[3].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4119 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.SM 0.00168f
C4120 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02762f
C4121 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Ien 0.00553f
C4122 XThR.Tn[1] XA.XIR[1].XIC[8].icell.PDM 0.00341f
C4123 XA.XIR[1].XIC[10].icell.Ien Iout 0.06417f
C4124 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C4125 XA.XIR[14].XIC[3].icell.PDM Iout 0.00117f
C4126 XA.XIR[2].XIC[2].icell.PUM VPWR 0.00937f
C4127 XThR.TB6 XThR.Tn[5] 0.20186f
C4128 XA.XIR[9].XIC[7].icell.PDM VPWR 0.00799f
C4129 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C4130 XThC.Tn[2] XThR.Tn[2] 0.28739f
C4131 XA.XIR[8].XIC[1].icell.Ien Vbias 0.21098f
C4132 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C4133 XA.XIR[13].XIC[7].icell.PDM Iout 0.00117f
C4134 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C4135 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Ien 0.00584f
C4136 XA.XIR[15].XIC_15.icell.PUM Vbias 0.0031f
C4137 XThR.Tn[5] XA.XIR[6].XIC[3].icell.SM 0.00121f
C4138 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PUM 0.00429f
C4139 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.03425f
C4140 XA.XIR[9].XIC[7].icell.Ien VPWR 0.1903f
C4141 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Ien 0.00232f
C4142 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00584f
C4143 XA.XIR[6].XIC_dummy_left.icell.SM VPWR 0.00269f
C4144 XThR.TBN XThR.TB3 0.17246f
C4145 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02762f
C4146 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00584f
C4147 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00584f
C4148 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C4149 XA.XIR[5].XIC[11].icell.SM Vbias 0.00701f
C4150 XA.XIR[15].XIC[9].icell.Ien Vbias 0.17899f
C4151 XA.XIR[9].XIC[3].icell.Ien Iout 0.06417f
C4152 XA.XIR[5].XIC[1].icell.PDM Vbias 0.04261f
C4153 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02762f
C4154 XA.XIR[3].XIC[13].icell.PDM Vbias 0.04261f
C4155 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.15202f
C4156 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C4157 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.SM 0.00168f
C4158 XA.XIR[7].XIC[0].icell.PDM VPWR 0.00799f
C4159 XThR.Tn[0] XA.XIR[1].XIC[8].icell.Ien 0.00338f
C4160 XA.XIR[8].XIC[3].icell.PDM Vbias 0.04261f
C4161 XA.XIR[4].XIC[3].icell.PUM VPWR 0.00937f
C4162 XThR.Tn[4] Vbias 3.74761f
C4163 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C4164 XA.XIR[2].XIC[7].icell.PUM VPWR 0.00937f
C4165 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14] 0.00341f
C4166 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.03425f
C4167 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.03425f
C4168 XThC.Tn[4] XThR.Tn[14] 0.28739f
C4169 XA.XIR[13].XIC[4].icell.PUM Vbias 0.0031f
C4170 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C4171 XA.XIR[8].XIC[6].icell.Ien Vbias 0.21098f
C4172 XA.XIR[7].XIC[3].icell.Ien VPWR 0.1903f
C4173 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04031f
C4174 XA.XIR[5].XIC[14].icell.Ien Iout 0.06417f
C4175 XA.XIR[0].XIC[12].icell.PDM VPWR 0.011f
C4176 XA.XIR[12].XIC[4].icell.SM Vbias 0.00701f
C4177 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02762f
C4178 XA.XIR[5].XIC[8].icell.PDM Iout 0.00117f
C4179 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C4180 XA.XIR[13].XIC_15.icell.Ien VPWR 0.25566f
C4181 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C4182 XA.XIR[14].XIC[7].icell.SM VPWR 0.00158f
C4183 XA.XIR[1].XIC[0].icell.PDM Vbias 0.04207f
C4184 XA.XIR[11].XIC[7].icell.PUM Vbias 0.0031f
C4185 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02762f
C4186 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Iout 0.00347f
C4187 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00584f
C4188 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C4189 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00584f
C4190 XA.XIR[6].XIC[1].icell.Ien Iout 0.06417f
C4191 XA.XIR[8].XIC[10].icell.PDM Iout 0.00117f
C4192 bias[1] bias[0] 0.13857f
C4193 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PUM 0.00465f
C4194 XA.XIR[14].XIC[3].icell.SM Iout 0.00388f
C4195 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00584f
C4196 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04031f
C4197 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00214f
C4198 XA.XIR[9].XIC_15.icell.Ien Vbias 0.21234f
C4199 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04031f
C4200 XThC.Tn[5] XThR.Tn[4] 0.28739f
C4201 XA.XIR[8].XIC[13].icell.PUM VPWR 0.00937f
C4202 XThR.Tn[2] XA.XIR[3].XIC[10].icell.SM 0.00121f
C4203 XA.XIR[10].XIC[9].icell.PUM Vbias 0.0031f
C4204 XThC.Tn[0] XA.XIR[14].XIC_dummy_left.icell.Iout 0.00109f
C4205 XA.XIR[15].XIC[10].icell.SM Vbias 0.00701f
C4206 XA.XIR[0].XIC[3].icell.PUM VPWR 0.00877f
C4207 XA.XIR[13].XIC[5].icell.SM Iout 0.00388f
C4208 XA.XIR[6].XIC[3].icell.SM Vbias 0.00701f
C4209 XThR.Tn[4] XA.XIR[4].XIC[11].icell.PDM 0.00341f
C4210 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C4211 XThC.TB3 a_7875_9569# 0.0061f
C4212 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.15202f
C4213 XA.XIR[12].XIC[7].icell.Ien Iout 0.06417f
C4214 XThR.TA1 VPWR 0.83112f
C4215 XA.XIR[10].XIC_dummy_right.icell.SM VPWR 0.00123f
C4216 XA.XIR[4].XIC[11].icell.PUM Vbias 0.0031f
C4217 XA.XIR[3].XIC[7].icell.SM VPWR 0.00158f
C4218 XA.XIR[1].XIC[7].icell.PDM Iout 0.00117f
C4219 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.SM 0.00168f
C4220 XA.XIR[2].XIC_15.icell.PUM Vbias 0.0031f
C4221 XA.XIR[11].XIC[8].icell.SM Iout 0.00388f
C4222 XA.XIR[12].XIC[10].icell.Ien Vbias 0.21098f
C4223 XA.XIR[2].XIC[8].icell.PDM Vbias 0.04261f
C4224 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C4225 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PUM 0.00465f
C4226 XA.XIR[6].XIC[10].icell.Ien VPWR 0.1903f
C4227 XA.XIR[3].XIC[3].icell.SM Iout 0.00388f
C4228 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.04036f
C4229 XA.XIR[7].XIC[11].icell.Ien Vbias 0.21098f
C4230 XA.XIR[4].XIC[7].icell.PDM VPWR 0.00799f
C4231 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.15202f
C4232 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C4233 XThC.Tn[7] XThR.Tn[0] 0.2882f
C4234 XA.XIR[6].XIC[6].icell.Ien Iout 0.06417f
C4235 XA.XIR[1].XIC[4].icell.SM VPWR 0.00158f
C4236 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7] 0.00341f
C4237 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02762f
C4238 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.SM 0.00168f
C4239 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00214f
C4240 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PUM 0.00465f
C4241 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02762f
C4242 a_2979_9615# Vbias 0.00736f
C4243 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.04036f
C4244 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00584f
C4245 XThR.TB3 a_n1049_5611# 0.009f
C4246 XA.XIR[4].XIC[12].icell.SM Iout 0.00388f
C4247 XA.XIR[15].XIC[13].icell.PUM Vbias 0.0031f
C4248 XThC.TAN XThC.Tn[13] 0.00276f
C4249 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.SM 0.00168f
C4250 XThC.TA3 data[1] 0.06544f
C4251 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.15202f
C4252 XThC.TB7 a_7875_9569# 0.00476f
C4253 XThR.Tn[8] Vbias 3.74624f
C4254 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.15202f
C4255 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Ien 0.00584f
C4256 XA.XIR[15].XIC[1].icell.Ien VPWR 0.32895f
C4257 XThR.TB5 a_n997_2667# 0.00427f
C4258 XA.XIR[2].XIC_15.icell.PDM Iout 0.00133f
C4259 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00214f
C4260 XA.XIR[0].XIC[11].icell.PUM Vbias 0.0031f
C4261 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C4262 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04031f
C4263 XA.XIR[4].XIC_15.icell.SM Vbias 0.00701f
C4264 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.SM 0.00168f
C4265 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.03425f
C4266 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C4267 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12] 0.00341f
C4268 XThC.Tn[6] XThR.Tn[13] 0.28739f
C4269 XThR.Tn[12] XA.XIR[13].XIC[8].icell.SM 0.00121f
C4270 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Iout 0.00347f
C4271 XA.XIR[11].XIC[2].icell.PDM VPWR 0.00799f
C4272 XA.XIR[11].XIC[1].icell.Ien Vbias 0.21098f
C4273 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.SM 0.0039f
C4274 XThR.Tn[4] XA.XIR[5].XIC[10].icell.Ien 0.00338f
C4275 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.03023f
C4276 XThR.Tn[1] XA.XIR[2].XIC[7].icell.SM 0.00121f
C4277 XA.XIR[5].XIC[3].icell.PUM Vbias 0.0031f
C4278 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PUM 0.00186f
C4279 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02774f
C4280 XThR.Tn[3] XA.XIR[4].XIC[12].icell.Ien 0.00338f
C4281 XThC.Tn[0] Iout 0.82523f
C4282 XThC.Tn[0] XThR.Tn[9] 0.28741f
C4283 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02762f
C4284 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PUM 0.00179f
C4285 XA.XIR[10].XIC[6].icell.PDM VPWR 0.00799f
C4286 XA.XIR[9].XIC[0].icell.SM Vbias 0.00675f
C4287 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.04036f
C4288 XA.XIR[1].XIC[0].icell.Ien Vbias 0.20957f
C4289 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C4290 XA.XIR[15].XIC[5].icell.PDM Vbias 0.04261f
C4291 XA.XIR[0].XIC[12].icell.SM Iout 0.00367f
C4292 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00214f
C4293 XThC.Tn[5] XThR.Tn[8] 0.28739f
C4294 XA.XIR[1].XIC[12].icell.SM Vbias 0.00704f
C4295 XThR.Tn[12] Iout 1.16233f
C4296 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.03425f
C4297 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.03425f
C4298 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C4299 a_7875_9569# VPWR 0.00639f
C4300 XThR.Tn[1] Vbias 3.74871f
C4301 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C4302 XA.XIR[5].XIC[8].icell.SM VPWR 0.00158f
C4303 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PUM 0.00465f
C4304 XA.XIR[15].XIC[6].icell.Ien VPWR 0.32895f
C4305 XA.XIR[15].XIC[14].icell.Ien Vbias 0.17899f
C4306 XA.XIR[0].XIC_15.icell.SM Vbias 0.00716f
C4307 XA.XIR[3].XIC[4].icell.PDM VPWR 0.00799f
C4308 XThR.TB1 XThR.TBN 0.20262f
C4309 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.15202f
C4310 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00214f
C4311 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.SM 0.0039f
C4312 XA.XIR[5].XIC[4].icell.SM Iout 0.00388f
C4313 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00584f
C4314 XA.XIR[15].XIC[2].icell.Ien Iout 0.06807f
C4315 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C4316 XA.XIR[9].XIC[3].icell.PDM Vbias 0.04261f
C4317 XThC.TB5 a_8963_9569# 0.00427f
C4318 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.03023f
C4319 XThR.TB5 XThR.Tn[11] 0.02067f
C4320 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6] 0.00341f
C4321 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PUM 0.00465f
C4322 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.SM 0.0039f
C4323 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C4324 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C4325 XThC.TB2 Vbias 0.0123f
C4326 XA.XIR[1].XIC_15.icell.Ien Iout 0.0642f
C4327 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02762f
C4328 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PUM 0.00465f
C4329 XA.XIR[9].XIC[5].icell.SM Vbias 0.00701f
C4330 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.SM 0.00168f
C4331 XA.XIR[8].XIC[3].icell.Ien VPWR 0.1903f
C4332 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.SM 0.0039f
C4333 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C4334 XThR.TA2 data[5] 0.37233f
C4335 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C4336 XThR.TA3 XThR.TB5 0.11935f
C4337 XA.XIR[12].XIC[1].icell.SM VPWR 0.00158f
C4338 XThC.Tn[5] XThR.Tn[1] 0.2874f
C4339 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.03535f
C4340 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C4341 XThR.TB2 VPWR 0.98816f
C4342 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Ien 0.00584f
C4343 a_8739_9569# XThC.Tn[10] 0.19671f
C4344 XA.XIR[11].XIC[4].icell.PUM VPWR 0.00937f
C4345 XThR.Tn[5] XA.XIR[6].XIC[8].icell.SM 0.00121f
C4346 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00214f
C4347 XA.XIR[9].XIC[10].icell.PDM Iout 0.00117f
C4348 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.SM 0.0039f
C4349 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9] 0.00341f
C4350 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.15202f
C4351 XA.XIR[2].XIC[5].icell.Ien Vbias 0.21098f
C4352 XA.XIR[9].XIC[12].icell.Ien VPWR 0.1903f
C4353 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11] 0.00341f
C4354 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02762f
C4355 XA.XIR[10].XIC[6].icell.PUM VPWR 0.00937f
C4356 XThR.Tn[2] XA.XIR[2].XIC[8].icell.PDM 0.00341f
C4357 XThR.Tn[14] XA.XIR[15].XIC[1].icell.SM 0.00121f
C4358 XA.XIR[9].XIC[8].icell.Ien Iout 0.06417f
C4359 XA.XIR[7].XIC[1].icell.SM Vbias 0.00701f
C4360 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.15202f
C4361 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00214f
C4362 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02762f
C4363 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04031f
C4364 XA.XIR[0].XIC[8].icell.PDM Vbias 0.04282f
C4365 XA.XIR[15].XIC[11].icell.PUM Vbias 0.0031f
C4366 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07214f
C4367 XThR.Tn[0] XA.XIR[1].XIC[13].icell.Ien 0.00338f
C4368 XThC.TB3 XThC.Tn[4] 0.00382f
C4369 XA.XIR[14].XIC[7].icell.PUM Vbias 0.0031f
C4370 XA.XIR[4].XIC[8].icell.PUM VPWR 0.00937f
C4371 XA.XIR[7].XIC[3].icell.PDM Iout 0.00117f
C4372 XA.XIR[11].XIC[13].icell.SM Iout 0.00388f
C4373 XA.XIR[2].XIC[12].icell.PUM VPWR 0.00937f
C4374 XThC.Tn[8] XThR.Tn[7] 0.28739f
C4375 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PUM 0.00465f
C4376 XA.XIR[12].XIC_15.icell.Ien Vbias 0.21234f
C4377 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C4378 XA.XIR[13].XIC[9].icell.PUM Vbias 0.0031f
C4379 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00584f
C4380 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00214f
C4381 XA.XIR[8].XIC[11].icell.Ien Vbias 0.21098f
C4382 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00584f
C4383 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C4384 XA.XIR[7].XIC[8].icell.Ien VPWR 0.1903f
C4385 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.03425f
C4386 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C4387 XThC.TB2 XThC.TA2 0.18237f
C4388 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00214f
C4389 data[2] data[3] 0.04128f
C4390 XA.XIR[7].XIC[4].icell.Ien Iout 0.06417f
C4391 XThC.TA1 XThC.TB2 0.02203f
C4392 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.SM 0.0039f
C4393 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.SM 0.00168f
C4394 XThR.TAN XThR.Tn[12] 0.00772f
C4395 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.04036f
C4396 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04031f
C4397 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00584f
C4398 XA.XIR[1].XIC_15.icell.PDM Vbias 0.04401f
C4399 XA.XIR[13].XIC_dummy_right.icell.SM VPWR 0.00123f
C4400 XA.XIR[3].XIC[1].icell.Ien VPWR 0.1903f
C4401 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.15202f
C4402 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00214f
C4403 XA.XIR[3].XIC[7].icell.PUM Vbias 0.0031f
C4404 XA.XIR[14].XIC[8].icell.SM Iout 0.00388f
C4405 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02762f
C4406 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[2].icell.SM 0.0039f
C4407 XThC.TA3 XThC.Tn[10] 0.00406f
C4408 XThR.Tn[3] XA.XIR[4].XIC[2].icell.SM 0.00121f
C4409 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.SM 0.0039f
C4410 XThR.Tn[7] XA.XIR[8].XIC[5].icell.Ien 0.00338f
C4411 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C4412 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00214f
C4413 XA.XIR[1].XIC[0].icell.SM Iout 0.00388f
C4414 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.SM 0.00168f
C4415 XA.XIR[6].XIC[8].icell.SM Vbias 0.00701f
C4416 XA.XIR[0].XIC[8].icell.PUM VPWR 0.00881f
C4417 XThC.Tn[10] XThC.Tn[11] 0.09949f
C4418 XA.XIR[15].XIC[12].icell.Ien Vbias 0.17899f
C4419 XThC.TA3 a_4861_9615# 0.02294f
C4420 XThC.TAN a_6243_10571# 0.00108f
C4421 XThR.TAN2 VPWR 0.90694f
C4422 XA.XIR[4].XIC[3].icell.PDM Vbias 0.04261f
C4423 XThR.Tn[12] XA.XIR[13].XIC[13].icell.SM 0.00121f
C4424 XThC.TBN XThC.Tn[12] 0.56523f
C4425 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00584f
C4426 XA.XIR[1].XIC[4].icell.PUM Vbias 0.0031f
C4427 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.15202f
C4428 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PUM 0.00465f
C4429 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.SM 0.00168f
C4430 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.SM 0.0039f
C4431 XThR.Tn[1] XThR.Tn[2] 0.10497f
C4432 XA.XIR[3].XIC[12].icell.SM VPWR 0.00158f
C4433 XA.XIR[4].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4434 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.03425f
C4435 XThR.Tn[6] VPWR 6.58002f
C4436 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12] 0.00341f
C4437 XThR.Tn[10] XA.XIR[11].XIC[6].icell.Ien 0.00338f
C4438 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C4439 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C4440 XA.XIR[10].XIC[0].icell.Ien VPWR 0.1903f
C4441 XA.XIR[6].XIC_15.icell.Ien VPWR 0.25566f
C4442 XThR.Tn[0] XA.XIR[0].XIC[9].icell.PDM 0.00341f
C4443 XA.XIR[6].XIC[11].icell.PDM VPWR 0.00799f
C4444 XA.XIR[3].XIC[8].icell.SM Iout 0.00388f
C4445 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02762f
C4446 XThR.TBN XA.XIR[11].XIC_dummy_left.icell.Iout 0.00401f
C4447 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.15202f
C4448 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C4449 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.SM 0.00168f
C4450 XThR.TB4 XThR.Tn[4] 0.00757f
C4451 XA.XIR[6].XIC[11].icell.Ien Iout 0.06417f
C4452 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.15202f
C4453 XA.XIR[1].XIC[9].icell.SM VPWR 0.00158f
C4454 XThR.TA2 XThR.Tn[9] 0.00838f
C4455 VPWR bias[0] 1.93694f
C4456 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C4457 XA.XIR[4].XIC[10].icell.PDM Iout 0.00117f
C4458 XA.XIR[14].XIC[1].icell.Ien Vbias 0.21098f
C4459 XA.XIR[14].XIC[2].icell.PDM VPWR 0.00799f
C4460 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.SM 0.00168f
C4461 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C4462 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02762f
C4463 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00584f
C4464 XThC.Tn[4] VPWR 5.88871f
C4465 XA.XIR[1].XIC[5].icell.SM Iout 0.00388f
C4466 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.SM 0.00168f
C4467 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.03425f
C4468 XA.XIR[13].XIC[6].icell.PDM VPWR 0.00799f
C4469 XThC.TB6 XThC.Tn[9] 0.0246f
C4470 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PUM 0.00465f
C4471 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00584f
C4472 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.15202f
C4473 XA.XIR[10].XIC[2].icell.PDM Vbias 0.04261f
C4474 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.15202f
C4475 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.SM 0.0039f
C4476 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.SM 0.00168f
C4477 XA.XIR[0].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4478 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00214f
C4479 XThC.TB6 XThC.TBN 0.18947f
C4480 a_8963_9569# XA.XIR[0].XIC[10].icell.PDM 0.0029f
C4481 XThR.TB3 XThR.TB7 0.03772f
C4482 XThR.TB4 XThR.TB6 0.04273f
C4483 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04031f
C4484 XThR.Tn[0] Iout 1.16239f
C4485 XA.XIR[9].XIC[2].icell.SM VPWR 0.00158f
C4486 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01432f
C4487 XThR.Tn[4] XA.XIR[5].XIC_15.icell.Ien 0.00117f
C4488 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C4489 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.15202f
C4490 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[10].icell.Ien 0.00214f
C4491 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04031f
C4492 XA.XIR[5].XIC[8].icell.PUM Vbias 0.0031f
C4493 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04031f
C4494 XA.XIR[15].XIC[4].icell.SM Vbias 0.00701f
C4495 XThR.Tn[1] XA.XIR[2].XIC[12].icell.SM 0.00121f
C4496 XA.XIR[11].XIC[5].icell.PDM Iout 0.00117f
C4497 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00214f
C4498 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C4499 XA.XIR[11].XIC[11].icell.SM Iout 0.00388f
C4500 XThR.Tn[7] XA.XIR[8].XIC[0].icell.Ien 0.00338f
C4501 XA.XIR[3].XIC[0].icell.PDM Vbias 0.04207f
C4502 XThC.TB2 XThC.TAN2 0.04716f
C4503 XThC.TAN XThC.Tn[2] 0.00273f
C4504 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.03425f
C4505 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.SM 0.0039f
C4506 XThR.Tn[0] XA.XIR[1].XIC[3].icell.SM 0.00121f
C4507 XA.XIR[10].XIC[9].icell.PDM Iout 0.00117f
C4508 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C4509 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00584f
C4510 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.11103f
C4511 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04031f
C4512 XA.XIR[2].XIC[2].icell.Ien VPWR 0.1903f
C4513 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00584f
C4514 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00214f
C4515 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PUM 0.00465f
C4516 XA.XIR[5].XIC[13].icell.SM VPWR 0.00158f
C4517 a_5155_9615# XThC.Tn[4] 0.26653f
C4518 XA.XIR[5].XIC[7].icell.PDM VPWR 0.00799f
C4519 XA.XIR[4].XIC[1].icell.Ien Vbias 0.21098f
C4520 XA.XIR[8].XIC[1].icell.SM Vbias 0.00701f
C4521 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.SM 0.00168f
C4522 XThR.Tn[10] XA.XIR[11].XIC[0].icell.SM 0.00121f
C4523 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C4524 XA.XIR[5].XIC[9].icell.SM Iout 0.00388f
C4525 XA.XIR[15].XIC[7].icell.Ien Iout 0.06807f
C4526 XA.XIR[6].XIC[0].icell.SM VPWR 0.00158f
C4527 XA.XIR[3].XIC[7].icell.PDM Iout 0.00117f
C4528 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.03425f
C4529 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C4530 XA.XIR[8].XIC[9].icell.PDM VPWR 0.00799f
C4531 XThC.TB3 a_6243_9615# 0.00899f
C4532 XA.XIR[14].XIC[4].icell.PUM VPWR 0.00937f
C4533 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C4534 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00584f
C4535 XA.XIR[11].XIC[2].icell.Ien Vbias 0.21098f
C4536 XA.XIR[15].XIC[10].icell.Ien Vbias 0.17899f
C4537 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PUM 0.00465f
C4538 XA.XIR[13].XIC[6].icell.PUM VPWR 0.00937f
C4539 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.SM 0.0039f
C4540 XA.XIR[9].XIC[10].icell.SM Vbias 0.00701f
C4541 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PUM 0.00465f
C4542 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04031f
C4543 XThR.Tn[12] XA.XIR[13].XIC[11].icell.SM 0.00121f
C4544 XA.XIR[8].XIC[8].icell.Ien VPWR 0.1903f
C4545 XA.XIR[10].XIC[4].icell.Ien Vbias 0.21098f
C4546 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.SM 0.00168f
C4547 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C4548 XThR.TB4 XThR.Tn[8] 0.01306f
C4549 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.SM 0.00168f
C4550 XA.XIR[12].XIC[6].icell.SM VPWR 0.00158f
C4551 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12] 0.00341f
C4552 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.02762f
C4553 XA.XIR[8].XIC[4].icell.Ien Iout 0.06417f
C4554 XThR.TAN XThR.TA2 1.47641f
C4555 XThR.TA1 XThR.TB2 0.02203f
C4556 XThR.Tn[8] XA.XIR[9].XIC[4].icell.Ien 0.00338f
C4557 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C4558 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07214f
C4559 XThR.Tn[3] XA.XIR[3].XIC[5].icell.PDM 0.00341f
C4560 XA.XIR[12].XIC[2].icell.SM Iout 0.00388f
C4561 XA.XIR[11].XIC[9].icell.PUM VPWR 0.00937f
C4562 XA.XIR[7].XIC[11].icell.PDM Vbias 0.04261f
C4563 XA.XIR[1].XIC[6].icell.PDM VPWR 0.00799f
C4564 XA.XIR[0].XIC[1].icell.Ien Vbias 0.2113f
C4565 XThR.Tn[5] XA.XIR[6].XIC[13].icell.SM 0.00121f
C4566 XA.XIR[4].XIC[6].icell.Ien Vbias 0.21098f
C4567 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04031f
C4568 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00214f
C4569 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.15202f
C4570 XA.XIR[14].XIC[13].icell.SM Iout 0.00388f
C4571 XA.XIR[3].XIC[4].icell.PUM VPWR 0.00937f
C4572 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00584f
C4573 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04031f
C4574 XA.XIR[2].XIC[10].icell.Ien Vbias 0.21098f
C4575 XThC.Tn[14] XThR.Tn[5] 0.28745f
C4576 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.PDM 0.00586f
C4577 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00584f
C4578 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00584f
C4579 XThR.Tn[14] XA.XIR[15].XIC[6].icell.SM 0.00121f
C4580 XA.XIR[6].XIC[5].icell.SM VPWR 0.00158f
C4581 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C4582 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00584f
C4583 XThC.TB7 a_6243_9615# 0.27822f
C4584 XThR.Tn[4] XA.XIR[5].XIC[0].icell.SM 0.00121f
C4585 XA.XIR[9].XIC[13].icell.Ien Iout 0.06417f
C4586 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.15202f
C4587 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02762f
C4588 XA.XIR[7].XIC[6].icell.SM Vbias 0.00701f
C4589 XA.XIR[6].XIC[1].icell.SM Iout 0.00388f
C4590 XA.XIR[9].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4591 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02762f
C4592 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02762f
C4593 XThC.TBN a_10915_9569# 0.21503f
C4594 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.SM 0.0039f
C4595 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C4596 XA.XIR[4].XIC[13].icell.PUM VPWR 0.00937f
C4597 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04035f
C4598 XA.XIR[2].XIC[14].icell.PDM VPWR 0.00809f
C4599 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.SM 0.00168f
C4600 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02762f
C4601 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8] 0.00341f
C4602 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.SM 0.0039f
C4603 XA.XIR[7].XIC[13].icell.Ien VPWR 0.1903f
C4604 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12] 0.00341f
C4605 XA.XIR[2].XIC[2].icell.PDM Iout 0.00117f
C4606 XA.XIR[5].XIC[0].icell.Ien VPWR 0.1903f
C4607 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.03425f
C4608 XA.XIR[0].XIC[6].icell.Ien Vbias 0.21134f
C4609 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.SM 0.00168f
C4610 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.15202f
C4611 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.SM 0.0039f
C4612 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PUM 0.00465f
C4613 XA.XIR[10].XIC_dummy_left.icell.SM VPWR 0.00269f
C4614 XA.XIR[7].XIC[9].icell.Ien Iout 0.06417f
C4615 XThR.Tn[6] XA.XIR[7].XIC[3].icell.Ien 0.00338f
C4616 XA.XIR[11].XIC[9].icell.SM Iout 0.00388f
C4617 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PDM 0.00172f
C4618 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00584f
C4619 a_6243_9615# VPWR 0.70553f
C4620 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00584f
C4621 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C4622 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00584f
C4623 XThR.Tn[4] XA.XIR[5].XIC[5].icell.SM 0.00121f
C4624 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.03425f
C4625 XA.XIR[3].XIC[12].icell.PUM Vbias 0.0031f
C4626 XThC.Tn[11] XThR.Tn[3] 0.28739f
C4627 XA.XIR[13].XIC[0].icell.Ien VPWR 0.1903f
C4628 XThR.Tn[3] XA.XIR[4].XIC[7].icell.SM 0.00121f
C4629 XThR.Tn[7] XA.XIR[8].XIC[10].icell.Ien 0.00338f
C4630 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02762f
C4631 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02762f
C4632 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.04036f
C4633 XA.XIR[0].XIC[13].icell.PUM VPWR 0.00877f
C4634 XA.XIR[6].XIC[13].icell.SM Vbias 0.00701f
C4635 XA.XIR[6].XIC[7].icell.PDM Vbias 0.04261f
C4636 XThR.TBN XA.XIR[14].XIC_dummy_left.icell.Iout 0.00116f
C4637 XA.XIR[12].XIC[2].icell.PUM VPWR 0.00937f
C4638 XThC.Tn[6] XThR.Tn[7] 0.28739f
C4639 XThC.Tn[14] Vbias 2.47342f
C4640 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.SM 0.00168f
C4641 XThR.TA1 XThR.TAN2 0.06303f
C4642 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5] 0.00341f
C4643 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00584f
C4644 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02762f
C4645 XA.XIR[1].XIC[9].icell.PUM Vbias 0.0031f
C4646 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Iout 0.00347f
C4647 XThC.Tn[5] XA.XIR[0].XIC[6].icell.Ien 0.0016f
C4648 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.15202f
C4649 XThR.TB3 XThR.Tn[10] 0.29462f
C4650 XA.XIR[5].XIC[5].icell.PUM VPWR 0.00937f
C4651 XA.XIR[15].XIC[1].icell.SM VPWR 0.00158f
C4652 XThR.TB1 XThR.TB7 0.05211f
C4653 XA.XIR[13].XIC[2].icell.PDM Vbias 0.04261f
C4654 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.03425f
C4655 XA.XIR[3].XIC[13].icell.SM Iout 0.00388f
C4656 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00584f
C4657 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.03425f
C4658 XThR.Tn[12] XA.XIR[13].XIC[9].icell.SM 0.00121f
C4659 XA.XIR[10].XIC[1].icell.Ien Iout 0.06417f
C4660 XThR.Tn[9] XA.XIR[10].XIC[1].icell.Ien 0.00338f
C4661 XA.XIR[6].XIC_dummy_right.icell.SM VPWR 0.00123f
C4662 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.15202f
C4663 XA.XIR[12].XIC[7].icell.PDM Vbias 0.04261f
C4664 XA.XIR[6].XIC[14].icell.PDM Iout 0.00117f
C4665 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02762f
C4666 XA.XIR[1].XIC[14].icell.SM VPWR 0.00207f
C4667 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C4668 XThC.TB1 a_7651_9569# 0.06353f
C4669 XThR.Tn[1] XA.XIR[1].XIC[10].icell.PDM 0.00341f
C4670 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00214f
C4671 XThC.TBN XThC.Tn[1] 0.7252f
C4672 XA.XIR[1].XIC[10].icell.SM Iout 0.00388f
C4673 XThR.TBN a_n1049_6699# 0.07601f
C4674 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00584f
C4675 XA.XIR[14].XIC[5].icell.PDM Iout 0.00117f
C4676 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02762f
C4677 XA.XIR[14].XIC[11].icell.SM Iout 0.00388f
C4678 XThC.Tn[10] XThR.Tn[12] 0.28739f
C4679 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.SM 0.00168f
C4680 XA.XIR[9].XIC[9].icell.PDM VPWR 0.00799f
C4681 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.15202f
C4682 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C4683 XA.XIR[13].XIC[9].icell.PDM Iout 0.00117f
C4684 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Ien 0.00584f
C4685 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.SM 0.0039f
C4686 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00584f
C4687 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.SM 0.0039f
C4688 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00214f
C4689 XA.XIR[10].XIC[12].icell.SM Vbias 0.00701f
C4690 XA.XIR[15].XIC_15.icell.Ien Vbias 0.17891f
C4691 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.SM 0.00168f
C4692 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C4693 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.03574f
C4694 XA.XIR[9].XIC[7].icell.SM VPWR 0.00158f
C4695 XThR.TB4 a_n997_3755# 0.00497f
C4696 XA.XIR[5].XIC[13].icell.PUM Vbias 0.0031f
C4697 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C4698 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C4699 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.15202f
C4700 XA.XIR[5].XIC[3].icell.PDM Vbias 0.04261f
C4701 XA.XIR[9].XIC[3].icell.SM Iout 0.00388f
C4702 XA.XIR[3].XIC_15.icell.PDM Vbias 0.04401f
C4703 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C4704 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.SM 0.0039f
C4705 XThC.Tn[0] XA.XIR[9].XIC_dummy_left.icell.Iout 0.00109f
C4706 XA.XIR[7].XIC[2].icell.PDM VPWR 0.00799f
C4707 XThR.Tn[0] XA.XIR[1].XIC[8].icell.SM 0.00121f
C4708 XThR.TBN XThR.Tn[9] 0.48048f
C4709 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00214f
C4710 XA.XIR[11].XIC[13].icell.Ien Iout 0.06417f
C4711 XThC.TB6 XThC.Tn[7] 0.01462f
C4712 XA.XIR[8].XIC[5].icell.PDM Vbias 0.04261f
C4713 XA.XIR[14].XIC[2].icell.Ien Vbias 0.21098f
C4714 XThC.Tn[9] XThR.Tn[10] 0.28739f
C4715 XA.XIR[4].XIC[3].icell.Ien VPWR 0.1903f
C4716 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10] 0.00341f
C4717 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C4718 XA.XIR[2].XIC[7].icell.Ien VPWR 0.1903f
C4719 XA.XIR[10].XIC[14].icell.PDM VPWR 0.00809f
C4720 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14] 0.00341f
C4721 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.SM 0.00168f
C4722 XA.XIR[13].XIC[4].icell.Ien Vbias 0.21098f
C4723 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.SM 0.00168f
C4724 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02852f
C4725 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02762f
C4726 XA.XIR[8].XIC[6].icell.SM Vbias 0.00701f
C4727 XA.XIR[2].XIC[3].icell.Ien Iout 0.06417f
C4728 XA.XIR[7].XIC[3].icell.SM VPWR 0.00158f
C4729 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04031f
C4730 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00214f
C4731 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C4732 XA.XIR[0].XIC[14].icell.PDM VPWR 0.00783f
C4733 XA.XIR[5].XIC[14].icell.SM Iout 0.00388f
C4734 XA.XIR[12].XIC[6].icell.PUM Vbias 0.0031f
C4735 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07214f
C4736 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00256f
C4737 XA.XIR[5].XIC[10].icell.PDM Iout 0.00117f
C4738 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.SM 0.00168f
C4739 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PUM 0.00465f
C4740 XA.XIR[14].XIC[9].icell.PUM VPWR 0.00937f
C4741 XA.XIR[10].XIC_15.icell.PUM Vbias 0.0031f
C4742 XA.XIR[1].XIC[2].icell.PDM Vbias 0.04261f
C4743 XA.XIR[11].XIC[7].icell.Ien Vbias 0.21098f
C4744 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.03425f
C4745 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.0353f
C4746 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.SM 0.00168f
C4747 XA.XIR[8].XIC[12].icell.PDM Iout 0.00117f
C4748 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.SM 0.0039f
C4749 XA.XIR[3].XIC[2].icell.Ien Vbias 0.21098f
C4750 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.04036f
C4751 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Ien 0.00584f
C4752 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02762f
C4753 XA.XIR[8].XIC[13].icell.Ien VPWR 0.1903f
C4754 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PUM 0.00465f
C4755 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00214f
C4756 XA.XIR[10].XIC[9].icell.Ien Vbias 0.21098f
C4757 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.SM 0.0039f
C4758 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.PDM 0.00578f
C4759 XA.XIR[6].XIC[5].icell.PUM Vbias 0.0031f
C4760 XThR.TB2 XThR.TAN2 0.04716f
C4761 XThC.TB5 a_5155_10571# 0.01188f
C4762 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18966f
C4763 XThC.TB5 Vbias 0.01581f
C4764 XA.XIR[8].XIC[9].icell.Ien Iout 0.06417f
C4765 XThR.Tn[4] XA.XIR[4].XIC[13].icell.PDM 0.00341f
C4766 XThR.Tn[12] XA.XIR[13].XIC[13].icell.Ien 0.00338f
C4767 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02762f
C4768 XThR.Tn[8] XA.XIR[9].XIC[9].icell.Ien 0.00338f
C4769 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.15202f
C4770 XA.XIR[11].XIC[14].icell.SM Iout 0.00388f
C4771 XThC.Tn[14] XThR.Tn[2] 0.28745f
C4772 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PUM 0.00465f
C4773 XA.XIR[12].XIC[7].icell.SM Iout 0.00388f
C4774 XThC.TB3 a_8963_9569# 0.002f
C4775 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12] 0.00341f
C4776 XA.XIR[12].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4777 XA.XIR[5].XIC_dummy_left.icell.SM VPWR 0.00269f
C4778 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C4779 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.SM 0.00168f
C4780 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.SM 0.0039f
C4781 XThR.TA3 XThR.Tn[5] 0.02751f
C4782 XA.XIR[4].XIC[11].icell.Ien Vbias 0.21098f
C4783 XA.XIR[3].XIC[9].icell.PUM VPWR 0.00937f
C4784 XA.XIR[2].XIC_15.icell.Ien Vbias 0.21234f
C4785 XA.XIR[1].XIC[9].icell.PDM Iout 0.00117f
C4786 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PUM 0.00465f
C4787 XA.XIR[2].XIC[10].icell.PDM Vbias 0.04261f
C4788 XA.XIR[15].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4789 XThR.Tn[10] XA.XIR[11].XIC[1].icell.SM 0.00121f
C4790 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C4791 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00214f
C4792 XA.XIR[6].XIC[10].icell.SM VPWR 0.00158f
C4793 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00214f
C4794 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.03425f
C4795 XA.XIR[7].XIC[11].icell.SM Vbias 0.00701f
C4796 XA.XIR[0].XIC[0].icell.PUM VPWR 0.00877f
C4797 XA.XIR[13].XIC_dummy_left.icell.SM VPWR 0.00269f
C4798 XA.XIR[4].XIC[9].icell.PDM VPWR 0.00799f
C4799 XThR.TB5 VPWR 1.0269f
C4800 XA.XIR[14].XIC[9].icell.SM Iout 0.00388f
C4801 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7] 0.00341f
C4802 XA.XIR[6].XIC[6].icell.SM Iout 0.00388f
C4803 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C4804 XA.XIR[1].XIC[6].icell.PUM VPWR 0.00937f
C4805 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.15202f
C4806 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PUM 0.00465f
C4807 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.PDM 0.00591f
C4808 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PUM 0.00465f
C4809 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.15202f
C4810 XThC.TB5 XThC.Tn[5] 0.01095f
C4811 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02762f
C4812 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PUM 0.00465f
C4813 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PDM 0.00172f
C4814 a_4067_9615# Vbias 0.00573f
C4815 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00584f
C4816 XThC.Tn[3] XThR.Tn[5] 0.28739f
C4817 XThR.Tn[13] XA.XIR[14].XIC[6].icell.Ien 0.00338f
C4818 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00584f
C4819 XA.XIR[10].XIC[10].icell.SM Vbias 0.00701f
C4820 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C4821 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C4822 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C4823 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02762f
C4824 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00584f
C4825 XThR.TAN XThR.TBN 0.3875f
C4826 XThC.TB7 a_8963_9569# 0.00474f
C4827 XThR.Tn[12] XA.XIR[13].XIC[14].icell.SM 0.00121f
C4828 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.25759f
C4829 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.SM 0.00168f
C4830 XA.XIR[0].XIC[11].icell.Ien Vbias 0.2113f
C4831 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.15202f
C4832 XA.XIR[12].XIC[0].icell.Ien Vbias 0.20951f
C4833 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00214f
C4834 a_n1049_8581# VPWR 0.71705f
C4835 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04031f
C4836 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C4837 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00214f
C4838 XA.XIR[7].XIC[14].icell.Ien Iout 0.06417f
C4839 XThR.Tn[6] XA.XIR[7].XIC[8].icell.Ien 0.00338f
C4840 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.SM 0.00168f
C4841 XThC.TB2 XThC.TAN 0.22599f
C4842 XThC.Tn[8] XThR.Tn[4] 0.28739f
C4843 XThC.TA2 XThC.TB5 0.01866f
C4844 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PUM 0.00465f
C4845 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C4846 XA.XIR[11].XIC[4].icell.PDM VPWR 0.00799f
C4847 XThR.Tn[11] Vbias 3.74874f
C4848 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C4849 XThC.TA1 XThC.TB5 0.0538f
C4850 XThR.Tn[4] XA.XIR[5].XIC[10].icell.SM 0.00121f
C4851 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00214f
C4852 XA.XIR[11].XIC[11].icell.Ien Iout 0.06417f
C4853 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[7].icell.SM 0.0039f
C4854 XA.XIR[5].XIC[3].icell.Ien Vbias 0.21098f
C4855 XThR.Tn[3] XA.XIR[4].XIC[12].icell.SM 0.00121f
C4856 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.SM 0.0039f
C4857 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02762f
C4858 XThR.Tn[7] XA.XIR[8].XIC_15.icell.Ien 0.00117f
C4859 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00584f
C4860 XA.XIR[10].XIC[8].icell.PDM VPWR 0.00799f
C4861 XA.XIR[9].XIC[2].icell.PUM Vbias 0.0031f
C4862 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C4863 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PDM 0.00172f
C4864 XA.XIR[13].XIC[1].icell.Ien Iout 0.06417f
C4865 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C4866 XA.XIR[15].XIC[7].icell.PDM Vbias 0.04261f
C4867 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.SM 0.00168f
C4868 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02762f
C4869 XA.XIR[1].XIC[14].icell.PUM Vbias 0.0031f
C4870 a_8963_9569# VPWR 0.0033f
C4871 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00584f
C4872 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C4873 XThR.Tn[6] XThR.TAN2 0.00131f
C4874 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.SM 0.00168f
C4875 XA.XIR[5].XIC[10].icell.PUM VPWR 0.00937f
C4876 XA.XIR[15].XIC[6].icell.SM VPWR 0.00158f
C4877 XA.XIR[10].XIC[13].icell.PUM Vbias 0.0031f
C4878 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.04498f
C4879 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02762f
C4880 XA.XIR[3].XIC[6].icell.PDM VPWR 0.00799f
C4881 XThC.Tn[0] XThR.Tn[3] 0.28747f
C4882 XThC.Tn[5] XThR.Tn[11] 0.28739f
C4883 XA.XIR[2].XIC[0].icell.SM Vbias 0.00675f
C4884 XThC.Tn[10] XThR.Tn[0] 0.28747f
C4885 XA.XIR[15].XIC[2].icell.SM Iout 0.00388f
C4886 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.SM 0.00168f
C4887 XA.XIR[9].XIC[5].icell.PDM Vbias 0.04261f
C4888 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00214f
C4889 XThC.TB5 a_10051_9569# 0.00133f
C4890 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C4891 XA.XIR[13].XIC[12].icell.SM Vbias 0.00701f
C4892 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.03425f
C4893 XThC.Tn[3] Vbias 2.45762f
C4894 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6] 0.00341f
C4895 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C4896 XThR.Tn[12] XA.XIR[13].XIC[11].icell.Ien 0.00338f
C4897 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.SM 0.0039f
C4898 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00584f
C4899 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C4900 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.03425f
C4901 XA.XIR[8].XIC[3].icell.SM VPWR 0.00158f
C4902 XA.XIR[9].XIC[7].icell.PUM Vbias 0.0031f
C4903 XThR.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.00338f
C4904 XA.XIR[10].XIC[13].icell.PDM VPWR 0.00799f
C4905 XThC.Tn[4] XThR.Tn[6] 0.28739f
C4906 XThR.Tn[13] XA.XIR[14].XIC[0].icell.SM 0.00127f
C4907 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02762f
C4908 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00584f
C4909 XA.XIR[12].XIC[3].icell.PUM VPWR 0.00937f
C4910 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C4911 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PUM 0.00465f
C4912 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00584f
C4913 XA.XIR[14].XIC[13].icell.Ien Iout 0.06417f
C4914 XThC.Tn[9] XThR.Tn[13] 0.28739f
C4915 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.SM 0.00168f
C4916 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04037f
C4917 XA.XIR[11].XIC[4].icell.Ien VPWR 0.1903f
C4918 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.SM 0.0039f
C4919 XA.XIR[9].XIC[12].icell.PDM Iout 0.00117f
C4920 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.SM 0.00168f
C4921 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9] 0.00341f
C4922 XA.XIR[13].XIC[14].icell.PDM VPWR 0.00809f
C4923 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.SM 0.0039f
C4924 XA.XIR[4].XIC[1].icell.SM Vbias 0.00701f
C4925 XA.XIR[9].XIC[12].icell.SM VPWR 0.00158f
C4926 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02762f
C4927 XA.XIR[2].XIC[5].icell.SM Vbias 0.00701f
C4928 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00214f
C4929 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.SM 0.0039f
C4930 XA.XIR[10].XIC[6].icell.Ien VPWR 0.1903f
C4931 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11] 0.00341f
C4932 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C4933 XA.XIR[10].XIC[14].icell.Ien Vbias 0.21098f
C4934 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC_15.icell.Ien 0.00214f
C4935 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.15202f
C4936 XThC.Tn[3] XThC.Tn[5] 0.00492f
C4937 XThR.Tn[2] XA.XIR[2].XIC[10].icell.PDM 0.00341f
C4938 XThC.Tn[12] Iout 0.84307f
C4939 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00214f
C4940 XA.XIR[9].XIC[8].icell.SM Iout 0.00388f
C4941 XA.XIR[10].XIC[2].icell.Ien Iout 0.06417f
C4942 XThC.Tn[12] XThR.Tn[9] 0.28739f
C4943 XA.XIR[7].XIC[3].icell.PUM Vbias 0.0031f
C4944 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C4945 XThR.Tn[9] XA.XIR[10].XIC[2].icell.Ien 0.00338f
C4946 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00584f
C4947 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PUM 0.00465f
C4948 XThR.TAN a_n1049_5611# 0.00927f
C4949 XThC.Tn[8] XThR.Tn[8] 0.28739f
C4950 XA.XIR[0].XIC[10].icell.PDM Vbias 0.04282f
C4951 XThR.Tn[7] XA.XIR[8].XIC[0].icell.SM 0.00121f
C4952 XThR.Tn[0] XA.XIR[1].XIC[13].icell.SM 0.00121f
C4953 XA.XIR[13].XIC_15.icell.PUM Vbias 0.0031f
C4954 XA.XIR[3].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4955 XA.XIR[14].XIC[7].icell.Ien Vbias 0.21098f
C4956 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00584f
C4957 XThC.TAN2 XThC.TB5 0.10854f
C4958 XA.XIR[4].XIC[8].icell.Ien VPWR 0.1903f
C4959 XA.XIR[7].XIC[5].icell.PDM Iout 0.00117f
C4960 XA.XIR[2].XIC[12].icell.Ien VPWR 0.1903f
C4961 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12] 0.00341f
C4962 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00584f
C4963 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.03425f
C4964 XA.XIR[2].XIC[1].icell.PDM VPWR 0.00799f
C4965 XA.XIR[13].XIC[9].icell.Ien Vbias 0.21098f
C4966 XA.XIR[4].XIC[4].icell.Ien Iout 0.06417f
C4967 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8] 0.00341f
C4968 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C4969 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02771f
C4970 XA.XIR[2].XIC[8].icell.Ien Iout 0.06417f
C4971 XA.XIR[8].XIC[11].icell.SM Vbias 0.00701f
C4972 XA.XIR[7].XIC[8].icell.SM VPWR 0.00158f
C4973 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00214f
C4974 XThC.TB4 XThC.Tn[2] 0.0021f
C4975 XA.XIR[0].XIC[1].icell.SM Vbias 0.00716f
C4976 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C4977 XA.XIR[14].XIC[14].icell.SM Iout 0.00388f
C4978 XA.XIR[7].XIC[4].icell.SM Iout 0.00388f
C4979 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04031f
C4980 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.SM 0.0039f
C4981 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C4982 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.15202f
C4983 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.38919f
C4984 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C4985 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11336f
C4986 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PUM 0.00465f
C4987 XA.XIR[3].XIC[7].icell.Ien Vbias 0.21098f
C4988 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PUM 0.00429f
C4989 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00214f
C4990 XThC.Tn[8] XThR.Tn[1] 0.28739f
C4991 XThC.Tn[7] XThR.Tn[10] 0.28739f
C4992 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.SM 0.00168f
C4993 XThR.Tn[7] XA.XIR[8].XIC[5].icell.SM 0.00121f
C4994 XA.XIR[6].XIC[10].icell.PUM Vbias 0.0031f
C4995 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C4996 XA.XIR[0].XIC[8].icell.Ien VPWR 0.19149f
C4997 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C4998 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.SM 0.0039f
C4999 XThC.TA3 a_5949_9615# 0.01824f
C5000 XA.XIR[8].XIC[14].icell.Ien Iout 0.06417f
C5001 XThR.TA3 XThR.Tn[2] 0.12549f
C5002 XThR.Tn[11] XA.XIR[12].XIC[3].icell.Ien 0.00338f
C5003 XA.XIR[10].XIC[11].icell.PUM Vbias 0.0031f
C5004 XThR.Tn[8] XA.XIR[9].XIC[14].icell.Ien 0.00338f
C5005 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.15202f
C5006 XA.XIR[4].XIC[5].icell.PDM Vbias 0.04261f
C5007 XA.XIR[0].XIC[4].icell.Ien Iout 0.06389f
C5008 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5009 XA.XIR[1].XIC[4].icell.Ien Vbias 0.21104f
C5010 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PUM 0.00465f
C5011 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02762f
C5012 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C5013 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00214f
C5014 XA.XIR[3].XIC[14].icell.PUM VPWR 0.00937f
C5015 XA.XIR[13].XIC[10].icell.SM Vbias 0.00701f
C5016 XThC.TB2 XThC.Tn[8] 0.00167f
C5017 XA.XIR[10].XIC[0].icell.SM VPWR 0.00158f
C5018 XThR.Tn[10] XA.XIR[11].XIC[6].icell.SM 0.00121f
C5019 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00584f
C5020 XThR.Tn[0] XA.XIR[0].XIC[11].icell.PDM 0.00341f
C5021 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.SM 0.0039f
C5022 a_3773_9615# XThC.Tn[1] 0.27139f
C5023 XA.XIR[6].XIC[13].icell.PDM VPWR 0.00799f
C5024 XA.XIR[15].XIC[1].icell.PUM Vbias 0.0031f
C5025 XThR.TA1 XThR.TB5 0.0538f
C5026 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.SM 0.00168f
C5027 XA.XIR[6].XIC[11].icell.SM Iout 0.00388f
C5028 XA.XIR[6].XIC[1].icell.PDM Iout 0.00117f
C5029 XA.XIR[1].XIC[11].icell.PUM VPWR 0.00937f
C5030 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.15202f
C5031 XA.XIR[4].XIC[12].icell.PDM Iout 0.00117f
C5032 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C5033 XThC.Tn[3] XThR.Tn[2] 0.28739f
C5034 XThR.Tn[14] Vbias 3.74893f
C5035 XA.XIR[14].XIC[4].icell.PDM VPWR 0.00799f
C5036 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.SM 0.0039f
C5037 XA.XIR[14].XIC[11].icell.Ien Iout 0.06417f
C5038 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02762f
C5039 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C5040 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Iout 0.00347f
C5041 XA.XIR[11].XIC[0].icell.PDM Vbias 0.04207f
C5042 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C5043 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C5044 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PUM 0.00465f
C5045 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.15202f
C5046 XA.XIR[13].XIC[8].icell.PDM VPWR 0.00799f
C5047 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.03425f
C5048 Vbias data[0] 0.00282f
C5049 XA.XIR[10].XIC[4].icell.PDM Vbias 0.04261f
C5050 XA.XIR[10].XIC[12].icell.Ien Vbias 0.21098f
C5051 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.15202f
C5052 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.SM 0.00168f
C5053 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C5054 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C5055 a_9827_9569# XA.XIR[0].XIC[11].icell.PDM 0.00136f
C5056 XA.XIR[2].XIC[0].icell.Ien VPWR 0.1903f
C5057 XThR.Tn[6] XA.XIR[7].XIC[13].icell.Ien 0.00338f
C5058 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.0284f
C5059 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PUM 0.00465f
C5060 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.03425f
C5061 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PUM 0.00465f
C5062 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.15202f
C5063 XA.XIR[9].XIC[4].icell.PUM VPWR 0.00937f
C5064 bias[1] Vbias 0.04991f
C5065 XA.XIR[12].XIC[1].icell.PDM Iout 0.00117f
C5066 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04031f
C5067 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00584f
C5068 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00584f
C5069 XA.XIR[13].XIC[13].icell.PUM Vbias 0.0031f
C5070 XA.XIR[5].XIC[8].icell.Ien Vbias 0.21098f
C5071 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.04036f
C5072 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.SM 0.00168f
C5073 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04031f
C5074 XA.XIR[15].XIC[6].icell.PUM Vbias 0.0031f
C5075 XThC.Tn[5] XThR.Tn[14] 0.28739f
C5076 XA.XIR[11].XIC[7].icell.PDM Iout 0.00117f
C5077 XA.XIR[3].XIC[2].icell.PDM Vbias 0.04261f
C5078 XA.XIR[11].XIC[12].icell.SM VPWR 0.00158f
C5079 XThR.TB7 XThR.Tn[9] 0.07413f
C5080 XA.XIR[1].XIC_15.icell.SM VPWR 0.00275f
C5081 XThR.TB4 a_n997_2667# 0.07199f
C5082 XA.XIR[10].XIC[12].icell.PDM VPWR 0.00799f
C5083 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.SM 0.0039f
C5084 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00584f
C5085 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Ien 0.00232f
C5086 XA.XIR[2].XIC[2].icell.SM VPWR 0.00158f
C5087 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02762f
C5088 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.03425f
C5089 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.15202f
C5090 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02762f
C5091 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PDM 0.0059f
C5092 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01577f
C5093 XA.XIR[5].XIC[9].icell.PDM VPWR 0.00799f
C5094 XA.XIR[8].XIC[3].icell.PUM Vbias 0.0031f
C5095 XA.XIR[13].XIC[13].icell.PDM VPWR 0.00799f
C5096 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C5097 XA.XIR[0].XIC[1].icell.PDM VPWR 0.00774f
C5098 XThC.Tn[6] XThR.Tn[4] 0.28739f
C5099 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.SM 0.0039f
C5100 XA.XIR[15].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5101 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00584f
C5102 XA.XIR[15].XIC[7].icell.SM Iout 0.00388f
C5103 XA.XIR[3].XIC[9].icell.PDM Iout 0.00117f
C5104 XA.XIR[6].XIC[2].icell.PUM VPWR 0.00937f
C5105 XA.XIR[8].XIC[11].icell.PDM VPWR 0.00799f
C5106 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00584f
C5107 XA.XIR[14].XIC[4].icell.Ien VPWR 0.19084f
C5108 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13] 0.00341f
C5109 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C5110 XA.XIR[11].XIC[2].icell.SM Vbias 0.00701f
C5111 XThC.TA2 data[0] 0.48493f
C5112 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.03425f
C5113 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.04036f
C5114 XA.XIR[13].XIC[6].icell.Ien VPWR 0.1903f
C5115 XThC.TA1 data[0] 0.14415f
C5116 XA.XIR[13].XIC[14].icell.Ien Vbias 0.21098f
C5117 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04031f
C5118 XA.XIR[9].XIC[12].icell.PUM Vbias 0.0031f
C5119 XThR.Tn[2] XA.XIR[3].XIC[7].icell.Ien 0.00338f
C5120 XA.XIR[8].XIC[8].icell.SM VPWR 0.00158f
C5121 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.SM 0.00168f
C5122 XA.XIR[10].XIC[4].icell.SM Vbias 0.00701f
C5123 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00584f
C5124 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C5125 XA.XIR[13].XIC[2].icell.Ien Iout 0.06417f
C5126 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C5127 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01577f
C5128 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12] 0.00341f
C5129 XA.XIR[12].XIC[8].icell.PUM VPWR 0.00937f
C5130 XThR.Tn[4] XA.XIR[4].XIC[0].icell.PDM 0.00346f
C5131 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02762f
C5132 XA.XIR[8].XIC[4].icell.SM Iout 0.00388f
C5133 XThR.TB3 a_n997_3979# 0.00604f
C5134 XThR.Tn[8] XA.XIR[9].XIC[4].icell.SM 0.00121f
C5135 XThR.Tn[3] XA.XIR[3].XIC[7].icell.PDM 0.00341f
C5136 XA.XIR[7].XIC[13].icell.PDM Vbias 0.04261f
C5137 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00584f
C5138 XA.XIR[1].XIC[8].icell.PDM VPWR 0.00799f
C5139 XA.XIR[11].XIC[9].icell.Ien VPWR 0.1903f
C5140 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.SM 0.0039f
C5141 XThR.TB4 XThR.Tn[11] 0.3042f
C5142 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PUM 0.00186f
C5143 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02762f
C5144 XA.XIR[4].XIC[6].icell.SM Vbias 0.00701f
C5145 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04031f
C5146 XA.XIR[3].XIC[4].icell.Ien VPWR 0.1903f
C5147 XA.XIR[2].XIC[10].icell.SM Vbias 0.00701f
C5148 XA.XIR[11].XIC[5].icell.Ien Iout 0.06417f
C5149 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C5150 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.SM 0.00168f
C5151 XA.XIR[5].XIC_15.icell.SM Iout 0.0047f
C5152 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C5153 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00214f
C5154 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.SM 0.0039f
C5155 XA.XIR[6].XIC[7].icell.PUM VPWR 0.00937f
C5156 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PUM 0.0047f
C5157 XA.XIR[9].XIC[13].icell.SM Iout 0.00388f
C5158 XA.XIR[7].XIC[8].icell.PUM Vbias 0.0031f
C5159 XThR.TA3 XThR.TB4 0.14536f
C5160 XThR.TB2 XThR.TB5 0.0451f
C5161 XA.XIR[10].XIC[7].icell.Ien Iout 0.06417f
C5162 XThR.Tn[9] XA.XIR[10].XIC[7].icell.Ien 0.00338f
C5163 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PUM 0.00465f
C5164 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C5165 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.SM 0.0039f
C5166 XThR.TBN XA.XIR[9].XIC_dummy_left.icell.Iout 0.00395f
C5167 XA.XIR[4].XIC[13].icell.Ien VPWR 0.1903f
C5168 XA.XIR[10].XIC[10].icell.Ien Vbias 0.21098f
C5169 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04031f
C5170 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PUM 0.00465f
C5171 XA.XIR[3].XIC[1].icell.PUM Vbias 0.0031f
C5172 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5173 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C5174 XA.XIR[4].XIC[9].icell.Ien Iout 0.06417f
C5175 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8] 0.00341f
C5176 XThR.Tn[13] XA.XIR[14].XIC[1].icell.SM 0.00121f
C5177 XThC.Tn[7] XThR.Tn[13] 0.28739f
C5178 XThR.TAN XThR.TB7 0.33493f
C5179 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C5180 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Iout 0.00347f
C5181 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PUM 0.00465f
C5182 XA.XIR[2].XIC[13].icell.Ien Iout 0.06417f
C5183 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PUM 0.00465f
C5184 XA.XIR[11].XIC_15.icell.SM Iout 0.0047f
C5185 XA.XIR[7].XIC[13].icell.SM VPWR 0.00158f
C5186 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02762f
C5187 a_n1319_5611# VPWR 0.00674f
C5188 XA.XIR[2].XIC[4].icell.PDM Iout 0.00117f
C5189 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.SM 0.00168f
C5190 XA.XIR[13].XIC[11].icell.PUM Vbias 0.0031f
C5191 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.03425f
C5192 XThC.Tn[1] Iout 0.84229f
C5193 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PUM 0.00465f
C5194 XA.XIR[0].XIC[6].icell.SM Vbias 0.00716f
C5195 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C5196 XThC.Tn[1] XThR.Tn[9] 0.28739f
C5197 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.SM 0.0039f
C5198 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C5199 XA.XIR[7].XIC[9].icell.SM Iout 0.00388f
C5200 XThR.Tn[6] XA.XIR[7].XIC[3].icell.SM 0.00121f
C5201 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.15202f
C5202 XA.XIR[2].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5203 XA.XIR[11].XIC[10].icell.SM VPWR 0.00158f
C5204 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.15202f
C5205 XThR.Tn[12] XA.XIR[13].XIC[5].icell.Ien 0.00338f
C5206 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C5207 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.SM 0.00168f
C5208 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.SM 0.0039f
C5209 XThC.Tn[6] XThR.Tn[8] 0.28739f
C5210 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Ien 0.00584f
C5211 XThR.Tn[1] XA.XIR[2].XIC[4].icell.Ien 0.00338f
C5212 XA.XIR[3].XIC[12].icell.Ien Vbias 0.21098f
C5213 XA.XIR[13].XIC[0].icell.SM VPWR 0.00158f
C5214 XThR.Tn[7] XA.XIR[8].XIC[10].icell.SM 0.00121f
C5215 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C5216 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11] 0.00341f
C5217 XA.XIR[6].XIC_15.icell.PUM Vbias 0.0031f
C5218 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04031f
C5219 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18966f
C5220 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C5221 XA.XIR[6].XIC[9].icell.PDM Vbias 0.04261f
C5222 XThR.Tn[11] XA.XIR[12].XIC[8].icell.Ien 0.00338f
C5223 XThR.TB3 XThR.Tn[7] 0.00819f
C5224 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.15202f
C5225 XThR.TB3 a_n997_2891# 0.07285f
C5226 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5] 0.00341f
C5227 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C5228 XA.XIR[0].XIC[9].icell.Ien Iout 0.06389f
C5229 XThC.TAN2 data[0] 0.02545f
C5230 XA.XIR[1].XIC[9].icell.Ien Vbias 0.21104f
C5231 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Iout 0.00347f
C5232 XA.XIR[14].XIC[0].icell.PDM Vbias 0.04207f
C5233 XA.XIR[5].XIC[5].icell.Ien VPWR 0.1903f
C5234 XA.XIR[2].XIC_dummy_left.icell.SM VPWR 0.00269f
C5235 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.15222f
C5236 XA.XIR[15].XIC[3].icell.PUM VPWR 0.00937f
C5237 XThR.Tn[5] XA.XIR[6].XIC[0].icell.Ien 0.00338f
C5238 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C5239 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00214f
C5240 XA.XIR[13].XIC[4].icell.PDM Vbias 0.04261f
C5241 XA.XIR[13].XIC[12].icell.Ien Vbias 0.21098f
C5242 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02799f
C5243 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.SM 0.0039f
C5244 XThC.TB3 Vbias 0.01225f
C5245 XThR.TB5 XThR.TAN2 0.10854f
C5246 XThR.Tn[10] Iout 1.16231f
C5247 XThC.TA3 a_8739_9569# 0.00342f
C5248 XA.XIR[11].XIC[13].icell.PUM VPWR 0.00937f
C5249 XThC.Tn[6] XThR.Tn[1] 0.2874f
C5250 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00584f
C5251 XThR.Tn[9] XThR.Tn[10] 0.07779f
C5252 XA.XIR[12].XIC[9].icell.PDM Vbias 0.04261f
C5253 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.SM 0.00168f
C5254 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PUM 0.00465f
C5255 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5256 XA.XIR[15].XIC[1].icell.PDM Iout 0.00117f
C5257 XA.XIR[10].XIC[11].icell.PDM VPWR 0.00799f
C5258 XThR.Tn[1] XA.XIR[1].XIC[12].icell.PDM 0.00341f
C5259 XThR.TB5 XThR.Tn[6] 0.00349f
C5260 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00584f
C5261 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.SM 0.00168f
C5262 XA.XIR[9].XIC[2].icell.Ien Vbias 0.21098f
C5263 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00214f
C5264 XThR.Tn[5] VPWR 6.61445f
C5265 XA.XIR[14].XIC[7].icell.PDM Iout 0.00117f
C5266 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00256f
C5267 XA.XIR[14].XIC[12].icell.SM VPWR 0.00158f
C5268 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C5269 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02762f
C5270 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00256f
C5271 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.15202f
C5272 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C5273 XA.XIR[9].XIC[11].icell.PDM VPWR 0.00799f
C5274 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C5275 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C5276 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02762f
C5277 XA.XIR[13].XIC[12].icell.PDM VPWR 0.00799f
C5278 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00214f
C5279 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02762f
C5280 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.15202f
C5281 XThR.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.00338f
C5282 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C5283 XThC.TB3 XThC.Tn[5] 0.00384f
C5284 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00584f
C5285 XA.XIR[9].XIC[9].icell.PUM VPWR 0.00937f
C5286 XA.XIR[10].XIC[1].icell.SM VPWR 0.00158f
C5287 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C5288 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C5289 XA.XIR[5].XIC[13].icell.Ien Vbias 0.21098f
C5290 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[12].icell.SM 0.0039f
C5291 XThC.TB7 Vbias 0.02353f
C5292 XThC.Tn[9] XThR.Tn[7] 0.28739f
C5293 XA.XIR[5].XIC[5].icell.PDM Vbias 0.04261f
C5294 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.SM 0.0039f
C5295 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.15202f
C5296 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.PDM 0.0059f
C5297 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00584f
C5298 XThC.TB5 XThC.TAN 0.30234f
C5299 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C5300 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.SM 0.00168f
C5301 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00214f
C5302 XA.XIR[7].XIC[4].icell.PDM VPWR 0.00799f
C5303 XA.XIR[11].XIC[14].icell.Ien VPWR 0.19036f
C5304 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04038f
C5305 XA.XIR[8].XIC[7].icell.PDM Vbias 0.04261f
C5306 XA.XIR[6].XIC[0].icell.Ien Vbias 0.20951f
C5307 XA.XIR[14].XIC[2].icell.SM Vbias 0.00701f
C5308 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C5309 XA.XIR[4].XIC[3].icell.SM VPWR 0.00158f
C5310 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10] 0.00341f
C5311 XThR.TB1 a_n997_3979# 0.06353f
C5312 XThC.TB2 XThC.TB4 0.04006f
C5313 XThC.TB1 a_3299_10575# 0.0097f
C5314 XThC.TA2 XThC.TB3 0.03869f
C5315 XA.XIR[2].XIC[7].icell.SM VPWR 0.00158f
C5316 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C5317 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14] 0.00341f
C5318 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.15202f
C5319 XThC.TB1 XThC.TA3 0.48957f
C5320 XThC.TA1 XThC.TB3 0.01156f
C5321 XA.XIR[13].XIC[4].icell.SM Vbias 0.00701f
C5322 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C5323 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PUM 0.00465f
C5324 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02762f
C5325 XA.XIR[8].XIC[8].icell.PUM Vbias 0.0031f
C5326 XA.XIR[7].XIC[5].icell.PUM VPWR 0.00937f
C5327 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01577f
C5328 XA.XIR[2].XIC[3].icell.SM Iout 0.00388f
C5329 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C5330 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02762f
C5331 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.SM 0.0039f
C5332 XA.XIR[5].XIC[12].icell.PDM Iout 0.00117f
C5333 XThC.Tn[0] XA.XIR[2].XIC_dummy_left.icell.Iout 0.00109f
C5334 XA.XIR[12].XIC[6].icell.Ien Vbias 0.21098f
C5335 XThR.TBN XThR.Tn[3] 0.62502f
C5336 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00214f
C5337 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.SM 0.0039f
C5338 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02762f
C5339 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.03425f
C5340 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C5341 a_5155_10571# VPWR 0.00653f
C5342 XA.XIR[14].XIC[9].icell.Ien VPWR 0.19084f
C5343 VPWR Vbias 0.21642p
C5344 XA.XIR[10].XIC_15.icell.Ien Vbias 0.21234f
C5345 XThC.Tn[10] XThC.Tn[12] 0.00453f
C5346 XA.XIR[11].XIC[7].icell.SM Vbias 0.00701f
C5347 XA.XIR[1].XIC[4].icell.PDM Vbias 0.04261f
C5348 XA.XIR[14].XIC[5].icell.Ien Iout 0.06417f
C5349 XThC.TBN XThC.Tn[13] 0.62331f
C5350 XA.XIR[8].XIC[14].icell.PDM Iout 0.00117f
C5351 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C5352 XA.XIR[1].XIC[1].icell.Ien VPWR 0.1903f
C5353 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PDM 0.00172f
C5354 XA.XIR[3].XIC[2].icell.SM Vbias 0.00701f
C5355 XA.XIR[8].XIC[13].icell.SM VPWR 0.00158f
C5356 XThR.Tn[2] XA.XIR[3].XIC[12].icell.Ien 0.00338f
C5357 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C5358 XThR.TAN XThR.Tn[10] 0.06102f
C5359 XA.XIR[13].XIC[7].icell.Ien Iout 0.06417f
C5360 XA.XIR[6].XIC[5].icell.Ien Vbias 0.21098f
C5361 XA.XIR[0].XIC[3].icell.SM VPWR 0.00158f
C5362 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C5363 XThR.Tn[4] XA.XIR[4].XIC_15.icell.PDM 0.00341f
C5364 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00256f
C5365 XA.XIR[8].XIC[9].icell.SM Iout 0.00388f
C5366 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C5367 XThR.Tn[8] XA.XIR[9].XIC[9].icell.SM 0.00121f
C5368 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C5369 XThC.TA2 XThC.TB7 0.01596f
C5370 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C5371 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.03426f
C5372 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PUM 0.00444f
C5373 XThC.TA1 XThC.TB7 0.00179f
C5374 XA.XIR[13].XIC[10].icell.Ien Vbias 0.21098f
C5375 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.SM 0.0039f
C5376 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PUM 0.00465f
C5377 XA.XIR[4].XIC[11].icell.SM Vbias 0.00701f
C5378 XA.XIR[3].XIC[9].icell.Ien VPWR 0.1903f
C5379 XA.XIR[11].XIC[11].icell.PUM VPWR 0.00937f
C5380 XA.XIR[1].XIC[11].icell.PDM Iout 0.00117f
C5381 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.03023f
C5382 XThC.Tn[5] VPWR 5.90052f
C5383 XA.XIR[2].XIC[12].icell.PDM Vbias 0.04261f
C5384 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C5385 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C5386 XA.XIR[14].XIC_15.icell.SM Iout 0.0047f
C5387 XA.XIR[3].XIC[5].icell.Ien Iout 0.06417f
C5388 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02762f
C5389 XA.XIR[6].XIC[12].icell.PUM VPWR 0.00937f
C5390 XA.XIR[7].XIC[13].icell.PUM Vbias 0.0031f
C5391 XA.XIR[6].XIC[0].icell.PDM VPWR 0.00799f
C5392 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00584f
C5393 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PUM 0.00465f
C5394 XThC.TB6 XThC.Tn[10] 0.02461f
C5395 XA.XIR[4].XIC[11].icell.PDM VPWR 0.00799f
C5396 XA.XIR[14].XIC[10].icell.SM VPWR 0.00158f
C5397 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7] 0.00341f
C5398 XA.XIR[1].XIC[6].icell.Ien VPWR 0.1903f
C5399 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.03425f
C5400 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.03425f
C5401 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11] 0.00341f
C5402 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C5403 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00584f
C5404 XThR.TBN XA.XIR[6].XIC_dummy_left.icell.Ien 0.00159f
C5405 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.SM 0.00168f
C5406 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.03425f
C5407 XThR.TB1 XThR.Tn[7] 0.00426f
C5408 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.03425f
C5409 a_5155_9615# Vbias 0.00695f
C5410 XA.XIR[1].XIC[2].icell.Ien Iout 0.06417f
C5411 XThR.Tn[13] XA.XIR[14].XIC[6].icell.SM 0.00121f
C5412 XA.XIR[4].XIC[14].icell.Ien Iout 0.06417f
C5413 XThC.TA2 VPWR 0.68179f
C5414 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.SM 0.00168f
C5415 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00584f
C5416 XThC.TB7 a_10051_9569# 0.013f
C5417 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00584f
C5418 XThC.TA1 VPWR 0.82807f
C5419 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00214f
C5420 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C5421 XA.XIR[0].XIC[11].icell.SM Vbias 0.00716f
C5422 XA.XIR[12].XIC[0].icell.PDM VPWR 0.00799f
C5423 XA.XIR[12].XIC[0].icell.SM Vbias 0.00675f
C5424 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04031f
C5425 XA.XIR[7].XIC[14].icell.SM Iout 0.00388f
C5426 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.SM 0.00168f
C5427 XThC.TAN XThC.Tn[3] 0.00532f
C5428 XThR.Tn[6] XA.XIR[7].XIC[8].icell.SM 0.00121f
C5429 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C5430 XA.XIR[5].XIC[1].icell.Ien Iout 0.06417f
C5431 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C5432 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PUM 0.00465f
C5433 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PUM 0.00465f
C5434 XThC.TB3 XThC.TAN2 0.03907f
C5435 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.03425f
C5436 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PUM 0.00465f
C5437 XA.XIR[11].XIC[6].icell.PDM VPWR 0.00799f
C5438 XA.XIR[11].XIC[12].icell.Ien VPWR 0.1903f
C5439 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PUM 0.00465f
C5440 XThR.Tn[1] XA.XIR[2].XIC[9].icell.Ien 0.00338f
C5441 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C5442 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00584f
C5443 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.04036f
C5444 XA.XIR[5].XIC[3].icell.SM Vbias 0.00701f
C5445 XA.XIR[14].XIC[0].icell.Ien Iout 0.06411f
C5446 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02762f
C5447 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02762f
C5448 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C5449 XA.XIR[10].XIC[10].icell.PDM VPWR 0.00799f
C5450 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.15202f
C5451 XThR.Tn[13] Iout 1.16236f
C5452 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C5453 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00214f
C5454 XA.XIR[15].XIC[9].icell.PDM Vbias 0.04261f
C5455 XA.XIR[14].XIC[13].icell.PUM VPWR 0.00937f
C5456 a_n1049_6405# XThR.Tn[4] 0.26564f
C5457 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PUM 0.00465f
C5458 XA.XIR[0].XIC[14].icell.Ien Iout 0.06389f
C5459 XA.XIR[1].XIC[14].icell.Ien Vbias 0.21104f
C5460 XA.XIR[13].XIC[11].icell.PDM VPWR 0.00799f
C5461 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C5462 a_10051_9569# VPWR 0.00319f
C5463 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C5464 XA.XIR[5].XIC[10].icell.Ien VPWR 0.1903f
C5465 XA.XIR[15].XIC[8].icell.PUM VPWR 0.00937f
C5466 XA.XIR[3].XIC[8].icell.PDM VPWR 0.00799f
C5467 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PUM 0.00102f
C5468 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11267f
C5469 XA.XIR[5].XIC[6].icell.Ien Iout 0.06417f
C5470 XA.XIR[2].XIC[2].icell.PUM Vbias 0.0031f
C5471 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.SM 0.00168f
C5472 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C5473 XA.XIR[9].XIC[7].icell.PDM Vbias 0.04261f
C5474 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C5475 XThC.TAN2 XThC.TB7 1.11562f
C5476 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00584f
C5477 XThC.TB5 XThC.Tn[8] 0.01728f
C5478 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.SM 0.0039f
C5479 XThC.Tn[12] XA.XIR[0].XIC[11].icell.PDM 0.00106f
C5480 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6] 0.00341f
C5481 XThR.Tn[2] VPWR 6.62952f
C5482 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C5483 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C5484 XThR.TAN a_n997_1803# 0.00228f
C5485 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00214f
C5486 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.SM 0.00168f
C5487 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PDM 0.00598f
C5488 XA.XIR[9].XIC[7].icell.Ien Vbias 0.21098f
C5489 XA.XIR[13].XIC[1].icell.SM VPWR 0.00158f
C5490 XA.XIR[8].XIC[5].icell.PUM VPWR 0.00937f
C5491 XThR.Tn[2] XA.XIR[3].XIC[2].icell.SM 0.00121f
C5492 XA.XIR[12].XIC[3].icell.Ien VPWR 0.1903f
C5493 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.15202f
C5494 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.SM 0.00168f
C5495 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.03425f
C5496 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.SM 0.0039f
C5497 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1909f
C5498 XA.XIR[11].XIC[4].icell.SM VPWR 0.00158f
C5499 XA.XIR[7].XIC[0].icell.PDM Vbias 0.04207f
C5500 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04031f
C5501 XA.XIR[9].XIC[14].icell.PDM Iout 0.00117f
C5502 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9] 0.00341f
C5503 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.15202f
C5504 XThR.Tn[5] XA.XIR[6].XIC[10].icell.Ien 0.00338f
C5505 XA.XIR[4].XIC[3].icell.PUM Vbias 0.0031f
C5506 XA.XIR[9].XIC[14].icell.PUM VPWR 0.00937f
C5507 XA.XIR[2].XIC[7].icell.PUM Vbias 0.0031f
C5508 XA.XIR[10].XIC[6].icell.SM VPWR 0.00158f
C5509 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02762f
C5510 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11] 0.00341f
C5511 XThR.Tn[2] XA.XIR[2].XIC[12].icell.PDM 0.00341f
C5512 XThC.TAN2 VPWR 0.88811f
C5513 XA.XIR[6].XIC[2].icell.Ien VPWR 0.1903f
C5514 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C5515 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.03023f
C5516 XThR.Tn[14] XA.XIR[15].XIC[3].icell.Ien 0.00338f
C5517 XA.XIR[7].XIC[3].icell.Ien Vbias 0.21098f
C5518 XA.XIR[10].XIC[2].icell.SM Iout 0.00388f
C5519 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Iout 0.00347f
C5520 XThR.Tn[9] XA.XIR[10].XIC[2].icell.SM 0.00121f
C5521 XA.XIR[0].XIC[12].icell.PDM Vbias 0.04282f
C5522 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00584f
C5523 XThR.TBN a_n1049_5317# 0.07731f
C5524 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.03425f
C5525 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C5526 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PUM 0.00186f
C5527 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.SM 0.0039f
C5528 XA.XIR[13].XIC_15.icell.Ien Vbias 0.21234f
C5529 XA.XIR[14].XIC[7].icell.SM Vbias 0.00701f
C5530 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00214f
C5531 XA.XIR[4].XIC[8].icell.SM VPWR 0.00158f
C5532 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C5533 XA.XIR[7].XIC[7].icell.PDM Iout 0.00117f
C5534 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.SM 0.0039f
C5535 XA.XIR[2].XIC[12].icell.SM VPWR 0.00158f
C5536 XA.XIR[2].XIC[3].icell.PDM VPWR 0.00799f
C5537 XThC.Tn[8] XThR.Tn[11] 0.28739f
C5538 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8] 0.00341f
C5539 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PUM 0.00465f
C5540 XA.XIR[4].XIC[4].icell.SM Iout 0.00388f
C5541 XA.XIR[8].XIC[13].icell.PUM Vbias 0.0031f
C5542 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02762f
C5543 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.15202f
C5544 XThR.TAN XThR.Tn[13] 0.00276f
C5545 XA.XIR[2].XIC[8].icell.SM Iout 0.00388f
C5546 XA.XIR[7].XIC[10].icell.PUM VPWR 0.00937f
C5547 XThC.Tn[12] XThR.Tn[3] 0.28739f
C5548 XA.XIR[11].XIC[10].icell.Ien VPWR 0.1903f
C5549 XA.XIR[0].XIC[3].icell.PUM Vbias 0.0031f
C5550 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04031f
C5551 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.SM 0.00168f
C5552 XThC.Tn[7] XThR.Tn[7] 0.28739f
C5553 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5554 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00584f
C5555 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00214f
C5556 XA.XIR[14].XIC[11].icell.PUM VPWR 0.00937f
C5557 XThR.Tn[4] XA.XIR[5].XIC[2].icell.Ien 0.00338f
C5558 XA.XIR[3].XIC[7].icell.SM Vbias 0.00701f
C5559 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11] 0.00341f
C5560 XThR.Tn[3] XA.XIR[4].XIC[4].icell.Ien 0.00338f
C5561 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.15202f
C5562 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.03511f
C5563 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C5564 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Ien 0.00232f
C5565 XThC.TAN data[0] 0.0138f
C5566 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.SM 0.00168f
C5567 XA.XIR[0].XIC[8].icell.SM VPWR 0.00158f
C5568 XA.XIR[6].XIC[10].icell.Ien Vbias 0.21098f
C5569 XThR.Tn[11] XA.XIR[12].XIC[3].icell.SM 0.00121f
C5570 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C5571 XA.XIR[8].XIC[14].icell.SM Iout 0.00388f
C5572 XThR.Tn[8] XA.XIR[9].XIC[14].icell.SM 0.00121f
C5573 XA.XIR[4].XIC[7].icell.PDM Vbias 0.04261f
C5574 XThC.TB1 XThC.Tn[0] 0.19116f
C5575 XA.XIR[0].XIC[4].icell.SM Iout 0.00367f
C5576 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.SM 0.00168f
C5577 XA.XIR[1].XIC[4].icell.SM Vbias 0.00704f
C5578 XA.XIR[11].XIC[0].icell.Ien VPWR 0.1903f
C5579 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Ien 0.00584f
C5580 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.03425f
C5581 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5582 XA.XIR[3].XIC[14].icell.Ien VPWR 0.19036f
C5583 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02762f
C5584 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C5585 XThC.TBN XThC.Tn[2] 0.64352f
C5586 XA.XIR[10].XIC[2].icell.PUM VPWR 0.00937f
C5587 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14] 0.00341f
C5588 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02762f
C5589 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.SM 0.0039f
C5590 XA.XIR[3].XIC[10].icell.Ien Iout 0.06417f
C5591 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C5592 XThR.Tn[0] XA.XIR[0].XIC[13].icell.PDM 0.00341f
C5593 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07214f
C5594 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.PDM 0.00591f
C5595 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C5596 XA.XIR[15].XIC[1].icell.Ien Vbias 0.17899f
C5597 XThC.Tn[11] XThR.Tn[12] 0.28739f
C5598 XA.XIR[15].XIC[0].icell.PDM VPWR 0.0114f
C5599 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00214f
C5600 XA.XIR[6].XIC[3].icell.PDM Iout 0.00117f
C5601 XA.XIR[1].XIC[11].icell.Ien VPWR 0.1903f
C5602 XA.XIR[4].XIC[14].icell.PDM Iout 0.00117f
C5603 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C5604 XA.XIR[14].XIC[6].icell.PDM VPWR 0.00799f
C5605 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C5606 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.SM 0.00168f
C5607 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PUM 0.00465f
C5608 XA.XIR[14].XIC[12].icell.Ien VPWR 0.19084f
C5609 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PUM 0.00465f
C5610 XA.XIR[11].XIC[2].icell.PDM Vbias 0.04261f
C5611 XA.XIR[1].XIC[7].icell.Ien Iout 0.06417f
C5612 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02762f
C5613 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.SM 0.0039f
C5614 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.03425f
C5615 XA.XIR[13].XIC[10].icell.PDM VPWR 0.00799f
C5616 XA.XIR[10].XIC[6].icell.PDM Vbias 0.04261f
C5617 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.SM 0.00168f
C5618 XThR.TB4 VPWR 0.92827f
C5619 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Ien 0.00595f
C5620 XThR.Tn[6] XA.XIR[7].XIC[13].icell.SM 0.00121f
C5621 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.SM 0.0039f
C5622 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.SM 0.00168f
C5623 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04031f
C5624 XThC.TB6 a_7651_9569# 0.0046f
C5625 XA.XIR[9].XIC[4].icell.Ien VPWR 0.1903f
C5626 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00584f
C5627 XA.XIR[12].XIC[3].icell.PDM Iout 0.00117f
C5628 a_7875_9569# Vbias 0.00315f
C5629 XThC.Tn[10] XThR.Tn[10] 0.28739f
C5630 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PDM 0.00172f
C5631 XThR.Tn[1] XA.XIR[2].XIC[14].icell.Ien 0.00338f
C5632 XA.XIR[5].XIC[8].icell.SM Vbias 0.00701f
C5633 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C5634 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04031f
C5635 XA.XIR[15].XIC[6].icell.Ien Vbias 0.17899f
C5636 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11153f
C5637 XA.XIR[11].XIC[9].icell.PDM Iout 0.00117f
C5638 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PUM 0.00465f
C5639 XA.XIR[3].XIC[4].icell.PDM Vbias 0.04261f
C5640 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00214f
C5641 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.15202f
C5642 XThR.Tn[0] XA.XIR[1].XIC[5].icell.Ien 0.00338f
C5643 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.03425f
C5644 XA.XIR[2].XIC[4].icell.PUM VPWR 0.00937f
C5645 XA.XIR[5].XIC_15.icell.Ien VPWR 0.25566f
C5646 XA.XIR[8].XIC[3].icell.Ien Vbias 0.21098f
C5647 XA.XIR[5].XIC[11].icell.PDM VPWR 0.00799f
C5648 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00584f
C5649 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00214f
C5650 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00584f
C5651 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C5652 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Iout 0.00347f
C5653 XA.XIR[0].XIC[3].icell.PDM VPWR 0.00774f
C5654 XThR.TB3 XThR.Tn[4] 0.00382f
C5655 XA.XIR[5].XIC[11].icell.Ien Iout 0.06417f
C5656 XThR.TBN XA.XIR[7].XIC_dummy_left.icell.Ien 0.00158f
C5657 XA.XIR[12].XIC[1].icell.SM Vbias 0.00701f
C5658 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.SM 0.0039f
C5659 XThR.TA3 a_n1331_2891# 0.00995f
C5660 XA.XIR[3].XIC[11].icell.PDM Iout 0.00117f
C5661 XA.XIR[8].XIC[13].icell.PDM VPWR 0.00799f
C5662 XA.XIR[14].XIC[4].icell.SM VPWR 0.00158f
C5663 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13] 0.00341f
C5664 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00584f
C5665 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[1].icell.Ien 0.00214f
C5666 XA.XIR[11].XIC[4].icell.PUM Vbias 0.0031f
C5667 XA.XIR[8].XIC[1].icell.PDM Iout 0.00117f
C5668 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.SM 0.00168f
C5669 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04031f
C5670 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00214f
C5671 XA.XIR[13].XIC[6].icell.SM VPWR 0.00158f
C5672 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04031f
C5673 XA.XIR[9].XIC[12].icell.Ien Vbias 0.21098f
C5674 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PUM 0.00465f
C5675 XA.XIR[10].XIC[6].icell.PUM Vbias 0.0031f
C5676 XA.XIR[8].XIC[10].icell.PUM VPWR 0.00937f
C5677 XThR.Tn[2] XA.XIR[3].XIC[7].icell.SM 0.00121f
C5678 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C5679 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07214f
C5680 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00214f
C5681 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C5682 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00256f
C5683 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.SM 0.00168f
C5684 XA.XIR[11].XIC_15.icell.Ien VPWR 0.25566f
C5685 XA.XIR[12].XIC[8].icell.Ien VPWR 0.1903f
C5686 XA.XIR[13].XIC[2].icell.SM Iout 0.00388f
C5687 XThR.Tn[4] XA.XIR[4].XIC[2].icell.PDM 0.00341f
C5688 XThC.TA2 a_7875_9569# 0.00149f
C5689 XThR.TB3 XThR.TB6 0.04428f
C5690 XThR.Tn[5] XThR.Tn[6] 0.06649f
C5691 XThR.Tn[3] XA.XIR[3].XIC[9].icell.PDM 0.00341f
C5692 XA.XIR[7].XIC_15.icell.PDM Vbias 0.04401f
C5693 XA.XIR[1].XIC[10].icell.PDM VPWR 0.00799f
C5694 XA.XIR[12].XIC[4].icell.Ien Iout 0.06417f
C5695 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00214f
C5696 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C5697 XThR.Tn[5] XA.XIR[6].XIC_15.icell.Ien 0.00117f
C5698 XA.XIR[4].XIC[8].icell.PUM Vbias 0.0031f
C5699 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04031f
C5700 XA.XIR[3].XIC[4].icell.SM VPWR 0.00158f
C5701 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C5702 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C5703 XA.XIR[11].XIC[5].icell.SM Iout 0.00388f
C5704 XThC.Tn[8] XThR.Tn[14] 0.28739f
C5705 XA.XIR[2].XIC[12].icell.PUM Vbias 0.0031f
C5706 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C5707 XThC.TB5 XThC.Tn[6] 0.00352f
C5708 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C5709 XThR.Tn[14] XA.XIR[15].XIC[8].icell.Ien 0.00338f
C5710 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.03425f
C5711 XA.XIR[6].XIC[7].icell.Ien VPWR 0.1903f
C5712 XA.XIR[14].XIC[10].icell.Ien VPWR 0.19084f
C5713 XA.XIR[7].XIC[8].icell.Ien Vbias 0.21098f
C5714 XA.XIR[10].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5715 XThC.Tn[4] XThR.Tn[5] 0.28739f
C5716 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11] 0.00341f
C5717 XA.XIR[10].XIC[7].icell.SM Iout 0.00388f
C5718 XThR.Tn[9] XA.XIR[10].XIC[7].icell.SM 0.00121f
C5719 XThC.Tn[8] data[0] 0.01643f
C5720 XA.XIR[6].XIC[3].icell.Ien Iout 0.06417f
C5721 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02803f
C5722 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.03023f
C5723 XA.XIR[1].XIC[1].icell.SM VPWR 0.00158f
C5724 XA.XIR[4].XIC[13].icell.SM VPWR 0.00158f
C5725 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04031f
C5726 XA.XIR[3].XIC[1].icell.Ien Vbias 0.21098f
C5727 XThC.Tn[9] XThR.Tn[4] 0.28739f
C5728 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.SM 0.00168f
C5729 XA.XIR[4].XIC[9].icell.SM Iout 0.00388f
C5730 XA.XIR[11].XIC_dummy_left.icell.SM VPWR 0.00269f
C5731 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C5732 XA.XIR[2].XIC[13].icell.SM Iout 0.00388f
C5733 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.03425f
C5734 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.15202f
C5735 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01577f
C5736 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00584f
C5737 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.03425f
C5738 XA.XIR[5].XIC[0].icell.SM VPWR 0.00158f
C5739 XA.XIR[2].XIC[6].icell.PDM Iout 0.00117f
C5740 XThC.TB4 XThC.TB5 2.06459f
C5741 XThC.TB3 XThC.TAN 0.23315f
C5742 XA.XIR[0].XIC[8].icell.PUM Vbias 0.0031f
C5743 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.SM 0.0039f
C5744 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.SM 0.00168f
C5745 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14] 0.00341f
C5746 XThR.Tn[12] XA.XIR[13].XIC[5].icell.SM 0.00121f
C5747 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02762f
C5748 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C5749 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C5750 XThR.Tn[4] XA.XIR[5].XIC[7].icell.Ien 0.00338f
C5751 XThR.TB3 XThR.Tn[8] 0.00178f
C5752 XA.XIR[3].XIC[12].icell.SM Vbias 0.00701f
C5753 XThR.Tn[1] XA.XIR[2].XIC[4].icell.SM 0.00121f
C5754 XA.XIR[13].XIC[2].icell.PUM VPWR 0.00937f
C5755 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[6].icell.Ien 0.00214f
C5756 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.15202f
C5757 XThR.Tn[6] Vbias 3.74624f
C5758 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00214f
C5759 XThR.Tn[3] XA.XIR[4].XIC[9].icell.Ien 0.00338f
C5760 XThR.Tn[1] a_n1049_7787# 0.26879f
C5761 XA.XIR[10].XIC[0].icell.Ien Vbias 0.20951f
C5762 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04031f
C5763 XA.XIR[6].XIC_15.icell.Ien Vbias 0.21234f
C5764 XA.XIR[0].XIC[13].icell.SM VPWR 0.00158f
C5765 XA.XIR[6].XIC[11].icell.PDM Vbias 0.04261f
C5766 XThC.Tn[1] XThR.Tn[3] 0.28739f
C5767 XThR.Tn[11] XA.XIR[12].XIC[8].icell.SM 0.00121f
C5768 XThC.Tn[6] XThR.Tn[11] 0.28739f
C5769 XThC.Tn[11] XThR.Tn[0] 0.28749f
C5770 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PUM 0.00465f
C5771 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00214f
C5772 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5] 0.00341f
C5773 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.SM 0.00168f
C5774 XA.XIR[0].XIC[9].icell.SM Iout 0.00367f
C5775 Vbias bias[0] 0.17404f
C5776 XA.XIR[1].XIC[9].icell.SM Vbias 0.00704f
C5777 bias[1] bias[2] 0.03172f
C5778 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.SM 0.0039f
C5779 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PUM 0.00176f
C5780 XThC.Tn[4] Vbias 2.48532f
C5781 XA.XIR[14].XIC[2].icell.PDM Vbias 0.04261f
C5782 XA.XIR[5].XIC[5].icell.SM VPWR 0.00158f
C5783 XThR.Tn[7] Iout 1.16233f
C5784 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PUM 0.00465f
C5785 XA.XIR[15].XIC[3].icell.Ien VPWR 0.32895f
C5786 XThC.TAN XThC.TB7 0.33493f
C5787 XThR.Tn[5] XA.XIR[6].XIC[0].icell.SM 0.00121f
C5788 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C5789 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.SM 0.0039f
C5790 XA.XIR[7].XIC_15.icell.SM Iout 0.0047f
C5791 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02762f
C5792 XA.XIR[5].XIC[1].icell.SM Iout 0.00388f
C5793 XA.XIR[3].XIC_15.icell.Ien Iout 0.0642f
C5794 XA.XIR[13].XIC[6].icell.PDM Vbias 0.04261f
C5795 XThC.TAN2 a_7875_9569# 0.01939f
C5796 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00584f
C5797 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01432f
C5798 XThC.Tn[5] XThR.Tn[6] 0.28739f
C5799 XThR.TB2 XThR.Tn[2] 0.00271f
C5800 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00214f
C5801 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.SM 0.0039f
C5802 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C5803 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6] 0.00341f
C5804 XThR.TAN a_n997_3979# 0.01152f
C5805 XA.XIR[15].XIC[3].icell.PDM Iout 0.00117f
C5806 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02762f
C5807 XThR.Tn[1] XA.XIR[1].XIC[14].icell.PDM 0.00341f
C5808 XThC.Tn[10] XThR.Tn[13] 0.28739f
C5809 XA.XIR[9].XIC[2].icell.SM Vbias 0.00701f
C5810 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.SM 0.0039f
C5811 XA.XIR[1].XIC[12].icell.Ien Iout 0.06417f
C5812 XA.XIR[14].XIC[9].icell.PDM Iout 0.00117f
C5813 XThC.Tn[4] XThC.Tn[5] 0.4169f
C5814 XA.XIR[9].XIC[13].icell.PDM VPWR 0.00799f
C5815 XThC.Tn[13] Iout 0.84238f
C5816 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PUM 0.00465f
C5817 XThC.Tn[13] XThR.Tn[9] 0.2874f
C5818 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.SM 0.0039f
C5819 XA.XIR[7].XIC[0].icell.Ien VPWR 0.1903f
C5820 XThC.TBN a_2979_9615# 0.0607f
C5821 XThC.Tn[0] XThR.Tn[12] 0.28741f
C5822 XThC.TAN VPWR 1.32988f
C5823 XA.XIR[9].XIC[1].icell.PDM Iout 0.00117f
C5824 XThR.TA1 XThR.TB4 0.02767f
C5825 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C5826 XThC.Tn[9] XThR.Tn[8] 0.28739f
C5827 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9] 0.00341f
C5828 XThR.Tn[5] XA.XIR[6].XIC[5].icell.SM 0.00121f
C5829 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.15202f
C5830 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00584f
C5831 XA.XIR[9].XIC[9].icell.Ien VPWR 0.1903f
C5832 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.SM 0.00168f
C5833 XA.XIR[10].XIC[3].icell.PUM VPWR 0.00937f
C5834 XA.XIR[2].XIC[2].icell.Ien Vbias 0.21098f
C5835 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00584f
C5836 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C5837 XA.XIR[5].XIC[13].icell.SM Vbias 0.00701f
C5838 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PUM 0.00465f
C5839 XA.XIR[5].XIC[7].icell.PDM Vbias 0.04261f
C5840 XA.XIR[9].XIC[5].icell.Ien Iout 0.06417f
C5841 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C5842 XA.XIR[12].XIC[12].icell.SM Iout 0.00388f
C5843 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.15202f
C5844 XThR.TB7 a_n1049_5317# 0.27822f
C5845 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04031f
C5846 XA.XIR[11].XIC[14].icell.PDM VPWR 0.00809f
C5847 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04031f
C5848 XThR.Tn[0] XA.XIR[1].XIC[10].icell.Ien 0.00338f
C5849 XA.XIR[7].XIC[6].icell.PDM VPWR 0.00799f
C5850 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PUM 0.00465f
C5851 XA.XIR[8].XIC[9].icell.PDM Vbias 0.04261f
C5852 XA.XIR[6].XIC[0].icell.SM Vbias 0.00675f
C5853 XThC.TB4 XThC.Tn[3] 0.18952f
C5854 XA.XIR[14].XIC[4].icell.PUM Vbias 0.0031f
C5855 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10] 0.00341f
C5856 XA.XIR[4].XIC[5].icell.PUM VPWR 0.00937f
C5857 XA.XIR[2].XIC[9].icell.PUM VPWR 0.00937f
C5858 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.15222f
C5859 XThR.TB1 XThR.TB6 0.05751f
C5860 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14] 0.00341f
C5861 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.SM 0.00168f
C5862 XThR.Tn[2] XA.XIR[3].XIC[1].icell.Ien 0.00338f
C5863 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C5864 XA.XIR[13].XIC[6].icell.PUM Vbias 0.0031f
C5865 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07214f
C5866 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.03425f
C5867 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.SM 0.00168f
C5868 XA.XIR[8].XIC[8].icell.Ien Vbias 0.21098f
C5869 XA.XIR[14].XIC_15.icell.Ien VPWR 0.25598f
C5870 XA.XIR[7].XIC[5].icell.Ien VPWR 0.1903f
C5871 XThC.Tn[9] XThR.Tn[1] 0.28739f
C5872 XA.XIR[5].XIC_dummy_right.icell.SM VPWR 0.00123f
C5873 XA.XIR[12].XIC[6].icell.SM Vbias 0.00701f
C5874 XA.XIR[5].XIC[14].icell.PDM Iout 0.00117f
C5875 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.SM 0.00168f
C5876 XA.XIR[10].XIC_15.icell.PDM Vbias 0.04401f
C5877 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PUM 0.00465f
C5878 XA.XIR[1].XIC[6].icell.PDM Vbias 0.04261f
C5879 XA.XIR[11].XIC[9].icell.PUM Vbias 0.0031f
C5880 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11] 0.00341f
C5881 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00584f
C5882 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_15.icell.SM 0.0039f
C5883 XThR.TAN XThR.Tn[7] 0.07415f
C5884 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.SM 0.0039f
C5885 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00584f
C5886 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.SM 0.00168f
C5887 XThC.TAN a_5155_9615# 0.00268f
C5888 XA.XIR[14].XIC[5].icell.SM Iout 0.00388f
C5889 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11154f
C5890 XThR.TAN a_n997_2891# 0.0168f
C5891 XA.XIR[3].XIC[4].icell.PUM Vbias 0.0031f
C5892 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.15202f
C5893 XThR.Tn[7] XA.XIR[8].XIC[2].icell.Ien 0.00338f
C5894 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01577f
C5895 XThR.Tn[2] XA.XIR[3].XIC[12].icell.SM 0.00121f
C5896 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.SM 0.00168f
C5897 XA.XIR[6].XIC[5].icell.SM Vbias 0.00701f
C5898 XA.XIR[13].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5899 XA.XIR[0].XIC[5].icell.PUM VPWR 0.00877f
C5900 XA.XIR[13].XIC[7].icell.SM Iout 0.00388f
C5901 XThC.TB2 XThC.Tn[9] 0.292f
C5902 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PUM 0.00465f
C5903 XA.XIR[11].XIC_dummy_right.icell.SM VPWR 0.00123f
C5904 a_3773_9615# XThC.Tn[2] 0.01175f
C5905 XThC.TB2 XThC.TBN 0.2075f
C5906 XThC.TB3 XThC.Tn[8] 0.00178f
C5907 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.03546f
C5908 XA.XIR[12].XIC[9].icell.Ien Iout 0.06417f
C5909 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.SM 0.0039f
C5910 XThR.TB3 a_n997_3755# 0.0061f
C5911 XA.XIR[4].XIC[13].icell.PUM Vbias 0.0031f
C5912 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C5913 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14] 0.00341f
C5914 XA.XIR[3].XIC[9].icell.SM VPWR 0.00158f
C5915 XThC.Tn[4] XThR.Tn[2] 0.28739f
C5916 XA.XIR[14].XIC[0].icell.PUM VPWR 0.00937f
C5917 XA.XIR[1].XIC[13].icell.PDM Iout 0.00117f
C5918 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C5919 XA.XIR[2].XIC[14].icell.PDM Vbias 0.04261f
C5920 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.SM 0.00168f
C5921 XThR.Tn[10] XA.XIR[11].XIC[3].icell.Ien 0.00338f
C5922 XThR.TB1 XThR.Tn[8] 0.29191f
C5923 XA.XIR[3].XIC[5].icell.SM Iout 0.00388f
C5924 XThR.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.00353f
C5925 XA.XIR[6].XIC[12].icell.Ien VPWR 0.1903f
C5926 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00584f
C5927 XA.XIR[7].XIC[13].icell.Ien Vbias 0.21098f
C5928 XA.XIR[9].XIC[0].icell.Ien Iout 0.06411f
C5929 XA.XIR[6].XIC[2].icell.PDM VPWR 0.00799f
C5930 XThR.Tn[11] XA.XIR[12].XIC[13].icell.SM 0.00121f
C5931 XA.XIR[5].XIC[0].icell.Ien Vbias 0.20951f
C5932 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.15202f
C5933 XA.XIR[4].XIC[13].icell.PDM VPWR 0.00799f
C5934 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PUM 0.00465f
C5935 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.15202f
C5936 XA.XIR[6].XIC[8].icell.Ien Iout 0.06417f
C5937 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.15202f
C5938 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7] 0.00341f
C5939 XA.XIR[1].XIC[6].icell.SM VPWR 0.00158f
C5940 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C5941 XA.XIR[4].XIC[1].icell.PDM Iout 0.00117f
C5942 XThC.TB6 a_5949_9615# 0.26831f
C5943 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00214f
C5944 a_6243_9615# Vbias 0.01019f
C5945 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C5946 XA.XIR[1].XIC[2].icell.SM Iout 0.00388f
C5947 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00584f
C5948 XA.XIR[8].XIC_15.icell.SM Iout 0.0047f
C5949 XA.XIR[4].XIC[14].icell.SM Iout 0.00388f
C5950 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C5951 XA.XIR[13].XIC[0].icell.Ien Vbias 0.20951f
C5952 XThC.TB7 XThC.Tn[8] 0.07806f
C5953 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.15202f
C5954 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.15202f
C5955 XThR.TB2 XThR.TB4 0.04006f
C5956 XA.XIR[0].XIC[13].icell.PUM Vbias 0.0031f
C5957 XA.XIR[12].XIC[2].icell.PUM Vbias 0.0031f
C5958 XA.XIR[12].XIC[2].icell.PDM VPWR 0.00799f
C5959 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PUM 0.00465f
C5960 XThC.Tn[6] XThR.Tn[14] 0.28739f
C5961 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04031f
C5962 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C5963 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.SM 0.00168f
C5964 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.0353f
C5965 XA.XIR[12].XIC[10].icell.SM Iout 0.00388f
C5966 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.03425f
C5967 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.03425f
C5968 XA.XIR[11].XIC[8].icell.PDM VPWR 0.00799f
C5969 XThR.Tn[4] XA.XIR[5].XIC[12].icell.Ien 0.00338f
C5970 XThR.TB1 XThR.Tn[1] 0.0099f
C5971 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.03425f
C5972 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.15202f
C5973 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C5974 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04031f
C5975 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C5976 XA.XIR[5].XIC[5].icell.PUM Vbias 0.0031f
C5977 XThR.Tn[1] XA.XIR[2].XIC[9].icell.SM 0.00121f
C5978 XThR.Tn[3] XA.XIR[4].XIC[14].icell.Ien 0.00338f
C5979 XA.XIR[15].XIC[1].icell.SM Vbias 0.00701f
C5980 a_6243_9615# XThC.Tn[5] 0.00158f
C5981 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02762f
C5982 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PUM 0.00465f
C5983 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C5984 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C5985 XA.XIR[10].XIC[0].icell.PDM Iout 0.00117f
C5986 XThC.Tn[7] XThR.Tn[4] 0.28739f
C5987 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04037f
C5988 XA.XIR[0].XIC[14].icell.SM Iout 0.00367f
C5989 XA.XIR[1].XIC[14].icell.SM Vbias 0.00704f
C5990 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PUM 0.00465f
C5991 XThC.Tn[8] VPWR 6.8418f
C5992 XA.XIR[7].XIC_dummy_left.icell.SM VPWR 0.00269f
C5993 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.SM 0.00168f
C5994 XA.XIR[15].XIC[8].icell.Ien VPWR 0.32895f
C5995 XA.XIR[5].XIC[10].icell.SM VPWR 0.00158f
C5996 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00214f
C5997 XA.XIR[3].XIC[10].icell.PDM VPWR 0.00799f
C5998 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00214f
C5999 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.SM 0.0039f
C6000 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C6001 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00584f
C6002 XA.XIR[5].XIC[6].icell.SM Iout 0.00388f
C6003 XA.XIR[15].XIC[4].icell.Ien Iout 0.06807f
C6004 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.15202f
C6005 XA.XIR[9].XIC[9].icell.PDM Vbias 0.04261f
C6006 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PUM 0.00465f
C6007 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.SM 0.00168f
C6008 XA.XIR[8].XIC[0].icell.PDM VPWR 0.00799f
C6009 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PUM 0.00465f
C6010 XThC.Tn[0] XThR.Tn[0] 0.28807f
C6011 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00214f
C6012 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6] 0.00341f
C6013 XA.XIR[11].XIC[13].icell.PDM VPWR 0.00799f
C6014 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.SM 0.0039f
C6015 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.03425f
C6016 XA.XIR[13].XIC[3].icell.PUM VPWR 0.00937f
C6017 XA.XIR[9].XIC[7].icell.SM Vbias 0.00701f
C6018 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C6019 XA.XIR[8].XIC[5].icell.Ien VPWR 0.1903f
C6020 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.SM 0.0039f
C6021 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.SM 0.0039f
C6022 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01745f
C6023 XA.XIR[12].XIC[3].icell.SM VPWR 0.00158f
C6024 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C6025 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00584f
C6026 XA.XIR[14].XIC[14].icell.PDM VPWR 0.00809f
C6027 XThR.TB4 XThR.TAN2 0.03415f
C6028 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00584f
C6029 a_n1335_4229# data[4] 0.00451f
C6030 VPWR bias[2] 1.5142f
C6031 XA.XIR[11].XIC[6].icell.PUM VPWR 0.00937f
C6032 XA.XIR[7].XIC[2].icell.PDM Vbias 0.04261f
C6033 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00214f
C6034 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6035 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04031f
C6036 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.SM 0.0039f
C6037 XThR.Tn[11] XA.XIR[12].XIC[11].icell.SM 0.00121f
C6038 XThR.Tn[5] XA.XIR[6].XIC[10].icell.SM 0.00121f
C6039 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.15202f
C6040 XA.XIR[7].XIC[1].icell.Ien Iout 0.06417f
C6041 XA.XIR[4].XIC[3].icell.Ien Vbias 0.21098f
C6042 XA.XIR[10].XIC[14].icell.PDM Vbias 0.04261f
C6043 XA.XIR[9].XIC[14].icell.Ien VPWR 0.19036f
C6044 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C6045 XA.XIR[10].XIC[8].icell.PUM VPWR 0.00937f
C6046 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PUM 0.00465f
C6047 XThR.TB4 XThR.Tn[6] 0.00605f
C6048 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00214f
C6049 XThR.TB5 XThR.Tn[5] 0.01094f
C6050 XA.XIR[2].XIC[7].icell.Ien Vbias 0.21098f
C6051 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11] 0.00341f
C6052 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00256f
C6053 XThR.Tn[2] XA.XIR[2].XIC[14].icell.PDM 0.00341f
C6054 XThR.Tn[14] XA.XIR[15].XIC[3].icell.SM 0.00121f
C6055 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Iout 0.00347f
C6056 XA.XIR[9].XIC[10].icell.Ien Iout 0.06417f
C6057 XA.XIR[6].XIC[2].icell.SM VPWR 0.00158f
C6058 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.15202f
C6059 XA.XIR[7].XIC[3].icell.SM Vbias 0.00701f
C6060 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00214f
C6061 XA.XIR[0].XIC[14].icell.PDM Vbias 0.04282f
C6062 XA.XIR[13].XIC_15.icell.PDM Vbias 0.04401f
C6063 XThR.Tn[0] XA.XIR[1].XIC_15.icell.Ien 0.00117f
C6064 XA.XIR[12].XIC[14].icell.Ien Iout 0.06417f
C6065 XThC.Tn[2] Iout 0.84806f
C6066 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C6067 XThC.Tn[2] XThR.Tn[9] 0.28739f
C6068 XA.XIR[4].XIC[10].icell.PUM VPWR 0.00937f
C6069 XA.XIR[14].XIC[9].icell.PUM Vbias 0.0031f
C6070 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6071 XA.XIR[2].XIC[14].icell.PUM VPWR 0.00937f
C6072 XThR.TAN a_n997_1579# 0.00209f
C6073 XA.XIR[7].XIC[9].icell.PDM Iout 0.00117f
C6074 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C6075 XA.XIR[2].XIC[5].icell.PDM VPWR 0.00799f
C6076 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00584f
C6077 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00584f
C6078 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8] 0.00341f
C6079 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.03425f
C6080 XThC.Tn[7] XThR.Tn[8] 0.28739f
C6081 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00584f
C6082 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C6083 XA.XIR[8].XIC[13].icell.Ien Vbias 0.21098f
C6084 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14] 0.00341f
C6085 XA.XIR[7].XIC[10].icell.Ien VPWR 0.1903f
C6086 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.389f
C6087 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C6088 XA.XIR[0].XIC[3].icell.Ien Vbias 0.21128f
C6089 XA.XIR[14].XIC_dummy_right.icell.SM VPWR 0.00123f
C6090 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00214f
C6091 XA.XIR[7].XIC[6].icell.Ien Iout 0.06417f
C6092 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C6093 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.SM 0.0039f
C6094 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.SM 0.00168f
C6095 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04031f
C6096 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00256f
C6097 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C6098 XThR.Tn[4] XA.XIR[5].XIC[2].icell.SM 0.00121f
C6099 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00214f
C6100 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.SM 0.0039f
C6101 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[3].icell.SM 0.0039f
C6102 XA.XIR[3].XIC[9].icell.PUM Vbias 0.0031f
C6103 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.SM 0.0039f
C6104 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.03425f
C6105 XThR.Tn[3] XA.XIR[4].XIC[4].icell.SM 0.00121f
C6106 XThR.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.00338f
C6107 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PUM 0.00465f
C6108 XA.XIR[8].XIC[0].icell.Ien VPWR 0.1903f
C6109 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00214f
C6110 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.SM 0.00168f
C6111 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C6112 XThR.TA3 a_n1049_6405# 0.02287f
C6113 XA.XIR[6].XIC[10].icell.SM Vbias 0.00701f
C6114 XA.XIR[0].XIC[10].icell.PUM VPWR 0.00877f
C6115 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C6116 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PUM 0.00465f
C6117 XA.XIR[4].XIC[9].icell.PDM Vbias 0.04261f
C6118 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.03425f
C6119 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Ien 0.00584f
C6120 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00584f
C6121 XA.XIR[1].XIC[6].icell.PUM Vbias 0.0031f
C6122 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C6123 XThC.Tn[7] XThR.Tn[1] 0.2877f
C6124 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.15202f
C6125 XA.XIR[3].XIC[14].icell.SM VPWR 0.00207f
C6126 XThC.TAN a_7875_9569# 0.01174f
C6127 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02762f
C6128 XThR.Tn[0] XA.XIR[0].XIC_15.icell.PDM 0.00341f
C6129 XThR.Tn[10] XA.XIR[11].XIC[8].icell.Ien 0.00338f
C6130 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C6131 XA.XIR[3].XIC[10].icell.SM Iout 0.00388f
C6132 XA.XIR[15].XIC[2].icell.PDM VPWR 0.0114f
C6133 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02762f
C6134 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.SM 0.00168f
C6135 XA.XIR[6].XIC[13].icell.Ien Iout 0.06417f
C6136 XA.XIR[1].XIC[11].icell.SM VPWR 0.00158f
C6137 XA.XIR[6].XIC[5].icell.PDM Iout 0.00117f
C6138 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.15202f
C6139 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C6140 XA.XIR[14].XIC[8].icell.PDM VPWR 0.00799f
C6141 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.03425f
C6142 XThR.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.00341f
C6143 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.03425f
C6144 XThR.Tn[0] XA.XIR[1].XIC[0].icell.SM 0.00121f
C6145 XA.XIR[11].XIC[4].icell.PDM Vbias 0.04261f
C6146 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C6147 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PDM 0.0059f
C6148 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C6149 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C6150 XA.XIR[6].XIC_dummy_right.icell.Ien Vbias 0.00288f
C6151 XA.XIR[15].XIC[12].icell.SM Iout 0.00388f
C6152 XA.XIR[1].XIC[7].icell.SM Iout 0.00388f
C6153 XThC.TB3 XThC.Tn[6] 0.00301f
C6154 XThR.Tn[11] XA.XIR[12].XIC[9].icell.SM 0.00121f
C6155 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00584f
C6156 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.15202f
C6157 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.15202f
C6158 XA.XIR[10].XIC[8].icell.PDM Vbias 0.04261f
C6159 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00214f
C6160 XA.XIR[9].XIC[0].icell.PDM VPWR 0.00799f
C6161 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.SM 0.0039f
C6162 XThC.Tn[10] XThR.Tn[7] 0.28739f
C6163 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C6164 XA.XIR[13].XIC[0].icell.PDM Iout 0.00117f
C6165 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PUM 0.00186f
C6166 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.03425f
C6167 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04052f
C6168 XA.XIR[12].XIC[5].icell.PDM Iout 0.00117f
C6169 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PUM 0.00465f
C6170 XThC.TB6 a_8739_9569# 0.00466f
C6171 XA.XIR[9].XIC[4].icell.SM VPWR 0.00158f
C6172 XThR.TB3 data[4] 0.03253f
C6173 XThR.TA3 data[6] 0.00197f
C6174 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6175 XA.XIR[12].XIC[12].icell.Ien Iout 0.06417f
C6176 a_8963_9569# Vbias 0.00243f
C6177 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.15202f
C6178 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Iout 0.00347f
C6179 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.SM 0.0039f
C6180 XA.XIR[5].XIC[10].icell.PUM Vbias 0.0031f
C6181 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[11].icell.Ien 0.00214f
C6182 XThR.Tn[1] XA.XIR[2].XIC[14].icell.SM 0.00121f
C6183 XA.XIR[15].XIC[6].icell.SM Vbias 0.00701f
C6184 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00214f
C6185 XA.XIR[11].XIC[12].icell.PDM VPWR 0.00799f
C6186 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04031f
C6187 XA.XIR[3].XIC[6].icell.PDM Vbias 0.04261f
C6188 XThC.TB3 XThC.TB4 2.13136f
C6189 a_n1049_6699# XThR.Tn[4] 0.00158f
C6190 XThR.Tn[0] XA.XIR[1].XIC[5].icell.SM 0.00121f
C6191 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PUM 0.00465f
C6192 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C6193 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00584f
C6194 XA.XIR[8].XIC[1].icell.Ien Iout 0.06417f
C6195 XThC.TB7 XThC.Tn[6] 0.2144f
C6196 XA.XIR[14].XIC[13].icell.PDM VPWR 0.00799f
C6197 XThR.Tn[8] XA.XIR[9].XIC[1].icell.Ien 0.00338f
C6198 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C6199 XA.XIR[2].XIC[4].icell.Ien VPWR 0.1903f
C6200 XThC.Tn[11] XThC.Tn[12] 0.22144f
C6201 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00584f
C6202 XA.XIR[5].XIC[13].icell.PDM VPWR 0.00799f
C6203 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PUM 0.00465f
C6204 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PUM 0.00465f
C6205 XA.XIR[8].XIC[3].icell.SM Vbias 0.00701f
C6206 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C6207 XThC.TBN XThC.Tn[14] 0.50214f
C6208 XA.XIR[10].XIC[13].icell.PDM Vbias 0.04261f
C6209 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04031f
C6210 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00214f
C6211 XA.XIR[12].XIC[3].icell.PUM Vbias 0.0031f
C6212 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PUM 0.00429f
C6213 XA.XIR[0].XIC[5].icell.PDM VPWR 0.00908f
C6214 XA.XIR[5].XIC[11].icell.SM Iout 0.00388f
C6215 XA.XIR[15].XIC[9].icell.Ien Iout 0.06807f
C6216 XA.XIR[5].XIC[1].icell.PDM Iout 0.00117f
C6217 XA.XIR[3].XIC[13].icell.PDM Iout 0.00117f
C6218 XA.XIR[14].XIC[6].icell.PUM VPWR 0.00937f
C6219 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07214f
C6220 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13] 0.00341f
C6221 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C6222 XA.XIR[11].XIC[4].icell.Ien Vbias 0.21098f
C6223 XA.XIR[8].XIC[3].icell.PDM Iout 0.00117f
C6224 XA.XIR[13].XIC[14].icell.PDM Vbias 0.04261f
C6225 XThR.Tn[4] Iout 1.16233f
C6226 XA.XIR[13].XIC[8].icell.PUM VPWR 0.00937f
C6227 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PUM 0.00465f
C6228 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04031f
C6229 XA.XIR[9].XIC[12].icell.SM Vbias 0.00701f
C6230 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02762f
C6231 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.03425f
C6232 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04031f
C6233 XThC.TB2 a_3773_9615# 0.2342f
C6234 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.SM 0.0039f
C6235 XA.XIR[8].XIC[10].icell.Ien VPWR 0.1903f
C6236 XA.XIR[10].XIC[6].icell.Ien Vbias 0.21098f
C6237 XThC.TB4 XThC.TB7 0.03475f
C6238 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.SM 0.00168f
C6239 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C6240 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C6241 XA.XIR[12].XIC[8].icell.SM VPWR 0.00158f
C6242 XThC.TA3 XThC.TB6 0.19112f
C6243 XA.XIR[8].XIC[6].icell.Ien Iout 0.06417f
C6244 XThC.Tn[6] VPWR 5.90436f
C6245 XThR.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.00341f
C6246 XThC.TB1 XThC.TB6 0.05752f
C6247 XThR.Tn[8] XA.XIR[9].XIC[6].icell.Ien 0.00338f
C6248 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14] 0.00341f
C6249 XThR.Tn[3] XA.XIR[3].XIC[11].icell.PDM 0.00341f
C6250 XA.XIR[12].XIC[4].icell.SM Iout 0.00388f
C6251 XThC.TB6 XThC.Tn[11] 0.02513f
C6252 XA.XIR[1].XIC[12].icell.PDM VPWR 0.008f
C6253 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C6254 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.04036f
C6255 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00214f
C6256 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.SM 0.0039f
C6257 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6258 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.15202f
C6259 XA.XIR[3].XIC[6].icell.PUM VPWR 0.00937f
C6260 XA.XIR[4].XIC[8].icell.Ien Vbias 0.21098f
C6261 XThR.TBN XThR.Tn[12] 0.50762f
C6262 XA.XIR[1].XIC[0].icell.PDM Iout 0.00117f
C6263 XThR.Tn[6] XA.XIR[7].XIC[0].icell.Ien 0.00338f
C6264 XA.XIR[2].XIC[12].icell.Ien Vbias 0.21098f
C6265 XA.XIR[2].XIC[1].icell.PDM Vbias 0.04261f
C6266 XThR.Tn[11] XA.XIR[12].XIC[13].icell.Ien 0.00338f
C6267 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C6268 XThR.TB6 XThR.Tn[9] 0.0246f
C6269 XA.XIR[6].XIC[7].icell.SM VPWR 0.00158f
C6270 XThR.Tn[14] XA.XIR[15].XIC[8].icell.SM 0.00121f
C6271 XThR.TB3 a_n997_2667# 0.002f
C6272 XA.XIR[9].XIC_15.icell.Ien Iout 0.0642f
C6273 XA.XIR[7].XIC[8].icell.SM Vbias 0.00701f
C6274 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C6275 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C6276 XA.XIR[15].XIC[10].icell.SM Iout 0.00388f
C6277 XA.XIR[4].XIC[0].icell.PDM VPWR 0.00799f
C6278 XA.XIR[8].XIC_dummy_left.icell.SM VPWR 0.00269f
C6279 XA.XIR[6].XIC[3].icell.SM Iout 0.00388f
C6280 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02762f
C6281 XA.XIR[1].XIC[3].icell.PUM VPWR 0.00937f
C6282 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.SM 0.0039f
C6283 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C6284 XThC.TB4 VPWR 0.91479f
C6285 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00214f
C6286 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C6287 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01577f
C6288 XA.XIR[0].XIC_dummy_left.icell.Ien Vbias 0.00348f
C6289 XThC.Tn[0] XA.XIR[6].XIC_dummy_left.icell.Iout 0.00109f
C6290 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.SM 0.0039f
C6291 XThC.TAN XThC.Tn[4] 0.00356f
C6292 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C6293 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04031f
C6294 XThR.Tn[13] XA.XIR[14].XIC[3].icell.Ien 0.00338f
C6295 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C6296 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.03425f
C6297 XA.XIR[12].XIC[10].icell.Ien Iout 0.06417f
C6298 XA.XIR[5].XIC[2].icell.PUM VPWR 0.00937f
C6299 XA.XIR[7].XIC_15.icell.Ien VPWR 0.25566f
C6300 XA.XIR[2].XIC[8].icell.PDM Iout 0.00117f
C6301 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C6302 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.15202f
C6303 XA.XIR[0].XIC[8].icell.Ien Vbias 0.2113f
C6304 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00214f
C6305 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C6306 XA.XIR[7].XIC[11].icell.Ien Iout 0.06417f
C6307 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.03425f
C6308 XThR.Tn[6] XA.XIR[7].XIC[5].icell.Ien 0.00338f
C6309 XA.XIR[14].XIC[1].icell.PUM VPWR 0.00937f
C6310 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00214f
C6311 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.SM 0.00168f
C6312 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00584f
C6313 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.SM 0.00168f
C6314 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Iout 0.00347f
C6315 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00584f
C6316 XThR.Tn[4] XA.XIR[5].XIC[7].icell.SM 0.00121f
C6317 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02762f
C6318 XA.XIR[3].XIC[14].icell.PUM Vbias 0.0031f
C6319 XThR.Tn[11] XA.XIR[12].XIC[14].icell.SM 0.00121f
C6320 XThR.Tn[7] XA.XIR[8].XIC[12].icell.Ien 0.00338f
C6321 XThR.Tn[3] XA.XIR[4].XIC[9].icell.SM 0.00121f
C6322 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.SM 0.00168f
C6323 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.SM 0.00168f
C6324 XA.XIR[10].XIC[0].icell.SM Vbias 0.00675f
C6325 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C6326 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C6327 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01499f
C6328 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04031f
C6329 XA.XIR[6].XIC[13].icell.PDM Vbias 0.04261f
C6330 a_5949_10571# VPWR 0.00653f
C6331 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.03425f
C6332 XThR.Tn[8] Iout 1.16233f
C6333 XThR.Tn[8] XThR.Tn[9] 0.05786f
C6334 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C6335 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5] 0.00341f
C6336 XThR.TAN XThR.Tn[4] 0.00356f
C6337 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6338 XA.XIR[1].XIC[11].icell.PUM Vbias 0.0031f
C6339 XA.XIR[4].XIC_15.icell.SM Iout 0.0047f
C6340 XThC.TB5 XThC.Tn[9] 0.01732f
C6341 XA.XIR[14].XIC[4].icell.PDM Vbias 0.04261f
C6342 XA.XIR[5].XIC[7].icell.PUM VPWR 0.00937f
C6343 XThC.TB4 a_5155_9615# 0.01546f
C6344 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.SM 0.0039f
C6345 XA.XIR[15].XIC[3].icell.SM VPWR 0.00158f
C6346 XThC.TB5 XThC.TBN 0.162f
C6347 XThR.TA3 XThR.TB3 0.57441f
C6348 XA.XIR[11].XIC[1].icell.Ien Iout 0.06417f
C6349 XThR.TB1 data[4] 0.06453f
C6350 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.SM 0.0039f
C6351 XA.XIR[13].XIC[8].icell.PDM Vbias 0.04261f
C6352 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6353 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01432f
C6354 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PUM 0.00465f
C6355 XThC.TAN2 a_8963_9569# 0.01679f
C6356 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00584f
C6357 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C6358 XA.XIR[11].XIC[11].icell.PDM VPWR 0.00799f
C6359 XA.XIR[9].XIC[0].icell.SM Iout 0.00388f
C6360 XA.XIR[1].XIC[0].icell.Ien Iout 0.06411f
C6361 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00584f
C6362 XA.XIR[2].XIC[0].icell.Ien Vbias 0.20951f
C6363 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6] 0.00341f
C6364 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.15202f
C6365 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.SM 0.00168f
C6366 XA.XIR[15].XIC[5].icell.PDM Iout 0.00117f
C6367 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00214f
C6368 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C6369 XThR.TAN XThR.TB6 0.30244f
C6370 XA.XIR[9].XIC[4].icell.PUM Vbias 0.0031f
C6371 XA.XIR[1].XIC[12].icell.SM Iout 0.00388f
C6372 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PUM 0.00465f
C6373 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PUM 0.00465f
C6374 XA.XIR[4].XIC[0].icell.Ien VPWR 0.1903f
C6375 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PUM 0.00465f
C6376 XA.XIR[14].XIC[12].icell.PDM VPWR 0.00799f
C6377 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00584f
C6378 XThR.Tn[1] Iout 1.16236f
C6379 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C6380 XA.XIR[15].XIC[14].icell.Ien Iout 0.06807f
C6381 XA.XIR[11].XIC[12].icell.SM Vbias 0.00701f
C6382 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C6383 XA.XIR[0].XIC_15.icell.SM Iout 0.00367f
C6384 XA.XIR[1].XIC_15.icell.SM Vbias 0.00704f
C6385 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07214f
C6386 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C6387 XA.XIR[7].XIC[0].icell.SM VPWR 0.00158f
C6388 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.03425f
C6389 XThR.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.00338f
C6390 XThC.TBN a_4067_9615# 0.08456f
C6391 XA.XIR[10].XIC[12].icell.PDM Vbias 0.04261f
C6392 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.SM 0.0039f
C6393 XA.XIR[9].XIC[3].icell.PDM Iout 0.00117f
C6394 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9] 0.00341f
C6395 XThR.Tn[12] XA.XIR[13].XIC[1].icell.Ien 0.00338f
C6396 XA.XIR[9].XIC[9].icell.SM VPWR 0.00158f
C6397 XA.XIR[2].XIC[2].icell.SM Vbias 0.00701f
C6398 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.SM 0.00168f
C6399 XA.XIR[10].XIC[3].icell.Ien VPWR 0.1903f
C6400 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Iout 0.00347f
C6401 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.15202f
C6402 XThR.Tn[2] XA.XIR[2].XIC[1].icell.PDM 0.00341f
C6403 XA.XIR[5].XIC_15.icell.PUM Vbias 0.0031f
C6404 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C6405 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00214f
C6406 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Ien 0.00232f
C6407 XA.XIR[9].XIC[5].icell.SM Iout 0.00388f
C6408 XA.XIR[12].XIC[13].icell.SM VPWR 0.00158f
C6409 XA.XIR[13].XIC[13].icell.PDM Vbias 0.04261f
C6410 XA.XIR[5].XIC[9].icell.PDM Vbias 0.04261f
C6411 XThC.Tn[9] XThR.Tn[11] 0.28739f
C6412 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04031f
C6413 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.SM 0.0039f
C6414 XA.XIR[0].XIC[1].icell.PDM Vbias 0.04282f
C6415 XThR.TB4 XThR.TB5 2.06459f
C6416 XThR.Tn[0] XA.XIR[1].XIC[10].icell.SM 0.00121f
C6417 XA.XIR[7].XIC[8].icell.PDM VPWR 0.00799f
C6418 XThC.Tn[13] XThR.Tn[3] 0.2874f
C6419 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00214f
C6420 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.03425f
C6421 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PUM 0.00429f
C6422 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04031f
C6423 XA.XIR[6].XIC[2].icell.PUM Vbias 0.0031f
C6424 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18966f
C6425 XA.XIR[8].XIC[11].icell.PDM Vbias 0.04261f
C6426 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C6427 XA.XIR[14].XIC[4].icell.Ien Vbias 0.21098f
C6428 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10] 0.00341f
C6429 XA.XIR[4].XIC[5].icell.Ien VPWR 0.1903f
C6430 XThR.TBN XThR.TA2 0.03867f
C6431 XA.XIR[2].XIC[9].icell.Ien VPWR 0.1903f
C6432 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14] 0.00341f
C6433 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C6434 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C6435 XA.XIR[13].XIC[6].icell.Ien Vbias 0.21098f
C6436 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C6437 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C6438 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Iout 0.00347f
C6439 XThR.Tn[14] XA.XIR[15].XIC[13].icell.SM 0.00121f
C6440 XA.XIR[7].XIC[5].icell.SM VPWR 0.00158f
C6441 XA.XIR[2].XIC[5].icell.Ien Iout 0.06417f
C6442 XA.XIR[8].XIC[8].icell.SM Vbias 0.00701f
C6443 XThC.Tn[8] XThR.Tn[6] 0.28739f
C6444 XA.XIR[11].XIC_15.icell.PUM Vbias 0.0031f
C6445 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00214f
C6446 XThR.TAN XThR.Tn[8] 0.05091f
C6447 XA.XIR[9].XIC[0].icell.PUM VPWR 0.00937f
C6448 XA.XIR[12].XIC[8].icell.PUM Vbias 0.0031f
C6449 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.SM 0.0039f
C6450 XA.XIR[7].XIC[1].icell.SM Iout 0.00388f
C6451 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C6452 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.15202f
C6453 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.03425f
C6454 XA.XIR[11].XIC[9].icell.Ien Vbias 0.21098f
C6455 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6456 XA.XIR[1].XIC[8].icell.PDM Vbias 0.04261f
C6457 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.PUM 0.00121f
C6458 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.SM 0.0039f
C6459 XThC.TAN a_6243_9615# 0.01743f
C6460 XThC.TB1 XThC.Tn[1] 0.01447f
C6461 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C6462 XA.XIR[3].XIC[4].icell.Ien Vbias 0.21098f
C6463 XThR.TBN XThR.Tn[0] 0.55717f
C6464 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02762f
C6465 XThR.Tn[7] XA.XIR[8].XIC[2].icell.SM 0.00121f
C6466 XA.XIR[8].XIC_15.icell.Ien VPWR 0.25566f
C6467 XA.XIR[12].XIC_15.icell.Ien Iout 0.0642f
C6468 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.SM 0.0039f
C6469 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C6470 XA.XIR[6].XIC[7].icell.PUM Vbias 0.0031f
C6471 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18987f
C6472 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02762f
C6473 XThC.TBN XThC.Tn[3] 0.62681f
C6474 XA.XIR[8].XIC[11].icell.Ien Iout 0.06417f
C6475 XThR.Tn[8] XA.XIR[9].XIC[11].icell.Ien 0.00338f
C6476 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.15202f
C6477 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C6478 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00584f
C6479 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.SM 0.0039f
C6480 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PUM 0.00465f
C6481 XThC.Tn[12] XThR.Tn[12] 0.28739f
C6482 XA.XIR[4].XIC[13].icell.Ien Vbias 0.21098f
C6483 XA.XIR[3].XIC[11].icell.PUM VPWR 0.00937f
C6484 XA.XIR[1].XIC_15.icell.PDM Iout 0.00133f
C6485 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Ien 0.00584f
C6486 XThR.Tn[10] XA.XIR[11].XIC[3].icell.SM 0.00121f
C6487 XA.XIR[6].XIC[12].icell.SM VPWR 0.00158f
C6488 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00214f
C6489 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C6490 XThR.Tn[0] XA.XIR[0].XIC[2].icell.PDM 0.00341f
C6491 XA.XIR[6].XIC[4].icell.PDM VPWR 0.00799f
C6492 XA.XIR[7].XIC[13].icell.SM Vbias 0.00701f
C6493 a_n997_3755# XThR.Tn[9] 0.19352f
C6494 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07214f
C6495 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02762f
C6496 XA.XIR[6].XIC[8].icell.SM Iout 0.00388f
C6497 XA.XIR[1].XIC[8].icell.PUM VPWR 0.00937f
C6498 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7] 0.00341f
C6499 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.SM 0.00168f
C6500 XA.XIR[11].XIC[10].icell.SM Vbias 0.00701f
C6501 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.15202f
C6502 XA.XIR[15].XIC[12].icell.Ien Iout 0.06807f
C6503 XA.XIR[4].XIC[3].icell.PDM Iout 0.00117f
C6504 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.15235f
C6505 XThR.Tn[13] XA.XIR[14].XIC[8].icell.Ien 0.00338f
C6506 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00584f
C6507 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6508 XThC.Tn[11] XThR.Tn[10] 0.28739f
C6509 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C6510 XA.XIR[13].XIC[0].icell.SM Vbias 0.00675f
C6511 XThR.TBN a_n1049_7493# 0.08456f
C6512 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.SM 0.00168f
C6513 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00584f
C6514 XThR.TB1 XThR.TA3 0.48957f
C6515 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C6516 XA.XIR[0].XIC[13].icell.Ien Vbias 0.2113f
C6517 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.03425f
C6518 XA.XIR[12].XIC[4].icell.PDM VPWR 0.00799f
C6519 XA.XIR[7].XIC_dummy_right.icell.SM VPWR 0.00123f
C6520 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04031f
C6521 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PUM 0.00465f
C6522 XA.XIR[3].XIC_15.icell.SM VPWR 0.00275f
C6523 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.SM 0.00168f
C6524 XA.XIR[12].XIC[11].icell.SM VPWR 0.00158f
C6525 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00214f
C6526 XThR.Tn[6] XA.XIR[7].XIC[10].icell.Ien 0.00338f
C6527 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C6528 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.SM 0.0039f
C6529 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04031f
C6530 XA.XIR[11].XIC[10].icell.PDM VPWR 0.00799f
C6531 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02762f
C6532 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Iout 0.00347f
C6533 XThR.Tn[4] XA.XIR[5].XIC[12].icell.SM 0.00121f
C6534 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04031f
C6535 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C6536 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[8].icell.SM 0.0039f
C6537 XA.XIR[15].XIC[3].icell.PUM Vbias 0.0031f
C6538 XA.XIR[5].XIC[5].icell.Ien Vbias 0.21098f
C6539 XA.XIR[14].XIC[1].icell.Ien Iout 0.06417f
C6540 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.SM 0.0039f
C6541 XThR.Tn[3] XA.XIR[4].XIC[14].icell.SM 0.00121f
C6542 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00584f
C6543 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.03425f
C6544 XA.XIR[8].XIC[0].icell.SM VPWR 0.00158f
C6545 XA.XIR[4].XIC_dummy_left.icell.SM VPWR 0.00269f
C6546 XThR.Tn[14] XA.XIR[15].XIC[11].icell.SM 0.00121f
C6547 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.SM 0.00168f
C6548 XA.XIR[14].XIC[11].icell.PDM VPWR 0.00799f
C6549 XA.XIR[10].XIC[2].icell.PDM Iout 0.00117f
C6550 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04031f
C6551 XA.XIR[11].XIC[13].icell.PUM Vbias 0.0031f
C6552 XA.XIR[1].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6553 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.03023f
C6554 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.SM 0.00168f
C6555 XA.XIR[5].XIC[12].icell.PUM VPWR 0.00937f
C6556 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C6557 XA.XIR[10].XIC[11].icell.PDM Vbias 0.04261f
C6558 XA.XIR[15].XIC[8].icell.SM VPWR 0.00158f
C6559 XA.XIR[5].XIC[0].icell.PDM VPWR 0.00799f
C6560 XA.XIR[3].XIC[12].icell.PDM VPWR 0.00799f
C6561 XThR.Tn[5] Vbias 3.74761f
C6562 XA.XIR[14].XIC[12].icell.SM Vbias 0.00701f
C6563 XA.XIR[15].XIC[4].icell.SM Iout 0.00388f
C6564 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.03425f
C6565 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C6566 XA.XIR[3].XIC[0].icell.PDM Iout 0.00117f
C6567 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.03425f
C6568 XA.XIR[8].XIC[2].icell.PDM VPWR 0.00799f
C6569 XA.XIR[9].XIC[11].icell.PDM Vbias 0.04261f
C6570 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00214f
C6571 XA.XIR[13].XIC[12].icell.PDM Vbias 0.04261f
C6572 a_n1049_6405# VPWR 0.72095f
C6573 XA.XIR[12].XIC[14].icell.PUM VPWR 0.00937f
C6574 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.03425f
C6575 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C6576 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.SM 0.0039f
C6577 XA.XIR[13].XIC[3].icell.Ien VPWR 0.1903f
C6578 XThC.TB4 a_7875_9569# 0.00497f
C6579 XA.XIR[0].XIC_dummy_left.icell.SM VPWR 0.00269f
C6580 XA.XIR[9].XIC[9].icell.PUM Vbias 0.0031f
C6581 XThR.Tn[2] XA.XIR[3].XIC[4].icell.Ien 0.00338f
C6582 XA.XIR[10].XIC[1].icell.SM Vbias 0.00701f
C6583 XA.XIR[8].XIC[5].icell.SM VPWR 0.00158f
C6584 XThR.TAN a_n997_3755# 0.01174f
C6585 XThC.Tn[9] XThR.Tn[14] 0.28739f
C6586 XThC.TB5 XThC.Tn[7] 0.00912f
C6587 XA.XIR[12].XIC[5].icell.PUM VPWR 0.00937f
C6588 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00584f
C6589 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12] 0.00341f
C6590 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00584f
C6591 XA.XIR[8].XIC[1].icell.SM Iout 0.00388f
C6592 XA.XIR[4].XIC[1].icell.Ien Iout 0.06417f
C6593 XThR.Tn[8] XA.XIR[9].XIC[1].icell.SM 0.00121f
C6594 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PUM 0.00465f
C6595 XThC.Tn[5] XThR.Tn[5] 0.28739f
C6596 XA.XIR[11].XIC[14].icell.Ien Vbias 0.21098f
C6597 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04031f
C6598 XA.XIR[7].XIC[4].icell.PDM Vbias 0.04261f
C6599 XA.XIR[11].XIC[6].icell.Ien VPWR 0.1903f
C6600 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38912f
C6601 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PUM 0.00465f
C6602 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.04036f
C6603 XA.XIR[4].XIC[3].icell.SM Vbias 0.00701f
C6604 XThR.TB7 XThR.Tn[12] 0.07066f
C6605 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.SM 0.0039f
C6606 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.0353f
C6607 XA.XIR[2].XIC[7].icell.SM Vbias 0.00701f
C6608 XA.XIR[11].XIC[2].icell.Ien Iout 0.06417f
C6609 XA.XIR[9].XIC[14].icell.SM VPWR 0.00207f
C6610 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.03425f
C6611 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.03591f
C6612 XA.XIR[10].XIC[8].icell.Ien VPWR 0.1903f
C6613 XA.XIR[15].XIC[10].icell.Ien Iout 0.06807f
C6614 XA.XIR[6].XIC[4].icell.PUM VPWR 0.00937f
C6615 XA.XIR[9].XIC[10].icell.SM Iout 0.00388f
C6616 XA.XIR[14].XIC_15.icell.PUM Vbias 0.0031f
C6617 XA.XIR[7].XIC[5].icell.PUM Vbias 0.0031f
C6618 XThC.Tn[10] XThR.Tn[4] 0.28739f
C6619 XA.XIR[10].XIC[4].icell.Ien Iout 0.06417f
C6620 XThR.Tn[9] XA.XIR[10].XIC[4].icell.Ien 0.00338f
C6621 XA.XIR[14].XIC[9].icell.Ien Vbias 0.21098f
C6622 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00584f
C6623 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02762f
C6624 XA.XIR[4].XIC[10].icell.Ien VPWR 0.1903f
C6625 XThC.TB2 data[1] 0.017f
C6626 data[5] data[4] 0.64735f
C6627 XA.XIR[7].XIC[11].icell.PDM Iout 0.00117f
C6628 XA.XIR[2].XIC[14].icell.Ien VPWR 0.19036f
C6629 XA.XIR[12].XIC[9].icell.SM VPWR 0.00158f
C6630 XA.XIR[0].XIC[1].icell.Ien Iout 0.06389f
C6631 XA.XIR[2].XIC[7].icell.PDM VPWR 0.00799f
C6632 XA.XIR[1].XIC[1].icell.Ien Vbias 0.21104f
C6633 XA.XIR[4].XIC[6].icell.Ien Iout 0.06417f
C6634 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8] 0.00341f
C6635 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.0404f
C6636 XA.XIR[7].XIC[10].icell.SM VPWR 0.00158f
C6637 XA.XIR[2].XIC[10].icell.Ien Iout 0.06417f
C6638 VPWR data[6] 0.21221f
C6639 XA.XIR[8].XIC[13].icell.SM Vbias 0.00701f
C6640 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00214f
C6641 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00214f
C6642 XA.XIR[0].XIC[3].icell.SM Vbias 0.00716f
C6643 XA.XIR[7].XIC[6].icell.SM Iout 0.00388f
C6644 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.SM 0.00168f
C6645 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C6646 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04031f
C6647 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.15202f
C6648 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PUM 0.00465f
C6649 XThC.Tn[2] XThR.Tn[3] 0.28739f
C6650 XThR.Tn[12] XA.XIR[13].XIC[2].icell.Ien 0.00338f
C6651 XThC.Tn[7] XThR.Tn[11] 0.28739f
C6652 XThC.Tn[12] XThR.Tn[0] 0.28786f
C6653 XThR.Tn[14] XA.XIR[15].XIC[9].icell.SM 0.00121f
C6654 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C6655 XA.XIR[3].XIC[9].icell.Ien Vbias 0.21098f
C6656 XA.XIR[11].XIC[11].icell.PUM Vbias 0.0031f
C6657 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.03425f
C6658 a_n1335_4229# VPWR 0.00633f
C6659 XThR.Tn[7] XA.XIR[8].XIC[7].icell.SM 0.00121f
C6660 XThC.Tn[5] Vbias 2.31635f
C6661 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C6662 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.SM 0.00168f
C6663 XA.XIR[6].XIC[0].icell.PDM Vbias 0.04207f
C6664 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18966f
C6665 XA.XIR[8].XIC_dummy_right.icell.SM VPWR 0.00123f
C6666 XA.XIR[6].XIC[12].icell.PUM Vbias 0.0031f
C6667 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C6668 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02762f
C6669 XThR.Tn[11] XA.XIR[12].XIC[5].icell.Ien 0.00338f
C6670 XA.XIR[4].XIC[11].icell.PDM Vbias 0.04261f
C6671 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.15202f
C6672 XA.XIR[0].XIC[6].icell.Ien Iout 0.06389f
C6673 XA.XIR[14].XIC[10].icell.SM Vbias 0.00701f
C6674 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PUM 0.00465f
C6675 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.03425f
C6676 XA.XIR[1].XIC[6].icell.Ien Vbias 0.21104f
C6677 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.SM 0.00168f
C6678 XThC.Tn[6] XThR.Tn[6] 0.28739f
C6679 XA.XIR[11].XIC[0].icell.SM VPWR 0.00158f
C6680 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6681 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00214f
C6682 XThC.TAN a_8963_9569# 0.02071f
C6683 XA.XIR[12].XIC[12].icell.PUM VPWR 0.00937f
C6684 XA.XIR[5].XIC[2].icell.Ien VPWR 0.1903f
C6685 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6686 XThC.Tn[11] XThR.Tn[13] 0.28739f
C6687 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C6688 a_9827_9569# XThC.Tn[12] 0.19481f
C6689 XThR.Tn[10] XA.XIR[11].XIC[8].icell.SM 0.00121f
C6690 XThC.TA2 a_5155_10571# 0.00306f
C6691 XThC.TA2 Vbias 0.00648f
C6692 XThC.Tn[0] XThC.Tn[1] 1.15401f
C6693 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.SM 0.0039f
C6694 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C6695 XThC.TA1 Vbias 0.00557f
C6696 XA.XIR[15].XIC[4].icell.PDM VPWR 0.0114f
C6697 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PUM 0.00465f
C6698 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C6699 XThC.Tn[4] XThC.Tn[6] 0.00202f
C6700 XA.XIR[12].XIC[0].icell.PDM Vbias 0.04207f
C6701 XA.XIR[6].XIC[13].icell.SM Iout 0.00388f
C6702 XA.XIR[6].XIC[7].icell.PDM Iout 0.00117f
C6703 XA.XIR[1].XIC[13].icell.PUM VPWR 0.00937f
C6704 XThC.Tn[14] Iout 0.84284f
C6705 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C6706 XThR.Tn[1] XA.XIR[1].XIC[3].icell.PDM 0.00341f
C6707 XA.XIR[14].XIC[10].icell.PDM VPWR 0.00799f
C6708 XThC.Tn[14] XThR.Tn[9] 0.28745f
C6709 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.SM 0.0039f
C6710 XThC.Tn[1] XThR.Tn[12] 0.28739f
C6711 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.SM 0.00168f
C6712 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02762f
C6713 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C6714 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PUM 0.00465f
C6715 XA.XIR[15].XIC[13].icell.SM VPWR 0.00158f
C6716 XA.XIR[11].XIC[6].icell.PDM Vbias 0.04261f
C6717 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01444f
C6718 XThC.Tn[10] XThR.Tn[8] 0.28739f
C6719 XA.XIR[11].XIC[12].icell.Ien Vbias 0.21098f
C6720 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.SM 0.0039f
C6721 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.15202f
C6722 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01432f
C6723 XA.XIR[10].XIC[10].icell.PDM Vbias 0.04261f
C6724 XA.XIR[9].XIC[2].icell.PDM VPWR 0.00799f
C6725 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6726 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.SM 0.00168f
C6727 XA.XIR[13].XIC[2].icell.PDM Iout 0.00117f
C6728 XA.XIR[14].XIC[13].icell.PUM Vbias 0.0031f
C6729 XThR.Tn[6] XA.XIR[7].XIC_15.icell.Ien 0.00117f
C6730 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.15202f
C6731 XThC.TA2 XThC.Tn[5] 0.00363f
C6732 XThR.Tn[5] XA.XIR[6].XIC[2].icell.Ien 0.00338f
C6733 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C6734 XA.XIR[12].XIC[7].icell.PDM Iout 0.00117f
C6735 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00256f
C6736 XThC.TB6 a_9827_9569# 0.00871f
C6737 XA.XIR[12].XIC[13].icell.Ien VPWR 0.1903f
C6738 XA.XIR[9].XIC[6].icell.PUM VPWR 0.00937f
C6739 XA.XIR[13].XIC[11].icell.PDM Vbias 0.04261f
C6740 a_10051_9569# Vbias 0.00827f
C6741 XThC.TB4 XThC.Tn[4] 0.00758f
C6742 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00584f
C6743 XA.XIR[5].XIC[10].icell.Ien Vbias 0.21098f
C6744 XA.XIR[15].XIC[8].icell.PUM Vbias 0.0031f
C6745 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04031f
C6746 XA.XIR[3].XIC[8].icell.PDM Vbias 0.04261f
C6747 XThC.Tn[0] XThR.Tn[10] 0.28736f
C6748 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C6749 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02762f
C6750 XThC.Tn[10] XThR.Tn[1] 0.28739f
C6751 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.03425f
C6752 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.SM 0.0039f
C6753 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.0353f
C6754 XThR.TA2 XThR.TB7 0.01596f
C6755 XThR.Tn[14] XA.XIR[15].XIC[13].icell.Ien 0.00338f
C6756 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C6757 XThR.Tn[2] Vbias 3.74868f
C6758 XA.XIR[2].XIC[4].icell.SM VPWR 0.00158f
C6759 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02762f
C6760 XThR.Tn[10] XThR.Tn[12] 0.00142f
C6761 XA.XIR[10].XIC[12].icell.SM Iout 0.00388f
C6762 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.SM 0.00168f
C6763 XThC.TA1 XThC.TA2 1.80461f
C6764 XA.XIR[13].XIC[1].icell.SM Vbias 0.00701f
C6765 XA.XIR[15].XIC_15.icell.Ien Iout 0.0681f
C6766 a_n1049_7787# VPWR 0.72173f
C6767 XThR.Tn[9] XA.XIR[10].XIC[12].icell.SM 0.00121f
C6768 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07214f
C6769 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.SM 0.00168f
C6770 XA.XIR[8].XIC[5].icell.PUM Vbias 0.0031f
C6771 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.03425f
C6772 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C6773 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.PDM 0.00591f
C6774 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04031f
C6775 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.SM 0.0039f
C6776 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00584f
C6777 XA.XIR[0].XIC[7].icell.PDM VPWR 0.00773f
C6778 XA.XIR[12].XIC[3].icell.Ien Vbias 0.21098f
C6779 XA.XIR[5].XIC[3].icell.PDM Iout 0.00117f
C6780 XA.XIR[3].XIC_15.icell.PDM Iout 0.00133f
C6781 XA.XIR[14].XIC[14].icell.Ien Vbias 0.21098f
C6782 XA.XIR[14].XIC[6].icell.Ien VPWR 0.19084f
C6783 XThC.TB2 XThC.Tn[10] 0.00106f
C6784 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00584f
C6785 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PUM 0.00465f
C6786 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13] 0.00341f
C6787 XA.XIR[11].XIC[4].icell.SM Vbias 0.00701f
C6788 XThR.TBN a_n1049_5611# 0.0768f
C6789 XA.XIR[12].XIC[14].icell.SM VPWR 0.00207f
C6790 XA.XIR[8].XIC[5].icell.PDM Iout 0.00117f
C6791 XA.XIR[14].XIC[2].icell.Ien Iout 0.06417f
C6792 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.03425f
C6793 XThC.TB3 XThC.Tn[9] 0.00285f
C6794 XA.XIR[13].XIC[8].icell.Ien VPWR 0.1903f
C6795 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04031f
C6796 XA.XIR[8].XIC[10].icell.SM VPWR 0.00158f
C6797 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02762f
C6798 XA.XIR[9].XIC[14].icell.PUM Vbias 0.0031f
C6799 XThC.TB2 a_4861_9615# 0.00851f
C6800 XA.XIR[10].XIC[6].icell.SM Vbias 0.00701f
C6801 XThR.TA3 data[5] 0.06538f
C6802 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C6803 XThR.Tn[2] XA.XIR[3].XIC[9].icell.Ien 0.00338f
C6804 XThC.TB3 XThC.TBN 0.17246f
C6805 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00584f
C6806 XA.XIR[13].XIC[4].icell.Ien Iout 0.06417f
C6807 XThC.TAN2 Vbias 0.01776f
C6808 XThC.Tn[5] XThR.Tn[2] 0.28739f
C6809 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.SM 0.00168f
C6810 XA.XIR[6].XIC[2].icell.Ien Vbias 0.21098f
C6811 XA.XIR[12].XIC[10].icell.PUM VPWR 0.00937f
C6812 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02762f
C6813 XA.XIR[8].XIC[6].icell.SM Iout 0.00388f
C6814 XThR.Tn[4] XA.XIR[4].XIC[6].icell.PDM 0.00341f
C6815 XThR.TB3 VPWR 1.07975f
C6816 XThR.Tn[8] XA.XIR[9].XIC[6].icell.SM 0.00121f
C6817 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PUM 0.00465f
C6818 XThR.Tn[3] XA.XIR[3].XIC[13].icell.PDM 0.00341f
C6819 XA.XIR[1].XIC[14].icell.PDM VPWR 0.00809f
C6820 XThR.Tn[14] XA.XIR[15].XIC[14].icell.SM 0.00121f
C6821 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PDM 0.00172f
C6822 XA.XIR[4].XIC[8].icell.SM Vbias 0.00701f
C6823 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.SM 0.00168f
C6824 XThR.Tn[6] XA.XIR[7].XIC[0].icell.SM 0.00121f
C6825 XA.XIR[3].XIC[6].icell.Ien VPWR 0.1903f
C6826 XThR.Tn[3] XThR.Tn[4] 0.06967f
C6827 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PUM 0.00186f
C6828 XA.XIR[1].XIC[2].icell.PDM Iout 0.00117f
C6829 XA.XIR[11].XIC[7].icell.Ien Iout 0.06417f
C6830 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C6831 XA.XIR[9].XIC[1].icell.PUM VPWR 0.00937f
C6832 XA.XIR[2].XIC[12].icell.SM Vbias 0.00701f
C6833 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PUM 0.00465f
C6834 XA.XIR[2].XIC[3].icell.PDM Vbias 0.04261f
C6835 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.SM 0.0039f
C6836 XA.XIR[3].XIC[2].icell.Ien Iout 0.06417f
C6837 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00584f
C6838 XA.XIR[6].XIC[9].icell.PUM VPWR 0.00937f
C6839 XA.XIR[15].XIC[11].icell.SM VPWR 0.00158f
C6840 XA.XIR[7].XIC[10].icell.PUM Vbias 0.0031f
C6841 XThR.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.00338f
C6842 XA.XIR[10].XIC[9].icell.Ien Iout 0.06417f
C6843 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00584f
C6844 XA.XIR[11].XIC[10].icell.Ien Vbias 0.21098f
C6845 XA.XIR[4].XIC[2].icell.PDM VPWR 0.00799f
C6846 XThR.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.00338f
C6847 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.SM 0.0039f
C6848 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02762f
C6849 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00214f
C6850 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7] 0.00341f
C6851 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PUM 0.00465f
C6852 XThC.TB7 XThC.Tn[9] 0.07413f
C6853 XA.XIR[1].XIC[3].icell.Ien VPWR 0.1903f
C6854 XThC.Tn[7] XThR.Tn[14] 0.28739f
C6855 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6856 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C6857 XA.XIR[4].XIC_15.icell.Ien VPWR 0.25566f
C6858 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.SM 0.00168f
C6859 XThC.TB7 XThC.TBN 0.50018f
C6860 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02762f
C6861 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04031f
C6862 XA.XIR[14].XIC[11].icell.PUM Vbias 0.0031f
C6863 XA.XIR[4].XIC[11].icell.Ien Iout 0.06417f
C6864 XThR.Tn[13] XA.XIR[14].XIC[3].icell.SM 0.00121f
C6865 XThR.Tn[10] XA.XIR[11].XIC[13].icell.SM 0.00121f
C6866 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.SM 0.00168f
C6867 XThR.TB4 XThR.Tn[5] 0.00751f
C6868 XThR.TAN data[4] 0.01382f
C6869 XA.XIR[2].XIC_15.icell.Ien Iout 0.0642f
C6870 XA.XIR[12].XIC[11].icell.Ien VPWR 0.1903f
C6871 XA.XIR[2].XIC[10].icell.PDM Iout 0.00117f
C6872 XA.XIR[0].XIC[8].icell.SM Vbias 0.00716f
C6873 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.SM 0.00168f
C6874 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.SM 0.0039f
C6875 a_6243_9615# XThC.Tn[6] 0.26142f
C6876 XThR.Tn[6] XA.XIR[7].XIC[5].icell.SM 0.00121f
C6877 XA.XIR[7].XIC[11].icell.SM Iout 0.00388f
C6878 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.15202f
C6879 XA.XIR[1].XIC[0].icell.PUM VPWR 0.00937f
C6880 XThC.TA2 XThC.TAN2 0.0513f
C6881 XA.XIR[14].XIC[0].icell.SM VPWR 0.00158f
C6882 XThC.TA1 XThC.TAN2 0.06305f
C6883 XThR.Tn[12] XA.XIR[13].XIC[7].icell.Ien 0.00338f
C6884 XA.XIR[11].XIC[0].icell.Ien Vbias 0.20951f
C6885 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C6886 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.SM 0.0039f
C6887 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00584f
C6888 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PDM 0.00172f
C6889 XA.XIR[3].XIC[14].icell.Ien Vbias 0.21098f
C6890 XThR.Tn[1] XA.XIR[2].XIC[6].icell.Ien 0.00338f
C6891 XThC.Tn[9] VPWR 6.83084f
C6892 XThR.Tn[14] XA.XIR[15].XIC[11].icell.Ien 0.00338f
C6893 XA.XIR[10].XIC[1].icell.PDM VPWR 0.00799f
C6894 XThR.Tn[7] XA.XIR[8].XIC[12].icell.SM 0.00121f
C6895 XThR.TA3 a_n1049_6699# 0.02294f
C6896 XA.XIR[10].XIC[2].icell.PUM Vbias 0.0031f
C6897 XThR.TA1 a_n1335_4229# 0.01243f
C6898 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.SM 0.0039f
C6899 XA.XIR[15].XIC[14].icell.PUM VPWR 0.00937f
C6900 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04031f
C6901 XA.XIR[10].XIC[10].icell.SM Iout 0.00388f
C6902 XThR.Tn[9] XA.XIR[10].XIC[10].icell.SM 0.00121f
C6903 XThC.TBN VPWR 4.08849f
C6904 XA.XIR[6].XIC_15.icell.PDM Vbias 0.04401f
C6905 XA.XIR[0].XIC_15.icell.Ien VPWR 0.2554f
C6906 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C6907 XA.XIR[15].XIC[0].icell.PDM Vbias 0.04207f
C6908 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5] 0.00341f
C6909 XThR.Tn[12] a_n997_1803# 0.18719f
C6910 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.SM 0.00168f
C6911 XA.XIR[0].XIC[11].icell.Ien Iout 0.06389f
C6912 XA.XIR[1].XIC[11].icell.Ien Vbias 0.21104f
C6913 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PUM 0.00465f
C6914 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6915 XA.XIR[12].XIC[0].icell.Ien Iout 0.06411f
C6916 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00214f
C6917 XA.XIR[14].XIC[6].icell.PDM Vbias 0.04261f
C6918 XThC.TB4 a_6243_9615# 0.00463f
C6919 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.02762f
C6920 XA.XIR[5].XIC[7].icell.Ien VPWR 0.1903f
C6921 XA.XIR[14].XIC[12].icell.Ien Vbias 0.21098f
C6922 XThC.Tn[1] XThR.Tn[0] 0.28784f
C6923 XA.XIR[15].XIC[5].icell.PUM VPWR 0.00937f
C6924 XThR.Tn[11] Iout 1.16235f
C6925 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C6926 XThR.Tn[9] XThR.Tn[11] 0.00252f
C6927 XA.XIR[13].XIC[10].icell.PDM Vbias 0.04261f
C6928 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00214f
C6929 XThR.TB2 a_n1049_6405# 0.00847f
C6930 XA.XIR[5].XIC[3].icell.Ien Iout 0.06417f
C6931 XThC.TAN2 a_10051_9569# 0.00199f
C6932 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.SM 0.0039f
C6933 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00584f
C6934 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6] 0.00341f
C6935 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C6936 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C6937 XA.XIR[15].XIC[7].icell.PDM Iout 0.00117f
C6938 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02762f
C6939 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.03425f
C6940 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PUM 0.00102f
C6941 XA.XIR[9].XIC[4].icell.Ien Vbias 0.21098f
C6942 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.03425f
C6943 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.03425f
C6944 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.03425f
C6945 XA.XIR[4].XIC[0].icell.SM VPWR 0.00158f
C6946 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00214f
C6947 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.15202f
C6948 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02762f
C6949 XThC.Tn[0] XThR.Tn[13] 0.28746f
C6950 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C6951 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02762f
C6952 XA.XIR[7].XIC[2].icell.PUM VPWR 0.00937f
C6953 XA.XIR[2].XIC[0].icell.SM Iout 0.00388f
C6954 XThR.TAN a_n997_2667# 0.02071f
C6955 XThC.TBN a_5155_9615# 0.07602f
C6956 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C6957 XA.XIR[11].XIC[1].icell.SM VPWR 0.00158f
C6958 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00214f
C6959 XA.XIR[15].XIC[9].icell.SM VPWR 0.00158f
C6960 XThR.Tn[5] XA.XIR[6].XIC[7].icell.Ien 0.00338f
C6961 XA.XIR[9].XIC[5].icell.PDM Iout 0.00117f
C6962 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.15202f
C6963 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9] 0.00341f
C6964 XThR.Tn[12] XThR.Tn[13] 0.06297f
C6965 XA.XIR[13].XIC[12].icell.SM Iout 0.00388f
C6966 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.SM 0.0039f
C6967 XA.XIR[9].XIC[11].icell.PUM VPWR 0.00937f
C6968 XThC.Tn[3] Iout 0.8384f
C6969 XA.XIR[10].XIC[3].icell.SM VPWR 0.00158f
C6970 XThR.TBN XA.XIR[11].XIC_dummy_left.icell.Ien 0.0016f
C6971 XA.XIR[2].XIC[4].icell.PUM Vbias 0.0031f
C6972 XThC.Tn[3] XThR.Tn[9] 0.28739f
C6973 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C6974 XA.XIR[5].XIC_15.icell.Ien Vbias 0.21234f
C6975 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[13].icell.SM 0.0039f
C6976 XThC.Tn[12] data[3] 0.00161f
C6977 XThR.Tn[2] XA.XIR[2].XIC[3].icell.PDM 0.00341f
C6978 XA.XIR[5].XIC[11].icell.PDM Vbias 0.04261f
C6979 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00214f
C6980 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.SM 0.0039f
C6981 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04031f
C6982 XA.XIR[0].XIC[3].icell.PDM Vbias 0.04278f
C6983 XThR.Tn[10] XA.XIR[11].XIC[11].icell.SM 0.00121f
C6984 XA.XIR[7].XIC[10].icell.PDM VPWR 0.00799f
C6985 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.03579f
C6986 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04031f
C6987 XA.XIR[0].XIC[0].icell.SM VPWR 0.00158f
C6988 XThR.TB1 VPWR 1.12978f
C6989 XA.XIR[8].XIC[13].icell.PDM Vbias 0.04261f
C6990 XA.XIR[14].XIC[4].icell.SM Vbias 0.00701f
C6991 XA.XIR[4].XIC[5].icell.SM VPWR 0.00158f
C6992 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00584f
C6993 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10] 0.00341f
C6994 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02762f
C6995 XA.XIR[2].XIC[9].icell.SM VPWR 0.00158f
C6996 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02762f
C6997 XA.XIR[13].XIC[6].icell.SM Vbias 0.00701f
C6998 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.SM 0.00168f
C6999 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.SM 0.00168f
C7000 XA.XIR[4].XIC[1].icell.SM Iout 0.00388f
C7001 XA.XIR[7].XIC[7].icell.PUM VPWR 0.00937f
C7002 XA.XIR[2].XIC[5].icell.SM Iout 0.00388f
C7003 XA.XIR[8].XIC[10].icell.PUM Vbias 0.0031f
C7004 VPWR data[2] 0.21031f
C7005 XA.XIR[11].XIC_15.icell.PDM Vbias 0.04401f
C7006 XA.XIR[10].XIC[14].icell.Ien Iout 0.06417f
C7007 XThR.Tn[9] XA.XIR[10].XIC[14].icell.Ien 0.00338f
C7008 XA.XIR[11].XIC_15.icell.Ien Vbias 0.21234f
C7009 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.SM 0.0039f
C7010 XA.XIR[12].XIC[8].icell.Ien Vbias 0.21098f
C7011 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.03023f
C7012 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00214f
C7013 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.SM 0.00168f
C7014 XA.XIR[9].XIC_15.icell.SM VPWR 0.00275f
C7015 XA.XIR[15].XIC[12].icell.PUM VPWR 0.00937f
C7016 XA.XIR[1].XIC[10].icell.PDM Vbias 0.04261f
C7017 XA.XIR[14].XIC[7].icell.Ien Iout 0.06417f
C7018 XThR.TAN XThR.Tn[11] 0.03888f
C7019 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.SM 0.00168f
C7020 XA.XIR[3].XIC[4].icell.SM Vbias 0.00701f
C7021 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PUM 0.00465f
C7022 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0404f
C7023 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.SM 0.0039f
C7024 XThR.Tn[2] XA.XIR[3].XIC[14].icell.Ien 0.00338f
C7025 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02762f
C7026 XA.XIR[13].XIC[9].icell.Ien Iout 0.06417f
C7027 XA.XIR[6].XIC[7].icell.Ien Vbias 0.21098f
C7028 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00214f
C7029 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PUM 0.00465f
C7030 XA.XIR[0].XIC[5].icell.SM VPWR 0.00158f
C7031 XA.XIR[14].XIC[10].icell.Ien Vbias 0.21098f
C7032 XThR.TA1 XThR.TB3 0.01152f
C7033 XA.XIR[8].XIC[11].icell.SM Iout 0.00388f
C7034 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02762f
C7035 XThR.TAN XThR.TA3 0.35833f
C7036 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PUM 0.00465f
C7037 XThR.TBN XThR.TB7 0.50018f
C7038 XThR.Tn[8] XA.XIR[9].XIC[11].icell.SM 0.00121f
C7039 XA.XIR[0].XIC[1].icell.SM Iout 0.00367f
C7040 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.03425f
C7041 XA.XIR[1].XIC[1].icell.SM Vbias 0.00704f
C7042 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.SM 0.0039f
C7043 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02762f
C7044 XA.XIR[4].XIC[13].icell.SM Vbias 0.00701f
C7045 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.SM 0.0039f
C7046 XA.XIR[3].XIC[11].icell.Ien VPWR 0.1903f
C7047 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39036f
C7048 XThC.TB2 a_7651_9569# 0.00191f
C7049 XThR.TB6 a_n1049_5317# 0.01199f
C7050 XThR.Tn[0] XA.XIR[0].XIC[4].icell.PDM 0.00341f
C7051 XA.XIR[6].XIC[14].icell.PUM VPWR 0.00937f
C7052 XA.XIR[3].XIC[7].icell.Ien Iout 0.06417f
C7053 XA.XIR[6].XIC[6].icell.PDM VPWR 0.00799f
C7054 XA.XIR[7].XIC_15.icell.PUM Vbias 0.0031f
C7055 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04052f
C7056 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PUM 0.00465f
C7057 XThC.TB3 XThC.Tn[7] 0.00819f
C7058 XA.XIR[5].XIC[0].icell.SM Vbias 0.00675f
C7059 XThR.TB2 a_n1335_8107# 0.01006f
C7060 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.SM 0.00168f
C7061 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C7062 XA.XIR[15].XIC[13].icell.Ien VPWR 0.32895f
C7063 XA.XIR[1].XIC[8].icell.Ien VPWR 0.1903f
C7064 XThC.Tn[11] XThR.Tn[7] 0.28739f
C7065 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00584f
C7066 XThR.Tn[2] XThR.TB4 0.0021f
C7067 XA.XIR[4].XIC[5].icell.PDM Iout 0.00117f
C7068 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.SM 0.0039f
C7069 XA.XIR[1].XIC[4].icell.Ien Iout 0.06417f
C7070 XThR.Tn[13] XA.XIR[14].XIC[8].icell.SM 0.00121f
C7071 XA.XIR[4].XIC_dummy_right.icell.SM VPWR 0.00123f
C7072 XA.XIR[13].XIC[1].icell.PDM VPWR 0.00799f
C7073 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C7074 XA.XIR[13].XIC[2].icell.PUM Vbias 0.0031f
C7075 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.SM 0.0039f
C7076 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.SM 0.0039f
C7077 XA.XIR[13].XIC[10].icell.SM Iout 0.00388f
C7078 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PUM 0.00465f
C7079 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00214f
C7080 XA.XIR[0].XIC[13].icell.SM Vbias 0.00716f
C7081 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PUM 0.00465f
C7082 XA.XIR[12].XIC[6].icell.PDM VPWR 0.00799f
C7083 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04031f
C7084 XThR.Tn[6] XA.XIR[7].XIC[10].icell.SM 0.00121f
C7085 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.03425f
C7086 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C7087 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PUM 0.00465f
C7088 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.SM 0.00168f
C7089 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02762f
C7090 XThR.Tn[10] XA.XIR[11].XIC[9].icell.SM 0.00121f
C7091 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04031f
C7092 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00214f
C7093 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C7094 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04031f
C7095 XThR.Tn[14] Iout 1.16234f
C7096 XThC.TB7 XThC.Tn[7] 0.0835f
C7097 XThR.Tn[1] XA.XIR[2].XIC[11].icell.Ien 0.00338f
C7098 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00584f
C7099 XA.XIR[5].XIC[5].icell.SM Vbias 0.00701f
C7100 XA.XIR[15].XIC[3].icell.Ien Vbias 0.17899f
C7101 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Ien 0.00584f
C7102 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.SM 0.00168f
C7103 XThC.Tn[11] XThC.Tn[13] 0.00226f
C7104 XA.XIR[11].XIC[0].icell.PDM Iout 0.00117f
C7105 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00214f
C7106 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Ien 0.00549f
C7107 XA.XIR[8].XIC[2].icell.PUM VPWR 0.00937f
C7108 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C7109 XThR.Tn[0] XA.XIR[1].XIC[2].icell.Ien 0.00338f
C7110 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PUM 0.00465f
C7111 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02762f
C7112 XA.XIR[10].XIC[4].icell.PDM Iout 0.00117f
C7113 XA.XIR[10].XIC[12].icell.Ien Iout 0.06417f
C7114 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04031f
C7115 XA.XIR[15].XIC[14].icell.SM VPWR 0.00207f
C7116 XA.XIR[0].XIC_dummy_right.icell.SM VPWR 0.00123f
C7117 XThR.Tn[9] XA.XIR[10].XIC[12].icell.Ien 0.00338f
C7118 XThR.TB2 a_n1049_7787# 0.2342f
C7119 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C7120 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02771f
C7121 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02762f
C7122 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.1106f
C7123 XA.XIR[5].XIC[12].icell.Ien VPWR 0.1903f
C7124 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.SM 0.00168f
C7125 XA.XIR[5].XIC[2].icell.PDM VPWR 0.00799f
C7126 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PUM 0.00465f
C7127 XA.XIR[15].XIC[10].icell.PUM VPWR 0.00937f
C7128 XA.XIR[3].XIC[14].icell.PDM VPWR 0.00809f
C7129 XA.XIR[5].XIC[8].icell.Ien Iout 0.06417f
C7130 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C7131 XThC.TB3 a_3773_9615# 0.00124f
C7132 XA.XIR[9].XIC[13].icell.PDM Vbias 0.04261f
C7133 XA.XIR[3].XIC[2].icell.PDM Iout 0.00117f
C7134 XA.XIR[8].XIC[4].icell.PDM VPWR 0.00799f
C7135 XThR.Tn[14] XA.XIR[15].XIC[0].icell.Ien 0.00377f
C7136 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.SM 0.00168f
C7137 XA.XIR[7].XIC[0].icell.Ien Vbias 0.20951f
C7138 XThC.Tn[7] VPWR 6.29093f
C7139 XA.XIR[14].XIC[1].icell.SM VPWR 0.00158f
C7140 a_n1049_5611# XThR.TB7 0.00153f
C7141 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.15202f
C7142 XThC.TAN Vbias 0.09241f
C7143 XThC.TB4 a_8963_9569# 0.07199f
C7144 XA.XIR[13].XIC[3].icell.SM VPWR 0.00158f
C7145 XThC.TB6 XThC.Tn[12] 0.02863f
C7146 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00214f
C7147 XThR.Tn[2] XA.XIR[3].XIC[4].icell.SM 0.00121f
C7148 XA.XIR[9].XIC[9].icell.Ien Vbias 0.21098f
C7149 XA.XIR[8].XIC[7].icell.PUM VPWR 0.00937f
C7150 XA.XIR[10].XIC[3].icell.PUM Vbias 0.0031f
C7151 XThR.TB2 XThR.TB3 2.04808f
C7152 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.15202f
C7153 XA.XIR[12].XIC[5].icell.Ien VPWR 0.1903f
C7154 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12] 0.00341f
C7155 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.0353f
C7156 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.03425f
C7157 XThR.Tn[3] XA.XIR[3].XIC[0].icell.PDM 0.00347f
C7158 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C7159 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PUM 0.00465f
C7160 XA.XIR[11].XIC[14].icell.PDM Vbias 0.04261f
C7161 XA.XIR[7].XIC[6].icell.PDM Vbias 0.04261f
C7162 XA.XIR[11].XIC[6].icell.SM VPWR 0.00158f
C7163 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04031f
C7164 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02762f
C7165 XA.XIR[1].XIC[1].icell.PDM VPWR 0.00799f
C7166 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.03425f
C7167 XThR.Tn[5] XA.XIR[6].XIC[12].icell.Ien 0.00338f
C7168 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.15202f
C7169 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C7170 XA.XIR[4].XIC[5].icell.PUM Vbias 0.0031f
C7171 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04031f
C7172 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7173 XA.XIR[3].XIC[1].icell.SM VPWR 0.00158f
C7174 XA.XIR[10].XIC[8].icell.SM VPWR 0.00158f
C7175 XA.XIR[11].XIC[2].icell.SM Iout 0.00388f
C7176 XA.XIR[2].XIC[9].icell.PUM Vbias 0.0031f
C7177 XA.XIR[15].XIC[11].icell.Ien VPWR 0.32895f
C7178 XThC.TAN XThC.Tn[5] 0.00714f
C7179 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PUM 0.00465f
C7180 XA.XIR[13].XIC[14].icell.Ien Iout 0.06417f
C7181 XA.XIR[14].XIC_15.icell.PDM Vbias 0.04401f
C7182 XA.XIR[6].XIC[4].icell.Ien VPWR 0.1903f
C7183 XThR.Tn[14] XA.XIR[15].XIC[5].icell.Ien 0.00338f
C7184 XA.XIR[7].XIC[5].icell.Ien Vbias 0.21098f
C7185 XA.XIR[14].XIC_15.icell.Ien Vbias 0.21234f
C7186 XA.XIR[10].XIC[4].icell.SM Iout 0.00388f
C7187 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[2].icell.Ien 0.00214f
C7188 XThR.Tn[9] XA.XIR[10].XIC[4].icell.SM 0.00121f
C7189 a_7875_9569# XThC.Tn[9] 0.19329f
C7190 XThR.Tn[3] XA.XIR[4].XIC[1].icell.Ien 0.00338f
C7191 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00214f
C7192 XA.XIR[12].XIC_15.icell.SM VPWR 0.00275f
C7193 XThR.TBN XThR.Tn[10] 0.46535f
C7194 XThC.TBN a_7875_9569# 0.229f
C7195 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02762f
C7196 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00214f
C7197 XThR.Tn[10] XA.XIR[11].XIC[13].icell.Ien 0.00338f
C7198 XA.XIR[4].XIC[10].icell.SM VPWR 0.00158f
C7199 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00214f
C7200 XThR.TA1 XThR.TB1 0.1098f
C7201 XA.XIR[2].XIC[14].icell.SM VPWR 0.00207f
C7202 XA.XIR[7].XIC[13].icell.PDM Iout 0.00117f
C7203 XA.XIR[2].XIC[9].icell.PDM VPWR 0.00799f
C7204 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.0353f
C7205 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C7206 XA.XIR[4].XIC[6].icell.SM Iout 0.00388f
C7207 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8] 0.00341f
C7208 XA.XIR[8].XIC_15.icell.PUM Vbias 0.0031f
C7209 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C7210 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02762f
C7211 XThC.TA2 XThC.TAN 1.47641f
C7212 XA.XIR[7].XIC[12].icell.PUM VPWR 0.00937f
C7213 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PUM 0.00465f
C7214 XA.XIR[2].XIC[10].icell.SM Iout 0.00388f
C7215 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7216 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00214f
C7217 XThC.TA1 XThC.TAN 0.30355f
C7218 XA.XIR[0].XIC[5].icell.PUM Vbias 0.0031f
C7219 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C7220 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04031f
C7221 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.03425f
C7222 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.04036f
C7223 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.SM 0.00168f
C7224 XThR.Tn[12] XA.XIR[13].XIC[2].icell.SM 0.00121f
C7225 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C7226 a_3773_9615# VPWR 0.70508f
C7227 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C7228 XThR.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.00338f
C7229 XA.XIR[10].XIC[10].icell.Ien Iout 0.06417f
C7230 XA.XIR[3].XIC[9].icell.SM Vbias 0.00701f
C7231 XThR.Tn[13] XA.XIR[14].XIC[13].icell.SM 0.00121f
C7232 XThC.TB5 XThC.Tn[10] 0.01742f
C7233 XThR.Tn[1] XA.XIR[2].XIC[1].icell.SM 0.00121f
C7234 XThR.Tn[9] XA.XIR[10].XIC[10].icell.Ien 0.00338f
C7235 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PUM 0.00465f
C7236 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.15202f
C7237 XThR.Tn[3] XA.XIR[4].XIC[6].icell.Ien 0.00338f
C7238 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C7239 XThR.TB3 XThR.TAN2 0.03907f
C7240 XA.XIR[0].XIC[10].icell.SM VPWR 0.00158f
C7241 XA.XIR[6].XIC[12].icell.Ien Vbias 0.21098f
C7242 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C7243 XA.XIR[6].XIC[2].icell.PDM Vbias 0.04261f
C7244 XThC.Tn[8] XThR.Tn[5] 0.28739f
C7245 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C7246 XThR.Tn[11] XA.XIR[12].XIC[5].icell.SM 0.00121f
C7247 XThC.TB5 a_4861_9615# 0.0021f
C7248 XA.XIR[4].XIC[13].icell.PDM Vbias 0.04261f
C7249 XA.XIR[0].XIC[6].icell.SM Iout 0.00367f
C7250 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C7251 XA.XIR[11].XIC[2].icell.PUM VPWR 0.00937f
C7252 XA.XIR[1].XIC[6].icell.SM Vbias 0.00704f
C7253 XThR.Tn[10] XA.XIR[11].XIC[14].icell.SM 0.00121f
C7254 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02762f
C7255 XThR.TB3 XThR.Tn[6] 0.00298f
C7256 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C7257 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PUM 0.00429f
C7258 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.SM 0.00168f
C7259 XThC.TAN a_10051_9569# 0.00209f
C7260 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PDM 0.00172f
C7261 XA.XIR[5].XIC[2].icell.SM VPWR 0.00158f
C7262 XThC.TA3 a_6243_10571# 0.0017f
C7263 XA.XIR[9].XIC[1].icell.Ien VPWR 0.1903f
C7264 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.SM 0.0039f
C7265 XA.XIR[3].XIC[12].icell.Ien Iout 0.06417f
C7266 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.SM 0.0039f
C7267 XA.XIR[1].XIC[1].icell.PUM VPWR 0.00937f
C7268 VPWR data[5] 0.4402f
C7269 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02762f
C7270 XA.XIR[15].XIC[6].icell.PDM VPWR 0.0114f
C7271 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.SM 0.00168f
C7272 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.03425f
C7273 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PUM 0.00465f
C7274 XA.XIR[6].XIC[9].icell.PDM Iout 0.00117f
C7275 XA.XIR[12].XIC[2].icell.PDM Vbias 0.04261f
C7276 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PUM 0.00179f
C7277 XA.XIR[1].XIC[13].icell.Ien VPWR 0.1903f
C7278 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C7279 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C7280 XThR.Tn[1] XA.XIR[1].XIC[5].icell.PDM 0.00341f
C7281 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00214f
C7282 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.SM 0.00168f
C7283 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.03425f
C7284 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C7285 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C7286 XA.XIR[11].XIC[8].icell.PDM Vbias 0.04261f
C7287 XA.XIR[1].XIC[9].icell.Ien Iout 0.06417f
C7288 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.SM 0.0039f
C7289 XA.XIR[14].XIC[0].icell.PDM Iout 0.00117f
C7290 XA.XIR[9].XIC[4].icell.PDM VPWR 0.00799f
C7291 XA.XIR[13].XIC[4].icell.PDM Iout 0.00117f
C7292 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C7293 XA.XIR[13].XIC[12].icell.Ien Iout 0.06417f
C7294 XThC.Tn[10] XThR.Tn[11] 0.28739f
C7295 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00214f
C7296 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PUM 0.00102f
C7297 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.SM 0.0039f
C7298 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02762f
C7299 XThR.Tn[5] XA.XIR[6].XIC[2].icell.SM 0.00121f
C7300 XThC.Tn[14] XThR.Tn[3] 0.28745f
C7301 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PUM 0.00465f
C7302 XThC.Tn[0] XThR.Tn[7] 0.2874f
C7303 XA.XIR[9].XIC[6].icell.Ien VPWR 0.1903f
C7304 XA.XIR[12].XIC[9].icell.PDM Iout 0.00117f
C7305 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PUM 0.00465f
C7306 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.1106f
C7307 XThC.Tn[8] Vbias 2.30271f
C7308 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.03425f
C7309 XA.XIR[5].XIC[10].icell.SM Vbias 0.00701f
C7310 XThC.TAN2 XThC.TAN 0.35142f
C7311 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.04036f
C7312 XThR.Tn[10] XA.XIR[11].XIC[11].icell.Ien 0.00338f
C7313 XA.XIR[15].XIC[8].icell.Ien Vbias 0.17899f
C7314 XThR.TBN a_n997_1803# 0.22873f
C7315 XA.XIR[9].XIC[2].icell.Ien Iout 0.06417f
C7316 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.15202f
C7317 XA.XIR[3].XIC[10].icell.PDM Vbias 0.04261f
C7318 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.SM 0.00168f
C7319 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00214f
C7320 XThC.Tn[9] XThR.Tn[6] 0.28739f
C7321 XThR.Tn[0] XA.XIR[1].XIC[7].icell.Ien 0.00338f
C7322 XThR.TB1 XThR.TB2 2.14864f
C7323 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00584f
C7324 XA.XIR[8].XIC[0].icell.PDM Vbias 0.04207f
C7325 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.SM 0.0039f
C7326 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C7327 XA.XIR[10].XIC[13].icell.SM VPWR 0.00158f
C7328 XA.XIR[2].XIC[6].icell.PUM VPWR 0.00937f
C7329 XThC.TA3 XThC.Tn[2] 0.12602f
C7330 XA.XIR[11].XIC[13].icell.PDM Vbias 0.04261f
C7331 XA.XIR[13].XIC[3].icell.PUM Vbias 0.0031f
C7332 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00584f
C7333 XA.XIR[8].XIC[5].icell.Ien Vbias 0.21098f
C7334 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C7335 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00214f
C7336 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00584f
C7337 data[1] data[0] 0.64735f
C7338 XA.XIR[7].XIC[2].icell.Ien VPWR 0.1903f
C7339 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04031f
C7340 XA.XIR[5].XIC[13].icell.Ien Iout 0.06417f
C7341 XThR.Tn[13] XA.XIR[14].XIC[11].icell.SM 0.00121f
C7342 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01093f
C7343 XA.XIR[12].XIC[3].icell.SM Vbias 0.00701f
C7344 XA.XIR[5].XIC[5].icell.PDM Iout 0.00117f
C7345 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.SM 0.0039f
C7346 a_n1049_6699# VPWR 0.72162f
C7347 XA.XIR[14].XIC[14].icell.PDM Vbias 0.04261f
C7348 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13] 0.00341f
C7349 XA.XIR[14].XIC[6].icell.SM VPWR 0.00158f
C7350 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00584f
C7351 XThC.TBN XThC.Tn[4] 0.61061f
C7352 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.03425f
C7353 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C7354 XA.XIR[5].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7355 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07214f
C7356 Vbias bias[2] 0.05684f
C7357 XA.XIR[11].XIC[6].icell.PUM Vbias 0.0031f
C7358 a_4861_9615# XThC.Tn[3] 0.27012f
C7359 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C7360 XA.XIR[6].XIC[0].icell.Ien Iout 0.06411f
C7361 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7362 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00214f
C7363 XA.XIR[14].XIC[2].icell.SM Iout 0.00388f
C7364 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04031f
C7365 XA.XIR[8].XIC[7].icell.PDM Iout 0.00117f
C7366 XThC.TB2 a_5949_9615# 0.00844f
C7367 XThC.Tn[13] XThR.Tn[12] 0.2874f
C7368 XA.XIR[13].XIC[8].icell.SM VPWR 0.00158f
C7369 XThR.Tn[2] XA.XIR[3].XIC[9].icell.SM 0.00121f
C7370 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.SM 0.0039f
C7371 XA.XIR[9].XIC[14].icell.Ien Vbias 0.21098f
C7372 XA.XIR[8].XIC[12].icell.PUM VPWR 0.00937f
C7373 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00214f
C7374 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.SM 0.00168f
C7375 XThR.TAN a_n1319_5317# 0.00108f
C7376 XA.XIR[10].XIC[8].icell.PUM Vbias 0.0031f
C7377 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C7378 XA.XIR[13].XIC[4].icell.SM Iout 0.00388f
C7379 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C7380 XThR.TA2 a_n1319_6405# 0.00306f
C7381 XA.XIR[6].XIC[2].icell.SM Vbias 0.00701f
C7382 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C7383 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02762f
C7384 XThR.Tn[4] XA.XIR[4].XIC[8].icell.PDM 0.00341f
C7385 XThR.TB5 a_n1049_6405# 0.24821f
C7386 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.03425f
C7387 XThR.TBN XThR.Tn[13] 0.56841f
C7388 XThR.Tn[3] XA.XIR[3].XIC_15.icell.PDM 0.00341f
C7389 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PUM 0.00465f
C7390 XThC.TA1 XThC.Tn[8] 0.00205f
C7391 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C7392 XA.XIR[12].XIC[6].icell.Ien Iout 0.06417f
C7393 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC[0].icell.Ien 0.00214f
C7394 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00214f
C7395 XA.XIR[4].XIC[10].icell.PUM Vbias 0.0031f
C7396 XA.XIR[10].XIC_15.icell.Ien Iout 0.0642f
C7397 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.SM 0.0039f
C7398 VPWR Iout 54.1536f
C7399 XA.XIR[3].XIC[6].icell.SM VPWR 0.00158f
C7400 XA.XIR[11].XIC[7].icell.SM Iout 0.00388f
C7401 XA.XIR[1].XIC[4].icell.PDM Iout 0.00117f
C7402 XThR.Tn[9] VPWR 7.55029f
C7403 XThR.Tn[9] XA.XIR[10].XIC_15.icell.Ien 0.00117f
C7404 XA.XIR[11].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7405 XA.XIR[2].XIC[14].icell.PUM Vbias 0.0031f
C7406 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04031f
C7407 XA.XIR[2].XIC[5].icell.PDM Vbias 0.04261f
C7408 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02762f
C7409 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C7410 XA.XIR[6].XIC[9].icell.Ien VPWR 0.1903f
C7411 XA.XIR[3].XIC[2].icell.SM Iout 0.00388f
C7412 XA.XIR[7].XIC[10].icell.Ien Vbias 0.21098f
C7413 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00214f
C7414 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C7415 XA.XIR[4].XIC[4].icell.PDM VPWR 0.00799f
C7416 XThC.Tn[12] XThR.Tn[10] 0.28739f
C7417 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.15202f
C7418 XA.XIR[6].XIC[5].icell.Ien Iout 0.06417f
C7419 XA.XIR[14].XIC_dummy_left.icell.Ien Vbias 0.00329f
C7420 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7] 0.00341f
C7421 XThR.TB1 XThR.TAN2 0.12307f
C7422 XA.XIR[1].XIC[3].icell.SM VPWR 0.00158f
C7423 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PUM 0.00465f
C7424 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C7425 XA.XIR[12].XIC[0].icell.PUM VPWR 0.00937f
C7426 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C7427 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04031f
C7428 XA.XIR[13].XIC[10].icell.Ien Iout 0.06417f
C7429 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PUM 0.00471f
C7430 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02762f
C7431 XA.XIR[4].XIC[11].icell.SM Iout 0.00388f
C7432 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C7433 XA.XIR[8].XIC[0].icell.Ien Vbias 0.20951f
C7434 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.15202f
C7435 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.15202f
C7436 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04052f
C7437 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00584f
C7438 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02762f
C7439 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PUM 0.00465f
C7440 XA.XIR[2].XIC[12].icell.PDM Iout 0.00117f
C7441 XA.XIR[15].XIC[0].icell.Ien VPWR 0.32895f
C7442 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.SM 0.0039f
C7443 XA.XIR[0].XIC[10].icell.PUM Vbias 0.0031f
C7444 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02762f
C7445 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02762f
C7446 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C7447 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C7448 XA.XIR[14].XIC[2].icell.PUM VPWR 0.00937f
C7449 XThR.Tn[12] XA.XIR[13].XIC[7].icell.SM 0.00121f
C7450 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02762f
C7451 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C7452 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.SM 0.00168f
C7453 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PUM 0.00465f
C7454 XThR.Tn[4] XA.XIR[5].XIC[9].icell.Ien 0.00338f
C7455 XA.XIR[3].XIC[14].icell.SM Vbias 0.00701f
C7456 XThR.Tn[1] XA.XIR[2].XIC[6].icell.SM 0.00121f
C7457 XThC.Tn[8] XThR.Tn[2] 0.28739f
C7458 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[7].icell.Ien 0.00214f
C7459 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.15202f
C7460 XThR.Tn[3] XA.XIR[4].XIC[11].icell.Ien 0.00338f
C7461 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PUM 0.00465f
C7462 XA.XIR[10].XIC[3].icell.PDM VPWR 0.00799f
C7463 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00214f
C7464 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.03425f
C7465 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C7466 XA.XIR[10].XIC[11].icell.SM VPWR 0.00158f
C7467 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04031f
C7468 XA.XIR[15].XIC[2].icell.PDM Vbias 0.04261f
C7469 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C7470 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5] 0.00341f
C7471 XThR.Tn[13] XA.XIR[14].XIC[9].icell.SM 0.00121f
C7472 XA.XIR[0].XIC[11].icell.SM Iout 0.00367f
C7473 XA.XIR[12].XIC[0].icell.SM Iout 0.00388f
C7474 XA.XIR[1].XIC[11].icell.SM Vbias 0.00704f
C7475 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.SM 0.0039f
C7476 XA.XIR[14].XIC[8].icell.PDM Vbias 0.04261f
C7477 XA.XIR[5].XIC[7].icell.SM VPWR 0.00158f
C7478 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02762f
C7479 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Ien 0.00309f
C7480 XA.XIR[15].XIC[5].icell.Ien VPWR 0.32895f
C7481 XA.XIR[3].XIC[1].icell.PDM VPWR 0.00799f
C7482 XA.XIR[5].XIC[3].icell.SM Iout 0.00388f
C7483 XThC.TAN2 XThC.Tn[8] 0.1369f
C7484 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02762f
C7485 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00584f
C7486 XA.XIR[9].XIC[0].icell.PDM Vbias 0.04207f
C7487 XThR.TA1 data[5] 0.11096f
C7488 XThC.Tn[10] XThR.Tn[14] 0.28739f
C7489 XThC.Tn[0] XA.XIR[5].XIC_dummy_left.icell.Iout 0.00109f
C7490 XThC.TB5 a_7651_9569# 0.00418f
C7491 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.SM 0.00168f
C7492 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6] 0.00341f
C7493 XThR.TAN VPWR 1.67379f
C7494 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.SM 0.00168f
C7495 XA.XIR[15].XIC[9].icell.PDM Iout 0.00117f
C7496 XThC.Tn[6] XThR.Tn[5] 0.28739f
C7497 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.SM 0.0039f
C7498 XA.XIR[9].XIC[4].icell.SM Vbias 0.00701f
C7499 XA.XIR[8].XIC[2].icell.Ien VPWR 0.1903f
C7500 XA.XIR[1].XIC[14].icell.Ien Iout 0.06417f
C7501 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.SM 0.00168f
C7502 XA.XIR[4].XIC[2].icell.PUM VPWR 0.00937f
C7503 XA.XIR[10].XIC[14].icell.PUM VPWR 0.00937f
C7504 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C7505 XA.XIR[11].XIC[12].icell.PDM Vbias 0.04261f
C7506 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C7507 XA.XIR[15].XIC_15.icell.SM VPWR 0.00275f
C7508 XThR.TBN XA.XIR[8].XIC_dummy_left.icell.Ien 0.00243f
C7509 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02762f
C7510 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.SM 0.00168f
C7511 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C7512 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.15202f
C7513 XThC.Tn[11] XThR.Tn[4] 0.28739f
C7514 XA.XIR[11].XIC[3].icell.PUM VPWR 0.00937f
C7515 XThC.TBN a_6243_9615# 0.07731f
C7516 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00214f
C7517 XThR.TA3 XThR.Tn[3] 0.0306f
C7518 XThR.Tn[5] XA.XIR[6].XIC[7].icell.SM 0.00121f
C7519 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9] 0.00341f
C7520 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00214f
C7521 XA.XIR[9].XIC[7].icell.PDM Iout 0.00117f
C7522 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.15202f
C7523 XA.XIR[9].XIC[11].icell.Ien VPWR 0.1903f
C7524 XA.XIR[13].XIC[13].icell.SM VPWR 0.00158f
C7525 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7526 XA.XIR[14].XIC[13].icell.PDM Vbias 0.04261f
C7527 XA.XIR[10].XIC[5].icell.PUM VPWR 0.00937f
C7528 XA.XIR[2].XIC[4].icell.Ien Vbias 0.21098f
C7529 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Ien 0.00232f
C7530 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11] 0.00341f
C7531 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00584f
C7532 XA.XIR[12].XIC[14].icell.PDM VPWR 0.00809f
C7533 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C7534 XThR.Tn[2] XA.XIR[2].XIC[5].icell.PDM 0.00341f
C7535 XA.XIR[5].XIC[13].icell.PDM Vbias 0.04261f
C7536 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00584f
C7537 XA.XIR[9].XIC[7].icell.Ien Iout 0.06417f
C7538 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.15202f
C7539 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04031f
C7540 XA.XIR[0].XIC[5].icell.PDM Vbias 0.04275f
C7541 XThR.TB7 XThR.Tn[10] 0.07406f
C7542 XA.XIR[7].XIC[12].icell.PDM VPWR 0.00799f
C7543 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04031f
C7544 XThR.Tn[0] XA.XIR[1].XIC[12].icell.Ien 0.00338f
C7545 XA.XIR[0].XIC[2].icell.PUM VPWR 0.00877f
C7546 XA.XIR[8].XIC_15.icell.PDM Vbias 0.04401f
C7547 XA.XIR[14].XIC[6].icell.PUM Vbias 0.0031f
C7548 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.SM 0.0039f
C7549 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07555f
C7550 XA.XIR[4].XIC[7].icell.PUM VPWR 0.00937f
C7551 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C7552 XA.XIR[7].XIC[0].icell.PDM Iout 0.00117f
C7553 XA.XIR[2].XIC[11].icell.PUM VPWR 0.00937f
C7554 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C7555 XThC.Tn[3] XThR.Tn[3] 0.28739f
C7556 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C7557 XA.XIR[13].XIC[8].icell.PUM Vbias 0.0031f
C7558 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.SM 0.0039f
C7559 XThC.Tn[13] XThR.Tn[0] 0.28789f
C7560 XA.XIR[8].XIC[10].icell.Ien Vbias 0.21098f
C7561 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C7562 XA.XIR[7].XIC[7].icell.Ien VPWR 0.1903f
C7563 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04031f
C7564 XThC.Tn[6] Vbias 2.22871f
C7565 XA.XIR[12].XIC[8].icell.SM Vbias 0.00701f
C7566 XA.XIR[7].XIC[3].icell.Ien Iout 0.06417f
C7567 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C7568 XThR.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.00338f
C7569 XA.XIR[10].XIC[9].icell.SM VPWR 0.00158f
C7570 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Iout 0.00347f
C7571 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PUM 0.00465f
C7572 XA.XIR[1].XIC[12].icell.PDM Vbias 0.04261f
C7573 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00584f
C7574 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PUM 0.00465f
C7575 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02827f
C7576 XA.XIR[3].XIC[0].icell.Ien VPWR 0.1903f
C7577 XA.XIR[13].XIC_15.icell.Ien Iout 0.0642f
C7578 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00584f
C7579 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02762f
C7580 XA.XIR[14].XIC[7].icell.SM Iout 0.00388f
C7581 XA.XIR[14].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7582 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C7583 XA.XIR[3].XIC[6].icell.PUM Vbias 0.0031f
C7584 XThC.Tn[7] XThR.Tn[6] 0.28739f
C7585 XThR.Tn[2] XA.XIR[3].XIC[14].icell.SM 0.00121f
C7586 XThR.Tn[3] XA.XIR[4].XIC[1].icell.SM 0.00121f
C7587 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38919f
C7588 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.SM 0.0039f
C7589 XThR.Tn[7] XA.XIR[8].XIC[4].icell.Ien 0.00338f
C7590 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.03425f
C7591 XA.XIR[6].XIC[7].icell.SM Vbias 0.00701f
C7592 XA.XIR[0].XIC[7].icell.PUM VPWR 0.00877f
C7593 XThC.Tn[12] XThR.Tn[13] 0.28739f
C7594 a_9827_9569# XThC.Tn[13] 0.00173f
C7595 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C7596 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.04036f
C7597 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C7598 XThC.Tn[0] XThC.Tn[2] 0.1179f
C7599 XA.XIR[4].XIC[0].icell.PDM Vbias 0.04207f
C7600 XA.XIR[2].XIC_15.icell.SM VPWR 0.00275f
C7601 XThC.TB1 a_2979_9615# 0.21263f
C7602 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02762f
C7603 XA.XIR[15].XIC_dummy_left.icell.SM VPWR 0.00269f
C7604 XA.XIR[1].XIC[3].icell.PUM Vbias 0.0031f
C7605 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.15202f
C7606 XThC.Tn[5] XThC.Tn[6] 0.30991f
C7607 XThC.TB4 Vbias 0.01548f
C7608 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01785f
C7609 XA.XIR[4].XIC_15.icell.PUM Vbias 0.0031f
C7610 XA.XIR[3].XIC[11].icell.SM VPWR 0.00158f
C7611 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.15202f
C7612 XThR.Tn[10] XA.XIR[11].XIC[5].icell.Ien 0.00338f
C7613 XThC.Tn[11] XThR.Tn[8] 0.28739f
C7614 XThC.Tn[2] XThR.Tn[12] 0.28739f
C7615 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02762f
C7616 XThR.TB3 XThR.TB5 0.04438f
C7617 XA.XIR[3].XIC[7].icell.SM Iout 0.00388f
C7618 XA.XIR[6].XIC[14].icell.Ien VPWR 0.19036f
C7619 XThR.Tn[0] XA.XIR[0].XIC[6].icell.PDM 0.00341f
C7620 XThR.TB2 data[5] 0.017f
C7621 XA.XIR[6].XIC[8].icell.PDM VPWR 0.00799f
C7622 XA.XIR[7].XIC_15.icell.Ien Vbias 0.21234f
C7623 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00584f
C7624 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PUM 0.00444f
C7625 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.03425f
C7626 XA.XIR[5].XIC[2].icell.PUM Vbias 0.0031f
C7627 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.03425f
C7628 VPWR data[1] 0.44103f
C7629 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.15202f
C7630 XA.XIR[6].XIC[10].icell.Ien Iout 0.06417f
C7631 XA.XIR[10].XIC[12].icell.PUM VPWR 0.00937f
C7632 XA.XIR[1].XIC[8].icell.SM VPWR 0.00158f
C7633 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.15202f
C7634 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C7635 XThR.Tn[13] XA.XIR[14].XIC[14].icell.SM 0.00121f
C7636 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.SM 0.00168f
C7637 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.SM 0.00168f
C7638 XA.XIR[4].XIC[7].icell.PDM Iout 0.00117f
C7639 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.03023f
C7640 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00214f
C7641 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C7642 XA.XIR[14].XIC[1].icell.PUM Vbias 0.0031f
C7643 XA.XIR[1].XIC[4].icell.SM Iout 0.00388f
C7644 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C7645 XThR.TB3 a_n1335_7243# 0.00941f
C7646 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00214f
C7647 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Iout 0.00347f
C7648 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PUM 0.00465f
C7649 XA.XIR[13].XIC[3].icell.PDM VPWR 0.00799f
C7650 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00584f
C7651 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.SM 0.00168f
C7652 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PUM 0.00465f
C7653 XThC.TB4 XThC.Tn[5] 0.00814f
C7654 XA.XIR[13].XIC[11].icell.SM VPWR 0.00158f
C7655 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.15202f
C7656 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.15202f
C7657 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PUM 0.00268f
C7658 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.03425f
C7659 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C7660 XA.XIR[0].XIC_15.icell.PUM Vbias 0.0031f
C7661 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.03425f
C7662 XA.XIR[12].XIC[8].icell.PDM VPWR 0.00799f
C7663 XThC.Tn[1] XThR.Tn[10] 0.28739f
C7664 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.04036f
C7665 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C7666 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02762f
C7667 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C7668 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C7669 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.03425f
C7670 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.SM 0.00168f
C7671 XA.XIR[15].XIC[1].icell.Ien Iout 0.06807f
C7672 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04031f
C7673 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00214f
C7674 XA.XIR[9].XIC[1].icell.SM VPWR 0.00158f
C7675 XThC.Tn[11] XThR.Tn[1] 0.28739f
C7676 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02762f
C7677 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C7678 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.15202f
C7679 XThR.Tn[4] XA.XIR[5].XIC[14].icell.Ien 0.00338f
C7680 XThR.Tn[1] XA.XIR[2].XIC[11].icell.SM 0.00121f
C7681 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02762f
C7682 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04031f
C7683 XA.XIR[5].XIC[7].icell.PUM Vbias 0.0031f
C7684 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.04036f
C7685 XThR.TB7 a_n997_1803# 0.00571f
C7686 XA.XIR[15].XIC[3].icell.SM Vbias 0.00701f
C7687 XThR.TBN a_n997_3979# 0.23021f
C7688 XA.XIR[11].XIC[2].icell.PDM Iout 0.00117f
C7689 XThC.TA2 XThC.TB4 0.04137f
C7690 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.SM 0.0039f
C7691 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PUM 0.00465f
C7692 XThC.TB2 XThC.TA3 0.2319f
C7693 XThC.TA1 XThC.TB4 0.02767f
C7694 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PUM 0.00465f
C7695 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00214f
C7696 XThR.Tn[0] XA.XIR[1].XIC[2].icell.SM 0.00121f
C7697 XA.XIR[10].XIC[13].icell.Ien VPWR 0.1903f
C7698 XA.XIR[10].XIC[6].icell.PDM Iout 0.00117f
C7699 XThC.TB1 XThC.TB2 2.14864f
C7700 XA.XIR[11].XIC[11].icell.PDM Vbias 0.04261f
C7701 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.03425f
C7702 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04031f
C7703 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7704 XThR.TB1 a_n1335_8331# 0.0097f
C7705 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C7706 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02762f
C7707 XA.XIR[5].XIC[12].icell.SM VPWR 0.00158f
C7708 XThR.Tn[13] XA.XIR[14].XIC[11].icell.Ien 0.00338f
C7709 XA.XIR[5].XIC[4].icell.PDM VPWR 0.00799f
C7710 XThC.TB3 XThC.Tn[10] 0.29462f
C7711 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00214f
C7712 XA.XIR[13].XIC[14].icell.PUM VPWR 0.00937f
C7713 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C7714 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00214f
C7715 XA.XIR[4].XIC[0].icell.Ien Vbias 0.20951f
C7716 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.SM 0.0039f
C7717 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00214f
C7718 XA.XIR[14].XIC[12].icell.PDM Vbias 0.04261f
C7719 XA.XIR[5].XIC[8].icell.SM Iout 0.00388f
C7720 XThR.TAN2 data[5] 0.0148f
C7721 XThR.TB2 a_n1049_6699# 0.00851f
C7722 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02762f
C7723 XA.XIR[15].XIC[6].icell.Ien Iout 0.06807f
C7724 XA.XIR[9].XIC_15.icell.PDM Vbias 0.04401f
C7725 XThR.Tn[14] XA.XIR[15].XIC[0].icell.SM 0.00128f
C7726 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C7727 XA.XIR[12].XIC[13].icell.PDM VPWR 0.00799f
C7728 XA.XIR[3].XIC[4].icell.PDM Iout 0.00117f
C7729 XThC.TB3 a_4861_9615# 0.0093f
C7730 XA.XIR[8].XIC[6].icell.PDM VPWR 0.00799f
C7731 XThC.Tn[6] XThR.Tn[2] 0.28739f
C7732 XA.XIR[7].XIC[0].icell.SM Vbias 0.00675f
C7733 XA.XIR[14].XIC[3].icell.PUM VPWR 0.00937f
C7734 XThR.TA3 a_n1049_5317# 0.02018f
C7735 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.SM 0.0039f
C7736 XThR.TA1 XThR.TAN 0.30355f
C7737 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C7738 XA.XIR[13].XIC[5].icell.PUM VPWR 0.00937f
C7739 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.SM 0.00168f
C7740 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.SM 0.0039f
C7741 XThC.TA2 a_5949_10571# 0.00467f
C7742 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04037f
C7743 XA.XIR[9].XIC[9].icell.SM Vbias 0.00701f
C7744 XA.XIR[10].XIC[3].icell.Ien Vbias 0.21098f
C7745 XA.XIR[8].XIC[7].icell.Ien VPWR 0.1903f
C7746 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.SM 0.0039f
C7747 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01149f
C7748 XA.XIR[12].XIC[5].icell.SM VPWR 0.00158f
C7749 XA.XIR[8].XIC[3].icell.Ien Iout 0.06417f
C7750 XA.XIR[12].XIC[13].icell.SM Vbias 0.00701f
C7751 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12] 0.00341f
C7752 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PUM 0.00465f
C7753 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.15202f
C7754 XThR.Tn[8] XA.XIR[9].XIC[3].icell.Ien 0.00338f
C7755 XThR.TB7 XThR.Tn[13] 0.10781f
C7756 XThR.Tn[3] XA.XIR[3].XIC[2].icell.PDM 0.00341f
C7757 XA.XIR[10].XIC[14].icell.SM VPWR 0.00207f
C7758 XA.XIR[12].XIC[1].icell.SM Iout 0.00388f
C7759 XA.XIR[11].XIC[8].icell.PUM VPWR 0.00937f
C7760 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C7761 XA.XIR[7].XIC[8].icell.PDM Vbias 0.04261f
C7762 XA.XIR[1].XIC[3].icell.PDM VPWR 0.00799f
C7763 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04031f
C7764 XA.XIR[0].XIC[0].icell.Ien Vbias 0.20983f
C7765 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.SM 0.0039f
C7766 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00214f
C7767 XThC.TB7 XThC.Tn[10] 0.07406f
C7768 XThR.Tn[5] XA.XIR[6].XIC[12].icell.SM 0.00121f
C7769 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.15202f
C7770 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04031f
C7771 XA.XIR[4].XIC[5].icell.Ien Vbias 0.21098f
C7772 XA.XIR[3].XIC[3].icell.PUM VPWR 0.00937f
C7773 XThC.TAN2 XThC.Tn[6] 0.00131f
C7774 XThR.TB2 XThR.Tn[9] 0.292f
C7775 XA.XIR[2].XIC[9].icell.Ien Vbias 0.21098f
C7776 XA.XIR[10].XIC[10].icell.PUM VPWR 0.00937f
C7777 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C7778 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.03425f
C7779 XThR.Tn[14] XA.XIR[15].XIC[5].icell.SM 0.00121f
C7780 XA.XIR[3].XIC_dummy_left.icell.SM VPWR 0.00269f
C7781 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00214f
C7782 XThR.TBN XThR.Tn[7] 0.8998f
C7783 XA.XIR[6].XIC[4].icell.SM VPWR 0.00158f
C7784 XA.XIR[9].XIC[12].icell.Ien Iout 0.06417f
C7785 XThR.TBN a_n997_2891# 0.22804f
C7786 XA.XIR[7].XIC[5].icell.SM Vbias 0.00701f
C7787 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.15202f
C7788 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7789 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C7790 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00214f
C7791 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02762f
C7792 XA.XIR[13].XIC[9].icell.SM VPWR 0.00158f
C7793 XThC.TBN a_8963_9569# 0.22784f
C7794 XA.XIR[4].XIC[12].icell.PUM VPWR 0.00937f
C7795 XThC.Tn[0] XThR.Tn[4] 0.28743f
C7796 XA.XIR[7].XIC_15.icell.PDM Iout 0.00133f
C7797 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7798 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04031f
C7799 XA.XIR[2].XIC[11].icell.PDM VPWR 0.00799f
C7800 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00584f
C7801 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8] 0.00341f
C7802 XA.XIR[8].XIC_15.icell.Ien Vbias 0.21234f
C7803 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00214f
C7804 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00584f
C7805 XA.XIR[7].XIC[12].icell.Ien VPWR 0.1903f
C7806 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.03425f
C7807 XThC.TB4 XThC.TAN2 0.03415f
C7808 XThC.Tn[10] VPWR 6.83631f
C7809 XA.XIR[0].XIC[5].icell.Ien Vbias 0.2113f
C7810 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.15202f
C7811 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00214f
C7812 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.SM 0.0039f
C7813 XA.XIR[7].XIC[8].icell.Ien Iout 0.06417f
C7814 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.SM 0.00168f
C7815 XThR.Tn[6] XA.XIR[7].XIC[2].icell.Ien 0.00338f
C7816 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C7817 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04031f
C7818 XThR.TB1 XThR.TB5 0.05054f
C7819 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PUM 0.00465f
C7820 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02764f
C7821 a_4861_9615# VPWR 0.70525f
C7822 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.03425f
C7823 XThR.Tn[4] XA.XIR[5].XIC[4].icell.SM 0.00121f
C7824 XA.XIR[10].XIC[11].icell.Ien VPWR 0.1903f
C7825 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00214f
C7826 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[4].icell.SM 0.0039f
C7827 XA.XIR[3].XIC[11].icell.PUM Vbias 0.0031f
C7828 XThR.Tn[3] XA.XIR[4].XIC[6].icell.SM 0.00121f
C7829 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.SM 0.0039f
C7830 XThR.Tn[7] XA.XIR[8].XIC[9].icell.Ien 0.00338f
C7831 XA.XIR[3].XIC[1].icell.Ien Iout 0.06417f
C7832 XThC.Tn[2] XThR.Tn[0] 0.28882f
C7833 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.SM 0.00168f
C7834 XA.XIR[0].XIC[12].icell.PUM VPWR 0.00878f
C7835 XA.XIR[6].XIC[12].icell.SM Vbias 0.00701f
C7836 XA.XIR[6].XIC[4].icell.PDM Vbias 0.04261f
C7837 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C7838 XA.XIR[12].XIC[1].icell.PUM VPWR 0.00937f
C7839 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.03425f
C7840 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C7841 XThC.TB5 a_5949_9615# 0.0093f
C7842 XA.XIR[4].XIC_15.icell.PDM Vbias 0.04401f
C7843 XThR.TB6 XThR.Tn[12] 0.02431f
C7844 XA.XIR[13].XIC[12].icell.PUM VPWR 0.00937f
C7845 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5] 0.00346f
C7846 XThR.TB1 a_n1049_8581# 0.21263f
C7847 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.0352f
C7848 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.SM 0.00168f
C7849 XA.XIR[1].XIC[8].icell.PUM Vbias 0.0031f
C7850 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.03425f
C7851 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.15202f
C7852 XThC.TAN XThC.Tn[8] 0.09736f
C7853 XThR.TAN2 XThR.Tn[9] 0.12398f
C7854 XA.XIR[5].XIC[4].icell.PUM VPWR 0.00937f
C7855 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C7856 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.1106f
C7857 XA.XIR[3].XIC[12].icell.SM Iout 0.00388f
C7858 XThR.Tn[6] Iout 1.1623f
C7859 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00214f
C7860 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C7861 XA.XIR[10].XIC[0].icell.Ien Iout 0.06411f
C7862 XA.XIR[15].XIC[8].icell.PDM VPWR 0.0114f
C7863 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C7864 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C7865 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.PDM 0.00591f
C7866 XThR.Tn[9] XA.XIR[10].XIC[0].icell.Ien 0.0037f
C7867 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C7868 XThR.TAN XThR.TB2 0.22599f
C7869 XThC.Tn[1] XThR.Tn[13] 0.28739f
C7870 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02762f
C7871 XA.XIR[6].XIC_15.icell.Ien Iout 0.0642f
C7872 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.03425f
C7873 XA.XIR[12].XIC[4].icell.PDM Vbias 0.04261f
C7874 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.15202f
C7875 XA.XIR[1].XIC[13].icell.SM VPWR 0.00158f
C7876 XA.XIR[6].XIC[11].icell.PDM Iout 0.00117f
C7877 XA.XIR[12].XIC[11].icell.SM Vbias 0.00701f
C7878 XA.XIR[3].XIC_15.icell.SM Vbias 0.00701f
C7879 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C7880 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.15202f
C7881 XThR.Tn[1] XA.XIR[1].XIC[7].icell.PDM 0.00341f
C7882 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C7883 XA.XIR[11].XIC[10].icell.PDM Vbias 0.04261f
C7884 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.SM 0.00168f
C7885 XA.XIR[1].XIC[9].icell.SM Iout 0.00388f
C7886 a_2979_9615# XThC.Tn[0] 0.28426f
C7887 XThC.Tn[4] Iout 0.83918f
C7888 XA.XIR[14].XIC[2].icell.PDM Iout 0.00117f
C7889 XA.XIR[2].XIC[1].icell.Ien VPWR 0.1903f
C7890 XThC.Tn[4] XThR.Tn[9] 0.28739f
C7891 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.15202f
C7892 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00584f
C7893 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00584f
C7894 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.15202f
C7895 XA.XIR[9].XIC[6].icell.PDM VPWR 0.00799f
C7896 XThC.Tn[0] XThR.Tn[8] 0.2874f
C7897 XA.XIR[8].XIC[0].icell.SM Vbias 0.00675f
C7898 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.SM 0.00168f
C7899 XA.XIR[13].XIC[13].icell.Ien VPWR 0.1903f
C7900 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.SM 0.00168f
C7901 XA.XIR[13].XIC[6].icell.PDM Iout 0.00117f
C7902 XA.XIR[14].XIC[11].icell.PDM Vbias 0.04261f
C7903 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02762f
C7904 XA.XIR[12].XIC[12].icell.PDM VPWR 0.00799f
C7905 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.03425f
C7906 XA.XIR[9].XIC[6].icell.SM VPWR 0.00158f
C7907 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.03426f
C7908 XA.XIR[6].XIC[0].icell.PUM VPWR 0.00937f
C7909 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.15202f
C7910 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[12].icell.Ien 0.00214f
C7911 XA.XIR[5].XIC[12].icell.PUM Vbias 0.0031f
C7912 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PDM 0.00172f
C7913 XA.XIR[15].XIC[8].icell.SM Vbias 0.00701f
C7914 XA.XIR[5].XIC[0].icell.PDM Vbias 0.04207f
C7915 XA.XIR[9].XIC[2].icell.SM Iout 0.00388f
C7916 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00214f
C7917 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00214f
C7918 XA.XIR[3].XIC[12].icell.PDM Vbias 0.04261f
C7919 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PDM 0.00587f
C7920 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C7921 XA.XIR[15].XIC[13].icell.PDM VPWR 0.0114f
C7922 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.03425f
C7923 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C7924 XThR.Tn[0] XA.XIR[1].XIC[7].icell.SM 0.00121f
C7925 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00214f
C7926 XThR.Tn[11] XA.XIR[12].XIC[1].icell.Ien 0.00338f
C7927 XA.XIR[8].XIC[2].icell.PDM Vbias 0.04261f
C7928 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00584f
C7929 XA.XIR[4].XIC[2].icell.Ien VPWR 0.1903f
C7930 XA.XIR[12].XIC[14].icell.PUM Vbias 0.0031f
C7931 XA.XIR[2].XIC[6].icell.Ien VPWR 0.1903f
C7932 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00584f
C7933 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14] 0.00341f
C7934 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PUM 0.00465f
C7935 XThC.Tn[0] XThR.Tn[1] 0.28748f
C7936 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.0353f
C7937 XA.XIR[13].XIC[3].icell.Ien Vbias 0.21098f
C7938 XA.XIR[8].XIC[5].icell.SM Vbias 0.00701f
C7939 XA.XIR[2].XIC[2].icell.Ien Iout 0.06417f
C7940 XA.XIR[7].XIC[2].icell.SM VPWR 0.00158f
C7941 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04031f
C7942 XA.XIR[12].XIC[5].icell.PUM Vbias 0.0031f
C7943 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00214f
C7944 XA.XIR[0].XIC[11].icell.PDM VPWR 0.00774f
C7945 XA.XIR[5].XIC[13].icell.SM Iout 0.00388f
C7946 XA.XIR[5].XIC[7].icell.PDM Iout 0.00117f
C7947 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.SM 0.0039f
C7948 XA.XIR[13].XIC[14].icell.SM VPWR 0.00207f
C7949 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02762f
C7950 XA.XIR[14].XIC[8].icell.PUM VPWR 0.00937f
C7951 XThR.TAN XThR.TAN2 0.35142f
C7952 XA.XIR[11].XIC[6].icell.Ien Vbias 0.21098f
C7953 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02762f
C7954 XA.XIR[9].XIC_dummy_left.icell.Ien Vbias 0.00329f
C7955 XA.XIR[8].XIC[9].icell.PDM Iout 0.00117f
C7956 XA.XIR[6].XIC[0].icell.SM Iout 0.00388f
C7957 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04031f
C7958 XA.XIR[13].XIC[10].icell.PUM VPWR 0.00937f
C7959 XA.XIR[9].XIC[14].icell.SM Vbias 0.00701f
C7960 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.SM 0.00168f
C7961 XThC.TB2 XThC.Tn[0] 0.00125f
C7962 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.SM 0.0039f
C7963 XA.XIR[8].XIC[12].icell.Ien VPWR 0.1903f
C7964 XA.XIR[10].XIC[8].icell.Ien Vbias 0.21098f
C7965 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00584f
C7966 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C7967 XThR.TAN XThR.Tn[6] 0.04822f
C7968 XThR.TBN a_n997_1579# 0.23006f
C7969 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04031f
C7970 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.SM 0.00168f
C7971 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18966f
C7972 XA.XIR[6].XIC[4].icell.PUM Vbias 0.0031f
C7973 XA.XIR[8].XIC[8].icell.Ien Iout 0.06417f
C7974 XThR.Tn[4] XA.XIR[4].XIC[10].icell.PDM 0.00341f
C7975 XThR.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.00338f
C7976 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.15202f
C7977 XThC.TB3 a_7651_9569# 0.00604f
C7978 XA.XIR[12].XIC[6].icell.SM Iout 0.00388f
C7979 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00214f
C7980 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PUM 0.00465f
C7981 XA.XIR[10].XIC_15.icell.PDM Iout 0.00133f
C7982 XA.XIR[3].XIC[8].icell.PUM VPWR 0.00937f
C7983 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C7984 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PDM 0.00172f
C7985 XA.XIR[4].XIC[10].icell.Ien Vbias 0.21098f
C7986 XThC.Tn[12] XThR.Tn[7] 0.28739f
C7987 XA.XIR[12].XIC[9].icell.SM Vbias 0.00701f
C7988 XA.XIR[2].XIC[14].icell.Ien Vbias 0.21098f
C7989 XA.XIR[2].XIC[7].icell.PDM Vbias 0.04261f
C7990 XA.XIR[1].XIC[6].icell.PDM Iout 0.00117f
C7991 data[7] VGND 0.49949f
C7992 data[6] VGND 0.47974f
C7993 data[4] VGND 0.59317f
C7994 data[5] VGND 1.17814f
C7995 Iout VGND 0.32054p
C7996 data[3] VGND 0.49953f
C7997 data[2] VGND 0.48064f
C7998 data[0] VGND 0.59421f
C7999 data[1] VGND 1.17844f
C8000 bias[2] VGND 0.77552f
C8001 bias[0] VGND 1.22004f
C8002 Vbias VGND 0.23106p
C8003 bias[1] VGND 0.62458f
C8004 VPWR VGND 0.34108p
C8005 a_n997_715# VGND 0.5638f
C8006 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.75246f
C8007 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C8008 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64516f
C8009 XA.XIR[15].XIC_15.icell.SM VGND 0.00474f
C8010 XA.XIR[15].XIC_dummy_right.icell.PUM VGND 0.00215f
C8011 XA.XIR[15].XIC_15.icell.Ien VGND 0.44292f
C8012 XA.XIR[15].XIC[14].icell.SM VGND 0.00502f
C8013 XA.XIR[15].XIC_15.icell.PUM VGND 0.00282f
C8014 XA.XIR[15].XIC[14].icell.Ien VGND 0.44322f
C8015 XA.XIR[15].XIC[13].icell.SM VGND 0.00502f
C8016 XA.XIR[15].XIC[14].icell.PUM VGND 0.00293f
C8017 XA.XIR[15].XIC[13].icell.Ien VGND 0.44322f
C8018 XA.XIR[15].XIC[12].icell.SM VGND 0.00502f
C8019 XA.XIR[15].XIC[13].icell.PUM VGND 0.00293f
C8020 XA.XIR[15].XIC[12].icell.Ien VGND 0.44322f
C8021 XA.XIR[15].XIC[11].icell.SM VGND 0.00502f
C8022 XA.XIR[15].XIC[12].icell.PUM VGND 0.00293f
C8023 XA.XIR[15].XIC[11].icell.Ien VGND 0.44322f
C8024 XA.XIR[15].XIC[10].icell.SM VGND 0.00502f
C8025 XA.XIR[15].XIC[11].icell.PUM VGND 0.00293f
C8026 XA.XIR[15].XIC[10].icell.Ien VGND 0.44322f
C8027 XA.XIR[15].XIC[9].icell.SM VGND 0.00502f
C8028 XA.XIR[15].XIC[10].icell.PUM VGND 0.00293f
C8029 XA.XIR[15].XIC[9].icell.Ien VGND 0.44322f
C8030 XA.XIR[15].XIC[8].icell.SM VGND 0.00502f
C8031 XA.XIR[15].XIC[9].icell.PUM VGND 0.00293f
C8032 XA.XIR[15].XIC[8].icell.Ien VGND 0.44322f
C8033 XA.XIR[15].XIC[7].icell.SM VGND 0.00502f
C8034 XA.XIR[15].XIC[8].icell.PUM VGND 0.00293f
C8035 XA.XIR[15].XIC[7].icell.Ien VGND 0.44322f
C8036 XA.XIR[15].XIC[6].icell.SM VGND 0.00502f
C8037 XA.XIR[15].XIC[7].icell.PUM VGND 0.00293f
C8038 XA.XIR[15].XIC[6].icell.Ien VGND 0.44322f
C8039 XA.XIR[15].XIC[5].icell.SM VGND 0.00502f
C8040 XA.XIR[15].XIC[6].icell.PUM VGND 0.00293f
C8041 XA.XIR[15].XIC[5].icell.Ien VGND 0.44322f
C8042 XA.XIR[15].XIC[4].icell.SM VGND 0.00502f
C8043 XA.XIR[15].XIC[5].icell.PUM VGND 0.00293f
C8044 XA.XIR[15].XIC[4].icell.Ien VGND 0.44322f
C8045 XA.XIR[15].XIC[3].icell.SM VGND 0.00502f
C8046 XA.XIR[15].XIC[4].icell.PUM VGND 0.00293f
C8047 XA.XIR[15].XIC[3].icell.Ien VGND 0.44322f
C8048 XA.XIR[15].XIC[2].icell.SM VGND 0.00502f
C8049 XA.XIR[15].XIC[3].icell.PUM VGND 0.00293f
C8050 XA.XIR[15].XIC[2].icell.Ien VGND 0.44322f
C8051 XA.XIR[15].XIC[1].icell.SM VGND 0.00502f
C8052 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70718f
C8053 XA.XIR[15].XIC[2].icell.PUM VGND 0.00293f
C8054 XA.XIR[15].XIC[1].icell.Ien VGND 0.44322f
C8055 XA.XIR[15].XIC[0].icell.SM VGND 0.00502f
C8056 XA.XIR[15].XIC[1].icell.PUM VGND 0.00293f
C8057 XA.XIR[15].XIC[0].icell.Ien VGND 0.44356f
C8058 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01044f
C8059 XA.XIR[15].XIC[0].icell.PUM VGND 0.00516f
C8060 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.61163f
C8061 XA.XIR[15].XIC_dummy_left.icell.PUM VGND 0.00215f
C8062 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23279f
C8063 XA.XIR[15].XIC_15.icell.PDM VGND 0.18779f
C8064 XA.XIR[15].XIC[14].icell.PDM VGND 0.18733f
C8065 XA.XIR[15].XIC[13].icell.PDM VGND 0.18733f
C8066 XA.XIR[15].XIC[12].icell.PDM VGND 0.18733f
C8067 XA.XIR[15].XIC[11].icell.PDM VGND 0.18733f
C8068 XA.XIR[15].XIC[10].icell.PDM VGND 0.18733f
C8069 XA.XIR[15].XIC[9].icell.PDM VGND 0.18733f
C8070 XA.XIR[15].XIC[8].icell.PDM VGND 0.18733f
C8071 XA.XIR[15].XIC[7].icell.PDM VGND 0.18733f
C8072 XA.XIR[15].XIC[6].icell.PDM VGND 0.18733f
C8073 XA.XIR[15].XIC[5].icell.PDM VGND 0.18733f
C8074 XA.XIR[15].XIC[4].icell.PDM VGND 0.18733f
C8075 XA.XIR[15].XIC[3].icell.PDM VGND 0.18733f
C8076 XA.XIR[15].XIC[2].icell.PDM VGND 0.18733f
C8077 XA.XIR[15].XIC[1].icell.PDM VGND 0.18733f
C8078 XA.XIR[15].XIC[0].icell.PDM VGND 0.18741f
C8079 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C8080 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85795f
C8081 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C8082 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60802f
C8083 XA.XIR[14].XIC_15.icell.SM VGND 0.00474f
C8084 XA.XIR[14].XIC_dummy_right.icell.PUM VGND 0.00215f
C8085 XA.XIR[14].XIC_15.icell.Ien VGND 0.37063f
C8086 XA.XIR[14].XIC[14].icell.SM VGND 0.00502f
C8087 XA.XIR[14].XIC_15.icell.PUM VGND 0.00282f
C8088 XA.XIR[14].XIC[14].icell.Ien VGND 0.37144f
C8089 XA.XIR[14].XIC[13].icell.SM VGND 0.00502f
C8090 XA.XIR[14].XIC[14].icell.PUM VGND 0.00293f
C8091 XA.XIR[14].XIC[13].icell.Ien VGND 0.37144f
C8092 XA.XIR[14].XIC[12].icell.SM VGND 0.00502f
C8093 XA.XIR[14].XIC[13].icell.PUM VGND 0.00293f
C8094 XA.XIR[14].XIC[12].icell.Ien VGND 0.37144f
C8095 XA.XIR[14].XIC[11].icell.SM VGND 0.00502f
C8096 XA.XIR[14].XIC[12].icell.PUM VGND 0.00293f
C8097 XA.XIR[14].XIC[11].icell.Ien VGND 0.37144f
C8098 XA.XIR[14].XIC[10].icell.SM VGND 0.00502f
C8099 XA.XIR[14].XIC[11].icell.PUM VGND 0.00293f
C8100 XA.XIR[14].XIC[10].icell.Ien VGND 0.37144f
C8101 XA.XIR[14].XIC[9].icell.SM VGND 0.00502f
C8102 XA.XIR[14].XIC[10].icell.PUM VGND 0.00293f
C8103 XA.XIR[14].XIC[9].icell.Ien VGND 0.37144f
C8104 XA.XIR[14].XIC[8].icell.SM VGND 0.00502f
C8105 XA.XIR[14].XIC[9].icell.PUM VGND 0.00293f
C8106 XA.XIR[14].XIC[8].icell.Ien VGND 0.37144f
C8107 XA.XIR[14].XIC[7].icell.SM VGND 0.00502f
C8108 XA.XIR[14].XIC[8].icell.PUM VGND 0.00293f
C8109 XA.XIR[14].XIC[7].icell.Ien VGND 0.37144f
C8110 XA.XIR[14].XIC[6].icell.SM VGND 0.00502f
C8111 XA.XIR[14].XIC[7].icell.PUM VGND 0.00293f
C8112 XA.XIR[14].XIC[6].icell.Ien VGND 0.37144f
C8113 XA.XIR[14].XIC[5].icell.SM VGND 0.00502f
C8114 XA.XIR[14].XIC[6].icell.PUM VGND 0.00293f
C8115 XA.XIR[14].XIC[5].icell.Ien VGND 0.37144f
C8116 XA.XIR[14].XIC[4].icell.SM VGND 0.00502f
C8117 XA.XIR[14].XIC[5].icell.PUM VGND 0.00293f
C8118 XA.XIR[14].XIC[4].icell.Ien VGND 0.37144f
C8119 XA.XIR[14].XIC[3].icell.SM VGND 0.00502f
C8120 XA.XIR[14].XIC[4].icell.PUM VGND 0.00293f
C8121 XA.XIR[14].XIC[3].icell.Ien VGND 0.37144f
C8122 XA.XIR[14].XIC[2].icell.SM VGND 0.00502f
C8123 XA.XIR[14].XIC[3].icell.PUM VGND 0.00293f
C8124 XA.XIR[14].XIC[2].icell.Ien VGND 0.37144f
C8125 XA.XIR[14].XIC[1].icell.SM VGND 0.00502f
C8126 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80696f
C8127 XThR.Tn[14] VGND 14.14128f
C8128 XA.XIR[14].XIC[2].icell.PUM VGND 0.00293f
C8129 XA.XIR[14].XIC[1].icell.Ien VGND 0.37144f
C8130 XA.XIR[14].XIC[0].icell.SM VGND 0.00502f
C8131 a_n997_1579# VGND 0.54776f
C8132 XA.XIR[14].XIC[1].icell.PUM VGND 0.00293f
C8133 XA.XIR[14].XIC[0].icell.Ien VGND 0.37178f
C8134 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01044f
C8135 XA.XIR[14].XIC[0].icell.PUM VGND 0.00516f
C8136 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57579f
C8137 XA.XIR[14].XIC_dummy_left.icell.PUM VGND 0.00215f
C8138 a_n997_1803# VGND 0.53619f
C8139 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C8140 XA.XIR[14].XIC_15.icell.PDM VGND 0.18855f
C8141 XA.XIR[14].XIC[14].icell.PDM VGND 0.18809f
C8142 XA.XIR[14].XIC[13].icell.PDM VGND 0.18809f
C8143 XA.XIR[14].XIC[12].icell.PDM VGND 0.18809f
C8144 XA.XIR[14].XIC[11].icell.PDM VGND 0.18809f
C8145 XA.XIR[14].XIC[10].icell.PDM VGND 0.18809f
C8146 XA.XIR[14].XIC[9].icell.PDM VGND 0.18809f
C8147 XA.XIR[14].XIC[8].icell.PDM VGND 0.18809f
C8148 XA.XIR[14].XIC[7].icell.PDM VGND 0.18809f
C8149 XA.XIR[14].XIC[6].icell.PDM VGND 0.18809f
C8150 XA.XIR[14].XIC[5].icell.PDM VGND 0.18809f
C8151 XA.XIR[14].XIC[4].icell.PDM VGND 0.18809f
C8152 XA.XIR[14].XIC[3].icell.PDM VGND 0.18809f
C8153 XA.XIR[14].XIC[2].icell.PDM VGND 0.18809f
C8154 XA.XIR[14].XIC[1].icell.PDM VGND 0.18809f
C8155 XA.XIR[14].XIC[0].icell.PDM VGND 0.18817f
C8156 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C8157 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85795f
C8158 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C8159 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60802f
C8160 XA.XIR[13].XIC_15.icell.SM VGND 0.00474f
C8161 XA.XIR[13].XIC_dummy_right.icell.PUM VGND 0.00215f
C8162 XA.XIR[13].XIC_15.icell.Ien VGND 0.37063f
C8163 XA.XIR[13].XIC[14].icell.SM VGND 0.00502f
C8164 XA.XIR[13].XIC_15.icell.PUM VGND 0.00282f
C8165 XA.XIR[13].XIC[14].icell.Ien VGND 0.37144f
C8166 XA.XIR[13].XIC[13].icell.SM VGND 0.00502f
C8167 XA.XIR[13].XIC[14].icell.PUM VGND 0.00293f
C8168 XA.XIR[13].XIC[13].icell.Ien VGND 0.37144f
C8169 XA.XIR[13].XIC[12].icell.SM VGND 0.00502f
C8170 XA.XIR[13].XIC[13].icell.PUM VGND 0.00293f
C8171 XA.XIR[13].XIC[12].icell.Ien VGND 0.37144f
C8172 XA.XIR[13].XIC[11].icell.SM VGND 0.00502f
C8173 XA.XIR[13].XIC[12].icell.PUM VGND 0.00293f
C8174 XA.XIR[13].XIC[11].icell.Ien VGND 0.37144f
C8175 XA.XIR[13].XIC[10].icell.SM VGND 0.00502f
C8176 XA.XIR[13].XIC[11].icell.PUM VGND 0.00293f
C8177 XA.XIR[13].XIC[10].icell.Ien VGND 0.37144f
C8178 XA.XIR[13].XIC[9].icell.SM VGND 0.00502f
C8179 XA.XIR[13].XIC[10].icell.PUM VGND 0.00293f
C8180 XA.XIR[13].XIC[9].icell.Ien VGND 0.37144f
C8181 XA.XIR[13].XIC[8].icell.SM VGND 0.00502f
C8182 XA.XIR[13].XIC[9].icell.PUM VGND 0.00293f
C8183 XA.XIR[13].XIC[8].icell.Ien VGND 0.37144f
C8184 XA.XIR[13].XIC[7].icell.SM VGND 0.00502f
C8185 XA.XIR[13].XIC[8].icell.PUM VGND 0.00293f
C8186 XA.XIR[13].XIC[7].icell.Ien VGND 0.37144f
C8187 XA.XIR[13].XIC[6].icell.SM VGND 0.00502f
C8188 XA.XIR[13].XIC[7].icell.PUM VGND 0.00293f
C8189 XA.XIR[13].XIC[6].icell.Ien VGND 0.37144f
C8190 XA.XIR[13].XIC[5].icell.SM VGND 0.00502f
C8191 XA.XIR[13].XIC[6].icell.PUM VGND 0.00293f
C8192 XA.XIR[13].XIC[5].icell.Ien VGND 0.37144f
C8193 XA.XIR[13].XIC[4].icell.SM VGND 0.00502f
C8194 XA.XIR[13].XIC[5].icell.PUM VGND 0.00293f
C8195 XA.XIR[13].XIC[4].icell.Ien VGND 0.37144f
C8196 XA.XIR[13].XIC[3].icell.SM VGND 0.00502f
C8197 XA.XIR[13].XIC[4].icell.PUM VGND 0.00293f
C8198 XA.XIR[13].XIC[3].icell.Ien VGND 0.37144f
C8199 XA.XIR[13].XIC[2].icell.SM VGND 0.00502f
C8200 XA.XIR[13].XIC[3].icell.PUM VGND 0.00293f
C8201 XA.XIR[13].XIC[2].icell.Ien VGND 0.37144f
C8202 XA.XIR[13].XIC[1].icell.SM VGND 0.00502f
C8203 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.807f
C8204 XThR.Tn[13] VGND 14.01892f
C8205 XA.XIR[13].XIC[2].icell.PUM VGND 0.00293f
C8206 XA.XIR[13].XIC[1].icell.Ien VGND 0.37144f
C8207 XA.XIR[13].XIC[0].icell.SM VGND 0.00502f
C8208 XA.XIR[13].XIC[1].icell.PUM VGND 0.00293f
C8209 XA.XIR[13].XIC[0].icell.Ien VGND 0.37178f
C8210 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01044f
C8211 XA.XIR[13].XIC[0].icell.PUM VGND 0.00516f
C8212 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57425f
C8213 XA.XIR[13].XIC_dummy_left.icell.PUM VGND 0.00215f
C8214 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C8215 XA.XIR[13].XIC_15.icell.PDM VGND 0.18855f
C8216 XA.XIR[13].XIC[14].icell.PDM VGND 0.18809f
C8217 XA.XIR[13].XIC[13].icell.PDM VGND 0.18809f
C8218 XA.XIR[13].XIC[12].icell.PDM VGND 0.18809f
C8219 XA.XIR[13].XIC[11].icell.PDM VGND 0.18809f
C8220 XA.XIR[13].XIC[10].icell.PDM VGND 0.18809f
C8221 XA.XIR[13].XIC[9].icell.PDM VGND 0.18809f
C8222 XA.XIR[13].XIC[8].icell.PDM VGND 0.18809f
C8223 XA.XIR[13].XIC[7].icell.PDM VGND 0.18809f
C8224 XA.XIR[13].XIC[6].icell.PDM VGND 0.18809f
C8225 XA.XIR[13].XIC[5].icell.PDM VGND 0.18809f
C8226 XA.XIR[13].XIC[4].icell.PDM VGND 0.18809f
C8227 XA.XIR[13].XIC[3].icell.PDM VGND 0.18809f
C8228 XA.XIR[13].XIC[2].icell.PDM VGND 0.18809f
C8229 XA.XIR[13].XIC[1].icell.PDM VGND 0.18809f
C8230 XA.XIR[13].XIC[0].icell.PDM VGND 0.18817f
C8231 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C8232 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85795f
C8233 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C8234 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60802f
C8235 XA.XIR[12].XIC_15.icell.SM VGND 0.00474f
C8236 XA.XIR[12].XIC_dummy_right.icell.PUM VGND 0.00215f
C8237 XA.XIR[12].XIC_15.icell.Ien VGND 0.37063f
C8238 XA.XIR[12].XIC[14].icell.SM VGND 0.00502f
C8239 XA.XIR[12].XIC_15.icell.PUM VGND 0.00282f
C8240 XA.XIR[12].XIC[14].icell.Ien VGND 0.37144f
C8241 XA.XIR[12].XIC[13].icell.SM VGND 0.00502f
C8242 XA.XIR[12].XIC[14].icell.PUM VGND 0.00293f
C8243 XA.XIR[12].XIC[13].icell.Ien VGND 0.37144f
C8244 XA.XIR[12].XIC[12].icell.SM VGND 0.00502f
C8245 XA.XIR[12].XIC[13].icell.PUM VGND 0.00293f
C8246 XA.XIR[12].XIC[12].icell.Ien VGND 0.37144f
C8247 XA.XIR[12].XIC[11].icell.SM VGND 0.00502f
C8248 XA.XIR[12].XIC[12].icell.PUM VGND 0.00293f
C8249 XA.XIR[12].XIC[11].icell.Ien VGND 0.37144f
C8250 XA.XIR[12].XIC[10].icell.SM VGND 0.00502f
C8251 XA.XIR[12].XIC[11].icell.PUM VGND 0.00293f
C8252 XA.XIR[12].XIC[10].icell.Ien VGND 0.37144f
C8253 XA.XIR[12].XIC[9].icell.SM VGND 0.00502f
C8254 XA.XIR[12].XIC[10].icell.PUM VGND 0.00293f
C8255 XA.XIR[12].XIC[9].icell.Ien VGND 0.37144f
C8256 XA.XIR[12].XIC[8].icell.SM VGND 0.00502f
C8257 XA.XIR[12].XIC[9].icell.PUM VGND 0.00293f
C8258 XA.XIR[12].XIC[8].icell.Ien VGND 0.37144f
C8259 XA.XIR[12].XIC[7].icell.SM VGND 0.00502f
C8260 XA.XIR[12].XIC[8].icell.PUM VGND 0.00293f
C8261 XA.XIR[12].XIC[7].icell.Ien VGND 0.37144f
C8262 XA.XIR[12].XIC[6].icell.SM VGND 0.00502f
C8263 XA.XIR[12].XIC[7].icell.PUM VGND 0.00293f
C8264 XA.XIR[12].XIC[6].icell.Ien VGND 0.37144f
C8265 XA.XIR[12].XIC[5].icell.SM VGND 0.00502f
C8266 XA.XIR[12].XIC[6].icell.PUM VGND 0.00293f
C8267 XA.XIR[12].XIC[5].icell.Ien VGND 0.37144f
C8268 XA.XIR[12].XIC[4].icell.SM VGND 0.00502f
C8269 XA.XIR[12].XIC[5].icell.PUM VGND 0.00293f
C8270 XA.XIR[12].XIC[4].icell.Ien VGND 0.37144f
C8271 XA.XIR[12].XIC[3].icell.SM VGND 0.00502f
C8272 XA.XIR[12].XIC[4].icell.PUM VGND 0.00293f
C8273 XA.XIR[12].XIC[3].icell.Ien VGND 0.37144f
C8274 XA.XIR[12].XIC[2].icell.SM VGND 0.00502f
C8275 XA.XIR[12].XIC[3].icell.PUM VGND 0.00293f
C8276 XA.XIR[12].XIC[2].icell.Ien VGND 0.37144f
C8277 XA.XIR[12].XIC[1].icell.SM VGND 0.00502f
C8278 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80565f
C8279 XThR.Tn[12] VGND 13.90987f
C8280 XA.XIR[12].XIC[2].icell.PUM VGND 0.00293f
C8281 XA.XIR[12].XIC[1].icell.Ien VGND 0.37144f
C8282 XA.XIR[12].XIC[0].icell.SM VGND 0.00502f
C8283 XA.XIR[12].XIC[1].icell.PUM VGND 0.00293f
C8284 XA.XIR[12].XIC[0].icell.Ien VGND 0.37178f
C8285 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01044f
C8286 XA.XIR[12].XIC[0].icell.PUM VGND 0.00516f
C8287 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.57283f
C8288 XA.XIR[12].XIC_dummy_left.icell.PUM VGND 0.00215f
C8289 a_n997_2667# VGND 0.5457f
C8290 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C8291 XA.XIR[12].XIC_15.icell.PDM VGND 0.18855f
C8292 XA.XIR[12].XIC[14].icell.PDM VGND 0.18809f
C8293 XA.XIR[12].XIC[13].icell.PDM VGND 0.18809f
C8294 XA.XIR[12].XIC[12].icell.PDM VGND 0.18809f
C8295 XA.XIR[12].XIC[11].icell.PDM VGND 0.18809f
C8296 XA.XIR[12].XIC[10].icell.PDM VGND 0.18809f
C8297 XA.XIR[12].XIC[9].icell.PDM VGND 0.18809f
C8298 XA.XIR[12].XIC[8].icell.PDM VGND 0.18809f
C8299 XA.XIR[12].XIC[7].icell.PDM VGND 0.18809f
C8300 XA.XIR[12].XIC[6].icell.PDM VGND 0.18809f
C8301 XA.XIR[12].XIC[5].icell.PDM VGND 0.18809f
C8302 XA.XIR[12].XIC[4].icell.PDM VGND 0.18809f
C8303 XA.XIR[12].XIC[3].icell.PDM VGND 0.18809f
C8304 XA.XIR[12].XIC[2].icell.PDM VGND 0.18809f
C8305 XA.XIR[12].XIC[1].icell.PDM VGND 0.18809f
C8306 XA.XIR[12].XIC[0].icell.PDM VGND 0.18817f
C8307 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C8308 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85795f
C8309 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C8310 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60802f
C8311 XA.XIR[11].XIC_15.icell.SM VGND 0.00474f
C8312 XA.XIR[11].XIC_dummy_right.icell.PUM VGND 0.00215f
C8313 XA.XIR[11].XIC_15.icell.Ien VGND 0.37063f
C8314 XA.XIR[11].XIC[14].icell.SM VGND 0.00502f
C8315 XA.XIR[11].XIC_15.icell.PUM VGND 0.00282f
C8316 XA.XIR[11].XIC[14].icell.Ien VGND 0.37144f
C8317 XA.XIR[11].XIC[13].icell.SM VGND 0.00502f
C8318 XA.XIR[11].XIC[14].icell.PUM VGND 0.00293f
C8319 XA.XIR[11].XIC[13].icell.Ien VGND 0.37144f
C8320 XA.XIR[11].XIC[12].icell.SM VGND 0.00502f
C8321 XA.XIR[11].XIC[13].icell.PUM VGND 0.00293f
C8322 XA.XIR[11].XIC[12].icell.Ien VGND 0.37144f
C8323 XA.XIR[11].XIC[11].icell.SM VGND 0.00502f
C8324 XA.XIR[11].XIC[12].icell.PUM VGND 0.00293f
C8325 XA.XIR[11].XIC[11].icell.Ien VGND 0.37144f
C8326 XA.XIR[11].XIC[10].icell.SM VGND 0.00502f
C8327 XA.XIR[11].XIC[11].icell.PUM VGND 0.00293f
C8328 XA.XIR[11].XIC[10].icell.Ien VGND 0.37144f
C8329 XA.XIR[11].XIC[9].icell.SM VGND 0.00502f
C8330 XA.XIR[11].XIC[10].icell.PUM VGND 0.00293f
C8331 XA.XIR[11].XIC[9].icell.Ien VGND 0.37144f
C8332 XA.XIR[11].XIC[8].icell.SM VGND 0.00502f
C8333 XA.XIR[11].XIC[9].icell.PUM VGND 0.00293f
C8334 XA.XIR[11].XIC[8].icell.Ien VGND 0.37144f
C8335 XA.XIR[11].XIC[7].icell.SM VGND 0.00502f
C8336 XA.XIR[11].XIC[8].icell.PUM VGND 0.00293f
C8337 XA.XIR[11].XIC[7].icell.Ien VGND 0.37144f
C8338 XA.XIR[11].XIC[6].icell.SM VGND 0.00502f
C8339 XA.XIR[11].XIC[7].icell.PUM VGND 0.00293f
C8340 XA.XIR[11].XIC[6].icell.Ien VGND 0.37144f
C8341 XA.XIR[11].XIC[5].icell.SM VGND 0.00502f
C8342 XA.XIR[11].XIC[6].icell.PUM VGND 0.00293f
C8343 XA.XIR[11].XIC[5].icell.Ien VGND 0.37144f
C8344 XA.XIR[11].XIC[4].icell.SM VGND 0.00502f
C8345 XA.XIR[11].XIC[5].icell.PUM VGND 0.00293f
C8346 XA.XIR[11].XIC[4].icell.Ien VGND 0.37144f
C8347 XA.XIR[11].XIC[3].icell.SM VGND 0.00502f
C8348 XA.XIR[11].XIC[4].icell.PUM VGND 0.00293f
C8349 XA.XIR[11].XIC[3].icell.Ien VGND 0.37144f
C8350 XA.XIR[11].XIC[2].icell.SM VGND 0.00502f
C8351 XA.XIR[11].XIC[3].icell.PUM VGND 0.00293f
C8352 XA.XIR[11].XIC[2].icell.Ien VGND 0.37144f
C8353 XA.XIR[11].XIC[1].icell.SM VGND 0.00502f
C8354 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.808f
C8355 XThR.Tn[11] VGND 13.97038f
C8356 XA.XIR[11].XIC[2].icell.PUM VGND 0.00293f
C8357 XA.XIR[11].XIC[1].icell.Ien VGND 0.37144f
C8358 XA.XIR[11].XIC[0].icell.SM VGND 0.00502f
C8359 a_n997_2891# VGND 0.54795f
C8360 a_n1331_2891# VGND 0.00194f
C8361 XA.XIR[11].XIC[1].icell.PUM VGND 0.00293f
C8362 XA.XIR[11].XIC[0].icell.Ien VGND 0.37178f
C8363 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01044f
C8364 XA.XIR[11].XIC[0].icell.PUM VGND 0.00516f
C8365 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57297f
C8366 XA.XIR[11].XIC_dummy_left.icell.PUM VGND 0.00215f
C8367 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C8368 XA.XIR[11].XIC_15.icell.PDM VGND 0.18855f
C8369 XA.XIR[11].XIC[14].icell.PDM VGND 0.18809f
C8370 XA.XIR[11].XIC[13].icell.PDM VGND 0.18809f
C8371 XA.XIR[11].XIC[12].icell.PDM VGND 0.18809f
C8372 XA.XIR[11].XIC[11].icell.PDM VGND 0.18809f
C8373 XA.XIR[11].XIC[10].icell.PDM VGND 0.18809f
C8374 XA.XIR[11].XIC[9].icell.PDM VGND 0.18809f
C8375 XA.XIR[11].XIC[8].icell.PDM VGND 0.18809f
C8376 XA.XIR[11].XIC[7].icell.PDM VGND 0.18809f
C8377 XA.XIR[11].XIC[6].icell.PDM VGND 0.18809f
C8378 XA.XIR[11].XIC[5].icell.PDM VGND 0.18809f
C8379 XA.XIR[11].XIC[4].icell.PDM VGND 0.18809f
C8380 XA.XIR[11].XIC[3].icell.PDM VGND 0.18809f
C8381 XA.XIR[11].XIC[2].icell.PDM VGND 0.18809f
C8382 XA.XIR[11].XIC[1].icell.PDM VGND 0.18809f
C8383 XA.XIR[11].XIC[0].icell.PDM VGND 0.18817f
C8384 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C8385 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85795f
C8386 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C8387 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60802f
C8388 XA.XIR[10].XIC_15.icell.SM VGND 0.00474f
C8389 XA.XIR[10].XIC_dummy_right.icell.PUM VGND 0.00215f
C8390 XA.XIR[10].XIC_15.icell.Ien VGND 0.37063f
C8391 XA.XIR[10].XIC[14].icell.SM VGND 0.00502f
C8392 XA.XIR[10].XIC_15.icell.PUM VGND 0.00282f
C8393 XA.XIR[10].XIC[14].icell.Ien VGND 0.37144f
C8394 XA.XIR[10].XIC[13].icell.SM VGND 0.00502f
C8395 XA.XIR[10].XIC[14].icell.PUM VGND 0.00293f
C8396 XA.XIR[10].XIC[13].icell.Ien VGND 0.37144f
C8397 XA.XIR[10].XIC[12].icell.SM VGND 0.00502f
C8398 XA.XIR[10].XIC[13].icell.PUM VGND 0.00293f
C8399 XA.XIR[10].XIC[12].icell.Ien VGND 0.37144f
C8400 XA.XIR[10].XIC[11].icell.SM VGND 0.00502f
C8401 XA.XIR[10].XIC[12].icell.PUM VGND 0.00293f
C8402 XA.XIR[10].XIC[11].icell.Ien VGND 0.37144f
C8403 XA.XIR[10].XIC[10].icell.SM VGND 0.00502f
C8404 XA.XIR[10].XIC[11].icell.PUM VGND 0.00293f
C8405 XA.XIR[10].XIC[10].icell.Ien VGND 0.37144f
C8406 XA.XIR[10].XIC[9].icell.SM VGND 0.00502f
C8407 XA.XIR[10].XIC[10].icell.PUM VGND 0.00293f
C8408 XA.XIR[10].XIC[9].icell.Ien VGND 0.37144f
C8409 XA.XIR[10].XIC[8].icell.SM VGND 0.00502f
C8410 XA.XIR[10].XIC[9].icell.PUM VGND 0.00293f
C8411 XA.XIR[10].XIC[8].icell.Ien VGND 0.37144f
C8412 XA.XIR[10].XIC[7].icell.SM VGND 0.00502f
C8413 XA.XIR[10].XIC[8].icell.PUM VGND 0.00293f
C8414 XA.XIR[10].XIC[7].icell.Ien VGND 0.37144f
C8415 XA.XIR[10].XIC[6].icell.SM VGND 0.00502f
C8416 XA.XIR[10].XIC[7].icell.PUM VGND 0.00293f
C8417 XA.XIR[10].XIC[6].icell.Ien VGND 0.37144f
C8418 XA.XIR[10].XIC[5].icell.SM VGND 0.00502f
C8419 XA.XIR[10].XIC[6].icell.PUM VGND 0.00293f
C8420 XA.XIR[10].XIC[5].icell.Ien VGND 0.37144f
C8421 XA.XIR[10].XIC[4].icell.SM VGND 0.00502f
C8422 XA.XIR[10].XIC[5].icell.PUM VGND 0.00293f
C8423 XA.XIR[10].XIC[4].icell.Ien VGND 0.37144f
C8424 XA.XIR[10].XIC[3].icell.SM VGND 0.00502f
C8425 XA.XIR[10].XIC[4].icell.PUM VGND 0.00293f
C8426 XA.XIR[10].XIC[3].icell.Ien VGND 0.37144f
C8427 XA.XIR[10].XIC[2].icell.SM VGND 0.00502f
C8428 XA.XIR[10].XIC[3].icell.PUM VGND 0.00293f
C8429 XA.XIR[10].XIC[2].icell.Ien VGND 0.37144f
C8430 XA.XIR[10].XIC[1].icell.SM VGND 0.00502f
C8431 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80684f
C8432 XThR.Tn[10] VGND 13.91105f
C8433 XA.XIR[10].XIC[2].icell.PUM VGND 0.00293f
C8434 XA.XIR[10].XIC[1].icell.Ien VGND 0.37144f
C8435 XA.XIR[10].XIC[0].icell.SM VGND 0.00502f
C8436 XA.XIR[10].XIC[1].icell.PUM VGND 0.00293f
C8437 XA.XIR[10].XIC[0].icell.Ien VGND 0.37178f
C8438 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01044f
C8439 XA.XIR[10].XIC[0].icell.PUM VGND 0.00516f
C8440 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57425f
C8441 XA.XIR[10].XIC_dummy_left.icell.PUM VGND 0.00215f
C8442 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C8443 XA.XIR[10].XIC_15.icell.PDM VGND 0.18855f
C8444 XA.XIR[10].XIC[14].icell.PDM VGND 0.18809f
C8445 XA.XIR[10].XIC[13].icell.PDM VGND 0.18809f
C8446 XA.XIR[10].XIC[12].icell.PDM VGND 0.18809f
C8447 XA.XIR[10].XIC[11].icell.PDM VGND 0.18809f
C8448 XA.XIR[10].XIC[10].icell.PDM VGND 0.18809f
C8449 XA.XIR[10].XIC[9].icell.PDM VGND 0.18809f
C8450 XA.XIR[10].XIC[8].icell.PDM VGND 0.18809f
C8451 XA.XIR[10].XIC[7].icell.PDM VGND 0.18809f
C8452 XA.XIR[10].XIC[6].icell.PDM VGND 0.18809f
C8453 XA.XIR[10].XIC[5].icell.PDM VGND 0.18809f
C8454 XA.XIR[10].XIC[4].icell.PDM VGND 0.18809f
C8455 XA.XIR[10].XIC[3].icell.PDM VGND 0.18809f
C8456 XA.XIR[10].XIC[2].icell.PDM VGND 0.18809f
C8457 XA.XIR[10].XIC[1].icell.PDM VGND 0.18809f
C8458 XA.XIR[10].XIC[0].icell.PDM VGND 0.18817f
C8459 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C8460 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85795f
C8461 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C8462 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60802f
C8463 XA.XIR[9].XIC_15.icell.SM VGND 0.00474f
C8464 XA.XIR[9].XIC_dummy_right.icell.PUM VGND 0.00215f
C8465 XA.XIR[9].XIC_15.icell.Ien VGND 0.37063f
C8466 XA.XIR[9].XIC[14].icell.SM VGND 0.00502f
C8467 XA.XIR[9].XIC_15.icell.PUM VGND 0.00282f
C8468 XA.XIR[9].XIC[14].icell.Ien VGND 0.37144f
C8469 XA.XIR[9].XIC[13].icell.SM VGND 0.00502f
C8470 XA.XIR[9].XIC[14].icell.PUM VGND 0.00293f
C8471 XA.XIR[9].XIC[13].icell.Ien VGND 0.37144f
C8472 XA.XIR[9].XIC[12].icell.SM VGND 0.00502f
C8473 XA.XIR[9].XIC[13].icell.PUM VGND 0.00293f
C8474 XA.XIR[9].XIC[12].icell.Ien VGND 0.37144f
C8475 XA.XIR[9].XIC[11].icell.SM VGND 0.00502f
C8476 XA.XIR[9].XIC[12].icell.PUM VGND 0.00293f
C8477 XA.XIR[9].XIC[11].icell.Ien VGND 0.37144f
C8478 XA.XIR[9].XIC[10].icell.SM VGND 0.00502f
C8479 XA.XIR[9].XIC[11].icell.PUM VGND 0.00293f
C8480 XA.XIR[9].XIC[10].icell.Ien VGND 0.37144f
C8481 XA.XIR[9].XIC[9].icell.SM VGND 0.00502f
C8482 XA.XIR[9].XIC[10].icell.PUM VGND 0.00293f
C8483 XA.XIR[9].XIC[9].icell.Ien VGND 0.37144f
C8484 XA.XIR[9].XIC[8].icell.SM VGND 0.00502f
C8485 XA.XIR[9].XIC[9].icell.PUM VGND 0.00293f
C8486 XA.XIR[9].XIC[8].icell.Ien VGND 0.37144f
C8487 XA.XIR[9].XIC[7].icell.SM VGND 0.00502f
C8488 XA.XIR[9].XIC[8].icell.PUM VGND 0.00293f
C8489 XA.XIR[9].XIC[7].icell.Ien VGND 0.37144f
C8490 XA.XIR[9].XIC[6].icell.SM VGND 0.00502f
C8491 XA.XIR[9].XIC[7].icell.PUM VGND 0.00293f
C8492 XA.XIR[9].XIC[6].icell.Ien VGND 0.37144f
C8493 XA.XIR[9].XIC[5].icell.SM VGND 0.00502f
C8494 XA.XIR[9].XIC[6].icell.PUM VGND 0.00293f
C8495 XA.XIR[9].XIC[5].icell.Ien VGND 0.37144f
C8496 XA.XIR[9].XIC[4].icell.SM VGND 0.00502f
C8497 XA.XIR[9].XIC[5].icell.PUM VGND 0.00293f
C8498 XA.XIR[9].XIC[4].icell.Ien VGND 0.37144f
C8499 XA.XIR[9].XIC[3].icell.SM VGND 0.00502f
C8500 XA.XIR[9].XIC[4].icell.PUM VGND 0.00293f
C8501 XA.XIR[9].XIC[3].icell.Ien VGND 0.37144f
C8502 XA.XIR[9].XIC[2].icell.SM VGND 0.00502f
C8503 XA.XIR[9].XIC[3].icell.PUM VGND 0.00293f
C8504 XA.XIR[9].XIC[2].icell.Ien VGND 0.37144f
C8505 XA.XIR[9].XIC[1].icell.SM VGND 0.00502f
C8506 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.8087f
C8507 XA.XIR[9].XIC[2].icell.PUM VGND 0.00293f
C8508 XA.XIR[9].XIC[1].icell.Ien VGND 0.37144f
C8509 XA.XIR[9].XIC[0].icell.SM VGND 0.00502f
C8510 XThR.Tn[9] VGND 13.95272f
C8511 a_n997_3755# VGND 0.54861f
C8512 XA.XIR[9].XIC[1].icell.PUM VGND 0.00293f
C8513 XA.XIR[9].XIC[0].icell.Ien VGND 0.37178f
C8514 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01044f
C8515 XA.XIR[9].XIC[0].icell.PUM VGND 0.00516f
C8516 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.57323f
C8517 a_n997_3979# VGND 0.54721f
C8518 XA.XIR[9].XIC_dummy_left.icell.PUM VGND 0.00215f
C8519 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C8520 XA.XIR[9].XIC_15.icell.PDM VGND 0.18855f
C8521 XA.XIR[9].XIC[14].icell.PDM VGND 0.18809f
C8522 XA.XIR[9].XIC[13].icell.PDM VGND 0.18809f
C8523 XA.XIR[9].XIC[12].icell.PDM VGND 0.18809f
C8524 XA.XIR[9].XIC[11].icell.PDM VGND 0.18809f
C8525 XA.XIR[9].XIC[10].icell.PDM VGND 0.18809f
C8526 XA.XIR[9].XIC[9].icell.PDM VGND 0.18809f
C8527 XA.XIR[9].XIC[8].icell.PDM VGND 0.18809f
C8528 XA.XIR[9].XIC[7].icell.PDM VGND 0.18809f
C8529 XA.XIR[9].XIC[6].icell.PDM VGND 0.18809f
C8530 XA.XIR[9].XIC[5].icell.PDM VGND 0.18809f
C8531 XA.XIR[9].XIC[4].icell.PDM VGND 0.18809f
C8532 XA.XIR[9].XIC[3].icell.PDM VGND 0.18809f
C8533 XA.XIR[9].XIC[2].icell.PDM VGND 0.18809f
C8534 XA.XIR[9].XIC[1].icell.PDM VGND 0.18809f
C8535 XA.XIR[9].XIC[0].icell.PDM VGND 0.18817f
C8536 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C8537 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85795f
C8538 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C8539 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60802f
C8540 XA.XIR[8].XIC_15.icell.SM VGND 0.00474f
C8541 XA.XIR[8].XIC_dummy_right.icell.PUM VGND 0.00215f
C8542 XA.XIR[8].XIC_15.icell.Ien VGND 0.37063f
C8543 XA.XIR[8].XIC[14].icell.SM VGND 0.00502f
C8544 XA.XIR[8].XIC_15.icell.PUM VGND 0.00282f
C8545 XA.XIR[8].XIC[14].icell.Ien VGND 0.37144f
C8546 XA.XIR[8].XIC[13].icell.SM VGND 0.00502f
C8547 XA.XIR[8].XIC[14].icell.PUM VGND 0.00293f
C8548 XA.XIR[8].XIC[13].icell.Ien VGND 0.37144f
C8549 XA.XIR[8].XIC[12].icell.SM VGND 0.00502f
C8550 XA.XIR[8].XIC[13].icell.PUM VGND 0.00293f
C8551 XA.XIR[8].XIC[12].icell.Ien VGND 0.37144f
C8552 XA.XIR[8].XIC[11].icell.SM VGND 0.00502f
C8553 XA.XIR[8].XIC[12].icell.PUM VGND 0.00293f
C8554 XA.XIR[8].XIC[11].icell.Ien VGND 0.37144f
C8555 XA.XIR[8].XIC[10].icell.SM VGND 0.00502f
C8556 XA.XIR[8].XIC[11].icell.PUM VGND 0.00293f
C8557 XA.XIR[8].XIC[10].icell.Ien VGND 0.37144f
C8558 XA.XIR[8].XIC[9].icell.SM VGND 0.00502f
C8559 XA.XIR[8].XIC[10].icell.PUM VGND 0.00293f
C8560 XA.XIR[8].XIC[9].icell.Ien VGND 0.37144f
C8561 XA.XIR[8].XIC[8].icell.SM VGND 0.00502f
C8562 XA.XIR[8].XIC[9].icell.PUM VGND 0.00293f
C8563 XA.XIR[8].XIC[8].icell.Ien VGND 0.37144f
C8564 XA.XIR[8].XIC[7].icell.SM VGND 0.00502f
C8565 XA.XIR[8].XIC[8].icell.PUM VGND 0.00293f
C8566 XA.XIR[8].XIC[7].icell.Ien VGND 0.37144f
C8567 XA.XIR[8].XIC[6].icell.SM VGND 0.00502f
C8568 XA.XIR[8].XIC[7].icell.PUM VGND 0.00293f
C8569 XA.XIR[8].XIC[6].icell.Ien VGND 0.37144f
C8570 XA.XIR[8].XIC[5].icell.SM VGND 0.00502f
C8571 XA.XIR[8].XIC[6].icell.PUM VGND 0.00293f
C8572 XA.XIR[8].XIC[5].icell.Ien VGND 0.37144f
C8573 XA.XIR[8].XIC[4].icell.SM VGND 0.00502f
C8574 XA.XIR[8].XIC[5].icell.PUM VGND 0.00293f
C8575 XA.XIR[8].XIC[4].icell.Ien VGND 0.37144f
C8576 XA.XIR[8].XIC[3].icell.SM VGND 0.00502f
C8577 XA.XIR[8].XIC[4].icell.PUM VGND 0.00293f
C8578 XA.XIR[8].XIC[3].icell.Ien VGND 0.37144f
C8579 XA.XIR[8].XIC[2].icell.SM VGND 0.00502f
C8580 XA.XIR[8].XIC[3].icell.PUM VGND 0.00293f
C8581 XA.XIR[8].XIC[2].icell.Ien VGND 0.37144f
C8582 XA.XIR[8].XIC[1].icell.SM VGND 0.00502f
C8583 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80602f
C8584 XA.XIR[8].XIC[2].icell.PUM VGND 0.00293f
C8585 XA.XIR[8].XIC[1].icell.Ien VGND 0.37144f
C8586 XA.XIR[8].XIC[0].icell.SM VGND 0.00502f
C8587 XThR.Tn[8] VGND 13.89711f
C8588 XA.XIR[8].XIC[1].icell.PUM VGND 0.00293f
C8589 XA.XIR[8].XIC[0].icell.Ien VGND 0.37178f
C8590 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01044f
C8591 XA.XIR[8].XIC[0].icell.PUM VGND 0.00516f
C8592 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57311f
C8593 XA.XIR[8].XIC_dummy_left.icell.PUM VGND 0.00215f
C8594 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C8595 XA.XIR[8].XIC_15.icell.PDM VGND 0.18855f
C8596 XA.XIR[8].XIC[14].icell.PDM VGND 0.18809f
C8597 XA.XIR[8].XIC[13].icell.PDM VGND 0.18809f
C8598 XA.XIR[8].XIC[12].icell.PDM VGND 0.18809f
C8599 XA.XIR[8].XIC[11].icell.PDM VGND 0.18809f
C8600 XA.XIR[8].XIC[10].icell.PDM VGND 0.18809f
C8601 XA.XIR[8].XIC[9].icell.PDM VGND 0.18809f
C8602 XA.XIR[8].XIC[8].icell.PDM VGND 0.18809f
C8603 XA.XIR[8].XIC[7].icell.PDM VGND 0.18809f
C8604 XA.XIR[8].XIC[6].icell.PDM VGND 0.18809f
C8605 XA.XIR[8].XIC[5].icell.PDM VGND 0.18809f
C8606 XA.XIR[8].XIC[4].icell.PDM VGND 0.18809f
C8607 XA.XIR[8].XIC[3].icell.PDM VGND 0.18809f
C8608 XA.XIR[8].XIC[2].icell.PDM VGND 0.18809f
C8609 XA.XIR[8].XIC[1].icell.PDM VGND 0.18809f
C8610 XA.XIR[8].XIC[0].icell.PDM VGND 0.18817f
C8611 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C8612 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85795f
C8613 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C8614 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60802f
C8615 XA.XIR[7].XIC_15.icell.SM VGND 0.00474f
C8616 XA.XIR[7].XIC_dummy_right.icell.PUM VGND 0.00215f
C8617 XA.XIR[7].XIC_15.icell.Ien VGND 0.37063f
C8618 XA.XIR[7].XIC[14].icell.SM VGND 0.00502f
C8619 XA.XIR[7].XIC_15.icell.PUM VGND 0.00282f
C8620 XA.XIR[7].XIC[14].icell.Ien VGND 0.37144f
C8621 XA.XIR[7].XIC[13].icell.SM VGND 0.00502f
C8622 XA.XIR[7].XIC[14].icell.PUM VGND 0.00293f
C8623 XA.XIR[7].XIC[13].icell.Ien VGND 0.37144f
C8624 XA.XIR[7].XIC[12].icell.SM VGND 0.00502f
C8625 XA.XIR[7].XIC[13].icell.PUM VGND 0.00293f
C8626 XA.XIR[7].XIC[12].icell.Ien VGND 0.37144f
C8627 XA.XIR[7].XIC[11].icell.SM VGND 0.00502f
C8628 XA.XIR[7].XIC[12].icell.PUM VGND 0.00293f
C8629 XA.XIR[7].XIC[11].icell.Ien VGND 0.37144f
C8630 XA.XIR[7].XIC[10].icell.SM VGND 0.00502f
C8631 XA.XIR[7].XIC[11].icell.PUM VGND 0.00293f
C8632 XA.XIR[7].XIC[10].icell.Ien VGND 0.37144f
C8633 XA.XIR[7].XIC[9].icell.SM VGND 0.00502f
C8634 XA.XIR[7].XIC[10].icell.PUM VGND 0.00293f
C8635 XA.XIR[7].XIC[9].icell.Ien VGND 0.37144f
C8636 XA.XIR[7].XIC[8].icell.SM VGND 0.00502f
C8637 XA.XIR[7].XIC[9].icell.PUM VGND 0.00293f
C8638 XA.XIR[7].XIC[8].icell.Ien VGND 0.37144f
C8639 XA.XIR[7].XIC[7].icell.SM VGND 0.00502f
C8640 XA.XIR[7].XIC[8].icell.PUM VGND 0.00293f
C8641 XA.XIR[7].XIC[7].icell.Ien VGND 0.37144f
C8642 XA.XIR[7].XIC[6].icell.SM VGND 0.00502f
C8643 XA.XIR[7].XIC[7].icell.PUM VGND 0.00293f
C8644 XA.XIR[7].XIC[6].icell.Ien VGND 0.37144f
C8645 XA.XIR[7].XIC[5].icell.SM VGND 0.00502f
C8646 XA.XIR[7].XIC[6].icell.PUM VGND 0.00293f
C8647 XA.XIR[7].XIC[5].icell.Ien VGND 0.37144f
C8648 XA.XIR[7].XIC[4].icell.SM VGND 0.00502f
C8649 XA.XIR[7].XIC[5].icell.PUM VGND 0.00293f
C8650 XA.XIR[7].XIC[4].icell.Ien VGND 0.37144f
C8651 XA.XIR[7].XIC[3].icell.SM VGND 0.00502f
C8652 XA.XIR[7].XIC[4].icell.PUM VGND 0.00293f
C8653 XA.XIR[7].XIC[3].icell.Ien VGND 0.37144f
C8654 XA.XIR[7].XIC[2].icell.SM VGND 0.00502f
C8655 XA.XIR[7].XIC[3].icell.PUM VGND 0.00293f
C8656 XA.XIR[7].XIC[2].icell.Ien VGND 0.37144f
C8657 XA.XIR[7].XIC[1].icell.SM VGND 0.00502f
C8658 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80634f
C8659 XA.XIR[7].XIC[2].icell.PUM VGND 0.00293f
C8660 XA.XIR[7].XIC[1].icell.Ien VGND 0.37144f
C8661 XA.XIR[7].XIC[0].icell.SM VGND 0.00502f
C8662 XA.XIR[7].XIC[1].icell.PUM VGND 0.00293f
C8663 XA.XIR[7].XIC[0].icell.Ien VGND 0.37178f
C8664 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01044f
C8665 XThR.Tn[7] VGND 14.38144f
C8666 XThR.TAN2 VGND 1.22814f
C8667 XA.XIR[7].XIC[0].icell.PUM VGND 0.00516f
C8668 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57579f
C8669 XA.XIR[7].XIC_dummy_left.icell.PUM VGND 0.00222f
C8670 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C8671 XA.XIR[7].XIC_15.icell.PDM VGND 0.18855f
C8672 XA.XIR[7].XIC[14].icell.PDM VGND 0.18809f
C8673 XA.XIR[7].XIC[13].icell.PDM VGND 0.18809f
C8674 XA.XIR[7].XIC[12].icell.PDM VGND 0.18809f
C8675 XA.XIR[7].XIC[11].icell.PDM VGND 0.18809f
C8676 XA.XIR[7].XIC[10].icell.PDM VGND 0.18809f
C8677 XA.XIR[7].XIC[9].icell.PDM VGND 0.18809f
C8678 XA.XIR[7].XIC[8].icell.PDM VGND 0.18809f
C8679 XA.XIR[7].XIC[7].icell.PDM VGND 0.18809f
C8680 XA.XIR[7].XIC[6].icell.PDM VGND 0.18809f
C8681 XA.XIR[7].XIC[5].icell.PDM VGND 0.18809f
C8682 XA.XIR[7].XIC[4].icell.PDM VGND 0.18809f
C8683 XA.XIR[7].XIC[3].icell.PDM VGND 0.18809f
C8684 XA.XIR[7].XIC[2].icell.PDM VGND 0.18809f
C8685 XA.XIR[7].XIC[1].icell.PDM VGND 0.18809f
C8686 XA.XIR[7].XIC[0].icell.PDM VGND 0.18817f
C8687 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C8688 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85795f
C8689 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C8690 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60802f
C8691 XA.XIR[6].XIC_15.icell.SM VGND 0.00474f
C8692 XA.XIR[6].XIC_dummy_right.icell.PUM VGND 0.00215f
C8693 XA.XIR[6].XIC_15.icell.Ien VGND 0.37063f
C8694 XA.XIR[6].XIC[14].icell.SM VGND 0.00502f
C8695 XA.XIR[6].XIC_15.icell.PUM VGND 0.00282f
C8696 XA.XIR[6].XIC[14].icell.Ien VGND 0.37144f
C8697 XA.XIR[6].XIC[13].icell.SM VGND 0.00502f
C8698 XA.XIR[6].XIC[14].icell.PUM VGND 0.00293f
C8699 XA.XIR[6].XIC[13].icell.Ien VGND 0.37144f
C8700 XA.XIR[6].XIC[12].icell.SM VGND 0.00502f
C8701 XA.XIR[6].XIC[13].icell.PUM VGND 0.00293f
C8702 XA.XIR[6].XIC[12].icell.Ien VGND 0.37144f
C8703 XA.XIR[6].XIC[11].icell.SM VGND 0.00502f
C8704 XA.XIR[6].XIC[12].icell.PUM VGND 0.00293f
C8705 XA.XIR[6].XIC[11].icell.Ien VGND 0.37144f
C8706 XA.XIR[6].XIC[10].icell.SM VGND 0.00502f
C8707 XA.XIR[6].XIC[11].icell.PUM VGND 0.00293f
C8708 XA.XIR[6].XIC[10].icell.Ien VGND 0.37144f
C8709 XA.XIR[6].XIC[9].icell.SM VGND 0.00502f
C8710 XA.XIR[6].XIC[10].icell.PUM VGND 0.00293f
C8711 XA.XIR[6].XIC[9].icell.Ien VGND 0.37144f
C8712 XA.XIR[6].XIC[8].icell.SM VGND 0.00502f
C8713 XA.XIR[6].XIC[9].icell.PUM VGND 0.00293f
C8714 XA.XIR[6].XIC[8].icell.Ien VGND 0.37144f
C8715 XA.XIR[6].XIC[7].icell.SM VGND 0.00502f
C8716 XA.XIR[6].XIC[8].icell.PUM VGND 0.00293f
C8717 XA.XIR[6].XIC[7].icell.Ien VGND 0.37144f
C8718 XA.XIR[6].XIC[6].icell.SM VGND 0.00502f
C8719 XA.XIR[6].XIC[7].icell.PUM VGND 0.00293f
C8720 XA.XIR[6].XIC[6].icell.Ien VGND 0.37144f
C8721 XA.XIR[6].XIC[5].icell.SM VGND 0.00502f
C8722 XA.XIR[6].XIC[6].icell.PUM VGND 0.00293f
C8723 XA.XIR[6].XIC[5].icell.Ien VGND 0.37144f
C8724 XA.XIR[6].XIC[4].icell.SM VGND 0.00502f
C8725 XA.XIR[6].XIC[5].icell.PUM VGND 0.00293f
C8726 XA.XIR[6].XIC[4].icell.Ien VGND 0.37144f
C8727 XA.XIR[6].XIC[3].icell.SM VGND 0.00502f
C8728 XA.XIR[6].XIC[4].icell.PUM VGND 0.00293f
C8729 XA.XIR[6].XIC[3].icell.Ien VGND 0.37144f
C8730 XA.XIR[6].XIC[2].icell.SM VGND 0.00502f
C8731 XA.XIR[6].XIC[3].icell.PUM VGND 0.00293f
C8732 XA.XIR[6].XIC[2].icell.Ien VGND 0.37144f
C8733 XA.XIR[6].XIC[1].icell.SM VGND 0.00502f
C8734 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80729f
C8735 XA.XIR[6].XIC[2].icell.PUM VGND 0.00293f
C8736 XA.XIR[6].XIC[1].icell.Ien VGND 0.37144f
C8737 XA.XIR[6].XIC[0].icell.SM VGND 0.00502f
C8738 XA.XIR[6].XIC[1].icell.PUM VGND 0.00293f
C8739 XA.XIR[6].XIC[0].icell.Ien VGND 0.37178f
C8740 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01044f
C8741 XA.XIR[6].XIC[0].icell.PUM VGND 0.00516f
C8742 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57425f
C8743 XThR.Tn[6] VGND 13.98754f
C8744 a_n1049_5317# VGND 0.02283f
C8745 XA.XIR[6].XIC_dummy_left.icell.PUM VGND 0.00215f
C8746 XThR.TB7 VGND 1.36132f
C8747 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C8748 XA.XIR[6].XIC_15.icell.PDM VGND 0.18855f
C8749 XA.XIR[6].XIC[14].icell.PDM VGND 0.18809f
C8750 XA.XIR[6].XIC[13].icell.PDM VGND 0.18809f
C8751 XA.XIR[6].XIC[12].icell.PDM VGND 0.18809f
C8752 XA.XIR[6].XIC[11].icell.PDM VGND 0.18809f
C8753 XA.XIR[6].XIC[10].icell.PDM VGND 0.18809f
C8754 XA.XIR[6].XIC[9].icell.PDM VGND 0.18809f
C8755 XA.XIR[6].XIC[8].icell.PDM VGND 0.18809f
C8756 XA.XIR[6].XIC[7].icell.PDM VGND 0.18809f
C8757 XA.XIR[6].XIC[6].icell.PDM VGND 0.18809f
C8758 XA.XIR[6].XIC[5].icell.PDM VGND 0.18809f
C8759 XA.XIR[6].XIC[4].icell.PDM VGND 0.18809f
C8760 XA.XIR[6].XIC[3].icell.PDM VGND 0.18809f
C8761 XA.XIR[6].XIC[2].icell.PDM VGND 0.18809f
C8762 XA.XIR[6].XIC[1].icell.PDM VGND 0.18809f
C8763 XA.XIR[6].XIC[0].icell.PDM VGND 0.18817f
C8764 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C8765 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85795f
C8766 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C8767 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60802f
C8768 XA.XIR[5].XIC_15.icell.SM VGND 0.00474f
C8769 XA.XIR[5].XIC_dummy_right.icell.PUM VGND 0.00215f
C8770 XA.XIR[5].XIC_15.icell.Ien VGND 0.37063f
C8771 XA.XIR[5].XIC[14].icell.SM VGND 0.00502f
C8772 XA.XIR[5].XIC_15.icell.PUM VGND 0.00282f
C8773 XA.XIR[5].XIC[14].icell.Ien VGND 0.37144f
C8774 XA.XIR[5].XIC[13].icell.SM VGND 0.00502f
C8775 XA.XIR[5].XIC[14].icell.PUM VGND 0.00293f
C8776 XA.XIR[5].XIC[13].icell.Ien VGND 0.37144f
C8777 XA.XIR[5].XIC[12].icell.SM VGND 0.00502f
C8778 XA.XIR[5].XIC[13].icell.PUM VGND 0.00293f
C8779 XA.XIR[5].XIC[12].icell.Ien VGND 0.37144f
C8780 XA.XIR[5].XIC[11].icell.SM VGND 0.00502f
C8781 XA.XIR[5].XIC[12].icell.PUM VGND 0.00293f
C8782 XA.XIR[5].XIC[11].icell.Ien VGND 0.37144f
C8783 XA.XIR[5].XIC[10].icell.SM VGND 0.00502f
C8784 XA.XIR[5].XIC[11].icell.PUM VGND 0.00293f
C8785 XA.XIR[5].XIC[10].icell.Ien VGND 0.37144f
C8786 XA.XIR[5].XIC[9].icell.SM VGND 0.00502f
C8787 XA.XIR[5].XIC[10].icell.PUM VGND 0.00293f
C8788 XA.XIR[5].XIC[9].icell.Ien VGND 0.37144f
C8789 XA.XIR[5].XIC[8].icell.SM VGND 0.00502f
C8790 XA.XIR[5].XIC[9].icell.PUM VGND 0.00293f
C8791 XA.XIR[5].XIC[8].icell.Ien VGND 0.37144f
C8792 XA.XIR[5].XIC[7].icell.SM VGND 0.00502f
C8793 XA.XIR[5].XIC[8].icell.PUM VGND 0.00293f
C8794 XA.XIR[5].XIC[7].icell.Ien VGND 0.37144f
C8795 XA.XIR[5].XIC[6].icell.SM VGND 0.00502f
C8796 XA.XIR[5].XIC[7].icell.PUM VGND 0.00293f
C8797 XA.XIR[5].XIC[6].icell.Ien VGND 0.37144f
C8798 XA.XIR[5].XIC[5].icell.SM VGND 0.00502f
C8799 XA.XIR[5].XIC[6].icell.PUM VGND 0.00293f
C8800 XA.XIR[5].XIC[5].icell.Ien VGND 0.37144f
C8801 XA.XIR[5].XIC[4].icell.SM VGND 0.00502f
C8802 XA.XIR[5].XIC[5].icell.PUM VGND 0.00293f
C8803 XA.XIR[5].XIC[4].icell.Ien VGND 0.37144f
C8804 XA.XIR[5].XIC[3].icell.SM VGND 0.00502f
C8805 XA.XIR[5].XIC[4].icell.PUM VGND 0.00293f
C8806 XA.XIR[5].XIC[3].icell.Ien VGND 0.37144f
C8807 XA.XIR[5].XIC[2].icell.SM VGND 0.00502f
C8808 XA.XIR[5].XIC[3].icell.PUM VGND 0.00293f
C8809 XA.XIR[5].XIC[2].icell.Ien VGND 0.37144f
C8810 XA.XIR[5].XIC[1].icell.SM VGND 0.00502f
C8811 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80598f
C8812 XA.XIR[5].XIC[2].icell.PUM VGND 0.00293f
C8813 XA.XIR[5].XIC[1].icell.Ien VGND 0.37144f
C8814 XA.XIR[5].XIC[0].icell.SM VGND 0.00502f
C8815 a_n1049_5611# VGND 0.02888f
C8816 XA.XIR[5].XIC[1].icell.PUM VGND 0.00293f
C8817 XA.XIR[5].XIC[0].icell.Ien VGND 0.37178f
C8818 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01044f
C8819 XA.XIR[5].XIC[0].icell.PUM VGND 0.00516f
C8820 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57291f
C8821 XA.XIR[5].XIC_dummy_left.icell.PUM VGND 0.00215f
C8822 XThR.Tn[5] VGND 13.96673f
C8823 XThR.TB6 VGND 1.38212f
C8824 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C8825 XA.XIR[5].XIC_15.icell.PDM VGND 0.18855f
C8826 XA.XIR[5].XIC[14].icell.PDM VGND 0.18809f
C8827 XA.XIR[5].XIC[13].icell.PDM VGND 0.18809f
C8828 XA.XIR[5].XIC[12].icell.PDM VGND 0.18809f
C8829 XA.XIR[5].XIC[11].icell.PDM VGND 0.18809f
C8830 XA.XIR[5].XIC[10].icell.PDM VGND 0.18809f
C8831 XA.XIR[5].XIC[9].icell.PDM VGND 0.18809f
C8832 XA.XIR[5].XIC[8].icell.PDM VGND 0.18809f
C8833 XA.XIR[5].XIC[7].icell.PDM VGND 0.18809f
C8834 XA.XIR[5].XIC[6].icell.PDM VGND 0.18809f
C8835 XA.XIR[5].XIC[5].icell.PDM VGND 0.18809f
C8836 XA.XIR[5].XIC[4].icell.PDM VGND 0.18809f
C8837 XA.XIR[5].XIC[3].icell.PDM VGND 0.18809f
C8838 XA.XIR[5].XIC[2].icell.PDM VGND 0.18809f
C8839 XA.XIR[5].XIC[1].icell.PDM VGND 0.18809f
C8840 XA.XIR[5].XIC[0].icell.PDM VGND 0.18817f
C8841 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C8842 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85795f
C8843 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C8844 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60802f
C8845 XA.XIR[4].XIC_15.icell.SM VGND 0.00474f
C8846 XA.XIR[4].XIC_dummy_right.icell.PUM VGND 0.00215f
C8847 XA.XIR[4].XIC_15.icell.Ien VGND 0.37063f
C8848 XA.XIR[4].XIC[14].icell.SM VGND 0.00502f
C8849 XA.XIR[4].XIC_15.icell.PUM VGND 0.00282f
C8850 XA.XIR[4].XIC[14].icell.Ien VGND 0.37144f
C8851 XA.XIR[4].XIC[13].icell.SM VGND 0.00502f
C8852 XA.XIR[4].XIC[14].icell.PUM VGND 0.00293f
C8853 XA.XIR[4].XIC[13].icell.Ien VGND 0.37144f
C8854 XA.XIR[4].XIC[12].icell.SM VGND 0.00502f
C8855 XA.XIR[4].XIC[13].icell.PUM VGND 0.00293f
C8856 XA.XIR[4].XIC[12].icell.Ien VGND 0.37144f
C8857 XA.XIR[4].XIC[11].icell.SM VGND 0.00502f
C8858 XA.XIR[4].XIC[12].icell.PUM VGND 0.00293f
C8859 XA.XIR[4].XIC[11].icell.Ien VGND 0.37144f
C8860 XA.XIR[4].XIC[10].icell.SM VGND 0.00502f
C8861 XA.XIR[4].XIC[11].icell.PUM VGND 0.00293f
C8862 XA.XIR[4].XIC[10].icell.Ien VGND 0.37144f
C8863 XA.XIR[4].XIC[9].icell.SM VGND 0.00502f
C8864 XA.XIR[4].XIC[10].icell.PUM VGND 0.00293f
C8865 XA.XIR[4].XIC[9].icell.Ien VGND 0.37144f
C8866 XA.XIR[4].XIC[8].icell.SM VGND 0.00502f
C8867 XA.XIR[4].XIC[9].icell.PUM VGND 0.00293f
C8868 XA.XIR[4].XIC[8].icell.Ien VGND 0.37144f
C8869 XA.XIR[4].XIC[7].icell.SM VGND 0.00502f
C8870 XA.XIR[4].XIC[8].icell.PUM VGND 0.00293f
C8871 XA.XIR[4].XIC[7].icell.Ien VGND 0.37144f
C8872 XA.XIR[4].XIC[6].icell.SM VGND 0.00502f
C8873 XA.XIR[4].XIC[7].icell.PUM VGND 0.00293f
C8874 XA.XIR[4].XIC[6].icell.Ien VGND 0.37144f
C8875 XA.XIR[4].XIC[5].icell.SM VGND 0.00502f
C8876 XA.XIR[4].XIC[6].icell.PUM VGND 0.00293f
C8877 XA.XIR[4].XIC[5].icell.Ien VGND 0.37144f
C8878 XA.XIR[4].XIC[4].icell.SM VGND 0.00502f
C8879 XA.XIR[4].XIC[5].icell.PUM VGND 0.00293f
C8880 XA.XIR[4].XIC[4].icell.Ien VGND 0.37144f
C8881 XA.XIR[4].XIC[3].icell.SM VGND 0.00502f
C8882 XA.XIR[4].XIC[4].icell.PUM VGND 0.00293f
C8883 XA.XIR[4].XIC[3].icell.Ien VGND 0.37144f
C8884 XA.XIR[4].XIC[2].icell.SM VGND 0.00502f
C8885 XA.XIR[4].XIC[3].icell.PUM VGND 0.00293f
C8886 XA.XIR[4].XIC[2].icell.Ien VGND 0.37144f
C8887 XA.XIR[4].XIC[1].icell.SM VGND 0.00502f
C8888 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.8077f
C8889 XA.XIR[4].XIC[2].icell.PUM VGND 0.00293f
C8890 XA.XIR[4].XIC[1].icell.Ien VGND 0.37144f
C8891 XA.XIR[4].XIC[0].icell.SM VGND 0.00502f
C8892 XA.XIR[4].XIC[1].icell.PUM VGND 0.00293f
C8893 XA.XIR[4].XIC[0].icell.Ien VGND 0.37178f
C8894 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01044f
C8895 XA.XIR[4].XIC[0].icell.PUM VGND 0.00516f
C8896 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57336f
C8897 XA.XIR[4].XIC_dummy_left.icell.PUM VGND 0.00215f
C8898 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C8899 XA.XIR[4].XIC_15.icell.PDM VGND 0.18855f
C8900 XA.XIR[4].XIC[14].icell.PDM VGND 0.18809f
C8901 XA.XIR[4].XIC[13].icell.PDM VGND 0.18809f
C8902 XA.XIR[4].XIC[12].icell.PDM VGND 0.18809f
C8903 XA.XIR[4].XIC[11].icell.PDM VGND 0.18809f
C8904 XA.XIR[4].XIC[10].icell.PDM VGND 0.18809f
C8905 XA.XIR[4].XIC[9].icell.PDM VGND 0.18809f
C8906 XA.XIR[4].XIC[8].icell.PDM VGND 0.18809f
C8907 XA.XIR[4].XIC[7].icell.PDM VGND 0.18809f
C8908 XA.XIR[4].XIC[6].icell.PDM VGND 0.18809f
C8909 XA.XIR[4].XIC[5].icell.PDM VGND 0.18809f
C8910 XA.XIR[4].XIC[4].icell.PDM VGND 0.18809f
C8911 XA.XIR[4].XIC[3].icell.PDM VGND 0.18809f
C8912 XA.XIR[4].XIC[2].icell.PDM VGND 0.18809f
C8913 XA.XIR[4].XIC[1].icell.PDM VGND 0.18809f
C8914 XA.XIR[4].XIC[0].icell.PDM VGND 0.18817f
C8915 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C8916 XThR.Tn[4] VGND 14.03736f
C8917 a_n1049_6405# VGND 0.02935f
C8918 a_n1319_6405# VGND 0.00166f
C8919 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85795f
C8920 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C8921 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60802f
C8922 XA.XIR[3].XIC_15.icell.SM VGND 0.00474f
C8923 XA.XIR[3].XIC_dummy_right.icell.PUM VGND 0.00215f
C8924 XA.XIR[3].XIC_15.icell.Ien VGND 0.37063f
C8925 XA.XIR[3].XIC[14].icell.SM VGND 0.00502f
C8926 XA.XIR[3].XIC_15.icell.PUM VGND 0.00282f
C8927 XA.XIR[3].XIC[14].icell.Ien VGND 0.37144f
C8928 XA.XIR[3].XIC[13].icell.SM VGND 0.00502f
C8929 XA.XIR[3].XIC[14].icell.PUM VGND 0.00293f
C8930 XA.XIR[3].XIC[13].icell.Ien VGND 0.37144f
C8931 XA.XIR[3].XIC[12].icell.SM VGND 0.00502f
C8932 XA.XIR[3].XIC[13].icell.PUM VGND 0.00293f
C8933 XA.XIR[3].XIC[12].icell.Ien VGND 0.37144f
C8934 XA.XIR[3].XIC[11].icell.SM VGND 0.00502f
C8935 XA.XIR[3].XIC[12].icell.PUM VGND 0.00293f
C8936 XA.XIR[3].XIC[11].icell.Ien VGND 0.37144f
C8937 XA.XIR[3].XIC[10].icell.SM VGND 0.00502f
C8938 XA.XIR[3].XIC[11].icell.PUM VGND 0.00293f
C8939 XA.XIR[3].XIC[10].icell.Ien VGND 0.37144f
C8940 XA.XIR[3].XIC[9].icell.SM VGND 0.00502f
C8941 XA.XIR[3].XIC[10].icell.PUM VGND 0.00293f
C8942 XA.XIR[3].XIC[9].icell.Ien VGND 0.37144f
C8943 XA.XIR[3].XIC[8].icell.SM VGND 0.00502f
C8944 XA.XIR[3].XIC[9].icell.PUM VGND 0.00293f
C8945 XA.XIR[3].XIC[8].icell.Ien VGND 0.37144f
C8946 XA.XIR[3].XIC[7].icell.SM VGND 0.00502f
C8947 XA.XIR[3].XIC[8].icell.PUM VGND 0.00293f
C8948 XA.XIR[3].XIC[7].icell.Ien VGND 0.37144f
C8949 XA.XIR[3].XIC[6].icell.SM VGND 0.00502f
C8950 XA.XIR[3].XIC[7].icell.PUM VGND 0.00293f
C8951 XA.XIR[3].XIC[6].icell.Ien VGND 0.37144f
C8952 XA.XIR[3].XIC[5].icell.SM VGND 0.00502f
C8953 XA.XIR[3].XIC[6].icell.PUM VGND 0.00293f
C8954 XA.XIR[3].XIC[5].icell.Ien VGND 0.37144f
C8955 XA.XIR[3].XIC[4].icell.SM VGND 0.00502f
C8956 XA.XIR[3].XIC[5].icell.PUM VGND 0.00293f
C8957 XA.XIR[3].XIC[4].icell.Ien VGND 0.37144f
C8958 XA.XIR[3].XIC[3].icell.SM VGND 0.00502f
C8959 XA.XIR[3].XIC[4].icell.PUM VGND 0.00293f
C8960 XA.XIR[3].XIC[3].icell.Ien VGND 0.37144f
C8961 XA.XIR[3].XIC[2].icell.SM VGND 0.00502f
C8962 XA.XIR[3].XIC[3].icell.PUM VGND 0.00293f
C8963 XA.XIR[3].XIC[2].icell.Ien VGND 0.37144f
C8964 XA.XIR[3].XIC[1].icell.SM VGND 0.00502f
C8965 XThR.TB5 VGND 1.32753f
C8966 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80611f
C8967 XA.XIR[3].XIC[2].icell.PUM VGND 0.00293f
C8968 XA.XIR[3].XIC[1].icell.Ien VGND 0.37144f
C8969 XA.XIR[3].XIC[0].icell.SM VGND 0.00502f
C8970 XA.XIR[3].XIC[1].icell.PUM VGND 0.00293f
C8971 XA.XIR[3].XIC[0].icell.Ien VGND 0.37178f
C8972 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01044f
C8973 XA.XIR[3].XIC[0].icell.PUM VGND 0.00516f
C8974 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57425f
C8975 a_n1049_6699# VGND 0.02979f
C8976 XA.XIR[3].XIC_dummy_left.icell.PUM VGND 0.00215f
C8977 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C8978 XA.XIR[3].XIC_15.icell.PDM VGND 0.18855f
C8979 XA.XIR[3].XIC[14].icell.PDM VGND 0.18809f
C8980 XA.XIR[3].XIC[13].icell.PDM VGND 0.18809f
C8981 XA.XIR[3].XIC[12].icell.PDM VGND 0.18809f
C8982 XA.XIR[3].XIC[11].icell.PDM VGND 0.18809f
C8983 XA.XIR[3].XIC[10].icell.PDM VGND 0.18809f
C8984 XA.XIR[3].XIC[9].icell.PDM VGND 0.18809f
C8985 XA.XIR[3].XIC[8].icell.PDM VGND 0.18809f
C8986 XA.XIR[3].XIC[7].icell.PDM VGND 0.18809f
C8987 XA.XIR[3].XIC[6].icell.PDM VGND 0.18809f
C8988 XA.XIR[3].XIC[5].icell.PDM VGND 0.18809f
C8989 XA.XIR[3].XIC[4].icell.PDM VGND 0.18809f
C8990 XA.XIR[3].XIC[3].icell.PDM VGND 0.18809f
C8991 XA.XIR[3].XIC[2].icell.PDM VGND 0.18809f
C8992 XA.XIR[3].XIC[1].icell.PDM VGND 0.18809f
C8993 XA.XIR[3].XIC[0].icell.PDM VGND 0.18817f
C8994 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C8995 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85795f
C8996 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C8997 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60802f
C8998 XA.XIR[2].XIC_15.icell.SM VGND 0.00474f
C8999 XA.XIR[2].XIC_dummy_right.icell.PUM VGND 0.00215f
C9000 XA.XIR[2].XIC_15.icell.Ien VGND 0.37063f
C9001 XA.XIR[2].XIC[14].icell.SM VGND 0.00502f
C9002 XA.XIR[2].XIC_15.icell.PUM VGND 0.00282f
C9003 XA.XIR[2].XIC[14].icell.Ien VGND 0.37144f
C9004 XA.XIR[2].XIC[13].icell.SM VGND 0.00502f
C9005 XA.XIR[2].XIC[14].icell.PUM VGND 0.00293f
C9006 XA.XIR[2].XIC[13].icell.Ien VGND 0.37144f
C9007 XA.XIR[2].XIC[12].icell.SM VGND 0.00502f
C9008 XA.XIR[2].XIC[13].icell.PUM VGND 0.00293f
C9009 XA.XIR[2].XIC[12].icell.Ien VGND 0.37144f
C9010 XA.XIR[2].XIC[11].icell.SM VGND 0.00502f
C9011 XA.XIR[2].XIC[12].icell.PUM VGND 0.00293f
C9012 XA.XIR[2].XIC[11].icell.Ien VGND 0.37144f
C9013 XA.XIR[2].XIC[10].icell.SM VGND 0.00502f
C9014 XA.XIR[2].XIC[11].icell.PUM VGND 0.00293f
C9015 XA.XIR[2].XIC[10].icell.Ien VGND 0.37144f
C9016 XA.XIR[2].XIC[9].icell.SM VGND 0.00502f
C9017 XA.XIR[2].XIC[10].icell.PUM VGND 0.00293f
C9018 XA.XIR[2].XIC[9].icell.Ien VGND 0.37144f
C9019 XA.XIR[2].XIC[8].icell.SM VGND 0.00502f
C9020 XA.XIR[2].XIC[9].icell.PUM VGND 0.00293f
C9021 XA.XIR[2].XIC[8].icell.Ien VGND 0.37144f
C9022 XA.XIR[2].XIC[7].icell.SM VGND 0.00502f
C9023 XA.XIR[2].XIC[8].icell.PUM VGND 0.00293f
C9024 XA.XIR[2].XIC[7].icell.Ien VGND 0.37144f
C9025 XA.XIR[2].XIC[6].icell.SM VGND 0.00502f
C9026 XA.XIR[2].XIC[7].icell.PUM VGND 0.00293f
C9027 XA.XIR[2].XIC[6].icell.Ien VGND 0.37144f
C9028 XA.XIR[2].XIC[5].icell.SM VGND 0.00502f
C9029 XA.XIR[2].XIC[6].icell.PUM VGND 0.00293f
C9030 XA.XIR[2].XIC[5].icell.Ien VGND 0.37144f
C9031 XA.XIR[2].XIC[4].icell.SM VGND 0.00502f
C9032 XA.XIR[2].XIC[5].icell.PUM VGND 0.00293f
C9033 XA.XIR[2].XIC[4].icell.Ien VGND 0.37144f
C9034 XA.XIR[2].XIC[3].icell.SM VGND 0.00502f
C9035 XA.XIR[2].XIC[4].icell.PUM VGND 0.00293f
C9036 XA.XIR[2].XIC[3].icell.Ien VGND 0.37144f
C9037 XA.XIR[2].XIC[2].icell.SM VGND 0.00502f
C9038 XA.XIR[2].XIC[3].icell.PUM VGND 0.00293f
C9039 XA.XIR[2].XIC[2].icell.Ien VGND 0.37144f
C9040 XA.XIR[2].XIC[1].icell.SM VGND 0.00502f
C9041 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80825f
C9042 XA.XIR[2].XIC[2].icell.PUM VGND 0.00293f
C9043 XA.XIR[2].XIC[1].icell.Ien VGND 0.37144f
C9044 XA.XIR[2].XIC[0].icell.SM VGND 0.00502f
C9045 XThR.Tn[3] VGND 13.98256f
C9046 XThR.TB4 VGND 1.48815f
C9047 XA.XIR[2].XIC[1].icell.PUM VGND 0.00293f
C9048 XA.XIR[2].XIC[0].icell.Ien VGND 0.37178f
C9049 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01044f
C9050 XA.XIR[2].XIC[0].icell.PUM VGND 0.00516f
C9051 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57559f
C9052 a_n1335_7243# VGND 0.00179f
C9053 XA.XIR[2].XIC_dummy_left.icell.PUM VGND 0.00215f
C9054 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C9055 XA.XIR[2].XIC_15.icell.PDM VGND 0.18855f
C9056 XA.XIR[2].XIC[14].icell.PDM VGND 0.18809f
C9057 XA.XIR[2].XIC[13].icell.PDM VGND 0.18809f
C9058 XA.XIR[2].XIC[12].icell.PDM VGND 0.18809f
C9059 XA.XIR[2].XIC[11].icell.PDM VGND 0.18809f
C9060 XA.XIR[2].XIC[10].icell.PDM VGND 0.18809f
C9061 XA.XIR[2].XIC[9].icell.PDM VGND 0.18809f
C9062 XA.XIR[2].XIC[8].icell.PDM VGND 0.18809f
C9063 XA.XIR[2].XIC[7].icell.PDM VGND 0.18809f
C9064 XA.XIR[2].XIC[6].icell.PDM VGND 0.18809f
C9065 XA.XIR[2].XIC[5].icell.PDM VGND 0.18809f
C9066 XA.XIR[2].XIC[4].icell.PDM VGND 0.18809f
C9067 XA.XIR[2].XIC[3].icell.PDM VGND 0.18809f
C9068 XA.XIR[2].XIC[2].icell.PDM VGND 0.18809f
C9069 XA.XIR[2].XIC[1].icell.PDM VGND 0.18809f
C9070 XA.XIR[2].XIC[0].icell.PDM VGND 0.18817f
C9071 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C9072 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85795f
C9073 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C9074 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60802f
C9075 XA.XIR[1].XIC_15.icell.SM VGND 0.00474f
C9076 XA.XIR[1].XIC_dummy_right.icell.PUM VGND 0.00215f
C9077 XA.XIR[1].XIC_15.icell.Ien VGND 0.37063f
C9078 XA.XIR[1].XIC[14].icell.SM VGND 0.00502f
C9079 XA.XIR[1].XIC_15.icell.PUM VGND 0.00282f
C9080 XA.XIR[1].XIC[14].icell.Ien VGND 0.37144f
C9081 XA.XIR[1].XIC[13].icell.SM VGND 0.00502f
C9082 XA.XIR[1].XIC[14].icell.PUM VGND 0.00293f
C9083 XA.XIR[1].XIC[13].icell.Ien VGND 0.37144f
C9084 XA.XIR[1].XIC[12].icell.SM VGND 0.00502f
C9085 XA.XIR[1].XIC[13].icell.PUM VGND 0.00293f
C9086 XA.XIR[1].XIC[12].icell.Ien VGND 0.37144f
C9087 XA.XIR[1].XIC[11].icell.SM VGND 0.00502f
C9088 XA.XIR[1].XIC[12].icell.PUM VGND 0.00293f
C9089 XA.XIR[1].XIC[11].icell.Ien VGND 0.37144f
C9090 XA.XIR[1].XIC[10].icell.SM VGND 0.00502f
C9091 XA.XIR[1].XIC[11].icell.PUM VGND 0.00293f
C9092 XA.XIR[1].XIC[10].icell.Ien VGND 0.37144f
C9093 XA.XIR[1].XIC[9].icell.SM VGND 0.00502f
C9094 XA.XIR[1].XIC[10].icell.PUM VGND 0.00293f
C9095 XA.XIR[1].XIC[9].icell.Ien VGND 0.37144f
C9096 XA.XIR[1].XIC[8].icell.SM VGND 0.00502f
C9097 XA.XIR[1].XIC[9].icell.PUM VGND 0.00293f
C9098 XA.XIR[1].XIC[8].icell.Ien VGND 0.37144f
C9099 XA.XIR[1].XIC[7].icell.SM VGND 0.00502f
C9100 XA.XIR[1].XIC[8].icell.PUM VGND 0.00293f
C9101 XA.XIR[1].XIC[7].icell.Ien VGND 0.37144f
C9102 XA.XIR[1].XIC[6].icell.SM VGND 0.00502f
C9103 XA.XIR[1].XIC[7].icell.PUM VGND 0.00293f
C9104 XA.XIR[1].XIC[6].icell.Ien VGND 0.37144f
C9105 XA.XIR[1].XIC[5].icell.SM VGND 0.00502f
C9106 XA.XIR[1].XIC[6].icell.PUM VGND 0.00293f
C9107 XA.XIR[1].XIC[5].icell.Ien VGND 0.37144f
C9108 XA.XIR[1].XIC[4].icell.SM VGND 0.00502f
C9109 XA.XIR[1].XIC[5].icell.PUM VGND 0.00293f
C9110 XA.XIR[1].XIC[4].icell.Ien VGND 0.37144f
C9111 XA.XIR[1].XIC[3].icell.SM VGND 0.00502f
C9112 XA.XIR[1].XIC[4].icell.PUM VGND 0.00293f
C9113 XA.XIR[1].XIC[3].icell.Ien VGND 0.37144f
C9114 XA.XIR[1].XIC[2].icell.SM VGND 0.00502f
C9115 XA.XIR[1].XIC[3].icell.PUM VGND 0.00293f
C9116 XA.XIR[1].XIC[2].icell.Ien VGND 0.37144f
C9117 XA.XIR[1].XIC[1].icell.SM VGND 0.00502f
C9118 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80611f
C9119 XA.XIR[1].XIC[2].icell.PUM VGND 0.00293f
C9120 XA.XIR[1].XIC[1].icell.Ien VGND 0.37144f
C9121 XA.XIR[1].XIC[0].icell.SM VGND 0.00502f
C9122 XThR.Tn[2] VGND 14.03476f
C9123 a_n1049_7493# VGND 0.02484f
C9124 XThR.TB3 VGND 3.11868f
C9125 XThR.TA3 VGND 1.95537f
C9126 XA.XIR[1].XIC[1].icell.PUM VGND 0.00293f
C9127 XA.XIR[1].XIC[0].icell.Ien VGND 0.37178f
C9128 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01044f
C9129 XA.XIR[1].XIC[0].icell.PUM VGND 0.00516f
C9130 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57378f
C9131 XA.XIR[1].XIC_dummy_left.icell.PUM VGND 0.00215f
C9132 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C9133 XA.XIR[1].XIC_15.icell.PDM VGND 0.18855f
C9134 XA.XIR[1].XIC[14].icell.PDM VGND 0.18809f
C9135 XA.XIR[1].XIC[13].icell.PDM VGND 0.18809f
C9136 XA.XIR[1].XIC[12].icell.PDM VGND 0.18809f
C9137 XA.XIR[1].XIC[11].icell.PDM VGND 0.18809f
C9138 XA.XIR[1].XIC[10].icell.PDM VGND 0.18809f
C9139 XA.XIR[1].XIC[9].icell.PDM VGND 0.18809f
C9140 XA.XIR[1].XIC[8].icell.PDM VGND 0.18809f
C9141 XA.XIR[1].XIC[7].icell.PDM VGND 0.18809f
C9142 XA.XIR[1].XIC[6].icell.PDM VGND 0.18809f
C9143 XA.XIR[1].XIC[5].icell.PDM VGND 0.18809f
C9144 XA.XIR[1].XIC[4].icell.PDM VGND 0.18809f
C9145 XA.XIR[1].XIC[3].icell.PDM VGND 0.18809f
C9146 XA.XIR[1].XIC[2].icell.PDM VGND 0.18809f
C9147 XA.XIR[1].XIC[1].icell.PDM VGND 0.18809f
C9148 XA.XIR[1].XIC[0].icell.PDM VGND 0.18817f
C9149 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C9150 a_n1049_7787# VGND 0.03396f
C9151 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87257f
C9152 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01019f
C9153 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61845f
C9154 XA.XIR[0].XIC_15.icell.SM VGND 0.00474f
C9155 XA.XIR[0].XIC_dummy_right.icell.PUM VGND 0.00216f
C9156 XA.XIR[0].XIC_15.icell.Ien VGND 0.37702f
C9157 XA.XIR[0].XIC[14].icell.SM VGND 0.00624f
C9158 XA.XIR[0].XIC_15.icell.PUM VGND 0.00475f
C9159 XA.XIR[0].XIC[14].icell.Ien VGND 0.38465f
C9160 XA.XIR[0].XIC[13].icell.SM VGND 0.00624f
C9161 XA.XIR[0].XIC[14].icell.PUM VGND 0.00392f
C9162 XA.XIR[0].XIC[13].icell.Ien VGND 0.38439f
C9163 XA.XIR[0].XIC[12].icell.SM VGND 0.00624f
C9164 XA.XIR[0].XIC[13].icell.PUM VGND 0.00397f
C9165 XA.XIR[0].XIC[12].icell.Ien VGND 0.381f
C9166 XA.XIR[0].XIC[11].icell.SM VGND 0.00624f
C9167 XA.XIR[0].XIC[12].icell.PUM VGND 0.00392f
C9168 XA.XIR[0].XIC[11].icell.Ien VGND 0.38167f
C9169 XA.XIR[0].XIC[10].icell.SM VGND 0.00624f
C9170 XA.XIR[0].XIC[11].icell.PUM VGND 0.00392f
C9171 XA.XIR[0].XIC[10].icell.Ien VGND 0.38301f
C9172 XA.XIR[0].XIC[9].icell.SM VGND 0.00624f
C9173 XA.XIR[0].XIC[10].icell.PUM VGND 0.00392f
C9174 XA.XIR[0].XIC[9].icell.Ien VGND 0.38128f
C9175 XA.XIR[0].XIC[8].icell.SM VGND 0.00624f
C9176 XA.XIR[0].XIC[9].icell.PUM VGND 0.00392f
C9177 XA.XIR[0].XIC[8].icell.Ien VGND 0.38176f
C9178 XA.XIR[0].XIC[7].icell.SM VGND 0.00624f
C9179 XA.XIR[0].XIC[8].icell.PUM VGND 0.00392f
C9180 XA.XIR[0].XIC[7].icell.Ien VGND 0.382f
C9181 XA.XIR[0].XIC[6].icell.SM VGND 0.00624f
C9182 XA.XIR[0].XIC[7].icell.PUM VGND 0.00392f
C9183 XA.XIR[0].XIC[6].icell.Ien VGND 0.38192f
C9184 XA.XIR[0].XIC[5].icell.SM VGND 0.00624f
C9185 XA.XIR[0].XIC[6].icell.PUM VGND 0.00403f
C9186 XA.XIR[0].XIC[5].icell.Ien VGND 0.38091f
C9187 XA.XIR[0].XIC[4].icell.SM VGND 0.00624f
C9188 XA.XIR[0].XIC[5].icell.PUM VGND 0.00392f
C9189 XA.XIR[0].XIC[4].icell.Ien VGND 0.38104f
C9190 XA.XIR[0].XIC[3].icell.SM VGND 0.00624f
C9191 XA.XIR[0].XIC[4].icell.PUM VGND 0.00392f
C9192 XA.XIR[0].XIC[3].icell.Ien VGND 0.38229f
C9193 XA.XIR[0].XIC[2].icell.SM VGND 0.00624f
C9194 XA.XIR[0].XIC[3].icell.PUM VGND 0.00392f
C9195 XA.XIR[0].XIC[2].icell.Ien VGND 0.38432f
C9196 XA.XIR[0].XIC[1].icell.SM VGND 0.00624f
C9197 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.841f
C9198 XA.XIR[0].XIC[2].icell.PUM VGND 0.00392f
C9199 XA.XIR[0].XIC[1].icell.Ien VGND 0.38432f
C9200 XA.XIR[0].XIC[0].icell.SM VGND 0.00624f
C9201 XA.XIR[0].XIC[1].icell.PUM VGND 0.00394f
C9202 XA.XIR[0].XIC[0].icell.Ien VGND 0.38446f
C9203 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01044f
C9204 XThR.Tn[1] VGND 14.06925f
C9205 a_n1335_8107# VGND 0.00163f
C9206 XThR.TB2 VGND 1.47668f
C9207 XThR.TA2 VGND 0.95641f
C9208 XA.XIR[0].XIC[0].icell.PUM VGND 0.00623f
C9209 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58675f
C9210 XA.XIR[0].XIC_dummy_left.icell.PUM VGND 0.0035f
C9211 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.25173f
C9212 XA.XIR[0].XIC_15.icell.PDM VGND 0.20835f
C9213 XA.XIR[0].XIC[14].icell.PDM VGND 0.24664f
C9214 XA.XIR[0].XIC[13].icell.PDM VGND 0.24612f
C9215 XA.XIR[0].XIC[12].icell.PDM VGND 0.24144f
C9216 XA.XIR[0].XIC[11].icell.PDM VGND 0.24182f
C9217 XA.XIR[0].XIC[10].icell.PDM VGND 0.24172f
C9218 XA.XIR[0].XIC[9].icell.PDM VGND 0.24144f
C9219 XA.XIR[0].XIC[8].icell.PDM VGND 0.24144f
C9220 XA.XIR[0].XIC[7].icell.PDM VGND 0.24388f
C9221 XA.XIR[0].XIC[6].icell.PDM VGND 0.24108f
C9222 XA.XIR[0].XIC[5].icell.PDM VGND 0.24297f
C9223 XA.XIR[0].XIC[4].icell.PDM VGND 0.24156f
C9224 XA.XIR[0].XIC[3].icell.PDM VGND 0.24455f
C9225 XA.XIR[0].XIC[2].icell.PDM VGND 0.24578f
C9226 XA.XIR[0].XIC[1].icell.PDM VGND 0.24578f
C9227 XA.XIR[0].XIC[0].icell.PDM VGND 0.24491f
C9228 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24713f
C9229 a_n1335_8331# VGND 0.00203f
C9230 XThR.Tn[0] VGND 14.40653f
C9231 a_n1049_8581# VGND 0.04324f
C9232 XThR.TBN VGND 7.8135f
C9233 XThR.TB1 VGND 2.41896f
C9234 XThR.TAN VGND 2.61156f
C9235 XThR.TA1 VGND 1.76044f
C9236 XThC.Tn[14] VGND 10.02286f
C9237 XThC.Tn[13] VGND 9.79583f
C9238 XThC.Tn[12] VGND 9.63554f
C9239 XThC.Tn[11] VGND 9.46598f
C9240 XThC.Tn[10] VGND 9.29745f
C9241 XThC.Tn[9] VGND 9.27278f
C9242 XThC.Tn[8] VGND 9.24802f
C9243 a_10915_9569# VGND 0.56659f
C9244 a_10051_9569# VGND 0.55927f
C9245 a_9827_9569# VGND 0.54559f
C9246 a_8963_9569# VGND 0.55448f
C9247 a_8739_9569# VGND 0.55288f
C9248 a_7875_9569# VGND 0.55432f
C9249 a_7651_9569# VGND 0.55717f
C9250 XThC.Tn[7] VGND 10.56205f
C9251 XThC.Tn[6] VGND 10.35711f
C9252 XThC.Tn[5] VGND 10.62787f
C9253 XThC.Tn[4] VGND 10.6808f
C9254 XThC.Tn[3] VGND 9.9249f
C9255 XThC.Tn[2] VGND 10.4557f
C9256 XThC.Tn[1] VGND 10.33149f
C9257 XThC.Tn[0] VGND 10.74903f
C9258 a_6243_9615# VGND 0.0299f
C9259 a_5949_9615# VGND 0.03432f
C9260 a_5155_9615# VGND 0.03615f
C9261 a_4861_9615# VGND 0.03632f
C9262 a_4067_9615# VGND 0.03071f
C9263 a_3773_9615# VGND 0.03867f
C9264 a_2979_9615# VGND 0.04107f
C9265 a_8739_10571# VGND 0.00194f
C9266 XThC.TBN VGND 7.91488f
C9267 XThC.TB7 VGND 1.38013f
C9268 XThC.TB6 VGND 1.38691f
C9269 a_5155_10571# VGND 0.00165f
C9270 XThC.TAN VGND 2.73083f
C9271 XThC.TB5 VGND 1.32648f
C9272 XThC.TAN2 VGND 1.2327f
C9273 a_4387_10575# VGND 0.00179f
C9274 a_3523_10575# VGND 0.00163f
C9275 a_3299_10575# VGND 0.00202f
C9276 XThC.TB4 VGND 2.79989f
C9277 XThC.TB3 VGND 3.08942f
C9278 XThC.TA3 VGND 1.96056f
C9279 XThC.TA2 VGND 0.95757f
C9280 XThC.TB2 VGND 1.47589f
C9281 XThC.TB1 VGND 2.409f
C9282 XThC.TA1 VGND 1.75974f
C9283 XThR.TB3.t2 VGND 0.06176f
C9284 XThR.TB3.n0 VGND 0.01521f
C9285 XThR.TB3.t8 VGND 0.04903f
C9286 XThR.TB3.t15 VGND 0.02889f
C9287 XThR.TB3.t13 VGND 0.04903f
C9288 XThR.TB3.t6 VGND 0.02889f
C9289 XThR.TB3.t9 VGND 0.04903f
C9290 XThR.TB3.t17 VGND 0.02889f
C9291 XThR.TB3.n1 VGND 0.08226f
C9292 XThR.TB3.n2 VGND 0.08688f
C9293 XThR.TB3.n3 VGND 0.03573f
C9294 XThR.TB3.n4 VGND 0.0707f
C9295 XThR.TB3.t12 VGND 0.04903f
C9296 XThR.TB3.t4 VGND 0.02889f
C9297 XThR.TB3.n5 VGND 0.06608f
C9298 XThR.TB3.n6 VGND 0.03236f
C9299 XThR.TB3.n7 VGND 0.02685f
C9300 XThR.TB3.t18 VGND 0.04903f
C9301 XThR.TB3.t5 VGND 0.02889f
C9302 XThR.TB3.n8 VGND 0.03005f
C9303 XThR.TB3.t7 VGND 0.04903f
C9304 XThR.TB3.t10 VGND 0.02889f
C9305 XThR.TB3.n9 VGND 0.05992f
C9306 XThR.TB3.t11 VGND 0.04903f
C9307 XThR.TB3.t16 VGND 0.02889f
C9308 XThR.TB3.n10 VGND 0.06454f
C9309 XThR.TB3.n11 VGND 0.03645f
C9310 XThR.TB3.n12 VGND 0.06034f
C9311 XThR.TB3.n13 VGND 0.03128f
C9312 XThR.TB3.n14 VGND 0.02851f
C9313 XThR.TB3.n15 VGND 0.06454f
C9314 XThR.TB3.t14 VGND 0.04903f
C9315 XThR.TB3.t3 VGND 0.02889f
C9316 XThR.TB3.n16 VGND 0.05838f
C9317 XThR.TB3.n17 VGND 0.03236f
C9318 XThR.TB3.n18 VGND 0.04707f
C9319 XThR.TB3.n19 VGND 0.28641f
C9320 XThR.TB3.t0 VGND 0.03152f
C9321 XThR.TB3.t1 VGND 0.03152f
C9322 XThR.TB3.n20 VGND 0.06766f
C9323 XThR.TB3.n21 VGND 0.157f
C9324 XThR.TB3.n22 VGND 0.03296f
C9325 XThR.TB1.t1 VGND 0.03165f
C9326 XThR.TB1.n0 VGND 0.0078f
C9327 XThR.TB1.t8 VGND 0.02512f
C9328 XThR.TB1.t15 VGND 0.0148f
C9329 XThR.TB1.t14 VGND 0.02512f
C9330 XThR.TB1.t7 VGND 0.0148f
C9331 XThR.TB1.t10 VGND 0.02512f
C9332 XThR.TB1.t18 VGND 0.0148f
C9333 XThR.TB1.n1 VGND 0.04215f
C9334 XThR.TB1.n2 VGND 0.04452f
C9335 XThR.TB1.n3 VGND 0.01831f
C9336 XThR.TB1.n4 VGND 0.03623f
C9337 XThR.TB1.t13 VGND 0.02512f
C9338 XThR.TB1.t4 VGND 0.0148f
C9339 XThR.TB1.n5 VGND 0.03386f
C9340 XThR.TB1.n6 VGND 0.01658f
C9341 XThR.TB1.n7 VGND 0.01376f
C9342 XThR.TB1.t6 VGND 0.02512f
C9343 XThR.TB1.t11 VGND 0.0148f
C9344 XThR.TB1.n8 VGND 0.0154f
C9345 XThR.TB1.t12 VGND 0.02512f
C9346 XThR.TB1.t16 VGND 0.0148f
C9347 XThR.TB1.n9 VGND 0.0307f
C9348 XThR.TB1.t17 VGND 0.02512f
C9349 XThR.TB1.t5 VGND 0.0148f
C9350 XThR.TB1.n10 VGND 0.03307f
C9351 XThR.TB1.n11 VGND 0.01868f
C9352 XThR.TB1.n12 VGND 0.03092f
C9353 XThR.TB1.n13 VGND 0.01603f
C9354 XThR.TB1.n14 VGND 0.01461f
C9355 XThR.TB1.n15 VGND 0.03307f
C9356 XThR.TB1.t3 VGND 0.02512f
C9357 XThR.TB1.t9 VGND 0.0148f
C9358 XThR.TB1.n16 VGND 0.02991f
C9359 XThR.TB1.n17 VGND 0.01658f
C9360 XThR.TB1.n18 VGND 0.02412f
C9361 XThR.TB1.n19 VGND 0.14588f
C9362 XThR.TB1.t2 VGND 0.01615f
C9363 XThR.TB1.t0 VGND 0.01615f
C9364 XThR.TB1.n20 VGND 0.03467f
C9365 XThR.TB1.n21 VGND 0.08068f
C9366 XThR.TB1.n22 VGND 0.01689f
C9367 XThR.Tn[13].t9 VGND 0.02397f
C9368 XThR.Tn[13].t11 VGND 0.02397f
C9369 XThR.Tn[13].n0 VGND 0.07277f
C9370 XThR.Tn[13].t10 VGND 0.02397f
C9371 XThR.Tn[13].t8 VGND 0.02397f
C9372 XThR.Tn[13].n1 VGND 0.05327f
C9373 XThR.Tn[13].n2 VGND 0.24224f
C9374 XThR.Tn[13].t7 VGND 0.01558f
C9375 XThR.Tn[13].t5 VGND 0.01558f
C9376 XThR.Tn[13].n3 VGND 0.03885f
C9377 XThR.Tn[13].t6 VGND 0.01558f
C9378 XThR.Tn[13].t4 VGND 0.01558f
C9379 XThR.Tn[13].n4 VGND 0.03116f
C9380 XThR.Tn[13].n5 VGND 0.07837f
C9381 XThR.Tn[13].t72 VGND 0.01873f
C9382 XThR.Tn[13].t64 VGND 0.02051f
C9383 XThR.Tn[13].n6 VGND 0.05008f
C9384 XThR.Tn[13].n7 VGND 0.09621f
C9385 XThR.Tn[13].t28 VGND 0.01873f
C9386 XThR.Tn[13].t21 VGND 0.02051f
C9387 XThR.Tn[13].n8 VGND 0.05008f
C9388 XThR.Tn[13].t44 VGND 0.01867f
C9389 XThR.Tn[13].t12 VGND 0.02044f
C9390 XThR.Tn[13].n9 VGND 0.05211f
C9391 XThR.Tn[13].n10 VGND 0.03661f
C9392 XThR.Tn[13].n11 VGND 0.00669f
C9393 XThR.Tn[13].n12 VGND 0.11748f
C9394 XThR.Tn[13].t65 VGND 0.01873f
C9395 XThR.Tn[13].t57 VGND 0.02051f
C9396 XThR.Tn[13].n13 VGND 0.05008f
C9397 XThR.Tn[13].t19 VGND 0.01867f
C9398 XThR.Tn[13].t52 VGND 0.02044f
C9399 XThR.Tn[13].n14 VGND 0.05211f
C9400 XThR.Tn[13].n15 VGND 0.03661f
C9401 XThR.Tn[13].n16 VGND 0.00669f
C9402 XThR.Tn[13].n17 VGND 0.11748f
C9403 XThR.Tn[13].t22 VGND 0.01873f
C9404 XThR.Tn[13].t14 VGND 0.02051f
C9405 XThR.Tn[13].n18 VGND 0.05008f
C9406 XThR.Tn[13].t34 VGND 0.01867f
C9407 XThR.Tn[13].t70 VGND 0.02044f
C9408 XThR.Tn[13].n19 VGND 0.05211f
C9409 XThR.Tn[13].n20 VGND 0.03661f
C9410 XThR.Tn[13].n21 VGND 0.00669f
C9411 XThR.Tn[13].n22 VGND 0.11748f
C9412 XThR.Tn[13].t49 VGND 0.01873f
C9413 XThR.Tn[13].t39 VGND 0.02051f
C9414 XThR.Tn[13].n23 VGND 0.05008f
C9415 XThR.Tn[13].t66 VGND 0.01867f
C9416 XThR.Tn[13].t35 VGND 0.02044f
C9417 XThR.Tn[13].n24 VGND 0.05211f
C9418 XThR.Tn[13].n25 VGND 0.03661f
C9419 XThR.Tn[13].n26 VGND 0.00669f
C9420 XThR.Tn[13].n27 VGND 0.11748f
C9421 XThR.Tn[13].t24 VGND 0.01873f
C9422 XThR.Tn[13].t16 VGND 0.02051f
C9423 XThR.Tn[13].n28 VGND 0.05008f
C9424 XThR.Tn[13].t37 VGND 0.01867f
C9425 XThR.Tn[13].t71 VGND 0.02044f
C9426 XThR.Tn[13].n29 VGND 0.05211f
C9427 XThR.Tn[13].n30 VGND 0.03661f
C9428 XThR.Tn[13].n31 VGND 0.00669f
C9429 XThR.Tn[13].n32 VGND 0.11748f
C9430 XThR.Tn[13].t60 VGND 0.01873f
C9431 XThR.Tn[13].t30 VGND 0.02051f
C9432 XThR.Tn[13].n33 VGND 0.05008f
C9433 XThR.Tn[13].t13 VGND 0.01867f
C9434 XThR.Tn[13].t26 VGND 0.02044f
C9435 XThR.Tn[13].n34 VGND 0.05211f
C9436 XThR.Tn[13].n35 VGND 0.03661f
C9437 XThR.Tn[13].n36 VGND 0.00669f
C9438 XThR.Tn[13].n37 VGND 0.11748f
C9439 XThR.Tn[13].t29 VGND 0.01873f
C9440 XThR.Tn[13].t25 VGND 0.02051f
C9441 XThR.Tn[13].n38 VGND 0.05008f
C9442 XThR.Tn[13].t43 VGND 0.01867f
C9443 XThR.Tn[13].t18 VGND 0.02044f
C9444 XThR.Tn[13].n39 VGND 0.05211f
C9445 XThR.Tn[13].n40 VGND 0.03661f
C9446 XThR.Tn[13].n41 VGND 0.00669f
C9447 XThR.Tn[13].n42 VGND 0.11748f
C9448 XThR.Tn[13].t32 VGND 0.01873f
C9449 XThR.Tn[13].t38 VGND 0.02051f
C9450 XThR.Tn[13].n43 VGND 0.05008f
C9451 XThR.Tn[13].t48 VGND 0.01867f
C9452 XThR.Tn[13].t33 VGND 0.02044f
C9453 XThR.Tn[13].n44 VGND 0.05211f
C9454 XThR.Tn[13].n45 VGND 0.03661f
C9455 XThR.Tn[13].n46 VGND 0.00669f
C9456 XThR.Tn[13].n47 VGND 0.11748f
C9457 XThR.Tn[13].t51 VGND 0.01873f
C9458 XThR.Tn[13].t59 VGND 0.02051f
C9459 XThR.Tn[13].n48 VGND 0.05008f
C9460 XThR.Tn[13].t68 VGND 0.01867f
C9461 XThR.Tn[13].t53 VGND 0.02044f
C9462 XThR.Tn[13].n49 VGND 0.05211f
C9463 XThR.Tn[13].n50 VGND 0.03661f
C9464 XThR.Tn[13].n51 VGND 0.00669f
C9465 XThR.Tn[13].n52 VGND 0.11748f
C9466 XThR.Tn[13].t41 VGND 0.01873f
C9467 XThR.Tn[13].t17 VGND 0.02051f
C9468 XThR.Tn[13].n53 VGND 0.05008f
C9469 XThR.Tn[13].t58 VGND 0.01867f
C9470 XThR.Tn[13].t73 VGND 0.02044f
C9471 XThR.Tn[13].n54 VGND 0.05211f
C9472 XThR.Tn[13].n55 VGND 0.03661f
C9473 XThR.Tn[13].n56 VGND 0.00669f
C9474 XThR.Tn[13].n57 VGND 0.11748f
C9475 XThR.Tn[13].t63 VGND 0.01873f
C9476 XThR.Tn[13].t55 VGND 0.02051f
C9477 XThR.Tn[13].n58 VGND 0.05008f
C9478 XThR.Tn[13].t15 VGND 0.01867f
C9479 XThR.Tn[13].t45 VGND 0.02044f
C9480 XThR.Tn[13].n59 VGND 0.05211f
C9481 XThR.Tn[13].n60 VGND 0.03661f
C9482 XThR.Tn[13].n61 VGND 0.00669f
C9483 XThR.Tn[13].n62 VGND 0.11748f
C9484 XThR.Tn[13].t31 VGND 0.01873f
C9485 XThR.Tn[13].t27 VGND 0.02051f
C9486 XThR.Tn[13].n63 VGND 0.05008f
C9487 XThR.Tn[13].t46 VGND 0.01867f
C9488 XThR.Tn[13].t20 VGND 0.02044f
C9489 XThR.Tn[13].n64 VGND 0.05211f
C9490 XThR.Tn[13].n65 VGND 0.03661f
C9491 XThR.Tn[13].n66 VGND 0.00669f
C9492 XThR.Tn[13].n67 VGND 0.11748f
C9493 XThR.Tn[13].t50 VGND 0.01873f
C9494 XThR.Tn[13].t40 VGND 0.02051f
C9495 XThR.Tn[13].n68 VGND 0.05008f
C9496 XThR.Tn[13].t67 VGND 0.01867f
C9497 XThR.Tn[13].t36 VGND 0.02044f
C9498 XThR.Tn[13].n69 VGND 0.05211f
C9499 XThR.Tn[13].n70 VGND 0.03661f
C9500 XThR.Tn[13].n71 VGND 0.00669f
C9501 XThR.Tn[13].n72 VGND 0.11748f
C9502 XThR.Tn[13].t69 VGND 0.01873f
C9503 XThR.Tn[13].t62 VGND 0.02051f
C9504 XThR.Tn[13].n73 VGND 0.05008f
C9505 XThR.Tn[13].t23 VGND 0.01867f
C9506 XThR.Tn[13].t54 VGND 0.02044f
C9507 XThR.Tn[13].n74 VGND 0.05211f
C9508 XThR.Tn[13].n75 VGND 0.03661f
C9509 XThR.Tn[13].n76 VGND 0.00669f
C9510 XThR.Tn[13].n77 VGND 0.11748f
C9511 XThR.Tn[13].t42 VGND 0.01873f
C9512 XThR.Tn[13].t56 VGND 0.02051f
C9513 XThR.Tn[13].n78 VGND 0.05008f
C9514 XThR.Tn[13].t61 VGND 0.01867f
C9515 XThR.Tn[13].t47 VGND 0.02044f
C9516 XThR.Tn[13].n79 VGND 0.05211f
C9517 XThR.Tn[13].n80 VGND 0.03661f
C9518 XThR.Tn[13].n81 VGND 0.00669f
C9519 XThR.Tn[13].n82 VGND 0.11748f
C9520 XThR.Tn[13].n83 VGND 0.10676f
C9521 XThR.Tn[13].n84 VGND 0.41858f
C9522 XThR.Tn[13].t2 VGND 0.02397f
C9523 XThR.Tn[13].t0 VGND 0.02397f
C9524 XThR.Tn[13].n85 VGND 0.05178f
C9525 XThR.Tn[13].t3 VGND 0.02397f
C9526 XThR.Tn[13].t1 VGND 0.02397f
C9527 XThR.Tn[13].n86 VGND 0.07881f
C9528 XThR.Tn[13].n87 VGND 0.21883f
C9529 XThR.Tn[13].n88 VGND 0.0293f
C9530 XThC.TB3.t1 VGND 0.06296f
C9531 XThC.TB3.n0 VGND 0.04069f
C9532 XThC.TB3.n1 VGND 0.05192f
C9533 XThC.TB3.t2 VGND 0.03159f
C9534 XThC.TB3.t0 VGND 0.03159f
C9535 XThC.TB3.n2 VGND 0.06782f
C9536 XThC.TB3.t10 VGND 0.04914f
C9537 XThC.TB3.t17 VGND 0.02896f
C9538 XThC.TB3.n3 VGND 0.05852f
C9539 XThC.TB3.t14 VGND 0.04914f
C9540 XThC.TB3.t5 VGND 0.02896f
C9541 XThC.TB3.n4 VGND 0.03012f
C9542 XThC.TB3.t15 VGND 0.04914f
C9543 XThC.TB3.t6 VGND 0.02896f
C9544 XThC.TB3.n5 VGND 0.06469f
C9545 XThC.TB3.t3 VGND 0.04914f
C9546 XThC.TB3.t9 VGND 0.02896f
C9547 XThC.TB3.n6 VGND 0.06006f
C9548 XThC.TB3.n7 VGND 0.03654f
C9549 XThC.TB3.n8 VGND 0.06049f
C9550 XThC.TB3.n9 VGND 0.0234f
C9551 XThC.TB3.n10 VGND 0.02857f
C9552 XThC.TB3.n11 VGND 0.06469f
C9553 XThC.TB3.n12 VGND 0.03243f
C9554 XThC.TB3.n13 VGND 0.05514f
C9555 XThC.TB3.t16 VGND 0.04914f
C9556 XThC.TB3.t7 VGND 0.02896f
C9557 XThC.TB3.n14 VGND 0.06624f
C9558 XThC.TB3.t4 VGND 0.04914f
C9559 XThC.TB3.t13 VGND 0.02896f
C9560 XThC.TB3.t12 VGND 0.04914f
C9561 XThC.TB3.t18 VGND 0.02896f
C9562 XThC.TB3.t11 VGND 0.04914f
C9563 XThC.TB3.t8 VGND 0.02896f
C9564 XThC.TB3.n15 VGND 0.08245f
C9565 XThC.TB3.n16 VGND 0.08709f
C9566 XThC.TB3.n17 VGND 0.03356f
C9567 XThC.TB3.n18 VGND 0.07087f
C9568 XThC.TB3.n19 VGND 0.03243f
C9569 XThC.TB3.n20 VGND 0.02691f
C9570 XThC.TB3.n21 VGND 0.27459f
C9571 XThC.TB3.n22 VGND 0.14933f
C9572 XThR.Tn[8].t10 VGND 0.02415f
C9573 XThR.Tn[8].t8 VGND 0.02415f
C9574 XThR.Tn[8].n0 VGND 0.07334f
C9575 XThR.Tn[8].t11 VGND 0.02415f
C9576 XThR.Tn[8].t9 VGND 0.02415f
C9577 XThR.Tn[8].n1 VGND 0.05369f
C9578 XThR.Tn[8].n2 VGND 0.24415f
C9579 XThR.Tn[8].t1 VGND 0.0157f
C9580 XThR.Tn[8].t3 VGND 0.0157f
C9581 XThR.Tn[8].n3 VGND 0.03916f
C9582 XThR.Tn[8].t2 VGND 0.0157f
C9583 XThR.Tn[8].t4 VGND 0.0157f
C9584 XThR.Tn[8].n4 VGND 0.0314f
C9585 XThR.Tn[8].n5 VGND 0.07241f
C9586 XThR.Tn[8].t39 VGND 0.01888f
C9587 XThR.Tn[8].t33 VGND 0.02067f
C9588 XThR.Tn[8].n6 VGND 0.05048f
C9589 XThR.Tn[8].n7 VGND 0.09697f
C9590 XThR.Tn[8].t59 VGND 0.01888f
C9591 XThR.Tn[8].t49 VGND 0.02067f
C9592 XThR.Tn[8].n8 VGND 0.05048f
C9593 XThR.Tn[8].t13 VGND 0.01882f
C9594 XThR.Tn[8].t45 VGND 0.02061f
C9595 XThR.Tn[8].n9 VGND 0.05252f
C9596 XThR.Tn[8].n10 VGND 0.0369f
C9597 XThR.Tn[8].n11 VGND 0.00675f
C9598 XThR.Tn[8].n12 VGND 0.11841f
C9599 XThR.Tn[8].t34 VGND 0.01888f
C9600 XThR.Tn[8].t26 VGND 0.02067f
C9601 XThR.Tn[8].n13 VGND 0.05048f
C9602 XThR.Tn[8].t53 VGND 0.01882f
C9603 XThR.Tn[8].t22 VGND 0.02061f
C9604 XThR.Tn[8].n14 VGND 0.05252f
C9605 XThR.Tn[8].n15 VGND 0.0369f
C9606 XThR.Tn[8].n16 VGND 0.00675f
C9607 XThR.Tn[8].n17 VGND 0.11841f
C9608 XThR.Tn[8].t50 VGND 0.01888f
C9609 XThR.Tn[8].t43 VGND 0.02067f
C9610 XThR.Tn[8].n18 VGND 0.05048f
C9611 XThR.Tn[8].t65 VGND 0.01882f
C9612 XThR.Tn[8].t40 VGND 0.02061f
C9613 XThR.Tn[8].n19 VGND 0.05252f
C9614 XThR.Tn[8].n20 VGND 0.0369f
C9615 XThR.Tn[8].n21 VGND 0.00675f
C9616 XThR.Tn[8].n22 VGND 0.11841f
C9617 XThR.Tn[8].t12 VGND 0.01888f
C9618 XThR.Tn[8].t70 VGND 0.02067f
C9619 XThR.Tn[8].n23 VGND 0.05048f
C9620 XThR.Tn[8].t36 VGND 0.01882f
C9621 XThR.Tn[8].t66 VGND 0.02061f
C9622 XThR.Tn[8].n24 VGND 0.05252f
C9623 XThR.Tn[8].n25 VGND 0.0369f
C9624 XThR.Tn[8].n26 VGND 0.00675f
C9625 XThR.Tn[8].n27 VGND 0.11841f
C9626 XThR.Tn[8].t52 VGND 0.01888f
C9627 XThR.Tn[8].t44 VGND 0.02067f
C9628 XThR.Tn[8].n28 VGND 0.05048f
C9629 XThR.Tn[8].t68 VGND 0.01882f
C9630 XThR.Tn[8].t41 VGND 0.02061f
C9631 XThR.Tn[8].n29 VGND 0.05252f
C9632 XThR.Tn[8].n30 VGND 0.0369f
C9633 XThR.Tn[8].n31 VGND 0.00675f
C9634 XThR.Tn[8].n32 VGND 0.11841f
C9635 XThR.Tn[8].t28 VGND 0.01888f
C9636 XThR.Tn[8].t61 VGND 0.02067f
C9637 XThR.Tn[8].n33 VGND 0.05048f
C9638 XThR.Tn[8].t47 VGND 0.01882f
C9639 XThR.Tn[8].t58 VGND 0.02061f
C9640 XThR.Tn[8].n34 VGND 0.05252f
C9641 XThR.Tn[8].n35 VGND 0.0369f
C9642 XThR.Tn[8].n36 VGND 0.00675f
C9643 XThR.Tn[8].n37 VGND 0.11841f
C9644 XThR.Tn[8].t60 VGND 0.01888f
C9645 XThR.Tn[8].t56 VGND 0.02067f
C9646 XThR.Tn[8].n38 VGND 0.05048f
C9647 XThR.Tn[8].t14 VGND 0.01882f
C9648 XThR.Tn[8].t51 VGND 0.02061f
C9649 XThR.Tn[8].n39 VGND 0.05252f
C9650 XThR.Tn[8].n40 VGND 0.0369f
C9651 XThR.Tn[8].n41 VGND 0.00675f
C9652 XThR.Tn[8].n42 VGND 0.11841f
C9653 XThR.Tn[8].t63 VGND 0.01888f
C9654 XThR.Tn[8].t69 VGND 0.02067f
C9655 XThR.Tn[8].n43 VGND 0.05048f
C9656 XThR.Tn[8].t20 VGND 0.01882f
C9657 XThR.Tn[8].t64 VGND 0.02061f
C9658 XThR.Tn[8].n44 VGND 0.05252f
C9659 XThR.Tn[8].n45 VGND 0.0369f
C9660 XThR.Tn[8].n46 VGND 0.00675f
C9661 XThR.Tn[8].n47 VGND 0.11841f
C9662 XThR.Tn[8].t17 VGND 0.01888f
C9663 XThR.Tn[8].t27 VGND 0.02067f
C9664 XThR.Tn[8].n48 VGND 0.05048f
C9665 XThR.Tn[8].t38 VGND 0.01882f
C9666 XThR.Tn[8].t24 VGND 0.02061f
C9667 XThR.Tn[8].n49 VGND 0.05252f
C9668 XThR.Tn[8].n50 VGND 0.0369f
C9669 XThR.Tn[8].n51 VGND 0.00675f
C9670 XThR.Tn[8].n52 VGND 0.11841f
C9671 XThR.Tn[8].t72 VGND 0.01888f
C9672 XThR.Tn[8].t46 VGND 0.02067f
C9673 XThR.Tn[8].n53 VGND 0.05048f
C9674 XThR.Tn[8].t31 VGND 0.01882f
C9675 XThR.Tn[8].t42 VGND 0.02061f
C9676 XThR.Tn[8].n54 VGND 0.05252f
C9677 XThR.Tn[8].n55 VGND 0.0369f
C9678 XThR.Tn[8].n56 VGND 0.00675f
C9679 XThR.Tn[8].n57 VGND 0.11841f
C9680 XThR.Tn[8].t30 VGND 0.01888f
C9681 XThR.Tn[8].t21 VGND 0.02067f
C9682 XThR.Tn[8].n58 VGND 0.05048f
C9683 XThR.Tn[8].t48 VGND 0.01882f
C9684 XThR.Tn[8].t16 VGND 0.02061f
C9685 XThR.Tn[8].n59 VGND 0.05252f
C9686 XThR.Tn[8].n60 VGND 0.0369f
C9687 XThR.Tn[8].n61 VGND 0.00675f
C9688 XThR.Tn[8].n62 VGND 0.11841f
C9689 XThR.Tn[8].t62 VGND 0.01888f
C9690 XThR.Tn[8].t57 VGND 0.02067f
C9691 XThR.Tn[8].n63 VGND 0.05048f
C9692 XThR.Tn[8].t18 VGND 0.01882f
C9693 XThR.Tn[8].t54 VGND 0.02061f
C9694 XThR.Tn[8].n64 VGND 0.05252f
C9695 XThR.Tn[8].n65 VGND 0.0369f
C9696 XThR.Tn[8].n66 VGND 0.00675f
C9697 XThR.Tn[8].n67 VGND 0.11841f
C9698 XThR.Tn[8].t15 VGND 0.01888f
C9699 XThR.Tn[8].t71 VGND 0.02067f
C9700 XThR.Tn[8].n68 VGND 0.05048f
C9701 XThR.Tn[8].t37 VGND 0.01882f
C9702 XThR.Tn[8].t67 VGND 0.02061f
C9703 XThR.Tn[8].n69 VGND 0.05252f
C9704 XThR.Tn[8].n70 VGND 0.0369f
C9705 XThR.Tn[8].n71 VGND 0.00675f
C9706 XThR.Tn[8].n72 VGND 0.11841f
C9707 XThR.Tn[8].t35 VGND 0.01888f
C9708 XThR.Tn[8].t29 VGND 0.02067f
C9709 XThR.Tn[8].n73 VGND 0.05048f
C9710 XThR.Tn[8].t55 VGND 0.01882f
C9711 XThR.Tn[8].t25 VGND 0.02061f
C9712 XThR.Tn[8].n74 VGND 0.05252f
C9713 XThR.Tn[8].n75 VGND 0.0369f
C9714 XThR.Tn[8].n76 VGND 0.00675f
C9715 XThR.Tn[8].n77 VGND 0.11841f
C9716 XThR.Tn[8].t73 VGND 0.01888f
C9717 XThR.Tn[8].t23 VGND 0.02067f
C9718 XThR.Tn[8].n78 VGND 0.05048f
C9719 XThR.Tn[8].t32 VGND 0.01882f
C9720 XThR.Tn[8].t19 VGND 0.02061f
C9721 XThR.Tn[8].n79 VGND 0.05252f
C9722 XThR.Tn[8].n80 VGND 0.0369f
C9723 XThR.Tn[8].n81 VGND 0.00675f
C9724 XThR.Tn[8].n82 VGND 0.11841f
C9725 XThR.Tn[8].n83 VGND 0.10761f
C9726 XThR.Tn[8].n84 VGND 0.32972f
C9727 XThR.Tn[8].t6 VGND 0.02415f
C9728 XThR.Tn[8].t0 VGND 0.02415f
C9729 XThR.Tn[8].n85 VGND 0.05219f
C9730 XThR.Tn[8].t5 VGND 0.02415f
C9731 XThR.Tn[8].t7 VGND 0.02415f
C9732 XThR.Tn[8].n86 VGND 0.07943f
C9733 XThR.Tn[8].n87 VGND 0.22055f
C9734 XThR.Tn[8].n88 VGND 0.01087f
C9735 XThR.Tn[0].t6 VGND 0.02293f
C9736 XThR.Tn[0].t7 VGND 0.02293f
C9737 XThR.Tn[0].n0 VGND 0.04628f
C9738 XThR.Tn[0].t5 VGND 0.02293f
C9739 XThR.Tn[0].t4 VGND 0.02293f
C9740 XThR.Tn[0].n1 VGND 0.05416f
C9741 XThR.Tn[0].n2 VGND 0.16245f
C9742 XThR.Tn[0].t9 VGND 0.0149f
C9743 XThR.Tn[0].t10 VGND 0.0149f
C9744 XThR.Tn[0].n3 VGND 0.03394f
C9745 XThR.Tn[0].t8 VGND 0.0149f
C9746 XThR.Tn[0].t11 VGND 0.0149f
C9747 XThR.Tn[0].n4 VGND 0.03394f
C9748 XThR.Tn[0].t3 VGND 0.0149f
C9749 XThR.Tn[0].t2 VGND 0.0149f
C9750 XThR.Tn[0].n5 VGND 0.05655f
C9751 XThR.Tn[0].t0 VGND 0.0149f
C9752 XThR.Tn[0].t1 VGND 0.0149f
C9753 XThR.Tn[0].n6 VGND 0.03394f
C9754 XThR.Tn[0].n7 VGND 0.16164f
C9755 XThR.Tn[0].n8 VGND 0.09992f
C9756 XThR.Tn[0].n9 VGND 0.11277f
C9757 XThR.Tn[0].t48 VGND 0.01792f
C9758 XThR.Tn[0].t40 VGND 0.01962f
C9759 XThR.Tn[0].n10 VGND 0.04792f
C9760 XThR.Tn[0].n11 VGND 0.09205f
C9761 XThR.Tn[0].t67 VGND 0.01792f
C9762 XThR.Tn[0].t58 VGND 0.01962f
C9763 XThR.Tn[0].n12 VGND 0.04792f
C9764 XThR.Tn[0].t24 VGND 0.01786f
C9765 XThR.Tn[0].t50 VGND 0.01956f
C9766 XThR.Tn[0].n13 VGND 0.04986f
C9767 XThR.Tn[0].n14 VGND 0.03503f
C9768 XThR.Tn[0].n15 VGND 0.0064f
C9769 XThR.Tn[0].n16 VGND 0.11241f
C9770 XThR.Tn[0].t41 VGND 0.01792f
C9771 XThR.Tn[0].t33 VGND 0.01962f
C9772 XThR.Tn[0].n17 VGND 0.04792f
C9773 XThR.Tn[0].t61 VGND 0.01786f
C9774 XThR.Tn[0].t26 VGND 0.01956f
C9775 XThR.Tn[0].n18 VGND 0.04986f
C9776 XThR.Tn[0].n19 VGND 0.03503f
C9777 XThR.Tn[0].n20 VGND 0.0064f
C9778 XThR.Tn[0].n21 VGND 0.11241f
C9779 XThR.Tn[0].t59 VGND 0.01792f
C9780 XThR.Tn[0].t51 VGND 0.01962f
C9781 XThR.Tn[0].n22 VGND 0.04792f
C9782 XThR.Tn[0].t12 VGND 0.01786f
C9783 XThR.Tn[0].t44 VGND 0.01956f
C9784 XThR.Tn[0].n23 VGND 0.04986f
C9785 XThR.Tn[0].n24 VGND 0.03503f
C9786 XThR.Tn[0].n25 VGND 0.0064f
C9787 XThR.Tn[0].n26 VGND 0.11241f
C9788 XThR.Tn[0].t21 VGND 0.01792f
C9789 XThR.Tn[0].t15 VGND 0.01962f
C9790 XThR.Tn[0].n27 VGND 0.04792f
C9791 XThR.Tn[0].t43 VGND 0.01786f
C9792 XThR.Tn[0].t72 VGND 0.01956f
C9793 XThR.Tn[0].n28 VGND 0.04986f
C9794 XThR.Tn[0].n29 VGND 0.03503f
C9795 XThR.Tn[0].n30 VGND 0.0064f
C9796 XThR.Tn[0].n31 VGND 0.11241f
C9797 XThR.Tn[0].t60 VGND 0.01792f
C9798 XThR.Tn[0].t52 VGND 0.01962f
C9799 XThR.Tn[0].n32 VGND 0.04792f
C9800 XThR.Tn[0].t13 VGND 0.01786f
C9801 XThR.Tn[0].t46 VGND 0.01956f
C9802 XThR.Tn[0].n33 VGND 0.04986f
C9803 XThR.Tn[0].n34 VGND 0.03503f
C9804 XThR.Tn[0].n35 VGND 0.0064f
C9805 XThR.Tn[0].n36 VGND 0.11241f
C9806 XThR.Tn[0].t35 VGND 0.01792f
C9807 XThR.Tn[0].t68 VGND 0.01962f
C9808 XThR.Tn[0].n37 VGND 0.04792f
C9809 XThR.Tn[0].t54 VGND 0.01786f
C9810 XThR.Tn[0].t64 VGND 0.01956f
C9811 XThR.Tn[0].n38 VGND 0.04986f
C9812 XThR.Tn[0].n39 VGND 0.03503f
C9813 XThR.Tn[0].n40 VGND 0.0064f
C9814 XThR.Tn[0].n41 VGND 0.11241f
C9815 XThR.Tn[0].t66 VGND 0.01792f
C9816 XThR.Tn[0].t63 VGND 0.01962f
C9817 XThR.Tn[0].n42 VGND 0.04792f
C9818 XThR.Tn[0].t23 VGND 0.01786f
C9819 XThR.Tn[0].t55 VGND 0.01956f
C9820 XThR.Tn[0].n43 VGND 0.04986f
C9821 XThR.Tn[0].n44 VGND 0.03503f
C9822 XThR.Tn[0].n45 VGND 0.0064f
C9823 XThR.Tn[0].n46 VGND 0.11241f
C9824 XThR.Tn[0].t70 VGND 0.01792f
C9825 XThR.Tn[0].t14 VGND 0.01962f
C9826 XThR.Tn[0].n47 VGND 0.04792f
C9827 XThR.Tn[0].t28 VGND 0.01786f
C9828 XThR.Tn[0].t71 VGND 0.01956f
C9829 XThR.Tn[0].n48 VGND 0.04986f
C9830 XThR.Tn[0].n49 VGND 0.03503f
C9831 XThR.Tn[0].n50 VGND 0.0064f
C9832 XThR.Tn[0].n51 VGND 0.11241f
C9833 XThR.Tn[0].t25 VGND 0.01792f
C9834 XThR.Tn[0].t34 VGND 0.01962f
C9835 XThR.Tn[0].n52 VGND 0.04792f
C9836 XThR.Tn[0].t47 VGND 0.01786f
C9837 XThR.Tn[0].t29 VGND 0.01956f
C9838 XThR.Tn[0].n53 VGND 0.04986f
C9839 XThR.Tn[0].n54 VGND 0.03503f
C9840 XThR.Tn[0].n55 VGND 0.0064f
C9841 XThR.Tn[0].n56 VGND 0.11241f
C9842 XThR.Tn[0].t17 VGND 0.01792f
C9843 XThR.Tn[0].t53 VGND 0.01962f
C9844 XThR.Tn[0].n57 VGND 0.04792f
C9845 XThR.Tn[0].t38 VGND 0.01786f
C9846 XThR.Tn[0].t49 VGND 0.01956f
C9847 XThR.Tn[0].n58 VGND 0.04986f
C9848 XThR.Tn[0].n59 VGND 0.03503f
C9849 XThR.Tn[0].n60 VGND 0.0064f
C9850 XThR.Tn[0].n61 VGND 0.11241f
C9851 XThR.Tn[0].t37 VGND 0.01792f
C9852 XThR.Tn[0].t31 VGND 0.01962f
C9853 XThR.Tn[0].n62 VGND 0.04792f
C9854 XThR.Tn[0].t56 VGND 0.01786f
C9855 XThR.Tn[0].t19 VGND 0.01956f
C9856 XThR.Tn[0].n63 VGND 0.04986f
C9857 XThR.Tn[0].n64 VGND 0.03503f
C9858 XThR.Tn[0].n65 VGND 0.0064f
C9859 XThR.Tn[0].n66 VGND 0.11241f
C9860 XThR.Tn[0].t69 VGND 0.01792f
C9861 XThR.Tn[0].t65 VGND 0.01962f
C9862 XThR.Tn[0].n67 VGND 0.04792f
C9863 XThR.Tn[0].t27 VGND 0.01786f
C9864 XThR.Tn[0].t57 VGND 0.01956f
C9865 XThR.Tn[0].n68 VGND 0.04986f
C9866 XThR.Tn[0].n69 VGND 0.03503f
C9867 XThR.Tn[0].n70 VGND 0.0064f
C9868 XThR.Tn[0].n71 VGND 0.11241f
C9869 XThR.Tn[0].t22 VGND 0.01792f
C9870 XThR.Tn[0].t16 VGND 0.01962f
C9871 XThR.Tn[0].n72 VGND 0.04792f
C9872 XThR.Tn[0].t45 VGND 0.01786f
C9873 XThR.Tn[0].t73 VGND 0.01956f
C9874 XThR.Tn[0].n73 VGND 0.04986f
C9875 XThR.Tn[0].n74 VGND 0.03503f
C9876 XThR.Tn[0].n75 VGND 0.0064f
C9877 XThR.Tn[0].n76 VGND 0.11241f
C9878 XThR.Tn[0].t42 VGND 0.01792f
C9879 XThR.Tn[0].t36 VGND 0.01962f
C9880 XThR.Tn[0].n77 VGND 0.04792f
C9881 XThR.Tn[0].t62 VGND 0.01786f
C9882 XThR.Tn[0].t30 VGND 0.01956f
C9883 XThR.Tn[0].n78 VGND 0.04986f
C9884 XThR.Tn[0].n79 VGND 0.03503f
C9885 XThR.Tn[0].n80 VGND 0.0064f
C9886 XThR.Tn[0].n81 VGND 0.11241f
C9887 XThR.Tn[0].t18 VGND 0.01792f
C9888 XThR.Tn[0].t32 VGND 0.01962f
C9889 XThR.Tn[0].n82 VGND 0.04792f
C9890 XThR.Tn[0].t39 VGND 0.01786f
C9891 XThR.Tn[0].t20 VGND 0.01956f
C9892 XThR.Tn[0].n83 VGND 0.04986f
C9893 XThR.Tn[0].n84 VGND 0.03503f
C9894 XThR.Tn[0].n85 VGND 0.0064f
C9895 XThR.Tn[0].n86 VGND 0.11241f
C9896 XThR.Tn[0].n87 VGND 0.10215f
C9897 XThR.Tn[0].n88 VGND 0.29249f
C9898 XThR.Tn[7].t2 VGND 0.01503f
C9899 XThR.Tn[7].t1 VGND 0.01503f
C9900 XThR.Tn[7].n0 VGND 0.03319f
C9901 XThR.Tn[7].t3 VGND 0.01503f
C9902 XThR.Tn[7].t0 VGND 0.01503f
C9903 XThR.Tn[7].n1 VGND 0.04638f
C9904 XThR.Tn[7].n2 VGND 0.17022f
C9905 XThR.Tn[7].t6 VGND 0.02312f
C9906 XThR.Tn[7].t7 VGND 0.02312f
C9907 XThR.Tn[7].n3 VGND 0.0704f
C9908 XThR.Tn[7].t5 VGND 0.02312f
C9909 XThR.Tn[7].t4 VGND 0.02312f
C9910 XThR.Tn[7].n4 VGND 0.05122f
C9911 XThR.Tn[7].n5 VGND 0.22538f
C9912 XThR.Tn[7].n6 VGND 0.02808f
C9913 XThR.Tn[7].t53 VGND 0.01807f
C9914 XThR.Tn[7].t45 VGND 0.01979f
C9915 XThR.Tn[7].n7 VGND 0.04832f
C9916 XThR.Tn[7].n8 VGND 0.09282f
C9917 XThR.Tn[7].t8 VGND 0.01807f
C9918 XThR.Tn[7].t60 VGND 0.01979f
C9919 XThR.Tn[7].n9 VGND 0.04832f
C9920 XThR.Tn[7].t26 VGND 0.01801f
C9921 XThR.Tn[7].t38 VGND 0.01972f
C9922 XThR.Tn[7].n10 VGND 0.05027f
C9923 XThR.Tn[7].n11 VGND 0.03532f
C9924 XThR.Tn[7].n12 VGND 0.00646f
C9925 XThR.Tn[7].n13 VGND 0.11334f
C9926 XThR.Tn[7].t47 VGND 0.01807f
C9927 XThR.Tn[7].t37 VGND 0.01979f
C9928 XThR.Tn[7].n14 VGND 0.04832f
C9929 XThR.Tn[7].t66 VGND 0.01801f
C9930 XThR.Tn[7].t15 VGND 0.01972f
C9931 XThR.Tn[7].n15 VGND 0.05027f
C9932 XThR.Tn[7].n16 VGND 0.03532f
C9933 XThR.Tn[7].n17 VGND 0.00646f
C9934 XThR.Tn[7].n18 VGND 0.11334f
C9935 XThR.Tn[7].t62 VGND 0.01807f
C9936 XThR.Tn[7].t55 VGND 0.01979f
C9937 XThR.Tn[7].n19 VGND 0.04832f
C9938 XThR.Tn[7].t18 VGND 0.01801f
C9939 XThR.Tn[7].t32 VGND 0.01972f
C9940 XThR.Tn[7].n20 VGND 0.05027f
C9941 XThR.Tn[7].n21 VGND 0.03532f
C9942 XThR.Tn[7].n22 VGND 0.00646f
C9943 XThR.Tn[7].n23 VGND 0.11334f
C9944 XThR.Tn[7].t25 VGND 0.01807f
C9945 XThR.Tn[7].t21 VGND 0.01979f
C9946 XThR.Tn[7].n24 VGND 0.04832f
C9947 XThR.Tn[7].t50 VGND 0.01801f
C9948 XThR.Tn[7].t63 VGND 0.01972f
C9949 XThR.Tn[7].n25 VGND 0.05027f
C9950 XThR.Tn[7].n26 VGND 0.03532f
C9951 XThR.Tn[7].n27 VGND 0.00646f
C9952 XThR.Tn[7].n28 VGND 0.11334f
C9953 XThR.Tn[7].t65 VGND 0.01807f
C9954 XThR.Tn[7].t56 VGND 0.01979f
C9955 XThR.Tn[7].n29 VGND 0.04832f
C9956 XThR.Tn[7].t19 VGND 0.01801f
C9957 XThR.Tn[7].t34 VGND 0.01972f
C9958 XThR.Tn[7].n30 VGND 0.05027f
C9959 XThR.Tn[7].n31 VGND 0.03532f
C9960 XThR.Tn[7].n32 VGND 0.00646f
C9961 XThR.Tn[7].n33 VGND 0.11334f
C9962 XThR.Tn[7].t40 VGND 0.01807f
C9963 XThR.Tn[7].t11 VGND 0.01979f
C9964 XThR.Tn[7].n34 VGND 0.04832f
C9965 XThR.Tn[7].t58 VGND 0.01801f
C9966 XThR.Tn[7].t54 VGND 0.01972f
C9967 XThR.Tn[7].n35 VGND 0.05027f
C9968 XThR.Tn[7].n36 VGND 0.03532f
C9969 XThR.Tn[7].n37 VGND 0.00646f
C9970 XThR.Tn[7].n38 VGND 0.11334f
C9971 XThR.Tn[7].t9 VGND 0.01807f
C9972 XThR.Tn[7].t68 VGND 0.01979f
C9973 XThR.Tn[7].n39 VGND 0.04832f
C9974 XThR.Tn[7].t27 VGND 0.01801f
C9975 XThR.Tn[7].t46 VGND 0.01972f
C9976 XThR.Tn[7].n40 VGND 0.05027f
C9977 XThR.Tn[7].n41 VGND 0.03532f
C9978 XThR.Tn[7].n42 VGND 0.00646f
C9979 XThR.Tn[7].n43 VGND 0.11334f
C9980 XThR.Tn[7].t14 VGND 0.01807f
C9981 XThR.Tn[7].t20 VGND 0.01979f
C9982 XThR.Tn[7].n44 VGND 0.04832f
C9983 XThR.Tn[7].t31 VGND 0.01801f
C9984 XThR.Tn[7].t61 VGND 0.01972f
C9985 XThR.Tn[7].n45 VGND 0.05027f
C9986 XThR.Tn[7].n46 VGND 0.03532f
C9987 XThR.Tn[7].n47 VGND 0.00646f
C9988 XThR.Tn[7].n48 VGND 0.11334f
C9989 XThR.Tn[7].t29 VGND 0.01807f
C9990 XThR.Tn[7].t39 VGND 0.01979f
C9991 XThR.Tn[7].n49 VGND 0.04832f
C9992 XThR.Tn[7].t52 VGND 0.01801f
C9993 XThR.Tn[7].t16 VGND 0.01972f
C9994 XThR.Tn[7].n50 VGND 0.05027f
C9995 XThR.Tn[7].n51 VGND 0.03532f
C9996 XThR.Tn[7].n52 VGND 0.00646f
C9997 XThR.Tn[7].n53 VGND 0.11334f
C9998 XThR.Tn[7].t23 VGND 0.01807f
C9999 XThR.Tn[7].t57 VGND 0.01979f
C10000 XThR.Tn[7].n54 VGND 0.04832f
C10001 XThR.Tn[7].t43 VGND 0.01801f
C10002 XThR.Tn[7].t36 VGND 0.01972f
C10003 XThR.Tn[7].n55 VGND 0.05027f
C10004 XThR.Tn[7].n56 VGND 0.03532f
C10005 XThR.Tn[7].n57 VGND 0.00646f
C10006 XThR.Tn[7].n58 VGND 0.11334f
C10007 XThR.Tn[7].t42 VGND 0.01807f
C10008 XThR.Tn[7].t33 VGND 0.01979f
C10009 XThR.Tn[7].n59 VGND 0.04832f
C10010 XThR.Tn[7].t59 VGND 0.01801f
C10011 XThR.Tn[7].t10 VGND 0.01972f
C10012 XThR.Tn[7].n60 VGND 0.05027f
C10013 XThR.Tn[7].n61 VGND 0.03532f
C10014 XThR.Tn[7].n62 VGND 0.00646f
C10015 XThR.Tn[7].n63 VGND 0.11334f
C10016 XThR.Tn[7].t12 VGND 0.01807f
C10017 XThR.Tn[7].t69 VGND 0.01979f
C10018 XThR.Tn[7].n64 VGND 0.04832f
C10019 XThR.Tn[7].t30 VGND 0.01801f
C10020 XThR.Tn[7].t48 VGND 0.01972f
C10021 XThR.Tn[7].n65 VGND 0.05027f
C10022 XThR.Tn[7].n66 VGND 0.03532f
C10023 XThR.Tn[7].n67 VGND 0.00646f
C10024 XThR.Tn[7].n68 VGND 0.11334f
C10025 XThR.Tn[7].t28 VGND 0.01807f
C10026 XThR.Tn[7].t22 VGND 0.01979f
C10027 XThR.Tn[7].n69 VGND 0.04832f
C10028 XThR.Tn[7].t51 VGND 0.01801f
C10029 XThR.Tn[7].t64 VGND 0.01972f
C10030 XThR.Tn[7].n70 VGND 0.05027f
C10031 XThR.Tn[7].n71 VGND 0.03532f
C10032 XThR.Tn[7].n72 VGND 0.00646f
C10033 XThR.Tn[7].n73 VGND 0.11334f
C10034 XThR.Tn[7].t49 VGND 0.01807f
C10035 XThR.Tn[7].t41 VGND 0.01979f
C10036 XThR.Tn[7].n74 VGND 0.04832f
C10037 XThR.Tn[7].t67 VGND 0.01801f
C10038 XThR.Tn[7].t17 VGND 0.01972f
C10039 XThR.Tn[7].n75 VGND 0.05027f
C10040 XThR.Tn[7].n76 VGND 0.03532f
C10041 XThR.Tn[7].n77 VGND 0.00646f
C10042 XThR.Tn[7].n78 VGND 0.11334f
C10043 XThR.Tn[7].t24 VGND 0.01807f
C10044 XThR.Tn[7].t35 VGND 0.01979f
C10045 XThR.Tn[7].n79 VGND 0.04832f
C10046 XThR.Tn[7].t44 VGND 0.01801f
C10047 XThR.Tn[7].t13 VGND 0.01972f
C10048 XThR.Tn[7].n80 VGND 0.05027f
C10049 XThR.Tn[7].n81 VGND 0.03532f
C10050 XThR.Tn[7].n82 VGND 0.00646f
C10051 XThR.Tn[7].n83 VGND 0.11334f
C10052 XThR.Tn[7].n84 VGND 0.103f
C10053 XThR.Tn[7].n85 VGND 0.41812f
C10054 XThR.Tn[11].t2 VGND 0.01567f
C10055 XThR.Tn[11].t0 VGND 0.01567f
C10056 XThR.Tn[11].n0 VGND 0.03134f
C10057 XThR.Tn[11].t3 VGND 0.01567f
C10058 XThR.Tn[11].t1 VGND 0.01567f
C10059 XThR.Tn[11].n1 VGND 0.03908f
C10060 XThR.Tn[11].n2 VGND 0.07883f
C10061 XThR.Tn[11].t8 VGND 0.0241f
C10062 XThR.Tn[11].t10 VGND 0.0241f
C10063 XThR.Tn[11].n3 VGND 0.07319f
C10064 XThR.Tn[11].t9 VGND 0.0241f
C10065 XThR.Tn[11].t11 VGND 0.0241f
C10066 XThR.Tn[11].n4 VGND 0.05358f
C10067 XThR.Tn[11].n5 VGND 0.24365f
C10068 XThR.Tn[11].t4 VGND 0.0241f
C10069 XThR.Tn[11].t6 VGND 0.0241f
C10070 XThR.Tn[11].n6 VGND 0.05208f
C10071 XThR.Tn[11].t5 VGND 0.0241f
C10072 XThR.Tn[11].t7 VGND 0.0241f
C10073 XThR.Tn[11].n7 VGND 0.07927f
C10074 XThR.Tn[11].n8 VGND 0.2201f
C10075 XThR.Tn[11].n9 VGND 0.02947f
C10076 XThR.Tn[11].t56 VGND 0.01884f
C10077 XThR.Tn[11].t48 VGND 0.02063f
C10078 XThR.Tn[11].n10 VGND 0.05037f
C10079 XThR.Tn[11].n11 VGND 0.09677f
C10080 XThR.Tn[11].t12 VGND 0.01884f
C10081 XThR.Tn[11].t67 VGND 0.02063f
C10082 XThR.Tn[11].n12 VGND 0.05037f
C10083 XThR.Tn[11].t27 VGND 0.01878f
C10084 XThR.Tn[11].t58 VGND 0.02056f
C10085 XThR.Tn[11].n13 VGND 0.05241f
C10086 XThR.Tn[11].n14 VGND 0.03682f
C10087 XThR.Tn[11].n15 VGND 0.00673f
C10088 XThR.Tn[11].n16 VGND 0.11816f
C10089 XThR.Tn[11].t49 VGND 0.01884f
C10090 XThR.Tn[11].t41 VGND 0.02063f
C10091 XThR.Tn[11].n17 VGND 0.05037f
C10092 XThR.Tn[11].t65 VGND 0.01878f
C10093 XThR.Tn[11].t36 VGND 0.02056f
C10094 XThR.Tn[11].n18 VGND 0.05241f
C10095 XThR.Tn[11].n19 VGND 0.03682f
C10096 XThR.Tn[11].n20 VGND 0.00673f
C10097 XThR.Tn[11].n21 VGND 0.11816f
C10098 XThR.Tn[11].t68 VGND 0.01884f
C10099 XThR.Tn[11].t60 VGND 0.02063f
C10100 XThR.Tn[11].n22 VGND 0.05037f
C10101 XThR.Tn[11].t18 VGND 0.01878f
C10102 XThR.Tn[11].t54 VGND 0.02056f
C10103 XThR.Tn[11].n23 VGND 0.05241f
C10104 XThR.Tn[11].n24 VGND 0.03682f
C10105 XThR.Tn[11].n25 VGND 0.00673f
C10106 XThR.Tn[11].n26 VGND 0.11816f
C10107 XThR.Tn[11].t33 VGND 0.01884f
C10108 XThR.Tn[11].t23 VGND 0.02063f
C10109 XThR.Tn[11].n27 VGND 0.05037f
C10110 XThR.Tn[11].t50 VGND 0.01878f
C10111 XThR.Tn[11].t19 VGND 0.02056f
C10112 XThR.Tn[11].n28 VGND 0.05241f
C10113 XThR.Tn[11].n29 VGND 0.03682f
C10114 XThR.Tn[11].n30 VGND 0.00673f
C10115 XThR.Tn[11].n31 VGND 0.11816f
C10116 XThR.Tn[11].t70 VGND 0.01884f
C10117 XThR.Tn[11].t62 VGND 0.02063f
C10118 XThR.Tn[11].n32 VGND 0.05037f
C10119 XThR.Tn[11].t21 VGND 0.01878f
C10120 XThR.Tn[11].t55 VGND 0.02056f
C10121 XThR.Tn[11].n33 VGND 0.05241f
C10122 XThR.Tn[11].n34 VGND 0.03682f
C10123 XThR.Tn[11].n35 VGND 0.00673f
C10124 XThR.Tn[11].n36 VGND 0.11816f
C10125 XThR.Tn[11].t44 VGND 0.01884f
C10126 XThR.Tn[11].t14 VGND 0.02063f
C10127 XThR.Tn[11].n37 VGND 0.05037f
C10128 XThR.Tn[11].t59 VGND 0.01878f
C10129 XThR.Tn[11].t72 VGND 0.02056f
C10130 XThR.Tn[11].n38 VGND 0.05241f
C10131 XThR.Tn[11].n39 VGND 0.03682f
C10132 XThR.Tn[11].n40 VGND 0.00673f
C10133 XThR.Tn[11].n41 VGND 0.11816f
C10134 XThR.Tn[11].t13 VGND 0.01884f
C10135 XThR.Tn[11].t71 VGND 0.02063f
C10136 XThR.Tn[11].n42 VGND 0.05037f
C10137 XThR.Tn[11].t28 VGND 0.01878f
C10138 XThR.Tn[11].t64 VGND 0.02056f
C10139 XThR.Tn[11].n43 VGND 0.05241f
C10140 XThR.Tn[11].n44 VGND 0.03682f
C10141 XThR.Tn[11].n45 VGND 0.00673f
C10142 XThR.Tn[11].n46 VGND 0.11816f
C10143 XThR.Tn[11].t16 VGND 0.01884f
C10144 XThR.Tn[11].t22 VGND 0.02063f
C10145 XThR.Tn[11].n47 VGND 0.05037f
C10146 XThR.Tn[11].t32 VGND 0.01878f
C10147 XThR.Tn[11].t17 VGND 0.02056f
C10148 XThR.Tn[11].n48 VGND 0.05241f
C10149 XThR.Tn[11].n49 VGND 0.03682f
C10150 XThR.Tn[11].n50 VGND 0.00673f
C10151 XThR.Tn[11].n51 VGND 0.11816f
C10152 XThR.Tn[11].t35 VGND 0.01884f
C10153 XThR.Tn[11].t43 VGND 0.02063f
C10154 XThR.Tn[11].n52 VGND 0.05037f
C10155 XThR.Tn[11].t52 VGND 0.01878f
C10156 XThR.Tn[11].t37 VGND 0.02056f
C10157 XThR.Tn[11].n53 VGND 0.05241f
C10158 XThR.Tn[11].n54 VGND 0.03682f
C10159 XThR.Tn[11].n55 VGND 0.00673f
C10160 XThR.Tn[11].n56 VGND 0.11816f
C10161 XThR.Tn[11].t25 VGND 0.01884f
C10162 XThR.Tn[11].t63 VGND 0.02063f
C10163 XThR.Tn[11].n57 VGND 0.05037f
C10164 XThR.Tn[11].t42 VGND 0.01878f
C10165 XThR.Tn[11].t57 VGND 0.02056f
C10166 XThR.Tn[11].n58 VGND 0.05241f
C10167 XThR.Tn[11].n59 VGND 0.03682f
C10168 XThR.Tn[11].n60 VGND 0.00673f
C10169 XThR.Tn[11].n61 VGND 0.11816f
C10170 XThR.Tn[11].t47 VGND 0.01884f
C10171 XThR.Tn[11].t39 VGND 0.02063f
C10172 XThR.Tn[11].n62 VGND 0.05037f
C10173 XThR.Tn[11].t61 VGND 0.01878f
C10174 XThR.Tn[11].t29 VGND 0.02056f
C10175 XThR.Tn[11].n63 VGND 0.05241f
C10176 XThR.Tn[11].n64 VGND 0.03682f
C10177 XThR.Tn[11].n65 VGND 0.00673f
C10178 XThR.Tn[11].n66 VGND 0.11816f
C10179 XThR.Tn[11].t15 VGND 0.01884f
C10180 XThR.Tn[11].t73 VGND 0.02063f
C10181 XThR.Tn[11].n67 VGND 0.05037f
C10182 XThR.Tn[11].t30 VGND 0.01878f
C10183 XThR.Tn[11].t66 VGND 0.02056f
C10184 XThR.Tn[11].n68 VGND 0.05241f
C10185 XThR.Tn[11].n69 VGND 0.03682f
C10186 XThR.Tn[11].n70 VGND 0.00673f
C10187 XThR.Tn[11].n71 VGND 0.11816f
C10188 XThR.Tn[11].t34 VGND 0.01884f
C10189 XThR.Tn[11].t24 VGND 0.02063f
C10190 XThR.Tn[11].n72 VGND 0.05037f
C10191 XThR.Tn[11].t51 VGND 0.01878f
C10192 XThR.Tn[11].t20 VGND 0.02056f
C10193 XThR.Tn[11].n73 VGND 0.05241f
C10194 XThR.Tn[11].n74 VGND 0.03682f
C10195 XThR.Tn[11].n75 VGND 0.00673f
C10196 XThR.Tn[11].n76 VGND 0.11816f
C10197 XThR.Tn[11].t53 VGND 0.01884f
C10198 XThR.Tn[11].t46 VGND 0.02063f
C10199 XThR.Tn[11].n77 VGND 0.05037f
C10200 XThR.Tn[11].t69 VGND 0.01878f
C10201 XThR.Tn[11].t38 VGND 0.02056f
C10202 XThR.Tn[11].n78 VGND 0.05241f
C10203 XThR.Tn[11].n79 VGND 0.03682f
C10204 XThR.Tn[11].n80 VGND 0.00673f
C10205 XThR.Tn[11].n81 VGND 0.11816f
C10206 XThR.Tn[11].t26 VGND 0.01884f
C10207 XThR.Tn[11].t40 VGND 0.02063f
C10208 XThR.Tn[11].n82 VGND 0.05037f
C10209 XThR.Tn[11].t45 VGND 0.01878f
C10210 XThR.Tn[11].t31 VGND 0.02056f
C10211 XThR.Tn[11].n83 VGND 0.05241f
C10212 XThR.Tn[11].n84 VGND 0.03682f
C10213 XThR.Tn[11].n85 VGND 0.00673f
C10214 XThR.Tn[11].n86 VGND 0.11816f
C10215 XThR.Tn[11].n87 VGND 0.10738f
C10216 XThR.Tn[11].n88 VGND 0.38486f
C10217 XThR.Tn[4].t5 VGND 0.02325f
C10218 XThR.Tn[4].t6 VGND 0.02325f
C10219 XThR.Tn[4].n0 VGND 0.04693f
C10220 XThR.Tn[4].t4 VGND 0.02325f
C10221 XThR.Tn[4].t7 VGND 0.02325f
C10222 XThR.Tn[4].n1 VGND 0.05491f
C10223 XThR.Tn[4].n2 VGND 0.16472f
C10224 XThR.Tn[4].t11 VGND 0.01511f
C10225 XThR.Tn[4].t8 VGND 0.01511f
C10226 XThR.Tn[4].n3 VGND 0.03442f
C10227 XThR.Tn[4].t10 VGND 0.01511f
C10228 XThR.Tn[4].t9 VGND 0.01511f
C10229 XThR.Tn[4].n4 VGND 0.03442f
C10230 XThR.Tn[4].t0 VGND 0.01511f
C10231 XThR.Tn[4].t1 VGND 0.01511f
C10232 XThR.Tn[4].n5 VGND 0.05735f
C10233 XThR.Tn[4].t3 VGND 0.01511f
C10234 XThR.Tn[4].t2 VGND 0.01511f
C10235 XThR.Tn[4].n6 VGND 0.03442f
C10236 XThR.Tn[4].n7 VGND 0.1639f
C10237 XThR.Tn[4].n8 VGND 0.10132f
C10238 XThR.Tn[4].n9 VGND 0.11435f
C10239 XThR.Tn[4].t44 VGND 0.01817f
C10240 XThR.Tn[4].t38 VGND 0.0199f
C10241 XThR.Tn[4].n10 VGND 0.04859f
C10242 XThR.Tn[4].n11 VGND 0.09334f
C10243 XThR.Tn[4].t65 VGND 0.01817f
C10244 XThR.Tn[4].t54 VGND 0.0199f
C10245 XThR.Tn[4].n12 VGND 0.04859f
C10246 XThR.Tn[4].t19 VGND 0.01811f
C10247 XThR.Tn[4].t50 VGND 0.01983f
C10248 XThR.Tn[4].n13 VGND 0.05056f
C10249 XThR.Tn[4].n14 VGND 0.03552f
C10250 XThR.Tn[4].n15 VGND 0.00649f
C10251 XThR.Tn[4].n16 VGND 0.11398f
C10252 XThR.Tn[4].t39 VGND 0.01817f
C10253 XThR.Tn[4].t31 VGND 0.0199f
C10254 XThR.Tn[4].n17 VGND 0.04859f
C10255 XThR.Tn[4].t58 VGND 0.01811f
C10256 XThR.Tn[4].t27 VGND 0.01983f
C10257 XThR.Tn[4].n18 VGND 0.05056f
C10258 XThR.Tn[4].n19 VGND 0.03552f
C10259 XThR.Tn[4].n20 VGND 0.00649f
C10260 XThR.Tn[4].n21 VGND 0.11398f
C10261 XThR.Tn[4].t55 VGND 0.01817f
C10262 XThR.Tn[4].t48 VGND 0.0199f
C10263 XThR.Tn[4].n22 VGND 0.04859f
C10264 XThR.Tn[4].t70 VGND 0.01811f
C10265 XThR.Tn[4].t45 VGND 0.01983f
C10266 XThR.Tn[4].n23 VGND 0.05056f
C10267 XThR.Tn[4].n24 VGND 0.03552f
C10268 XThR.Tn[4].n25 VGND 0.00649f
C10269 XThR.Tn[4].n26 VGND 0.11398f
C10270 XThR.Tn[4].t17 VGND 0.01817f
C10271 XThR.Tn[4].t13 VGND 0.0199f
C10272 XThR.Tn[4].n27 VGND 0.04859f
C10273 XThR.Tn[4].t41 VGND 0.01811f
C10274 XThR.Tn[4].t71 VGND 0.01983f
C10275 XThR.Tn[4].n28 VGND 0.05056f
C10276 XThR.Tn[4].n29 VGND 0.03552f
C10277 XThR.Tn[4].n30 VGND 0.00649f
C10278 XThR.Tn[4].n31 VGND 0.11398f
C10279 XThR.Tn[4].t57 VGND 0.01817f
C10280 XThR.Tn[4].t49 VGND 0.0199f
C10281 XThR.Tn[4].n32 VGND 0.04859f
C10282 XThR.Tn[4].t73 VGND 0.01811f
C10283 XThR.Tn[4].t46 VGND 0.01983f
C10284 XThR.Tn[4].n33 VGND 0.05056f
C10285 XThR.Tn[4].n34 VGND 0.03552f
C10286 XThR.Tn[4].n35 VGND 0.00649f
C10287 XThR.Tn[4].n36 VGND 0.11398f
C10288 XThR.Tn[4].t33 VGND 0.01817f
C10289 XThR.Tn[4].t66 VGND 0.0199f
C10290 XThR.Tn[4].n37 VGND 0.04859f
C10291 XThR.Tn[4].t52 VGND 0.01811f
C10292 XThR.Tn[4].t63 VGND 0.01983f
C10293 XThR.Tn[4].n38 VGND 0.05056f
C10294 XThR.Tn[4].n39 VGND 0.03552f
C10295 XThR.Tn[4].n40 VGND 0.00649f
C10296 XThR.Tn[4].n41 VGND 0.11398f
C10297 XThR.Tn[4].t64 VGND 0.01817f
C10298 XThR.Tn[4].t61 VGND 0.0199f
C10299 XThR.Tn[4].n42 VGND 0.04859f
C10300 XThR.Tn[4].t18 VGND 0.01811f
C10301 XThR.Tn[4].t56 VGND 0.01983f
C10302 XThR.Tn[4].n43 VGND 0.05056f
C10303 XThR.Tn[4].n44 VGND 0.03552f
C10304 XThR.Tn[4].n45 VGND 0.00649f
C10305 XThR.Tn[4].n46 VGND 0.11398f
C10306 XThR.Tn[4].t68 VGND 0.01817f
C10307 XThR.Tn[4].t12 VGND 0.0199f
C10308 XThR.Tn[4].n47 VGND 0.04859f
C10309 XThR.Tn[4].t25 VGND 0.01811f
C10310 XThR.Tn[4].t69 VGND 0.01983f
C10311 XThR.Tn[4].n48 VGND 0.05056f
C10312 XThR.Tn[4].n49 VGND 0.03552f
C10313 XThR.Tn[4].n50 VGND 0.00649f
C10314 XThR.Tn[4].n51 VGND 0.11398f
C10315 XThR.Tn[4].t22 VGND 0.01817f
C10316 XThR.Tn[4].t32 VGND 0.0199f
C10317 XThR.Tn[4].n52 VGND 0.04859f
C10318 XThR.Tn[4].t43 VGND 0.01811f
C10319 XThR.Tn[4].t29 VGND 0.01983f
C10320 XThR.Tn[4].n53 VGND 0.05056f
C10321 XThR.Tn[4].n54 VGND 0.03552f
C10322 XThR.Tn[4].n55 VGND 0.00649f
C10323 XThR.Tn[4].n56 VGND 0.11398f
C10324 XThR.Tn[4].t15 VGND 0.01817f
C10325 XThR.Tn[4].t51 VGND 0.0199f
C10326 XThR.Tn[4].n57 VGND 0.04859f
C10327 XThR.Tn[4].t36 VGND 0.01811f
C10328 XThR.Tn[4].t47 VGND 0.01983f
C10329 XThR.Tn[4].n58 VGND 0.05056f
C10330 XThR.Tn[4].n59 VGND 0.03552f
C10331 XThR.Tn[4].n60 VGND 0.00649f
C10332 XThR.Tn[4].n61 VGND 0.11398f
C10333 XThR.Tn[4].t35 VGND 0.01817f
C10334 XThR.Tn[4].t26 VGND 0.0199f
C10335 XThR.Tn[4].n62 VGND 0.04859f
C10336 XThR.Tn[4].t53 VGND 0.01811f
C10337 XThR.Tn[4].t21 VGND 0.01983f
C10338 XThR.Tn[4].n63 VGND 0.05056f
C10339 XThR.Tn[4].n64 VGND 0.03552f
C10340 XThR.Tn[4].n65 VGND 0.00649f
C10341 XThR.Tn[4].n66 VGND 0.11398f
C10342 XThR.Tn[4].t67 VGND 0.01817f
C10343 XThR.Tn[4].t62 VGND 0.0199f
C10344 XThR.Tn[4].n67 VGND 0.04859f
C10345 XThR.Tn[4].t23 VGND 0.01811f
C10346 XThR.Tn[4].t59 VGND 0.01983f
C10347 XThR.Tn[4].n68 VGND 0.05056f
C10348 XThR.Tn[4].n69 VGND 0.03552f
C10349 XThR.Tn[4].n70 VGND 0.00649f
C10350 XThR.Tn[4].n71 VGND 0.11398f
C10351 XThR.Tn[4].t20 VGND 0.01817f
C10352 XThR.Tn[4].t14 VGND 0.0199f
C10353 XThR.Tn[4].n72 VGND 0.04859f
C10354 XThR.Tn[4].t42 VGND 0.01811f
C10355 XThR.Tn[4].t72 VGND 0.01983f
C10356 XThR.Tn[4].n73 VGND 0.05056f
C10357 XThR.Tn[4].n74 VGND 0.03552f
C10358 XThR.Tn[4].n75 VGND 0.00649f
C10359 XThR.Tn[4].n76 VGND 0.11398f
C10360 XThR.Tn[4].t40 VGND 0.01817f
C10361 XThR.Tn[4].t34 VGND 0.0199f
C10362 XThR.Tn[4].n77 VGND 0.04859f
C10363 XThR.Tn[4].t60 VGND 0.01811f
C10364 XThR.Tn[4].t30 VGND 0.01983f
C10365 XThR.Tn[4].n78 VGND 0.05056f
C10366 XThR.Tn[4].n79 VGND 0.03552f
C10367 XThR.Tn[4].n80 VGND 0.00649f
C10368 XThR.Tn[4].n81 VGND 0.11398f
C10369 XThR.Tn[4].t16 VGND 0.01817f
C10370 XThR.Tn[4].t28 VGND 0.0199f
C10371 XThR.Tn[4].n82 VGND 0.04859f
C10372 XThR.Tn[4].t37 VGND 0.01811f
C10373 XThR.Tn[4].t24 VGND 0.01983f
C10374 XThR.Tn[4].n83 VGND 0.05056f
C10375 XThR.Tn[4].n84 VGND 0.03552f
C10376 XThR.Tn[4].n85 VGND 0.00649f
C10377 XThR.Tn[4].n86 VGND 0.11398f
C10378 XThR.Tn[4].n87 VGND 0.10358f
C10379 XThR.Tn[4].n88 VGND 0.19569f
C10380 XThC.Tn[7].t4 VGND 0.0189f
C10381 XThC.Tn[7].t7 VGND 0.0189f
C10382 XThC.Tn[7].n0 VGND 0.0407f
C10383 XThC.Tn[7].t6 VGND 0.0189f
C10384 XThC.Tn[7].t5 VGND 0.0189f
C10385 XThC.Tn[7].n1 VGND 0.06179f
C10386 XThC.Tn[7].n2 VGND 0.18167f
C10387 XThC.Tn[7].t8 VGND 0.01498f
C10388 XThC.Tn[7].t11 VGND 0.01636f
C10389 XThC.Tn[7].n3 VGND 0.03652f
C10390 XThC.Tn[7].n4 VGND 0.02502f
C10391 XThC.Tn[7].n5 VGND 0.08213f
C10392 XThC.Tn[7].t25 VGND 0.01498f
C10393 XThC.Tn[7].t30 VGND 0.01636f
C10394 XThC.Tn[7].n6 VGND 0.03652f
C10395 XThC.Tn[7].n7 VGND 0.02502f
C10396 XThC.Tn[7].n8 VGND 0.08235f
C10397 XThC.Tn[7].n9 VGND 0.13573f
C10398 XThC.Tn[7].t27 VGND 0.01498f
C10399 XThC.Tn[7].t34 VGND 0.01636f
C10400 XThC.Tn[7].n10 VGND 0.03652f
C10401 XThC.Tn[7].n11 VGND 0.02502f
C10402 XThC.Tn[7].n12 VGND 0.08235f
C10403 XThC.Tn[7].n13 VGND 0.13573f
C10404 XThC.Tn[7].t29 VGND 0.01498f
C10405 XThC.Tn[7].t35 VGND 0.01636f
C10406 XThC.Tn[7].n14 VGND 0.03652f
C10407 XThC.Tn[7].n15 VGND 0.02502f
C10408 XThC.Tn[7].n16 VGND 0.08235f
C10409 XThC.Tn[7].n17 VGND 0.13573f
C10410 XThC.Tn[7].t18 VGND 0.01498f
C10411 XThC.Tn[7].t22 VGND 0.01636f
C10412 XThC.Tn[7].n18 VGND 0.03652f
C10413 XThC.Tn[7].n19 VGND 0.02502f
C10414 XThC.Tn[7].n20 VGND 0.08235f
C10415 XThC.Tn[7].n21 VGND 0.13573f
C10416 XThC.Tn[7].t20 VGND 0.01498f
C10417 XThC.Tn[7].t23 VGND 0.01636f
C10418 XThC.Tn[7].n22 VGND 0.03652f
C10419 XThC.Tn[7].n23 VGND 0.02502f
C10420 XThC.Tn[7].n24 VGND 0.08235f
C10421 XThC.Tn[7].n25 VGND 0.13573f
C10422 XThC.Tn[7].t33 VGND 0.01498f
C10423 XThC.Tn[7].t39 VGND 0.01636f
C10424 XThC.Tn[7].n26 VGND 0.03652f
C10425 XThC.Tn[7].n27 VGND 0.02502f
C10426 XThC.Tn[7].n28 VGND 0.08235f
C10427 XThC.Tn[7].n29 VGND 0.13573f
C10428 XThC.Tn[7].t10 VGND 0.01498f
C10429 XThC.Tn[7].t14 VGND 0.01636f
C10430 XThC.Tn[7].n30 VGND 0.03652f
C10431 XThC.Tn[7].n31 VGND 0.02502f
C10432 XThC.Tn[7].n32 VGND 0.08235f
C10433 XThC.Tn[7].n33 VGND 0.13573f
C10434 XThC.Tn[7].t12 VGND 0.01498f
C10435 XThC.Tn[7].t16 VGND 0.01636f
C10436 XThC.Tn[7].n34 VGND 0.03652f
C10437 XThC.Tn[7].n35 VGND 0.02502f
C10438 XThC.Tn[7].n36 VGND 0.08235f
C10439 XThC.Tn[7].n37 VGND 0.13573f
C10440 XThC.Tn[7].t31 VGND 0.01498f
C10441 XThC.Tn[7].t36 VGND 0.01636f
C10442 XThC.Tn[7].n38 VGND 0.03652f
C10443 XThC.Tn[7].n39 VGND 0.02502f
C10444 XThC.Tn[7].n40 VGND 0.08235f
C10445 XThC.Tn[7].n41 VGND 0.13573f
C10446 XThC.Tn[7].t32 VGND 0.01498f
C10447 XThC.Tn[7].t38 VGND 0.01636f
C10448 XThC.Tn[7].n42 VGND 0.03652f
C10449 XThC.Tn[7].n43 VGND 0.02502f
C10450 XThC.Tn[7].n44 VGND 0.08235f
C10451 XThC.Tn[7].n45 VGND 0.13573f
C10452 XThC.Tn[7].t13 VGND 0.01498f
C10453 XThC.Tn[7].t17 VGND 0.01636f
C10454 XThC.Tn[7].n46 VGND 0.03652f
C10455 XThC.Tn[7].n47 VGND 0.02502f
C10456 XThC.Tn[7].n48 VGND 0.08235f
C10457 XThC.Tn[7].n49 VGND 0.13573f
C10458 XThC.Tn[7].t21 VGND 0.01498f
C10459 XThC.Tn[7].t26 VGND 0.01636f
C10460 XThC.Tn[7].n50 VGND 0.03652f
C10461 XThC.Tn[7].n51 VGND 0.02502f
C10462 XThC.Tn[7].n52 VGND 0.08235f
C10463 XThC.Tn[7].n53 VGND 0.13573f
C10464 XThC.Tn[7].t24 VGND 0.01498f
C10465 XThC.Tn[7].t28 VGND 0.01636f
C10466 XThC.Tn[7].n54 VGND 0.03652f
C10467 XThC.Tn[7].n55 VGND 0.02502f
C10468 XThC.Tn[7].n56 VGND 0.08235f
C10469 XThC.Tn[7].n57 VGND 0.13573f
C10470 XThC.Tn[7].t37 VGND 0.01498f
C10471 XThC.Tn[7].t9 VGND 0.01636f
C10472 XThC.Tn[7].n58 VGND 0.03652f
C10473 XThC.Tn[7].n59 VGND 0.02502f
C10474 XThC.Tn[7].n60 VGND 0.08235f
C10475 XThC.Tn[7].n61 VGND 0.13573f
C10476 XThC.Tn[7].t15 VGND 0.01498f
C10477 XThC.Tn[7].t19 VGND 0.01636f
C10478 XThC.Tn[7].n62 VGND 0.03652f
C10479 XThC.Tn[7].n63 VGND 0.02502f
C10480 XThC.Tn[7].n64 VGND 0.08235f
C10481 XThC.Tn[7].n65 VGND 0.13573f
C10482 XThC.Tn[7].n66 VGND 0.34086f
C10483 XThC.Tn[7].t2 VGND 0.01228f
C10484 XThC.Tn[7].t1 VGND 0.01228f
C10485 XThC.Tn[7].n67 VGND 0.03791f
C10486 XThC.Tn[7].t0 VGND 0.01228f
C10487 XThC.Tn[7].t3 VGND 0.01228f
C10488 XThC.Tn[7].n68 VGND 0.02713f
C10489 XThC.Tn[7].n69 VGND 0.13418f
C10490 XThC.Tn[7].n70 VGND 0.02261f
C10491 XThR.Tn[1].t11 VGND 0.01497f
C10492 XThR.Tn[1].t8 VGND 0.01497f
C10493 XThR.Tn[1].n0 VGND 0.05682f
C10494 XThR.Tn[1].t10 VGND 0.01497f
C10495 XThR.Tn[1].t9 VGND 0.01497f
C10496 XThR.Tn[1].n1 VGND 0.0341f
C10497 XThR.Tn[1].n2 VGND 0.16239f
C10498 XThR.Tn[1].t6 VGND 0.01497f
C10499 XThR.Tn[1].t5 VGND 0.01497f
C10500 XThR.Tn[1].n3 VGND 0.0341f
C10501 XThR.Tn[1].n4 VGND 0.10039f
C10502 XThR.Tn[1].t7 VGND 0.01497f
C10503 XThR.Tn[1].t4 VGND 0.01497f
C10504 XThR.Tn[1].n5 VGND 0.0341f
C10505 XThR.Tn[1].n6 VGND 0.11329f
C10506 XThR.Tn[1].t24 VGND 0.01801f
C10507 XThR.Tn[1].t18 VGND 0.01972f
C10508 XThR.Tn[1].n7 VGND 0.04814f
C10509 XThR.Tn[1].n8 VGND 0.09248f
C10510 XThR.Tn[1].t44 VGND 0.01801f
C10511 XThR.Tn[1].t34 VGND 0.01972f
C10512 XThR.Tn[1].n9 VGND 0.04814f
C10513 XThR.Tn[1].t61 VGND 0.01795f
C10514 XThR.Tn[1].t30 VGND 0.01965f
C10515 XThR.Tn[1].n10 VGND 0.05009f
C10516 XThR.Tn[1].n11 VGND 0.03519f
C10517 XThR.Tn[1].n12 VGND 0.00643f
C10518 XThR.Tn[1].n13 VGND 0.11293f
C10519 XThR.Tn[1].t19 VGND 0.01801f
C10520 XThR.Tn[1].t73 VGND 0.01972f
C10521 XThR.Tn[1].n14 VGND 0.04814f
C10522 XThR.Tn[1].t38 VGND 0.01795f
C10523 XThR.Tn[1].t69 VGND 0.01965f
C10524 XThR.Tn[1].n15 VGND 0.05009f
C10525 XThR.Tn[1].n16 VGND 0.03519f
C10526 XThR.Tn[1].n17 VGND 0.00643f
C10527 XThR.Tn[1].n18 VGND 0.11293f
C10528 XThR.Tn[1].t35 VGND 0.01801f
C10529 XThR.Tn[1].t28 VGND 0.01972f
C10530 XThR.Tn[1].n19 VGND 0.04814f
C10531 XThR.Tn[1].t50 VGND 0.01795f
C10532 XThR.Tn[1].t25 VGND 0.01965f
C10533 XThR.Tn[1].n20 VGND 0.05009f
C10534 XThR.Tn[1].n21 VGND 0.03519f
C10535 XThR.Tn[1].n22 VGND 0.00643f
C10536 XThR.Tn[1].n23 VGND 0.11293f
C10537 XThR.Tn[1].t59 VGND 0.01801f
C10538 XThR.Tn[1].t55 VGND 0.01972f
C10539 XThR.Tn[1].n24 VGND 0.04814f
C10540 XThR.Tn[1].t21 VGND 0.01795f
C10541 XThR.Tn[1].t51 VGND 0.01965f
C10542 XThR.Tn[1].n25 VGND 0.05009f
C10543 XThR.Tn[1].n26 VGND 0.03519f
C10544 XThR.Tn[1].n27 VGND 0.00643f
C10545 XThR.Tn[1].n28 VGND 0.11293f
C10546 XThR.Tn[1].t37 VGND 0.01801f
C10547 XThR.Tn[1].t29 VGND 0.01972f
C10548 XThR.Tn[1].n29 VGND 0.04814f
C10549 XThR.Tn[1].t53 VGND 0.01795f
C10550 XThR.Tn[1].t26 VGND 0.01965f
C10551 XThR.Tn[1].n30 VGND 0.05009f
C10552 XThR.Tn[1].n31 VGND 0.03519f
C10553 XThR.Tn[1].n32 VGND 0.00643f
C10554 XThR.Tn[1].n33 VGND 0.11293f
C10555 XThR.Tn[1].t13 VGND 0.01801f
C10556 XThR.Tn[1].t46 VGND 0.01972f
C10557 XThR.Tn[1].n34 VGND 0.04814f
C10558 XThR.Tn[1].t32 VGND 0.01795f
C10559 XThR.Tn[1].t43 VGND 0.01965f
C10560 XThR.Tn[1].n35 VGND 0.05009f
C10561 XThR.Tn[1].n36 VGND 0.03519f
C10562 XThR.Tn[1].n37 VGND 0.00643f
C10563 XThR.Tn[1].n38 VGND 0.11293f
C10564 XThR.Tn[1].t45 VGND 0.01801f
C10565 XThR.Tn[1].t41 VGND 0.01972f
C10566 XThR.Tn[1].n39 VGND 0.04814f
C10567 XThR.Tn[1].t60 VGND 0.01795f
C10568 XThR.Tn[1].t36 VGND 0.01965f
C10569 XThR.Tn[1].n40 VGND 0.05009f
C10570 XThR.Tn[1].n41 VGND 0.03519f
C10571 XThR.Tn[1].n42 VGND 0.00643f
C10572 XThR.Tn[1].n43 VGND 0.11293f
C10573 XThR.Tn[1].t48 VGND 0.01801f
C10574 XThR.Tn[1].t54 VGND 0.01972f
C10575 XThR.Tn[1].n44 VGND 0.04814f
C10576 XThR.Tn[1].t67 VGND 0.01795f
C10577 XThR.Tn[1].t49 VGND 0.01965f
C10578 XThR.Tn[1].n45 VGND 0.05009f
C10579 XThR.Tn[1].n46 VGND 0.03519f
C10580 XThR.Tn[1].n47 VGND 0.00643f
C10581 XThR.Tn[1].n48 VGND 0.11293f
C10582 XThR.Tn[1].t64 VGND 0.01801f
C10583 XThR.Tn[1].t12 VGND 0.01972f
C10584 XThR.Tn[1].n49 VGND 0.04814f
C10585 XThR.Tn[1].t23 VGND 0.01795f
C10586 XThR.Tn[1].t71 VGND 0.01965f
C10587 XThR.Tn[1].n50 VGND 0.05009f
C10588 XThR.Tn[1].n51 VGND 0.03519f
C10589 XThR.Tn[1].n52 VGND 0.00643f
C10590 XThR.Tn[1].n53 VGND 0.11293f
C10591 XThR.Tn[1].t57 VGND 0.01801f
C10592 XThR.Tn[1].t31 VGND 0.01972f
C10593 XThR.Tn[1].n54 VGND 0.04814f
C10594 XThR.Tn[1].t16 VGND 0.01795f
C10595 XThR.Tn[1].t27 VGND 0.01965f
C10596 XThR.Tn[1].n55 VGND 0.05009f
C10597 XThR.Tn[1].n56 VGND 0.03519f
C10598 XThR.Tn[1].n57 VGND 0.00643f
C10599 XThR.Tn[1].n58 VGND 0.11293f
C10600 XThR.Tn[1].t15 VGND 0.01801f
C10601 XThR.Tn[1].t68 VGND 0.01972f
C10602 XThR.Tn[1].n59 VGND 0.04814f
C10603 XThR.Tn[1].t33 VGND 0.01795f
C10604 XThR.Tn[1].t63 VGND 0.01965f
C10605 XThR.Tn[1].n60 VGND 0.05009f
C10606 XThR.Tn[1].n61 VGND 0.03519f
C10607 XThR.Tn[1].n62 VGND 0.00643f
C10608 XThR.Tn[1].n63 VGND 0.11293f
C10609 XThR.Tn[1].t47 VGND 0.01801f
C10610 XThR.Tn[1].t42 VGND 0.01972f
C10611 XThR.Tn[1].n64 VGND 0.04814f
C10612 XThR.Tn[1].t65 VGND 0.01795f
C10613 XThR.Tn[1].t39 VGND 0.01965f
C10614 XThR.Tn[1].n65 VGND 0.05009f
C10615 XThR.Tn[1].n66 VGND 0.03519f
C10616 XThR.Tn[1].n67 VGND 0.00643f
C10617 XThR.Tn[1].n68 VGND 0.11293f
C10618 XThR.Tn[1].t62 VGND 0.01801f
C10619 XThR.Tn[1].t56 VGND 0.01972f
C10620 XThR.Tn[1].n69 VGND 0.04814f
C10621 XThR.Tn[1].t22 VGND 0.01795f
C10622 XThR.Tn[1].t52 VGND 0.01965f
C10623 XThR.Tn[1].n70 VGND 0.05009f
C10624 XThR.Tn[1].n71 VGND 0.03519f
C10625 XThR.Tn[1].n72 VGND 0.00643f
C10626 XThR.Tn[1].n73 VGND 0.11293f
C10627 XThR.Tn[1].t20 VGND 0.01801f
C10628 XThR.Tn[1].t14 VGND 0.01972f
C10629 XThR.Tn[1].n74 VGND 0.04814f
C10630 XThR.Tn[1].t40 VGND 0.01795f
C10631 XThR.Tn[1].t72 VGND 0.01965f
C10632 XThR.Tn[1].n75 VGND 0.05009f
C10633 XThR.Tn[1].n76 VGND 0.03519f
C10634 XThR.Tn[1].n77 VGND 0.00643f
C10635 XThR.Tn[1].n78 VGND 0.11293f
C10636 XThR.Tn[1].t58 VGND 0.01801f
C10637 XThR.Tn[1].t70 VGND 0.01972f
C10638 XThR.Tn[1].n79 VGND 0.04814f
C10639 XThR.Tn[1].t17 VGND 0.01795f
C10640 XThR.Tn[1].t66 VGND 0.01965f
C10641 XThR.Tn[1].n80 VGND 0.05009f
C10642 XThR.Tn[1].n81 VGND 0.03519f
C10643 XThR.Tn[1].n82 VGND 0.00643f
C10644 XThR.Tn[1].n83 VGND 0.11293f
C10645 XThR.Tn[1].n84 VGND 0.10263f
C10646 XThR.Tn[1].n85 VGND 0.29541f
C10647 XThR.Tn[1].t0 VGND 0.02304f
C10648 XThR.Tn[1].t1 VGND 0.02304f
C10649 XThR.Tn[1].n86 VGND 0.0465f
C10650 XThR.Tn[1].t3 VGND 0.02304f
C10651 XThR.Tn[1].t2 VGND 0.02304f
C10652 XThR.Tn[1].n87 VGND 0.05441f
C10653 XThR.Tn[1].n88 VGND 0.15232f
C10654 XThR.Tn[1].n89 VGND 0.04821f
C10655 XThC.Tn[8].t5 VGND 0.01304f
C10656 XThC.Tn[8].t4 VGND 0.01304f
C10657 XThC.Tn[8].n0 VGND 0.03253f
C10658 XThC.Tn[8].t7 VGND 0.01304f
C10659 XThC.Tn[8].t6 VGND 0.01304f
C10660 XThC.Tn[8].n1 VGND 0.02608f
C10661 XThC.Tn[8].n2 VGND 0.06561f
C10662 XThC.Tn[8].n3 VGND 0.02453f
C10663 XThC.Tn[8].t43 VGND 0.0159f
C10664 XThC.Tn[8].t41 VGND 0.01737f
C10665 XThC.Tn[8].n4 VGND 0.03878f
C10666 XThC.Tn[8].n5 VGND 0.02657f
C10667 XThC.Tn[8].n6 VGND 0.0872f
C10668 XThC.Tn[8].t29 VGND 0.0159f
C10669 XThC.Tn[8].t26 VGND 0.01737f
C10670 XThC.Tn[8].n7 VGND 0.03878f
C10671 XThC.Tn[8].n8 VGND 0.02657f
C10672 XThC.Tn[8].n9 VGND 0.08744f
C10673 XThC.Tn[8].n10 VGND 0.1441f
C10674 XThC.Tn[8].t34 VGND 0.0159f
C10675 XThC.Tn[8].t28 VGND 0.01737f
C10676 XThC.Tn[8].n11 VGND 0.03878f
C10677 XThC.Tn[8].n12 VGND 0.02657f
C10678 XThC.Tn[8].n13 VGND 0.08744f
C10679 XThC.Tn[8].n14 VGND 0.1441f
C10680 XThC.Tn[8].t35 VGND 0.0159f
C10681 XThC.Tn[8].t30 VGND 0.01737f
C10682 XThC.Tn[8].n15 VGND 0.03878f
C10683 XThC.Tn[8].n16 VGND 0.02657f
C10684 XThC.Tn[8].n17 VGND 0.08744f
C10685 XThC.Tn[8].n18 VGND 0.1441f
C10686 XThC.Tn[8].t22 VGND 0.0159f
C10687 XThC.Tn[8].t19 VGND 0.01737f
C10688 XThC.Tn[8].n19 VGND 0.03878f
C10689 XThC.Tn[8].n20 VGND 0.02657f
C10690 XThC.Tn[8].n21 VGND 0.08744f
C10691 XThC.Tn[8].n22 VGND 0.1441f
C10692 XThC.Tn[8].t23 VGND 0.0159f
C10693 XThC.Tn[8].t20 VGND 0.01737f
C10694 XThC.Tn[8].n23 VGND 0.03878f
C10695 XThC.Tn[8].n24 VGND 0.02657f
C10696 XThC.Tn[8].n25 VGND 0.08744f
C10697 XThC.Tn[8].n26 VGND 0.1441f
C10698 XThC.Tn[8].t39 VGND 0.0159f
C10699 XThC.Tn[8].t33 VGND 0.01737f
C10700 XThC.Tn[8].n27 VGND 0.03878f
C10701 XThC.Tn[8].n28 VGND 0.02657f
C10702 XThC.Tn[8].n29 VGND 0.08744f
C10703 XThC.Tn[8].n30 VGND 0.1441f
C10704 XThC.Tn[8].t14 VGND 0.0159f
C10705 XThC.Tn[8].t42 VGND 0.01737f
C10706 XThC.Tn[8].n31 VGND 0.03878f
C10707 XThC.Tn[8].n32 VGND 0.02657f
C10708 XThC.Tn[8].n33 VGND 0.08744f
C10709 XThC.Tn[8].n34 VGND 0.1441f
C10710 XThC.Tn[8].t16 VGND 0.0159f
C10711 XThC.Tn[8].t12 VGND 0.01737f
C10712 XThC.Tn[8].n35 VGND 0.03878f
C10713 XThC.Tn[8].n36 VGND 0.02657f
C10714 XThC.Tn[8].n37 VGND 0.08744f
C10715 XThC.Tn[8].n38 VGND 0.1441f
C10716 XThC.Tn[8].t36 VGND 0.0159f
C10717 XThC.Tn[8].t31 VGND 0.01737f
C10718 XThC.Tn[8].n39 VGND 0.03878f
C10719 XThC.Tn[8].n40 VGND 0.02657f
C10720 XThC.Tn[8].n41 VGND 0.08744f
C10721 XThC.Tn[8].n42 VGND 0.1441f
C10722 XThC.Tn[8].t38 VGND 0.0159f
C10723 XThC.Tn[8].t32 VGND 0.01737f
C10724 XThC.Tn[8].n43 VGND 0.03878f
C10725 XThC.Tn[8].n44 VGND 0.02657f
C10726 XThC.Tn[8].n45 VGND 0.08744f
C10727 XThC.Tn[8].n46 VGND 0.1441f
C10728 XThC.Tn[8].t17 VGND 0.0159f
C10729 XThC.Tn[8].t13 VGND 0.01737f
C10730 XThC.Tn[8].n47 VGND 0.03878f
C10731 XThC.Tn[8].n48 VGND 0.02657f
C10732 XThC.Tn[8].n49 VGND 0.08744f
C10733 XThC.Tn[8].n50 VGND 0.1441f
C10734 XThC.Tn[8].t25 VGND 0.0159f
C10735 XThC.Tn[8].t21 VGND 0.01737f
C10736 XThC.Tn[8].n51 VGND 0.03878f
C10737 XThC.Tn[8].n52 VGND 0.02657f
C10738 XThC.Tn[8].n53 VGND 0.08744f
C10739 XThC.Tn[8].n54 VGND 0.1441f
C10740 XThC.Tn[8].t27 VGND 0.0159f
C10741 XThC.Tn[8].t24 VGND 0.01737f
C10742 XThC.Tn[8].n55 VGND 0.03878f
C10743 XThC.Tn[8].n56 VGND 0.02657f
C10744 XThC.Tn[8].n57 VGND 0.08744f
C10745 XThC.Tn[8].n58 VGND 0.1441f
C10746 XThC.Tn[8].t40 VGND 0.0159f
C10747 XThC.Tn[8].t37 VGND 0.01737f
C10748 XThC.Tn[8].n59 VGND 0.03878f
C10749 XThC.Tn[8].n60 VGND 0.02657f
C10750 XThC.Tn[8].n61 VGND 0.08744f
C10751 XThC.Tn[8].n62 VGND 0.1441f
C10752 XThC.Tn[8].t18 VGND 0.0159f
C10753 XThC.Tn[8].t15 VGND 0.01737f
C10754 XThC.Tn[8].n63 VGND 0.03878f
C10755 XThC.Tn[8].n64 VGND 0.02657f
C10756 XThC.Tn[8].n65 VGND 0.08744f
C10757 XThC.Tn[8].n66 VGND 0.1441f
C10758 XThC.Tn[8].n67 VGND 0.60346f
C10759 XThC.Tn[8].n68 VGND 0.23618f
C10760 XThC.Tn[8].t9 VGND 0.02006f
C10761 XThC.Tn[8].t10 VGND 0.02006f
C10762 XThC.Tn[8].n69 VGND 0.04335f
C10763 XThC.Tn[8].t8 VGND 0.02006f
C10764 XThC.Tn[8].t11 VGND 0.02006f
C10765 XThC.Tn[8].n70 VGND 0.06598f
C10766 XThC.Tn[8].n71 VGND 0.18333f
C10767 XThC.Tn[8].n72 VGND 0.02883f
C10768 XThC.Tn[8].t2 VGND 0.02006f
C10769 XThC.Tn[8].t1 VGND 0.02006f
C10770 XThC.Tn[8].n73 VGND 0.0446f
C10771 XThC.Tn[8].t0 VGND 0.02006f
C10772 XThC.Tn[8].t3 VGND 0.02006f
C10773 XThC.Tn[8].n74 VGND 0.06092f
C10774 XThC.Tn[8].n75 VGND 0.1985f
C10775 XThC.TB1.t1 VGND 0.03224f
C10776 XThC.TB1.n0 VGND 0.02084f
C10777 XThC.TB1.n1 VGND 0.02659f
C10778 XThC.TB1.t0 VGND 0.01618f
C10779 XThC.TB1.t2 VGND 0.01618f
C10780 XThC.TB1.n2 VGND 0.03473f
C10781 XThC.TB1.t17 VGND 0.02517f
C10782 XThC.TB1.t5 VGND 0.01483f
C10783 XThC.TB1.n3 VGND 0.02997f
C10784 XThC.TB1.t6 VGND 0.02517f
C10785 XThC.TB1.t12 VGND 0.01483f
C10786 XThC.TB1.n4 VGND 0.01542f
C10787 XThC.TB1.t8 VGND 0.02517f
C10788 XThC.TB1.t13 VGND 0.01483f
C10789 XThC.TB1.n5 VGND 0.03313f
C10790 XThC.TB1.t11 VGND 0.02517f
C10791 XThC.TB1.t16 VGND 0.01483f
C10792 XThC.TB1.n6 VGND 0.03076f
C10793 XThC.TB1.n7 VGND 0.01871f
C10794 XThC.TB1.n8 VGND 0.03098f
C10795 XThC.TB1.n9 VGND 0.01198f
C10796 XThC.TB1.n10 VGND 0.01463f
C10797 XThC.TB1.n11 VGND 0.03313f
C10798 XThC.TB1.n12 VGND 0.01661f
C10799 XThC.TB1.n13 VGND 0.02824f
C10800 XThC.TB1.t18 VGND 0.02517f
C10801 XThC.TB1.t9 VGND 0.01483f
C10802 XThC.TB1.n14 VGND 0.03392f
C10803 XThC.TB1.t7 VGND 0.02517f
C10804 XThC.TB1.t15 VGND 0.01483f
C10805 XThC.TB1.t14 VGND 0.02517f
C10806 XThC.TB1.t3 VGND 0.01483f
C10807 XThC.TB1.t10 VGND 0.02517f
C10808 XThC.TB1.t4 VGND 0.01483f
C10809 XThC.TB1.n15 VGND 0.04223f
C10810 XThC.TB1.n16 VGND 0.0446f
C10811 XThC.TB1.n17 VGND 0.01719f
C10812 XThC.TB1.n18 VGND 0.0363f
C10813 XThC.TB1.n19 VGND 0.01661f
C10814 XThC.TB1.n20 VGND 0.01378f
C10815 XThC.TB1.n21 VGND 0.13924f
C10816 XThC.TB1.n22 VGND 0.07634f
C10817 XThC.Tn[14].t0 VGND 0.01262f
C10818 XThC.Tn[14].t2 VGND 0.01262f
C10819 XThC.Tn[14].n0 VGND 0.03148f
C10820 XThC.Tn[14].t1 VGND 0.01262f
C10821 XThC.Tn[14].t3 VGND 0.01262f
C10822 XThC.Tn[14].n1 VGND 0.02524f
C10823 XThC.Tn[14].n2 VGND 0.06349f
C10824 XThC.Tn[14].t4 VGND 0.01942f
C10825 XThC.Tn[14].t5 VGND 0.01942f
C10826 XThC.Tn[14].n3 VGND 0.04195f
C10827 XThC.Tn[14].t7 VGND 0.01942f
C10828 XThC.Tn[14].t6 VGND 0.01942f
C10829 XThC.Tn[14].n4 VGND 0.06385f
C10830 XThC.Tn[14].n5 VGND 0.1774f
C10831 XThC.Tn[14].t11 VGND 0.01942f
C10832 XThC.Tn[14].t10 VGND 0.01942f
C10833 XThC.Tn[14].n6 VGND 0.05895f
C10834 XThC.Tn[14].t9 VGND 0.01942f
C10835 XThC.Tn[14].t8 VGND 0.01942f
C10836 XThC.Tn[14].n7 VGND 0.04316f
C10837 XThC.Tn[14].n8 VGND 0.19209f
C10838 XThC.Tn[14].n9 VGND 0.02789f
C10839 XThC.Tn[14].t43 VGND 0.01539f
C10840 XThC.Tn[14].t38 VGND 0.01681f
C10841 XThC.Tn[14].n10 VGND 0.03752f
C10842 XThC.Tn[14].n11 VGND 0.02571f
C10843 XThC.Tn[14].n12 VGND 0.08438f
C10844 XThC.Tn[14].t29 VGND 0.01539f
C10845 XThC.Tn[14].t22 VGND 0.01681f
C10846 XThC.Tn[14].n13 VGND 0.03752f
C10847 XThC.Tn[14].n14 VGND 0.02571f
C10848 XThC.Tn[14].n15 VGND 0.08461f
C10849 XThC.Tn[14].n16 VGND 0.13945f
C10850 XThC.Tn[14].t32 VGND 0.01539f
C10851 XThC.Tn[14].t25 VGND 0.01681f
C10852 XThC.Tn[14].n17 VGND 0.03752f
C10853 XThC.Tn[14].n18 VGND 0.02571f
C10854 XThC.Tn[14].n19 VGND 0.08461f
C10855 XThC.Tn[14].n20 VGND 0.13945f
C10856 XThC.Tn[14].t34 VGND 0.01539f
C10857 XThC.Tn[14].t26 VGND 0.01681f
C10858 XThC.Tn[14].n21 VGND 0.03752f
C10859 XThC.Tn[14].n22 VGND 0.02571f
C10860 XThC.Tn[14].n23 VGND 0.08461f
C10861 XThC.Tn[14].n24 VGND 0.13945f
C10862 XThC.Tn[14].t20 VGND 0.01539f
C10863 XThC.Tn[14].t14 VGND 0.01681f
C10864 XThC.Tn[14].n25 VGND 0.03752f
C10865 XThC.Tn[14].n26 VGND 0.02571f
C10866 XThC.Tn[14].n27 VGND 0.08461f
C10867 XThC.Tn[14].n28 VGND 0.13945f
C10868 XThC.Tn[14].t23 VGND 0.01539f
C10869 XThC.Tn[14].t17 VGND 0.01681f
C10870 XThC.Tn[14].n29 VGND 0.03752f
C10871 XThC.Tn[14].n30 VGND 0.02571f
C10872 XThC.Tn[14].n31 VGND 0.08461f
C10873 XThC.Tn[14].n32 VGND 0.13945f
C10874 XThC.Tn[14].t37 VGND 0.01539f
C10875 XThC.Tn[14].t31 VGND 0.01681f
C10876 XThC.Tn[14].n33 VGND 0.03752f
C10877 XThC.Tn[14].n34 VGND 0.02571f
C10878 XThC.Tn[14].n35 VGND 0.08461f
C10879 XThC.Tn[14].n36 VGND 0.13945f
C10880 XThC.Tn[14].t13 VGND 0.01539f
C10881 XThC.Tn[14].t39 VGND 0.01681f
C10882 XThC.Tn[14].n37 VGND 0.03752f
C10883 XThC.Tn[14].n38 VGND 0.02571f
C10884 XThC.Tn[14].n39 VGND 0.08461f
C10885 XThC.Tn[14].n40 VGND 0.13945f
C10886 XThC.Tn[14].t15 VGND 0.01539f
C10887 XThC.Tn[14].t41 VGND 0.01681f
C10888 XThC.Tn[14].n41 VGND 0.03752f
C10889 XThC.Tn[14].n42 VGND 0.02571f
C10890 XThC.Tn[14].n43 VGND 0.08461f
C10891 XThC.Tn[14].n44 VGND 0.13945f
C10892 XThC.Tn[14].t35 VGND 0.01539f
C10893 XThC.Tn[14].t27 VGND 0.01681f
C10894 XThC.Tn[14].n45 VGND 0.03752f
C10895 XThC.Tn[14].n46 VGND 0.02571f
C10896 XThC.Tn[14].n47 VGND 0.08461f
C10897 XThC.Tn[14].n48 VGND 0.13945f
C10898 XThC.Tn[14].t36 VGND 0.01539f
C10899 XThC.Tn[14].t30 VGND 0.01681f
C10900 XThC.Tn[14].n49 VGND 0.03752f
C10901 XThC.Tn[14].n50 VGND 0.02571f
C10902 XThC.Tn[14].n51 VGND 0.08461f
C10903 XThC.Tn[14].n52 VGND 0.13945f
C10904 XThC.Tn[14].t16 VGND 0.01539f
C10905 XThC.Tn[14].t42 VGND 0.01681f
C10906 XThC.Tn[14].n53 VGND 0.03752f
C10907 XThC.Tn[14].n54 VGND 0.02571f
C10908 XThC.Tn[14].n55 VGND 0.08461f
C10909 XThC.Tn[14].n56 VGND 0.13945f
C10910 XThC.Tn[14].t24 VGND 0.01539f
C10911 XThC.Tn[14].t19 VGND 0.01681f
C10912 XThC.Tn[14].n57 VGND 0.03752f
C10913 XThC.Tn[14].n58 VGND 0.02571f
C10914 XThC.Tn[14].n59 VGND 0.08461f
C10915 XThC.Tn[14].n60 VGND 0.13945f
C10916 XThC.Tn[14].t28 VGND 0.01539f
C10917 XThC.Tn[14].t21 VGND 0.01681f
C10918 XThC.Tn[14].n61 VGND 0.03752f
C10919 XThC.Tn[14].n62 VGND 0.02571f
C10920 XThC.Tn[14].n63 VGND 0.08461f
C10921 XThC.Tn[14].n64 VGND 0.13945f
C10922 XThC.Tn[14].t40 VGND 0.01539f
C10923 XThC.Tn[14].t33 VGND 0.01681f
C10924 XThC.Tn[14].n65 VGND 0.03752f
C10925 XThC.Tn[14].n66 VGND 0.02571f
C10926 XThC.Tn[14].n67 VGND 0.08461f
C10927 XThC.Tn[14].n68 VGND 0.13945f
C10928 XThC.Tn[14].t18 VGND 0.01539f
C10929 XThC.Tn[14].t12 VGND 0.01681f
C10930 XThC.Tn[14].n69 VGND 0.03752f
C10931 XThC.Tn[14].n70 VGND 0.02571f
C10932 XThC.Tn[14].n71 VGND 0.08461f
C10933 XThC.Tn[14].n72 VGND 0.13945f
C10934 XThC.Tn[14].n73 VGND 0.91462f
C10935 XThC.Tn[14].n74 VGND 0.26906f
C10936 XThR.Tn[10].t10 VGND 0.02415f
C10937 XThR.Tn[10].t8 VGND 0.02415f
C10938 XThR.Tn[10].n0 VGND 0.07333f
C10939 XThR.Tn[10].t11 VGND 0.02415f
C10940 XThR.Tn[10].t9 VGND 0.02415f
C10941 XThR.Tn[10].n1 VGND 0.05368f
C10942 XThR.Tn[10].n2 VGND 0.2441f
C10943 XThR.Tn[10].t1 VGND 0.0157f
C10944 XThR.Tn[10].t4 VGND 0.0157f
C10945 XThR.Tn[10].n3 VGND 0.03915f
C10946 XThR.Tn[10].t2 VGND 0.0157f
C10947 XThR.Tn[10].t7 VGND 0.0157f
C10948 XThR.Tn[10].n4 VGND 0.0314f
C10949 XThR.Tn[10].n5 VGND 0.07239f
C10950 XThR.Tn[10].t54 VGND 0.01887f
C10951 XThR.Tn[10].t47 VGND 0.02067f
C10952 XThR.Tn[10].n6 VGND 0.05047f
C10953 XThR.Tn[10].n7 VGND 0.09695f
C10954 XThR.Tn[10].t13 VGND 0.01887f
C10955 XThR.Tn[10].t63 VGND 0.02067f
C10956 XThR.Tn[10].n8 VGND 0.05047f
C10957 XThR.Tn[10].t50 VGND 0.01881f
C10958 XThR.Tn[10].t60 VGND 0.0206f
C10959 XThR.Tn[10].n9 VGND 0.05251f
C10960 XThR.Tn[10].n10 VGND 0.03689f
C10961 XThR.Tn[10].n11 VGND 0.00674f
C10962 XThR.Tn[10].n12 VGND 0.11838f
C10963 XThR.Tn[10].t48 VGND 0.01887f
C10964 XThR.Tn[10].t41 VGND 0.02067f
C10965 XThR.Tn[10].n13 VGND 0.05047f
C10966 XThR.Tn[10].t23 VGND 0.01881f
C10967 XThR.Tn[10].t36 VGND 0.0206f
C10968 XThR.Tn[10].n14 VGND 0.05251f
C10969 XThR.Tn[10].n15 VGND 0.03689f
C10970 XThR.Tn[10].n16 VGND 0.00674f
C10971 XThR.Tn[10].n17 VGND 0.11838f
C10972 XThR.Tn[10].t65 VGND 0.01887f
C10973 XThR.Tn[10].t58 VGND 0.02067f
C10974 XThR.Tn[10].n18 VGND 0.05047f
C10975 XThR.Tn[10].t40 VGND 0.01881f
C10976 XThR.Tn[10].t55 VGND 0.0206f
C10977 XThR.Tn[10].n19 VGND 0.05251f
C10978 XThR.Tn[10].n20 VGND 0.03689f
C10979 XThR.Tn[10].n21 VGND 0.00674f
C10980 XThR.Tn[10].n22 VGND 0.11838f
C10981 XThR.Tn[10].t30 VGND 0.01887f
C10982 XThR.Tn[10].t26 VGND 0.02067f
C10983 XThR.Tn[10].n23 VGND 0.05047f
C10984 XThR.Tn[10].t70 VGND 0.01881f
C10985 XThR.Tn[10].t21 VGND 0.0206f
C10986 XThR.Tn[10].n24 VGND 0.05251f
C10987 XThR.Tn[10].n25 VGND 0.03689f
C10988 XThR.Tn[10].n26 VGND 0.00674f
C10989 XThR.Tn[10].n27 VGND 0.11838f
C10990 XThR.Tn[10].t67 VGND 0.01887f
C10991 XThR.Tn[10].t59 VGND 0.02067f
C10992 XThR.Tn[10].n28 VGND 0.05047f
C10993 XThR.Tn[10].t42 VGND 0.01881f
C10994 XThR.Tn[10].t56 VGND 0.0206f
C10995 XThR.Tn[10].n29 VGND 0.05251f
C10996 XThR.Tn[10].n30 VGND 0.03689f
C10997 XThR.Tn[10].n31 VGND 0.00674f
C10998 XThR.Tn[10].n32 VGND 0.11838f
C10999 XThR.Tn[10].t44 VGND 0.01887f
C11000 XThR.Tn[10].t15 VGND 0.02067f
C11001 XThR.Tn[10].n33 VGND 0.05047f
C11002 XThR.Tn[10].t18 VGND 0.01881f
C11003 XThR.Tn[10].t12 VGND 0.0206f
C11004 XThR.Tn[10].n34 VGND 0.05251f
C11005 XThR.Tn[10].n35 VGND 0.03689f
C11006 XThR.Tn[10].n36 VGND 0.00674f
C11007 XThR.Tn[10].n37 VGND 0.11838f
C11008 XThR.Tn[10].t14 VGND 0.01887f
C11009 XThR.Tn[10].t69 VGND 0.02067f
C11010 XThR.Tn[10].n38 VGND 0.05047f
C11011 XThR.Tn[10].t51 VGND 0.01881f
C11012 XThR.Tn[10].t66 VGND 0.0206f
C11013 XThR.Tn[10].n39 VGND 0.05251f
C11014 XThR.Tn[10].n40 VGND 0.03689f
C11015 XThR.Tn[10].n41 VGND 0.00674f
C11016 XThR.Tn[10].n42 VGND 0.11838f
C11017 XThR.Tn[10].t17 VGND 0.01887f
C11018 XThR.Tn[10].t24 VGND 0.02067f
C11019 XThR.Tn[10].n43 VGND 0.05047f
C11020 XThR.Tn[10].t53 VGND 0.01881f
C11021 XThR.Tn[10].t20 VGND 0.0206f
C11022 XThR.Tn[10].n44 VGND 0.05251f
C11023 XThR.Tn[10].n45 VGND 0.03689f
C11024 XThR.Tn[10].n46 VGND 0.00674f
C11025 XThR.Tn[10].n47 VGND 0.11838f
C11026 XThR.Tn[10].t33 VGND 0.01887f
C11027 XThR.Tn[10].t43 VGND 0.02067f
C11028 XThR.Tn[10].n48 VGND 0.05047f
C11029 XThR.Tn[10].t73 VGND 0.01881f
C11030 XThR.Tn[10].t38 VGND 0.0206f
C11031 XThR.Tn[10].n49 VGND 0.05251f
C11032 XThR.Tn[10].n50 VGND 0.03689f
C11033 XThR.Tn[10].n51 VGND 0.00674f
C11034 XThR.Tn[10].n52 VGND 0.11838f
C11035 XThR.Tn[10].t28 VGND 0.01887f
C11036 XThR.Tn[10].t61 VGND 0.02067f
C11037 XThR.Tn[10].n53 VGND 0.05047f
C11038 XThR.Tn[10].t62 VGND 0.01881f
C11039 XThR.Tn[10].t57 VGND 0.0206f
C11040 XThR.Tn[10].n54 VGND 0.05251f
C11041 XThR.Tn[10].n55 VGND 0.03689f
C11042 XThR.Tn[10].n56 VGND 0.00674f
C11043 XThR.Tn[10].n57 VGND 0.11838f
C11044 XThR.Tn[10].t46 VGND 0.01887f
C11045 XThR.Tn[10].t35 VGND 0.02067f
C11046 XThR.Tn[10].n58 VGND 0.05047f
C11047 XThR.Tn[10].t19 VGND 0.01881f
C11048 XThR.Tn[10].t32 VGND 0.0206f
C11049 XThR.Tn[10].n59 VGND 0.05251f
C11050 XThR.Tn[10].n60 VGND 0.03689f
C11051 XThR.Tn[10].n61 VGND 0.00674f
C11052 XThR.Tn[10].n62 VGND 0.11838f
C11053 XThR.Tn[10].t16 VGND 0.01887f
C11054 XThR.Tn[10].t72 VGND 0.02067f
C11055 XThR.Tn[10].n63 VGND 0.05047f
C11056 XThR.Tn[10].t52 VGND 0.01881f
C11057 XThR.Tn[10].t68 VGND 0.0206f
C11058 XThR.Tn[10].n64 VGND 0.05251f
C11059 XThR.Tn[10].n65 VGND 0.03689f
C11060 XThR.Tn[10].n66 VGND 0.00674f
C11061 XThR.Tn[10].n67 VGND 0.11838f
C11062 XThR.Tn[10].t31 VGND 0.01887f
C11063 XThR.Tn[10].t27 VGND 0.02067f
C11064 XThR.Tn[10].n68 VGND 0.05047f
C11065 XThR.Tn[10].t71 VGND 0.01881f
C11066 XThR.Tn[10].t22 VGND 0.0206f
C11067 XThR.Tn[10].n69 VGND 0.05251f
C11068 XThR.Tn[10].n70 VGND 0.03689f
C11069 XThR.Tn[10].n71 VGND 0.00674f
C11070 XThR.Tn[10].n72 VGND 0.11838f
C11071 XThR.Tn[10].t49 VGND 0.01887f
C11072 XThR.Tn[10].t45 VGND 0.02067f
C11073 XThR.Tn[10].n73 VGND 0.05047f
C11074 XThR.Tn[10].t25 VGND 0.01881f
C11075 XThR.Tn[10].t39 VGND 0.0206f
C11076 XThR.Tn[10].n74 VGND 0.05251f
C11077 XThR.Tn[10].n75 VGND 0.03689f
C11078 XThR.Tn[10].n76 VGND 0.00674f
C11079 XThR.Tn[10].n77 VGND 0.11838f
C11080 XThR.Tn[10].t29 VGND 0.01887f
C11081 XThR.Tn[10].t37 VGND 0.02067f
C11082 XThR.Tn[10].n78 VGND 0.05047f
C11083 XThR.Tn[10].t64 VGND 0.01881f
C11084 XThR.Tn[10].t34 VGND 0.0206f
C11085 XThR.Tn[10].n79 VGND 0.05251f
C11086 XThR.Tn[10].n80 VGND 0.03689f
C11087 XThR.Tn[10].n81 VGND 0.00674f
C11088 XThR.Tn[10].n82 VGND 0.11838f
C11089 XThR.Tn[10].n83 VGND 0.10758f
C11090 XThR.Tn[10].n84 VGND 0.3312f
C11091 XThR.Tn[10].t5 VGND 0.02415f
C11092 XThR.Tn[10].t3 VGND 0.02415f
C11093 XThR.Tn[10].n85 VGND 0.05218f
C11094 XThR.Tn[10].t0 VGND 0.02415f
C11095 XThR.Tn[10].t6 VGND 0.02415f
C11096 XThR.Tn[10].n86 VGND 0.07942f
C11097 XThR.Tn[10].n87 VGND 0.22051f
C11098 XThR.Tn[10].n88 VGND 0.01087f
C11099 XThC.Tn[3].t1 VGND 0.01826f
C11100 XThC.Tn[3].t0 VGND 0.01826f
C11101 XThC.Tn[3].n0 VGND 0.03685f
C11102 XThC.Tn[3].t3 VGND 0.01826f
C11103 XThC.Tn[3].t2 VGND 0.01826f
C11104 XThC.Tn[3].n1 VGND 0.04312f
C11105 XThC.Tn[3].n2 VGND 0.12934f
C11106 XThC.Tn[3].t11 VGND 0.01187f
C11107 XThC.Tn[3].t10 VGND 0.01187f
C11108 XThC.Tn[3].n3 VGND 0.04503f
C11109 XThC.Tn[3].t9 VGND 0.01187f
C11110 XThC.Tn[3].t8 VGND 0.01187f
C11111 XThC.Tn[3].n4 VGND 0.02703f
C11112 XThC.Tn[3].n5 VGND 0.1287f
C11113 XThC.Tn[3].t7 VGND 0.01187f
C11114 XThC.Tn[3].t6 VGND 0.01187f
C11115 XThC.Tn[3].n6 VGND 0.02703f
C11116 XThC.Tn[3].n7 VGND 0.07956f
C11117 XThC.Tn[3].t5 VGND 0.01187f
C11118 XThC.Tn[3].t4 VGND 0.01187f
C11119 XThC.Tn[3].n8 VGND 0.02703f
C11120 XThC.Tn[3].n9 VGND 0.08979f
C11121 XThC.Tn[3].t12 VGND 0.01447f
C11122 XThC.Tn[3].t42 VGND 0.01581f
C11123 XThC.Tn[3].n10 VGND 0.03529f
C11124 XThC.Tn[3].n11 VGND 0.02417f
C11125 XThC.Tn[3].n12 VGND 0.07935f
C11126 XThC.Tn[3].t30 VGND 0.01447f
C11127 XThC.Tn[3].t27 VGND 0.01581f
C11128 XThC.Tn[3].n13 VGND 0.03529f
C11129 XThC.Tn[3].n14 VGND 0.02417f
C11130 XThC.Tn[3].n15 VGND 0.07957f
C11131 XThC.Tn[3].n16 VGND 0.13113f
C11132 XThC.Tn[3].t35 VGND 0.01447f
C11133 XThC.Tn[3].t29 VGND 0.01581f
C11134 XThC.Tn[3].n17 VGND 0.03529f
C11135 XThC.Tn[3].n18 VGND 0.02417f
C11136 XThC.Tn[3].n19 VGND 0.07957f
C11137 XThC.Tn[3].n20 VGND 0.13113f
C11138 XThC.Tn[3].t36 VGND 0.01447f
C11139 XThC.Tn[3].t31 VGND 0.01581f
C11140 XThC.Tn[3].n21 VGND 0.03529f
C11141 XThC.Tn[3].n22 VGND 0.02417f
C11142 XThC.Tn[3].n23 VGND 0.07957f
C11143 XThC.Tn[3].n24 VGND 0.13113f
C11144 XThC.Tn[3].t23 VGND 0.01447f
C11145 XThC.Tn[3].t20 VGND 0.01581f
C11146 XThC.Tn[3].n25 VGND 0.03529f
C11147 XThC.Tn[3].n26 VGND 0.02417f
C11148 XThC.Tn[3].n27 VGND 0.07957f
C11149 XThC.Tn[3].n28 VGND 0.13113f
C11150 XThC.Tn[3].t24 VGND 0.01447f
C11151 XThC.Tn[3].t21 VGND 0.01581f
C11152 XThC.Tn[3].n29 VGND 0.03529f
C11153 XThC.Tn[3].n30 VGND 0.02417f
C11154 XThC.Tn[3].n31 VGND 0.07957f
C11155 XThC.Tn[3].n32 VGND 0.13113f
C11156 XThC.Tn[3].t40 VGND 0.01447f
C11157 XThC.Tn[3].t34 VGND 0.01581f
C11158 XThC.Tn[3].n33 VGND 0.03529f
C11159 XThC.Tn[3].n34 VGND 0.02417f
C11160 XThC.Tn[3].n35 VGND 0.07957f
C11161 XThC.Tn[3].n36 VGND 0.13113f
C11162 XThC.Tn[3].t15 VGND 0.01447f
C11163 XThC.Tn[3].t43 VGND 0.01581f
C11164 XThC.Tn[3].n37 VGND 0.03529f
C11165 XThC.Tn[3].n38 VGND 0.02417f
C11166 XThC.Tn[3].n39 VGND 0.07957f
C11167 XThC.Tn[3].n40 VGND 0.13113f
C11168 XThC.Tn[3].t17 VGND 0.01447f
C11169 XThC.Tn[3].t13 VGND 0.01581f
C11170 XThC.Tn[3].n41 VGND 0.03529f
C11171 XThC.Tn[3].n42 VGND 0.02417f
C11172 XThC.Tn[3].n43 VGND 0.07957f
C11173 XThC.Tn[3].n44 VGND 0.13113f
C11174 XThC.Tn[3].t37 VGND 0.01447f
C11175 XThC.Tn[3].t32 VGND 0.01581f
C11176 XThC.Tn[3].n45 VGND 0.03529f
C11177 XThC.Tn[3].n46 VGND 0.02417f
C11178 XThC.Tn[3].n47 VGND 0.07957f
C11179 XThC.Tn[3].n48 VGND 0.13113f
C11180 XThC.Tn[3].t39 VGND 0.01447f
C11181 XThC.Tn[3].t33 VGND 0.01581f
C11182 XThC.Tn[3].n49 VGND 0.03529f
C11183 XThC.Tn[3].n50 VGND 0.02417f
C11184 XThC.Tn[3].n51 VGND 0.07957f
C11185 XThC.Tn[3].n52 VGND 0.13113f
C11186 XThC.Tn[3].t18 VGND 0.01447f
C11187 XThC.Tn[3].t14 VGND 0.01581f
C11188 XThC.Tn[3].n53 VGND 0.03529f
C11189 XThC.Tn[3].n54 VGND 0.02417f
C11190 XThC.Tn[3].n55 VGND 0.07957f
C11191 XThC.Tn[3].n56 VGND 0.13113f
C11192 XThC.Tn[3].t26 VGND 0.01447f
C11193 XThC.Tn[3].t22 VGND 0.01581f
C11194 XThC.Tn[3].n57 VGND 0.03529f
C11195 XThC.Tn[3].n58 VGND 0.02417f
C11196 XThC.Tn[3].n59 VGND 0.07957f
C11197 XThC.Tn[3].n60 VGND 0.13113f
C11198 XThC.Tn[3].t28 VGND 0.01447f
C11199 XThC.Tn[3].t25 VGND 0.01581f
C11200 XThC.Tn[3].n61 VGND 0.03529f
C11201 XThC.Tn[3].n62 VGND 0.02417f
C11202 XThC.Tn[3].n63 VGND 0.07957f
C11203 XThC.Tn[3].n64 VGND 0.13113f
C11204 XThC.Tn[3].t41 VGND 0.01447f
C11205 XThC.Tn[3].t38 VGND 0.01581f
C11206 XThC.Tn[3].n65 VGND 0.03529f
C11207 XThC.Tn[3].n66 VGND 0.02417f
C11208 XThC.Tn[3].n67 VGND 0.07957f
C11209 XThC.Tn[3].n68 VGND 0.13113f
C11210 XThC.Tn[3].t19 VGND 0.01447f
C11211 XThC.Tn[3].t16 VGND 0.01581f
C11212 XThC.Tn[3].n69 VGND 0.03529f
C11213 XThC.Tn[3].n70 VGND 0.02417f
C11214 XThC.Tn[3].n71 VGND 0.07957f
C11215 XThC.Tn[3].n72 VGND 0.13113f
C11216 XThC.Tn[3].n73 VGND 0.77119f
C11217 XThC.Tn[3].n74 VGND 0.1112f
C11218 XThC.Tn[1].t7 VGND 0.01715f
C11219 XThC.Tn[1].t6 VGND 0.01715f
C11220 XThC.Tn[1].n0 VGND 0.03462f
C11221 XThC.Tn[1].t5 VGND 0.01715f
C11222 XThC.Tn[1].t4 VGND 0.01715f
C11223 XThC.Tn[1].n1 VGND 0.04051f
C11224 XThC.Tn[1].n2 VGND 0.12152f
C11225 XThC.Tn[1].t9 VGND 0.01115f
C11226 XThC.Tn[1].t8 VGND 0.01115f
C11227 XThC.Tn[1].n3 VGND 0.02539f
C11228 XThC.Tn[1].t11 VGND 0.01115f
C11229 XThC.Tn[1].t10 VGND 0.01115f
C11230 XThC.Tn[1].n4 VGND 0.02539f
C11231 XThC.Tn[1].t1 VGND 0.01115f
C11232 XThC.Tn[1].t0 VGND 0.01115f
C11233 XThC.Tn[1].n5 VGND 0.02539f
C11234 XThC.Tn[1].t3 VGND 0.01115f
C11235 XThC.Tn[1].t2 VGND 0.01115f
C11236 XThC.Tn[1].n6 VGND 0.04231f
C11237 XThC.Tn[1].n7 VGND 0.12091f
C11238 XThC.Tn[1].n8 VGND 0.07475f
C11239 XThC.Tn[1].n9 VGND 0.08436f
C11240 XThC.Tn[1].t31 VGND 0.0136f
C11241 XThC.Tn[1].t29 VGND 0.01485f
C11242 XThC.Tn[1].n10 VGND 0.03315f
C11243 XThC.Tn[1].n11 VGND 0.02271f
C11244 XThC.Tn[1].n12 VGND 0.07455f
C11245 XThC.Tn[1].t17 VGND 0.0136f
C11246 XThC.Tn[1].t14 VGND 0.01485f
C11247 XThC.Tn[1].n13 VGND 0.03315f
C11248 XThC.Tn[1].n14 VGND 0.02271f
C11249 XThC.Tn[1].n15 VGND 0.07475f
C11250 XThC.Tn[1].n16 VGND 0.1232f
C11251 XThC.Tn[1].t22 VGND 0.0136f
C11252 XThC.Tn[1].t16 VGND 0.01485f
C11253 XThC.Tn[1].n17 VGND 0.03315f
C11254 XThC.Tn[1].n18 VGND 0.02271f
C11255 XThC.Tn[1].n19 VGND 0.07475f
C11256 XThC.Tn[1].n20 VGND 0.1232f
C11257 XThC.Tn[1].t23 VGND 0.0136f
C11258 XThC.Tn[1].t18 VGND 0.01485f
C11259 XThC.Tn[1].n21 VGND 0.03315f
C11260 XThC.Tn[1].n22 VGND 0.02271f
C11261 XThC.Tn[1].n23 VGND 0.07475f
C11262 XThC.Tn[1].n24 VGND 0.1232f
C11263 XThC.Tn[1].t42 VGND 0.0136f
C11264 XThC.Tn[1].t39 VGND 0.01485f
C11265 XThC.Tn[1].n25 VGND 0.03315f
C11266 XThC.Tn[1].n26 VGND 0.02271f
C11267 XThC.Tn[1].n27 VGND 0.07475f
C11268 XThC.Tn[1].n28 VGND 0.1232f
C11269 XThC.Tn[1].t43 VGND 0.0136f
C11270 XThC.Tn[1].t40 VGND 0.01485f
C11271 XThC.Tn[1].n29 VGND 0.03315f
C11272 XThC.Tn[1].n30 VGND 0.02271f
C11273 XThC.Tn[1].n31 VGND 0.07475f
C11274 XThC.Tn[1].n32 VGND 0.1232f
C11275 XThC.Tn[1].t27 VGND 0.0136f
C11276 XThC.Tn[1].t21 VGND 0.01485f
C11277 XThC.Tn[1].n33 VGND 0.03315f
C11278 XThC.Tn[1].n34 VGND 0.02271f
C11279 XThC.Tn[1].n35 VGND 0.07475f
C11280 XThC.Tn[1].n36 VGND 0.1232f
C11281 XThC.Tn[1].t34 VGND 0.0136f
C11282 XThC.Tn[1].t30 VGND 0.01485f
C11283 XThC.Tn[1].n37 VGND 0.03315f
C11284 XThC.Tn[1].n38 VGND 0.02271f
C11285 XThC.Tn[1].n39 VGND 0.07475f
C11286 XThC.Tn[1].n40 VGND 0.1232f
C11287 XThC.Tn[1].t36 VGND 0.0136f
C11288 XThC.Tn[1].t32 VGND 0.01485f
C11289 XThC.Tn[1].n41 VGND 0.03315f
C11290 XThC.Tn[1].n42 VGND 0.02271f
C11291 XThC.Tn[1].n43 VGND 0.07475f
C11292 XThC.Tn[1].n44 VGND 0.1232f
C11293 XThC.Tn[1].t24 VGND 0.0136f
C11294 XThC.Tn[1].t19 VGND 0.01485f
C11295 XThC.Tn[1].n45 VGND 0.03315f
C11296 XThC.Tn[1].n46 VGND 0.02271f
C11297 XThC.Tn[1].n47 VGND 0.07475f
C11298 XThC.Tn[1].n48 VGND 0.1232f
C11299 XThC.Tn[1].t26 VGND 0.0136f
C11300 XThC.Tn[1].t20 VGND 0.01485f
C11301 XThC.Tn[1].n49 VGND 0.03315f
C11302 XThC.Tn[1].n50 VGND 0.02271f
C11303 XThC.Tn[1].n51 VGND 0.07475f
C11304 XThC.Tn[1].n52 VGND 0.1232f
C11305 XThC.Tn[1].t37 VGND 0.0136f
C11306 XThC.Tn[1].t33 VGND 0.01485f
C11307 XThC.Tn[1].n53 VGND 0.03315f
C11308 XThC.Tn[1].n54 VGND 0.02271f
C11309 XThC.Tn[1].n55 VGND 0.07475f
C11310 XThC.Tn[1].n56 VGND 0.1232f
C11311 XThC.Tn[1].t13 VGND 0.0136f
C11312 XThC.Tn[1].t41 VGND 0.01485f
C11313 XThC.Tn[1].n57 VGND 0.03315f
C11314 XThC.Tn[1].n58 VGND 0.02271f
C11315 XThC.Tn[1].n59 VGND 0.07475f
C11316 XThC.Tn[1].n60 VGND 0.1232f
C11317 XThC.Tn[1].t15 VGND 0.0136f
C11318 XThC.Tn[1].t12 VGND 0.01485f
C11319 XThC.Tn[1].n61 VGND 0.03315f
C11320 XThC.Tn[1].n62 VGND 0.02271f
C11321 XThC.Tn[1].n63 VGND 0.07475f
C11322 XThC.Tn[1].n64 VGND 0.1232f
C11323 XThC.Tn[1].t28 VGND 0.0136f
C11324 XThC.Tn[1].t25 VGND 0.01485f
C11325 XThC.Tn[1].n65 VGND 0.03315f
C11326 XThC.Tn[1].n66 VGND 0.02271f
C11327 XThC.Tn[1].n67 VGND 0.07475f
C11328 XThC.Tn[1].n68 VGND 0.1232f
C11329 XThC.Tn[1].t38 VGND 0.0136f
C11330 XThC.Tn[1].t35 VGND 0.01485f
C11331 XThC.Tn[1].n69 VGND 0.03315f
C11332 XThC.Tn[1].n70 VGND 0.02271f
C11333 XThC.Tn[1].n71 VGND 0.07475f
C11334 XThC.Tn[1].n72 VGND 0.1232f
C11335 XThC.Tn[1].n73 VGND 0.62603f
C11336 XThC.Tn[1].n74 VGND 0.11896f
C11337 Vbias.t2 VGND 0.26877f
C11338 Vbias.t1 VGND 1.05767f
C11339 Vbias.n0 VGND 1.97597f
C11340 Vbias.t3 VGND 0.05767f
C11341 Vbias.t5 VGND 0.05767f
C11342 Vbias.n1 VGND 0.3885f
C11343 Vbias.t4 VGND 0.05767f
C11344 Vbias.t0 VGND 0.05767f
C11345 Vbias.n2 VGND 0.3885f
C11346 Vbias.n3 VGND 1.16485f
C11347 Vbias.n4 VGND 0.8158f
C11348 Vbias.n5 VGND 0.8811f
C11349 Vbias.t181 VGND 0.2822f
C11350 Vbias.n6 VGND 0.27871f
C11351 Vbias.t110 VGND 0.2822f
C11352 Vbias.n7 VGND 0.27871f
C11353 Vbias.n8 VGND 0.07848f
C11354 Vbias.n9 VGND 0.29662f
C11355 Vbias.t146 VGND 0.2822f
C11356 Vbias.n10 VGND 0.27871f
C11357 Vbias.t238 VGND 0.2822f
C11358 Vbias.n11 VGND 0.27871f
C11359 Vbias.n12 VGND 0.29662f
C11360 Vbias.t210 VGND 0.2822f
C11361 Vbias.n13 VGND 0.27871f
C11362 Vbias.n14 VGND 0.07848f
C11363 Vbias.t24 VGND 0.2822f
C11364 Vbias.n15 VGND 0.27871f
C11365 Vbias.t12 VGND 0.2822f
C11366 Vbias.n16 VGND 0.27871f
C11367 Vbias.n17 VGND 0.29662f
C11368 Vbias.t193 VGND 0.2822f
C11369 Vbias.n18 VGND 0.27871f
C11370 Vbias.n19 VGND 0.16575f
C11371 Vbias.n20 VGND 0.16575f
C11372 Vbias.t173 VGND 0.2822f
C11373 Vbias.n21 VGND 0.27871f
C11374 Vbias.n22 VGND 0.29662f
C11375 Vbias.t248 VGND 0.2822f
C11376 Vbias.n23 VGND 0.27871f
C11377 Vbias.t95 VGND 0.2822f
C11378 Vbias.n24 VGND 0.27871f
C11379 Vbias.n25 VGND 0.29662f
C11380 Vbias.t25 VGND 0.2822f
C11381 Vbias.n26 VGND 0.27871f
C11382 Vbias.t258 VGND 0.2822f
C11383 Vbias.n27 VGND 0.27871f
C11384 Vbias.n28 VGND 0.29662f
C11385 Vbias.t75 VGND 0.2822f
C11386 Vbias.n29 VGND 0.27871f
C11387 Vbias.t246 VGND 0.2822f
C11388 Vbias.n30 VGND 0.27871f
C11389 Vbias.n31 VGND 0.29662f
C11390 Vbias.t171 VGND 0.2822f
C11391 Vbias.n32 VGND 0.27871f
C11392 Vbias.t96 VGND 0.2822f
C11393 Vbias.n33 VGND 0.27871f
C11394 Vbias.n34 VGND 0.29662f
C11395 Vbias.t169 VGND 0.2822f
C11396 Vbias.n35 VGND 0.27871f
C11397 Vbias.t147 VGND 0.2822f
C11398 Vbias.n36 VGND 0.27871f
C11399 Vbias.n37 VGND 0.29662f
C11400 Vbias.t76 VGND 0.2822f
C11401 Vbias.n38 VGND 0.27871f
C11402 Vbias.t247 VGND 0.2822f
C11403 Vbias.n39 VGND 0.27871f
C11404 Vbias.n40 VGND 0.29662f
C11405 Vbias.t60 VGND 0.2822f
C11406 Vbias.n41 VGND 0.27871f
C11407 Vbias.t227 VGND 0.2822f
C11408 Vbias.n42 VGND 0.27871f
C11409 Vbias.n43 VGND 0.29662f
C11410 Vbias.t156 VGND 0.2822f
C11411 Vbias.n44 VGND 0.27871f
C11412 Vbias.t69 VGND 0.2822f
C11413 Vbias.n45 VGND 0.27871f
C11414 Vbias.n46 VGND 0.29662f
C11415 Vbias.t141 VGND 0.2822f
C11416 Vbias.n47 VGND 0.27871f
C11417 Vbias.t56 VGND 0.2822f
C11418 Vbias.n48 VGND 0.27871f
C11419 Vbias.n49 VGND 0.29662f
C11420 Vbias.t242 VGND 0.2822f
C11421 Vbias.n50 VGND 0.27871f
C11422 Vbias.t229 VGND 0.2822f
C11423 Vbias.n51 VGND 0.27871f
C11424 Vbias.n52 VGND 0.29662f
C11425 Vbias.t41 VGND 0.2822f
C11426 Vbias.n53 VGND 0.27871f
C11427 Vbias.t201 VGND 0.2822f
C11428 Vbias.n54 VGND 0.27871f
C11429 Vbias.n55 VGND 0.29662f
C11430 Vbias.t130 VGND 0.2822f
C11431 Vbias.n56 VGND 0.27871f
C11432 Vbias.t57 VGND 0.2822f
C11433 Vbias.n57 VGND 0.27871f
C11434 Vbias.t129 VGND 0.2822f
C11435 Vbias.n58 VGND 0.27871f
C11436 Vbias.n59 VGND 0.03744f
C11437 Vbias.t87 VGND 0.2822f
C11438 Vbias.n60 VGND 0.27871f
C11439 Vbias.t225 VGND 0.2822f
C11440 Vbias.n61 VGND 0.27871f
C11441 Vbias.n62 VGND 0.07848f
C11442 Vbias.n63 VGND 0.16575f
C11443 Vbias.t205 VGND 0.2822f
C11444 Vbias.n64 VGND 0.27871f
C11445 Vbias.n65 VGND 0.07848f
C11446 Vbias.n66 VGND 0.16575f
C11447 Vbias.t52 VGND 0.2822f
C11448 Vbias.n67 VGND 0.27871f
C11449 Vbias.n68 VGND 0.07848f
C11450 Vbias.n69 VGND 0.16575f
C11451 Vbias.t32 VGND 0.2822f
C11452 Vbias.n70 VGND 0.27871f
C11453 Vbias.n71 VGND 0.07848f
C11454 Vbias.n72 VGND 0.16575f
C11455 Vbias.t199 VGND 0.2822f
C11456 Vbias.n73 VGND 0.27871f
C11457 Vbias.n74 VGND 0.07848f
C11458 Vbias.n75 VGND 0.16575f
C11459 Vbias.t125 VGND 0.2822f
C11460 Vbias.n76 VGND 0.27871f
C11461 Vbias.n77 VGND 0.07848f
C11462 Vbias.n78 VGND 0.16575f
C11463 Vbias.t102 VGND 0.2822f
C11464 Vbias.n79 VGND 0.27871f
C11465 Vbias.n80 VGND 0.07848f
C11466 Vbias.n81 VGND 0.16575f
C11467 Vbias.t18 VGND 0.2822f
C11468 Vbias.n82 VGND 0.27871f
C11469 Vbias.n83 VGND 0.07848f
C11470 Vbias.n84 VGND 0.16575f
C11471 Vbias.t183 VGND 0.2822f
C11472 Vbias.n85 VGND 0.27871f
C11473 Vbias.n86 VGND 0.07848f
C11474 Vbias.n87 VGND 0.16575f
C11475 Vbias.t99 VGND 0.2822f
C11476 Vbias.n88 VGND 0.27871f
C11477 Vbias.n89 VGND 0.07848f
C11478 Vbias.n90 VGND 0.16575f
C11479 Vbias.t14 VGND 0.2822f
C11480 Vbias.n91 VGND 0.27871f
C11481 Vbias.n92 VGND 0.07848f
C11482 Vbias.n93 VGND 0.16575f
C11483 Vbias.t262 VGND 0.2822f
C11484 Vbias.n94 VGND 0.27871f
C11485 Vbias.n95 VGND 0.07848f
C11486 Vbias.n96 VGND 0.16575f
C11487 Vbias.t160 VGND 0.2822f
C11488 Vbias.n97 VGND 0.27871f
C11489 Vbias.n98 VGND 0.07848f
C11490 Vbias.n99 VGND 0.16575f
C11491 Vbias.n100 VGND 0.07618f
C11492 Vbias.n101 VGND 0.29662f
C11493 Vbias.t16 VGND 0.2822f
C11494 Vbias.n102 VGND 0.27871f
C11495 Vbias.t88 VGND 0.2822f
C11496 Vbias.n103 VGND 0.27871f
C11497 Vbias.n104 VGND 0.29662f
C11498 Vbias.t17 VGND 0.2822f
C11499 Vbias.n105 VGND 0.27871f
C11500 Vbias.t113 VGND 0.2822f
C11501 Vbias.n106 VGND 0.27871f
C11502 Vbias.n107 VGND 0.29662f
C11503 Vbias.t185 VGND 0.2822f
C11504 Vbias.n108 VGND 0.27871f
C11505 Vbias.t196 VGND 0.2822f
C11506 Vbias.n109 VGND 0.27871f
C11507 Vbias.n110 VGND 0.29662f
C11508 Vbias.t124 VGND 0.2822f
C11509 Vbias.n111 VGND 0.27871f
C11510 Vbias.t213 VGND 0.2822f
C11511 Vbias.n112 VGND 0.27871f
C11512 Vbias.n113 VGND 0.29662f
C11513 Vbias.t29 VGND 0.2822f
C11514 Vbias.n114 VGND 0.27871f
C11515 Vbias.t112 VGND 0.2822f
C11516 Vbias.n115 VGND 0.27871f
C11517 Vbias.n116 VGND 0.29662f
C11518 Vbias.t40 VGND 0.2822f
C11519 Vbias.n117 VGND 0.27871f
C11520 Vbias.t127 VGND 0.2822f
C11521 Vbias.n118 VGND 0.27871f
C11522 Vbias.n119 VGND 0.29662f
C11523 Vbias.t200 VGND 0.2822f
C11524 Vbias.n120 VGND 0.27871f
C11525 Vbias.t33 VGND 0.2822f
C11526 Vbias.n121 VGND 0.27871f
C11527 Vbias.n122 VGND 0.29662f
C11528 Vbias.t219 VGND 0.2822f
C11529 Vbias.n123 VGND 0.27871f
C11530 Vbias.t240 VGND 0.2822f
C11531 Vbias.n124 VGND 0.27871f
C11532 Vbias.n125 VGND 0.29662f
C11533 Vbias.t53 VGND 0.2822f
C11534 Vbias.n126 VGND 0.27871f
C11535 Vbias.t126 VGND 0.2822f
C11536 Vbias.n127 VGND 0.27871f
C11537 Vbias.n128 VGND 0.29662f
C11538 Vbias.t54 VGND 0.2822f
C11539 Vbias.n129 VGND 0.27871f
C11540 Vbias.t144 VGND 0.2822f
C11541 Vbias.n130 VGND 0.27871f
C11542 Vbias.n131 VGND 0.29662f
C11543 Vbias.t217 VGND 0.2822f
C11544 Vbias.n132 VGND 0.27871f
C11545 Vbias.t239 VGND 0.2822f
C11546 Vbias.n133 VGND 0.27871f
C11547 Vbias.n134 VGND 0.29662f
C11548 Vbias.t166 VGND 0.2822f
C11549 Vbias.n135 VGND 0.27871f
C11550 Vbias.t62 VGND 0.2822f
C11551 Vbias.n136 VGND 0.27871f
C11552 Vbias.n137 VGND 0.29662f
C11553 Vbias.t133 VGND 0.2822f
C11554 Vbias.n138 VGND 0.27871f
C11555 Vbias.t153 VGND 0.2822f
C11556 Vbias.n139 VGND 0.27871f
C11557 Vbias.n140 VGND 0.29662f
C11558 Vbias.t81 VGND 0.2822f
C11559 Vbias.n141 VGND 0.27871f
C11560 Vbias.t92 VGND 0.2822f
C11561 Vbias.n142 VGND 0.27871f
C11562 Vbias.n143 VGND 0.29662f
C11563 Vbias.t20 VGND 0.2822f
C11564 Vbias.n144 VGND 0.27871f
C11565 Vbias.t121 VGND 0.2822f
C11566 Vbias.n145 VGND 0.27871f
C11567 Vbias.t49 VGND 0.2822f
C11568 Vbias.n146 VGND 0.27871f
C11569 Vbias.n147 VGND 0.07618f
C11570 Vbias.n148 VGND 0.29662f
C11571 Vbias.t82 VGND 0.2822f
C11572 Vbias.n149 VGND 0.27871f
C11573 Vbias.t154 VGND 0.2822f
C11574 Vbias.n150 VGND 0.27871f
C11575 Vbias.n151 VGND 0.29662f
C11576 Vbias.t122 VGND 0.2822f
C11577 Vbias.n152 VGND 0.27871f
C11578 Vbias.t222 VGND 0.2822f
C11579 Vbias.n153 VGND 0.27871f
C11580 Vbias.n154 VGND 0.29662f
C11581 Vbias.t257 VGND 0.2822f
C11582 Vbias.n155 VGND 0.27871f
C11583 Vbias.t8 VGND 0.2822f
C11584 Vbias.n156 VGND 0.27871f
C11585 Vbias.n157 VGND 0.29662f
C11586 Vbias.t235 VGND 0.2822f
C11587 Vbias.n158 VGND 0.27871f
C11588 Vbias.t63 VGND 0.2822f
C11589 Vbias.n159 VGND 0.27871f
C11590 Vbias.n160 VGND 0.29662f
C11591 Vbias.t93 VGND 0.2822f
C11592 Vbias.n161 VGND 0.27871f
C11593 Vbias.t179 VGND 0.2822f
C11594 Vbias.n162 VGND 0.27871f
C11595 Vbias.n163 VGND 0.29662f
C11596 Vbias.t150 VGND 0.2822f
C11597 Vbias.n164 VGND 0.27871f
C11598 Vbias.t237 VGND 0.2822f
C11599 Vbias.n165 VGND 0.27871f
C11600 Vbias.n166 VGND 0.29662f
C11601 Vbias.t11 VGND 0.2822f
C11602 Vbias.n167 VGND 0.27871f
C11603 Vbias.t98 VGND 0.2822f
C11604 Vbias.n168 VGND 0.27871f
C11605 Vbias.n169 VGND 0.29662f
C11606 Vbias.t68 VGND 0.2822f
C11607 Vbias.n170 VGND 0.27871f
C11608 Vbias.t91 VGND 0.2822f
C11609 Vbias.n171 VGND 0.27871f
C11610 Vbias.n172 VGND 0.29662f
C11611 Vbias.t118 VGND 0.2822f
C11612 Vbias.n173 VGND 0.27871f
C11613 Vbias.t190 VGND 0.2822f
C11614 Vbias.n174 VGND 0.27871f
C11615 Vbias.n175 VGND 0.29662f
C11616 Vbias.t164 VGND 0.2822f
C11617 Vbias.n176 VGND 0.27871f
C11618 Vbias.t251 VGND 0.2822f
C11619 Vbias.n177 VGND 0.27871f
C11620 Vbias.n178 VGND 0.29662f
C11621 Vbias.t27 VGND 0.2822f
C11622 Vbias.n179 VGND 0.27871f
C11623 Vbias.t44 VGND 0.2822f
C11624 Vbias.n180 VGND 0.27871f
C11625 Vbias.n181 VGND 0.29662f
C11626 Vbias.t21 VGND 0.2822f
C11627 Vbias.n182 VGND 0.27871f
C11628 Vbias.t168 VGND 0.2822f
C11629 Vbias.n183 VGND 0.27871f
C11630 Vbias.n184 VGND 0.29662f
C11631 Vbias.t197 VGND 0.2822f
C11632 Vbias.n185 VGND 0.27871f
C11633 Vbias.t220 VGND 0.2822f
C11634 Vbias.n186 VGND 0.27871f
C11635 Vbias.n187 VGND 0.29662f
C11636 Vbias.t187 VGND 0.2822f
C11637 Vbias.n188 VGND 0.27871f
C11638 Vbias.t105 VGND 0.2822f
C11639 Vbias.n189 VGND 0.27871f
C11640 Vbias.n190 VGND 0.29662f
C11641 Vbias.t137 VGND 0.2822f
C11642 Vbias.n191 VGND 0.27871f
C11643 Vbias.n192 VGND 0.07848f
C11644 Vbias.n193 VGND 0.29662f
C11645 Vbias.t64 VGND 0.2822f
C11646 Vbias.n194 VGND 0.27871f
C11647 Vbias.t9 VGND 0.2822f
C11648 Vbias.n195 VGND 0.27871f
C11649 Vbias.n196 VGND 0.07618f
C11650 Vbias.t83 VGND 0.2822f
C11651 Vbias.n197 VGND 0.27871f
C11652 Vbias.n198 VGND 0.07848f
C11653 Vbias.n199 VGND 0.16575f
C11654 Vbias.t180 VGND 0.2822f
C11655 Vbias.n200 VGND 0.27871f
C11656 Vbias.n201 VGND 0.07848f
C11657 Vbias.n202 VGND 0.16575f
C11658 Vbias.t188 VGND 0.2822f
C11659 Vbias.n203 VGND 0.27871f
C11660 Vbias.n204 VGND 0.07848f
C11661 Vbias.n205 VGND 0.16575f
C11662 Vbias.t23 VGND 0.2822f
C11663 Vbias.n206 VGND 0.27871f
C11664 Vbias.n207 VGND 0.07848f
C11665 Vbias.n208 VGND 0.16575f
C11666 Vbias.t107 VGND 0.2822f
C11667 Vbias.n209 VGND 0.27871f
C11668 Vbias.n210 VGND 0.07848f
C11669 Vbias.n211 VGND 0.16575f
C11670 Vbias.t192 VGND 0.2822f
C11671 Vbias.n212 VGND 0.27871f
C11672 Vbias.n213 VGND 0.07848f
C11673 Vbias.n214 VGND 0.16575f
C11674 Vbias.t28 VGND 0.2822f
C11675 Vbias.n215 VGND 0.27871f
C11676 Vbias.n216 VGND 0.07848f
C11677 Vbias.n217 VGND 0.16575f
C11678 Vbias.t45 VGND 0.2822f
C11679 Vbias.n218 VGND 0.27871f
C11680 Vbias.n219 VGND 0.07848f
C11681 Vbias.n220 VGND 0.16575f
C11682 Vbias.t119 VGND 0.2822f
C11683 Vbias.n221 VGND 0.27871f
C11684 Vbias.n222 VGND 0.07848f
C11685 Vbias.n223 VGND 0.16575f
C11686 Vbias.t211 VGND 0.2822f
C11687 Vbias.n224 VGND 0.27871f
C11688 Vbias.n225 VGND 0.07848f
C11689 Vbias.n226 VGND 0.16575f
C11690 Vbias.t233 VGND 0.2822f
C11691 Vbias.n227 VGND 0.27871f
C11692 Vbias.n228 VGND 0.07848f
C11693 Vbias.n229 VGND 0.16575f
C11694 Vbias.t123 VGND 0.2822f
C11695 Vbias.n230 VGND 0.27871f
C11696 Vbias.n231 VGND 0.07848f
C11697 Vbias.n232 VGND 0.16575f
C11698 Vbias.t149 VGND 0.2822f
C11699 Vbias.n233 VGND 0.27871f
C11700 Vbias.n234 VGND 0.07848f
C11701 Vbias.n235 VGND 0.16575f
C11702 Vbias.t161 VGND 0.2822f
C11703 Vbias.n236 VGND 0.27871f
C11704 Vbias.n237 VGND 0.29662f
C11705 Vbias.t232 VGND 0.2822f
C11706 Vbias.n238 VGND 0.27871f
C11707 Vbias.n239 VGND 0.8811f
C11708 Vbias.t80 VGND 0.2822f
C11709 Vbias.n240 VGND 0.27871f
C11710 Vbias.n241 VGND 0.29662f
C11711 Vbias.t191 VGND 0.2822f
C11712 Vbias.n242 VGND 0.27871f
C11713 Vbias.t172 VGND 0.2822f
C11714 Vbias.n243 VGND 0.27871f
C11715 Vbias.n244 VGND 0.29662f
C11716 Vbias.t51 VGND 0.2822f
C11717 Vbias.n245 VGND 0.27871f
C11718 Vbias.t162 VGND 0.2822f
C11719 Vbias.n246 VGND 0.27871f
C11720 Vbias.n247 VGND 0.29662f
C11721 Vbias.t22 VGND 0.2822f
C11722 Vbias.n248 VGND 0.27871f
C11723 Vbias.t256 VGND 0.2822f
C11724 Vbias.n249 VGND 0.27871f
C11725 Vbias.n250 VGND 0.29662f
C11726 Vbias.t136 VGND 0.2822f
C11727 Vbias.n251 VGND 0.27871f
C11728 Vbias.t46 VGND 0.2822f
C11729 Vbias.n252 VGND 0.27871f
C11730 Vbias.n253 VGND 0.29662f
C11731 Vbias.t167 VGND 0.2822f
C11732 Vbias.n254 VGND 0.27871f
C11733 Vbias.t94 VGND 0.2822f
C11734 Vbias.n255 VGND 0.27871f
C11735 Vbias.n256 VGND 0.29662f
C11736 Vbias.t234 VGND 0.2822f
C11737 Vbias.n257 VGND 0.27871f
C11738 Vbias.t212 VGND 0.2822f
C11739 Vbias.n258 VGND 0.27871f
C11740 Vbias.n259 VGND 0.29662f
C11741 Vbias.t74 VGND 0.2822f
C11742 Vbias.n260 VGND 0.27871f
C11743 Vbias.t244 VGND 0.2822f
C11744 Vbias.n261 VGND 0.27871f
C11745 Vbias.n262 VGND 0.29662f
C11746 Vbias.t120 VGND 0.2822f
C11747 Vbias.n263 VGND 0.27871f
C11748 Vbias.t36 VGND 0.2822f
C11749 Vbias.n264 VGND 0.27871f
C11750 Vbias.n265 VGND 0.29662f
C11751 Vbias.t155 VGND 0.2822f
C11752 Vbias.n266 VGND 0.27871f
C11753 Vbias.t66 VGND 0.2822f
C11754 Vbias.n267 VGND 0.27871f
C11755 Vbias.n268 VGND 0.29662f
C11756 Vbias.t208 VGND 0.2822f
C11757 Vbias.n269 VGND 0.27871f
C11758 Vbias.t117 VGND 0.2822f
C11759 Vbias.n270 VGND 0.27871f
C11760 Vbias.n271 VGND 0.29662f
C11761 Vbias.t241 VGND 0.2822f
C11762 Vbias.n272 VGND 0.27871f
C11763 Vbias.t226 VGND 0.2822f
C11764 Vbias.n273 VGND 0.27871f
C11765 Vbias.n274 VGND 0.29662f
C11766 Vbias.t108 VGND 0.2822f
C11767 Vbias.n275 VGND 0.27871f
C11768 Vbias.t10 VGND 0.2822f
C11769 Vbias.n276 VGND 0.27871f
C11770 Vbias.n277 VGND 0.29662f
C11771 Vbias.t128 VGND 0.2822f
C11772 Vbias.n278 VGND 0.27871f
C11773 Vbias.t55 VGND 0.2822f
C11774 Vbias.n279 VGND 0.27871f
C11775 Vbias.t189 VGND 0.2822f
C11776 Vbias.n280 VGND 0.27871f
C11777 Vbias.n281 VGND 0.07618f
C11778 Vbias.n282 VGND 0.29662f
C11779 Vbias.n283 VGND 0.29662f
C11780 Vbias.t186 VGND 0.2822f
C11781 Vbias.n284 VGND 0.27871f
C11782 Vbias.t85 VGND 0.2822f
C11783 Vbias.n285 VGND 0.27871f
C11784 Vbias.n286 VGND 0.29662f
C11785 Vbias.t207 VGND 0.2822f
C11786 Vbias.n287 VGND 0.27871f
C11787 Vbias.t109 VGND 0.2822f
C11788 Vbias.n288 VGND 0.27871f
C11789 Vbias.t249 VGND 0.2822f
C11790 Vbias.n289 VGND 0.27871f
C11791 Vbias.n290 VGND 0.07848f
C11792 Vbias.n291 VGND 0.29662f
C11793 Vbias.t86 VGND 0.2822f
C11794 Vbias.n292 VGND 0.27871f
C11795 Vbias.t170 VGND 0.2822f
C11796 Vbias.n293 VGND 0.27871f
C11797 Vbias.n294 VGND 0.30595f
C11798 Vbias.t97 VGND 0.2822f
C11799 Vbias.n295 VGND 0.27871f
C11800 Vbias.t77 VGND 0.2822f
C11801 Vbias.n296 VGND 0.27871f
C11802 Vbias.n297 VGND 0.30595f
C11803 Vbias.t148 VGND 0.2822f
C11804 Vbias.n298 VGND 0.27871f
C11805 Vbias.t252 VGND 0.2822f
C11806 Vbias.n299 VGND 0.27871f
C11807 Vbias.n300 VGND 0.30595f
C11808 Vbias.t177 VGND 0.2822f
C11809 Vbias.n301 VGND 0.27871f
C11810 Vbias.t157 VGND 0.2822f
C11811 Vbias.n302 VGND 0.27871f
C11812 Vbias.n303 VGND 0.30595f
C11813 Vbias.t228 VGND 0.2822f
C11814 Vbias.n304 VGND 0.27871f
C11815 Vbias.t143 VGND 0.2822f
C11816 Vbias.n305 VGND 0.27871f
C11817 Vbias.n306 VGND 0.30595f
C11818 Vbias.t71 VGND 0.2822f
C11819 Vbias.n307 VGND 0.27871f
C11820 Vbias.t253 VGND 0.2822f
C11821 Vbias.n308 VGND 0.27871f
C11822 Vbias.n309 VGND 0.30595f
C11823 Vbias.t70 VGND 0.2822f
C11824 Vbias.n310 VGND 0.27871f
C11825 Vbias.t42 VGND 0.2822f
C11826 Vbias.n311 VGND 0.27871f
C11827 Vbias.n312 VGND 0.30595f
C11828 Vbias.t230 VGND 0.2822f
C11829 Vbias.n313 VGND 0.27871f
C11830 Vbias.t145 VGND 0.2822f
C11831 Vbias.n314 VGND 0.27871f
C11832 Vbias.n315 VGND 0.30595f
C11833 Vbias.t218 VGND 0.2822f
C11834 Vbias.n316 VGND 0.27871f
C11835 Vbias.t131 VGND 0.2822f
C11836 Vbias.n317 VGND 0.27871f
C11837 Vbias.n318 VGND 0.30595f
C11838 Vbias.t58 VGND 0.2822f
C11839 Vbias.n319 VGND 0.27871f
C11840 Vbias.t224 VGND 0.2822f
C11841 Vbias.n320 VGND 0.27871f
C11842 Vbias.n321 VGND 0.30595f
C11843 Vbias.t38 VGND 0.2822f
C11844 Vbias.n322 VGND 0.27871f
C11845 Vbias.t214 VGND 0.2822f
C11846 Vbias.n323 VGND 0.27871f
C11847 Vbias.n324 VGND 0.30595f
C11848 Vbias.t139 VGND 0.2822f
C11849 Vbias.n325 VGND 0.27871f
C11850 Vbias.t132 VGND 0.2822f
C11851 Vbias.n326 VGND 0.27871f
C11852 Vbias.n327 VGND 0.30595f
C11853 Vbias.t203 VGND 0.2822f
C11854 Vbias.n328 VGND 0.27871f
C11855 Vbias.t30 VGND 0.2822f
C11856 Vbias.n329 VGND 0.27871f
C11857 Vbias.n330 VGND 0.07618f
C11858 Vbias.t100 VGND 0.2822f
C11859 Vbias.n331 VGND 0.27871f
C11860 Vbias.n332 VGND 0.30595f
C11861 Vbias.t31 VGND 0.2822f
C11862 Vbias.n333 VGND 0.27871f
C11863 Vbias.t215 VGND 0.2822f
C11864 Vbias.n334 VGND 0.27871f
C11865 Vbias.t140 VGND 0.2822f
C11866 Vbias.n335 VGND 0.27871f
C11867 Vbias.n336 VGND 0.07618f
C11868 Vbias.t261 VGND 0.2822f
C11869 Vbias.n337 VGND 0.27871f
C11870 Vbias.t151 VGND 0.2822f
C11871 Vbias.n338 VGND 0.27871f
C11872 Vbias.t35 VGND 0.2822f
C11873 Vbias.n339 VGND 0.27871f
C11874 Vbias.n340 VGND 0.07848f
C11875 Vbias.t104 VGND 0.2822f
C11876 Vbias.n341 VGND 0.27871f
C11877 Vbias.t260 VGND 44.3836f
C11878 Vbias.n342 VGND 1.7799f
C11879 Vbias.t216 VGND 0.2822f
C11880 Vbias.n343 VGND 0.27871f
C11881 Vbias.n344 VGND 0.07848f
C11882 Vbias.n345 VGND 0.16575f
C11883 Vbias.t59 VGND 0.2822f
C11884 Vbias.n346 VGND 0.27871f
C11885 Vbias.n347 VGND 0.07848f
C11886 Vbias.n348 VGND 0.16575f
C11887 Vbias.t67 VGND 0.2822f
C11888 Vbias.n349 VGND 0.27871f
C11889 Vbias.n350 VGND 0.07848f
C11890 Vbias.n351 VGND 0.16575f
C11891 Vbias.t152 VGND 0.2822f
C11892 Vbias.n352 VGND 0.27871f
C11893 Vbias.n353 VGND 0.07848f
C11894 Vbias.n354 VGND 0.16575f
C11895 Vbias.t245 VGND 0.2822f
C11896 Vbias.n355 VGND 0.27871f
C11897 Vbias.n356 VGND 0.07848f
C11898 Vbias.n357 VGND 0.16575f
C11899 Vbias.t72 VGND 0.2822f
C11900 Vbias.n358 VGND 0.27871f
C11901 Vbias.n359 VGND 0.07848f
C11902 Vbias.n360 VGND 0.16575f
C11903 Vbias.t158 VGND 0.2822f
C11904 Vbias.n361 VGND 0.27871f
C11905 Vbias.n362 VGND 0.07848f
C11906 Vbias.n363 VGND 0.16575f
C11907 Vbias.t178 VGND 0.2822f
C11908 Vbias.n364 VGND 0.27871f
C11909 Vbias.n365 VGND 0.07848f
C11910 Vbias.n366 VGND 0.16575f
C11911 Vbias.t254 VGND 0.2822f
C11912 Vbias.n367 VGND 0.27871f
C11913 Vbias.n368 VGND 0.07848f
C11914 Vbias.n369 VGND 0.16575f
C11915 Vbias.t84 VGND 0.2822f
C11916 Vbias.n370 VGND 0.27871f
C11917 Vbias.n371 VGND 0.07848f
C11918 Vbias.n372 VGND 0.16575f
C11919 Vbias.t106 VGND 0.2822f
C11920 Vbias.n373 VGND 0.27871f
C11921 Vbias.n374 VGND 0.07848f
C11922 Vbias.n375 VGND 0.16575f
C11923 Vbias.t259 VGND 0.2822f
C11924 Vbias.n376 VGND 0.27871f
C11925 Vbias.n377 VGND 0.07848f
C11926 Vbias.n378 VGND 0.16575f
C11927 Vbias.t26 VGND 0.2822f
C11928 Vbias.n379 VGND 0.27871f
C11929 Vbias.n380 VGND 0.07848f
C11930 Vbias.n381 VGND 0.16575f
C11931 Vbias.n382 VGND 0.16575f
C11932 Vbias.t194 VGND 0.2822f
C11933 Vbias.n383 VGND 0.27871f
C11934 Vbias.t61 VGND 0.2822f
C11935 Vbias.n384 VGND 0.27871f
C11936 Vbias.n385 VGND 0.68957f
C11937 Vbias.n386 VGND 0.16575f
C11938 Vbias.n387 VGND 0.2262f
C11939 Vbias.n388 VGND 0.30595f
C11940 Vbias.n389 VGND 0.07848f
C11941 Vbias.n390 VGND 0.16575f
C11942 Vbias.n391 VGND 0.67535f
C11943 Vbias.n392 VGND 0.16575f
C11944 Vbias.n393 VGND 0.8811f
C11945 Vbias.n394 VGND 0.8811f
C11946 Vbias.n395 VGND 0.8811f
C11947 Vbias.t13 VGND 0.2822f
C11948 Vbias.n396 VGND 0.27871f
C11949 Vbias.n397 VGND 0.07848f
C11950 Vbias.n398 VGND 0.16575f
C11951 Vbias.n399 VGND 0.16575f
C11952 Vbias.n400 VGND 0.07848f
C11953 Vbias.n401 VGND 0.29662f
C11954 Vbias.n402 VGND 0.30595f
C11955 Vbias.n403 VGND 0.2262f
C11956 Vbias.n404 VGND 0.16575f
C11957 Vbias.t142 VGND 0.2822f
C11958 Vbias.n405 VGND 0.27871f
C11959 Vbias.n406 VGND 0.2262f
C11960 Vbias.n407 VGND 0.16575f
C11961 Vbias.t114 VGND 0.2822f
C11962 Vbias.n408 VGND 0.27871f
C11963 Vbias.n409 VGND 0.2262f
C11964 Vbias.n410 VGND 0.16575f
C11965 Vbias.t223 VGND 0.2822f
C11966 Vbias.n411 VGND 0.27871f
C11967 Vbias.n412 VGND 0.2262f
C11968 Vbias.n413 VGND 0.16575f
C11969 Vbias.t202 VGND 0.2822f
C11970 Vbias.n414 VGND 0.27871f
C11971 Vbias.n415 VGND 0.2262f
C11972 Vbias.n416 VGND 0.16575f
C11973 Vbias.t111 VGND 0.2822f
C11974 Vbias.n417 VGND 0.27871f
C11975 Vbias.n418 VGND 0.2262f
C11976 Vbias.n419 VGND 0.16575f
C11977 Vbias.t39 VGND 0.2822f
C11978 Vbias.n420 VGND 0.27871f
C11979 Vbias.n421 VGND 0.2262f
C11980 Vbias.n422 VGND 0.16575f
C11981 Vbias.t19 VGND 0.2822f
C11982 Vbias.n423 VGND 0.27871f
C11983 Vbias.n424 VGND 0.2262f
C11984 Vbias.n425 VGND 0.16575f
C11985 Vbias.t184 VGND 0.2822f
C11986 Vbias.n426 VGND 0.27871f
C11987 Vbias.n427 VGND 0.2262f
C11988 Vbias.n428 VGND 0.16575f
C11989 Vbias.t101 VGND 0.2822f
C11990 Vbias.n429 VGND 0.27871f
C11991 Vbias.n430 VGND 0.2262f
C11992 Vbias.n431 VGND 0.16575f
C11993 Vbias.t15 VGND 0.2822f
C11994 Vbias.n432 VGND 0.27871f
C11995 Vbias.n433 VGND 0.2262f
C11996 Vbias.n434 VGND 0.16575f
C11997 Vbias.t182 VGND 0.2822f
C11998 Vbias.n435 VGND 0.27871f
C11999 Vbias.n436 VGND 0.2262f
C12000 Vbias.n437 VGND 0.16575f
C12001 Vbias.t174 VGND 0.2822f
C12002 Vbias.n438 VGND 0.27871f
C12003 Vbias.n439 VGND 0.2262f
C12004 Vbias.n440 VGND 0.16575f
C12005 Vbias.t79 VGND 0.2822f
C12006 Vbias.n441 VGND 0.27871f
C12007 Vbias.n442 VGND 0.2262f
C12008 Vbias.n443 VGND 0.16575f
C12009 Vbias.n444 VGND 0.2239f
C12010 Vbias.n445 VGND 0.30595f
C12011 Vbias.n446 VGND 0.29662f
C12012 Vbias.n447 VGND 0.07618f
C12013 Vbias.n448 VGND 0.16575f
C12014 Vbias.n449 VGND 0.07848f
C12015 Vbias.n450 VGND 0.29662f
C12016 Vbias.n451 VGND 0.29662f
C12017 Vbias.n452 VGND 0.07848f
C12018 Vbias.n453 VGND 0.16575f
C12019 Vbias.n454 VGND 0.16575f
C12020 Vbias.n455 VGND 0.07848f
C12021 Vbias.n456 VGND 0.29662f
C12022 Vbias.n457 VGND 0.29662f
C12023 Vbias.n458 VGND 0.07848f
C12024 Vbias.n459 VGND 0.16575f
C12025 Vbias.n460 VGND 0.16575f
C12026 Vbias.n461 VGND 0.07848f
C12027 Vbias.n462 VGND 0.29662f
C12028 Vbias.n463 VGND 0.29662f
C12029 Vbias.n464 VGND 0.07848f
C12030 Vbias.n465 VGND 0.16575f
C12031 Vbias.n466 VGND 0.16575f
C12032 Vbias.n467 VGND 0.07848f
C12033 Vbias.n468 VGND 0.29662f
C12034 Vbias.n469 VGND 0.29662f
C12035 Vbias.n470 VGND 0.07848f
C12036 Vbias.n471 VGND 0.16575f
C12037 Vbias.n472 VGND 0.16575f
C12038 Vbias.n473 VGND 0.07848f
C12039 Vbias.n474 VGND 0.29662f
C12040 Vbias.n475 VGND 0.29662f
C12041 Vbias.n476 VGND 0.07848f
C12042 Vbias.n477 VGND 0.16575f
C12043 Vbias.n478 VGND 0.16575f
C12044 Vbias.n479 VGND 0.07848f
C12045 Vbias.n480 VGND 0.29662f
C12046 Vbias.n481 VGND 0.29662f
C12047 Vbias.n482 VGND 0.07848f
C12048 Vbias.n483 VGND 0.16575f
C12049 Vbias.n484 VGND 0.16575f
C12050 Vbias.n485 VGND 0.07848f
C12051 Vbias.n486 VGND 0.29662f
C12052 Vbias.n487 VGND 0.29662f
C12053 Vbias.n488 VGND 0.07848f
C12054 Vbias.n489 VGND 0.16575f
C12055 Vbias.n490 VGND 0.16575f
C12056 Vbias.n491 VGND 0.07848f
C12057 Vbias.n492 VGND 0.29662f
C12058 Vbias.n493 VGND 0.29662f
C12059 Vbias.n494 VGND 0.07848f
C12060 Vbias.n495 VGND 0.16575f
C12061 Vbias.n496 VGND 0.16575f
C12062 Vbias.n497 VGND 0.07848f
C12063 Vbias.n498 VGND 0.29662f
C12064 Vbias.n499 VGND 0.29662f
C12065 Vbias.n500 VGND 0.07848f
C12066 Vbias.n501 VGND 0.16575f
C12067 Vbias.n502 VGND 0.16575f
C12068 Vbias.n503 VGND 0.07848f
C12069 Vbias.n504 VGND 0.29662f
C12070 Vbias.n505 VGND 0.29662f
C12071 Vbias.n506 VGND 0.07848f
C12072 Vbias.n507 VGND 0.16575f
C12073 Vbias.n508 VGND 0.16575f
C12074 Vbias.n509 VGND 0.07848f
C12075 Vbias.n510 VGND 0.29662f
C12076 Vbias.n511 VGND 0.29662f
C12077 Vbias.n512 VGND 0.07848f
C12078 Vbias.n513 VGND 0.16575f
C12079 Vbias.n514 VGND 0.16575f
C12080 Vbias.n515 VGND 0.07848f
C12081 Vbias.n516 VGND 0.29662f
C12082 Vbias.n517 VGND 0.29662f
C12083 Vbias.n518 VGND 0.07848f
C12084 Vbias.n519 VGND 0.16575f
C12085 Vbias.n520 VGND 0.16575f
C12086 Vbias.n521 VGND 0.07848f
C12087 Vbias.n522 VGND 0.29662f
C12088 Vbias.n523 VGND 0.29662f
C12089 Vbias.n524 VGND 0.07848f
C12090 Vbias.n525 VGND 0.16575f
C12091 Vbias.t175 VGND 0.2822f
C12092 Vbias.n526 VGND 0.27871f
C12093 Vbias.n527 VGND 0.07848f
C12094 Vbias.n528 VGND 0.16575f
C12095 Vbias.n529 VGND 0.16575f
C12096 Vbias.n530 VGND 0.07848f
C12097 Vbias.n531 VGND 0.29662f
C12098 Vbias.n532 VGND 0.29662f
C12099 Vbias.n533 VGND 0.29662f
C12100 Vbias.n534 VGND 0.07848f
C12101 Vbias.n535 VGND 0.16575f
C12102 Vbias.n536 VGND 0.16575f
C12103 Vbias.n537 VGND 0.07848f
C12104 Vbias.n538 VGND 0.29662f
C12105 Vbias.n539 VGND 0.29662f
C12106 Vbias.n540 VGND 0.07848f
C12107 Vbias.n541 VGND 0.16575f
C12108 Vbias.t78 VGND 0.2822f
C12109 Vbias.n542 VGND 0.27871f
C12110 Vbias.n543 VGND 0.07848f
C12111 Vbias.n544 VGND 0.16575f
C12112 Vbias.t47 VGND 0.2822f
C12113 Vbias.n545 VGND 0.27871f
C12114 Vbias.n546 VGND 0.07848f
C12115 Vbias.n547 VGND 0.16575f
C12116 Vbias.t159 VGND 0.2822f
C12117 Vbias.n548 VGND 0.27871f
C12118 Vbias.n549 VGND 0.07848f
C12119 Vbias.n550 VGND 0.16575f
C12120 Vbias.t134 VGND 0.2822f
C12121 Vbias.n551 VGND 0.27871f
C12122 Vbias.n552 VGND 0.07848f
C12123 Vbias.n553 VGND 0.16575f
C12124 Vbias.t43 VGND 0.2822f
C12125 Vbias.n554 VGND 0.27871f
C12126 Vbias.n555 VGND 0.07848f
C12127 Vbias.n556 VGND 0.16575f
C12128 Vbias.t231 VGND 0.2822f
C12129 Vbias.n557 VGND 0.27871f
C12130 Vbias.n558 VGND 0.07848f
C12131 Vbias.n559 VGND 0.16575f
C12132 Vbias.t209 VGND 0.2822f
C12133 Vbias.n560 VGND 0.27871f
C12134 Vbias.n561 VGND 0.07848f
C12135 Vbias.n562 VGND 0.16575f
C12136 Vbias.t116 VGND 0.2822f
C12137 Vbias.n563 VGND 0.27871f
C12138 Vbias.n564 VGND 0.07848f
C12139 Vbias.n565 VGND 0.16575f
C12140 Vbias.t34 VGND 0.2822f
C12141 Vbias.n566 VGND 0.27871f
C12142 Vbias.n567 VGND 0.07848f
C12143 Vbias.n568 VGND 0.16575f
C12144 Vbias.t206 VGND 0.2822f
C12145 Vbias.n569 VGND 0.27871f
C12146 Vbias.n570 VGND 0.07848f
C12147 Vbias.n571 VGND 0.16575f
C12148 Vbias.t115 VGND 0.2822f
C12149 Vbias.n572 VGND 0.27871f
C12150 Vbias.n573 VGND 0.07848f
C12151 Vbias.n574 VGND 0.16575f
C12152 Vbias.t103 VGND 0.2822f
C12153 Vbias.n575 VGND 0.27871f
C12154 Vbias.n576 VGND 0.07848f
C12155 Vbias.n577 VGND 0.16575f
C12156 Vbias.t6 VGND 0.2822f
C12157 Vbias.n578 VGND 0.27871f
C12158 Vbias.n579 VGND 0.07848f
C12159 Vbias.n580 VGND 0.16575f
C12160 Vbias.n581 VGND 0.07618f
C12161 Vbias.n582 VGND 0.29662f
C12162 Vbias.n583 VGND 0.29662f
C12163 Vbias.n584 VGND 0.07618f
C12164 Vbias.n585 VGND 0.16575f
C12165 Vbias.n586 VGND 0.07848f
C12166 Vbias.n587 VGND 0.29662f
C12167 Vbias.n588 VGND 0.29662f
C12168 Vbias.n589 VGND 0.07848f
C12169 Vbias.n590 VGND 0.16575f
C12170 Vbias.n591 VGND 0.16575f
C12171 Vbias.n592 VGND 0.07848f
C12172 Vbias.n593 VGND 0.29662f
C12173 Vbias.n594 VGND 0.29662f
C12174 Vbias.n595 VGND 0.07848f
C12175 Vbias.n596 VGND 0.16575f
C12176 Vbias.n597 VGND 0.16575f
C12177 Vbias.n598 VGND 0.07848f
C12178 Vbias.n599 VGND 0.29662f
C12179 Vbias.n600 VGND 0.29662f
C12180 Vbias.n601 VGND 0.07848f
C12181 Vbias.n602 VGND 0.16575f
C12182 Vbias.n603 VGND 0.16575f
C12183 Vbias.n604 VGND 0.07848f
C12184 Vbias.n605 VGND 0.29662f
C12185 Vbias.n606 VGND 0.29662f
C12186 Vbias.n607 VGND 0.07848f
C12187 Vbias.n608 VGND 0.16575f
C12188 Vbias.n609 VGND 0.16575f
C12189 Vbias.n610 VGND 0.07848f
C12190 Vbias.n611 VGND 0.29662f
C12191 Vbias.n612 VGND 0.29662f
C12192 Vbias.n613 VGND 0.07848f
C12193 Vbias.n614 VGND 0.16575f
C12194 Vbias.n615 VGND 0.16575f
C12195 Vbias.n616 VGND 0.07848f
C12196 Vbias.n617 VGND 0.29662f
C12197 Vbias.n618 VGND 0.29662f
C12198 Vbias.n619 VGND 0.07848f
C12199 Vbias.n620 VGND 0.16575f
C12200 Vbias.n621 VGND 0.16575f
C12201 Vbias.n622 VGND 0.07848f
C12202 Vbias.n623 VGND 0.29662f
C12203 Vbias.n624 VGND 0.29662f
C12204 Vbias.n625 VGND 0.07848f
C12205 Vbias.n626 VGND 0.16575f
C12206 Vbias.n627 VGND 0.16575f
C12207 Vbias.n628 VGND 0.07848f
C12208 Vbias.n629 VGND 0.29662f
C12209 Vbias.n630 VGND 0.29662f
C12210 Vbias.n631 VGND 0.07848f
C12211 Vbias.n632 VGND 0.16575f
C12212 Vbias.n633 VGND 0.16575f
C12213 Vbias.n634 VGND 0.07848f
C12214 Vbias.n635 VGND 0.29662f
C12215 Vbias.n636 VGND 0.29662f
C12216 Vbias.n637 VGND 0.07848f
C12217 Vbias.n638 VGND 0.16575f
C12218 Vbias.n639 VGND 0.16575f
C12219 Vbias.n640 VGND 0.07848f
C12220 Vbias.n641 VGND 0.29662f
C12221 Vbias.n642 VGND 0.29662f
C12222 Vbias.n643 VGND 0.07848f
C12223 Vbias.n644 VGND 0.16575f
C12224 Vbias.n645 VGND 0.16575f
C12225 Vbias.n646 VGND 0.07848f
C12226 Vbias.n647 VGND 0.29662f
C12227 Vbias.n648 VGND 0.29662f
C12228 Vbias.n649 VGND 0.07848f
C12229 Vbias.n650 VGND 0.16575f
C12230 Vbias.n651 VGND 0.16575f
C12231 Vbias.n652 VGND 0.07848f
C12232 Vbias.n653 VGND 0.29662f
C12233 Vbias.n654 VGND 0.29662f
C12234 Vbias.n655 VGND 0.07848f
C12235 Vbias.n656 VGND 0.16575f
C12236 Vbias.n657 VGND 0.16575f
C12237 Vbias.n658 VGND 0.07848f
C12238 Vbias.n659 VGND 0.29662f
C12239 Vbias.n660 VGND 0.29662f
C12240 Vbias.n661 VGND 0.07848f
C12241 Vbias.n662 VGND 0.16575f
C12242 Vbias.t89 VGND 0.2822f
C12243 Vbias.n663 VGND 0.27871f
C12244 Vbias.n664 VGND 0.07848f
C12245 Vbias.n665 VGND 0.16575f
C12246 Vbias.t250 VGND 0.2822f
C12247 Vbias.n666 VGND 0.27871f
C12248 Vbias.n667 VGND 0.07848f
C12249 Vbias.n668 VGND 0.16575f
C12250 Vbias.n669 VGND 0.8811f
C12251 Vbias.n670 VGND 0.8811f
C12252 Vbias.n671 VGND 0.8811f
C12253 Vbias.t165 VGND 0.2822f
C12254 Vbias.n672 VGND 0.27871f
C12255 Vbias.n673 VGND 0.07848f
C12256 Vbias.n674 VGND 0.16575f
C12257 Vbias.t73 VGND 0.2822f
C12258 Vbias.n675 VGND 0.27871f
C12259 Vbias.n676 VGND 0.07848f
C12260 Vbias.n677 VGND 0.16575f
C12261 Vbias.n678 VGND 0.8811f
C12262 Vbias.t255 VGND 0.2822f
C12263 Vbias.n679 VGND 0.27871f
C12264 Vbias.n680 VGND 0.29662f
C12265 Vbias.n681 VGND 0.07848f
C12266 Vbias.n682 VGND 0.16575f
C12267 Vbias.n683 VGND 0.8811f
C12268 Vbias.t176 VGND 0.2822f
C12269 Vbias.n684 VGND 0.27871f
C12270 Vbias.n685 VGND 0.07848f
C12271 Vbias.n686 VGND 0.16575f
C12272 Vbias.n687 VGND 0.8811f
C12273 Vbias.n688 VGND 0.8811f
C12274 Vbias.n689 VGND 0.8811f
C12275 Vbias.n690 VGND 0.16575f
C12276 Vbias.n691 VGND 0.16575f
C12277 Vbias.n692 VGND 0.07848f
C12278 Vbias.n693 VGND 0.29662f
C12279 Vbias.n694 VGND 0.29662f
C12280 Vbias.n695 VGND 0.07848f
C12281 Vbias.n696 VGND 0.16575f
C12282 Vbias.n697 VGND 0.16575f
C12283 Vbias.n698 VGND 0.07848f
C12284 Vbias.n699 VGND 0.29662f
C12285 Vbias.n700 VGND 0.29662f
C12286 Vbias.n701 VGND 0.29662f
C12287 Vbias.n702 VGND 0.07848f
C12288 Vbias.n703 VGND 0.16575f
C12289 Vbias.t204 VGND 0.2822f
C12290 Vbias.n704 VGND 0.27871f
C12291 Vbias.n705 VGND 0.07848f
C12292 Vbias.n706 VGND 0.16575f
C12293 Vbias.n707 VGND 0.16575f
C12294 Vbias.n708 VGND 0.07848f
C12295 Vbias.n709 VGND 0.29662f
C12296 Vbias.n710 VGND 0.29662f
C12297 Vbias.n711 VGND 0.07848f
C12298 Vbias.n712 VGND 0.16575f
C12299 Vbias.n713 VGND 0.16575f
C12300 Vbias.n714 VGND 0.07848f
C12301 Vbias.n715 VGND 0.29662f
C12302 Vbias.n716 VGND 0.29662f
C12303 Vbias.n717 VGND 0.07848f
C12304 Vbias.n718 VGND 0.16575f
C12305 Vbias.n719 VGND 0.16575f
C12306 Vbias.n720 VGND 0.07848f
C12307 Vbias.n721 VGND 0.29662f
C12308 Vbias.n722 VGND 0.29662f
C12309 Vbias.n723 VGND 0.07848f
C12310 Vbias.n724 VGND 0.16575f
C12311 Vbias.n725 VGND 0.16575f
C12312 Vbias.n726 VGND 0.07848f
C12313 Vbias.n727 VGND 0.29662f
C12314 Vbias.n728 VGND 0.29662f
C12315 Vbias.n729 VGND 0.07848f
C12316 Vbias.n730 VGND 0.16575f
C12317 Vbias.n731 VGND 0.16575f
C12318 Vbias.n732 VGND 0.07848f
C12319 Vbias.n733 VGND 0.29662f
C12320 Vbias.n734 VGND 0.29662f
C12321 Vbias.n735 VGND 0.07848f
C12322 Vbias.n736 VGND 0.16575f
C12323 Vbias.n737 VGND 0.16575f
C12324 Vbias.n738 VGND 0.07848f
C12325 Vbias.n739 VGND 0.29662f
C12326 Vbias.n740 VGND 0.29662f
C12327 Vbias.n741 VGND 0.07848f
C12328 Vbias.n742 VGND 0.16575f
C12329 Vbias.n743 VGND 0.16575f
C12330 Vbias.n744 VGND 0.07848f
C12331 Vbias.n745 VGND 0.29662f
C12332 Vbias.n746 VGND 0.29662f
C12333 Vbias.n747 VGND 0.07848f
C12334 Vbias.n748 VGND 0.16575f
C12335 Vbias.n749 VGND 0.16575f
C12336 Vbias.n750 VGND 0.07848f
C12337 Vbias.n751 VGND 0.29662f
C12338 Vbias.n752 VGND 0.29662f
C12339 Vbias.n753 VGND 0.07848f
C12340 Vbias.n754 VGND 0.16575f
C12341 Vbias.n755 VGND 0.16575f
C12342 Vbias.n756 VGND 0.07848f
C12343 Vbias.n757 VGND 0.29662f
C12344 Vbias.n758 VGND 0.29662f
C12345 Vbias.n759 VGND 0.07848f
C12346 Vbias.n760 VGND 0.16575f
C12347 Vbias.n761 VGND 0.16575f
C12348 Vbias.n762 VGND 0.07848f
C12349 Vbias.n763 VGND 0.29662f
C12350 Vbias.n764 VGND 0.29662f
C12351 Vbias.n765 VGND 0.07848f
C12352 Vbias.n766 VGND 0.16575f
C12353 Vbias.n767 VGND 0.16575f
C12354 Vbias.n768 VGND 0.07848f
C12355 Vbias.n769 VGND 0.29662f
C12356 Vbias.n770 VGND 0.29662f
C12357 Vbias.n771 VGND 0.07848f
C12358 Vbias.n772 VGND 0.16575f
C12359 Vbias.n773 VGND 0.16575f
C12360 Vbias.n774 VGND 0.07848f
C12361 Vbias.n775 VGND 0.29662f
C12362 Vbias.n776 VGND 0.29662f
C12363 Vbias.n777 VGND 0.07848f
C12364 Vbias.n778 VGND 0.16575f
C12365 Vbias.n779 VGND 0.16575f
C12366 Vbias.n780 VGND 0.07848f
C12367 Vbias.n781 VGND 0.29662f
C12368 Vbias.n782 VGND 0.29662f
C12369 Vbias.n783 VGND 0.07848f
C12370 Vbias.n784 VGND 0.16575f
C12371 Vbias.n785 VGND 0.07618f
C12372 Vbias.n786 VGND 0.29662f
C12373 Vbias.n787 VGND 0.29662f
C12374 Vbias.n788 VGND 0.29662f
C12375 Vbias.n789 VGND 0.07618f
C12376 Vbias.t195 VGND 0.2822f
C12377 Vbias.n790 VGND 0.27871f
C12378 Vbias.n791 VGND 0.07848f
C12379 Vbias.n792 VGND 0.16575f
C12380 Vbias.t37 VGND 0.2822f
C12381 Vbias.n793 VGND 0.27871f
C12382 Vbias.n794 VGND 0.07848f
C12383 Vbias.n795 VGND 0.16575f
C12384 Vbias.t48 VGND 0.2822f
C12385 Vbias.n796 VGND 0.27871f
C12386 Vbias.n797 VGND 0.07848f
C12387 Vbias.n798 VGND 0.16575f
C12388 Vbias.t135 VGND 0.2822f
C12389 Vbias.n799 VGND 0.27871f
C12390 Vbias.n800 VGND 0.07848f
C12391 Vbias.n801 VGND 0.16575f
C12392 Vbias.t221 VGND 0.2822f
C12393 Vbias.n802 VGND 0.27871f
C12394 Vbias.n803 VGND 0.07848f
C12395 Vbias.n804 VGND 0.16575f
C12396 Vbias.t50 VGND 0.2822f
C12397 Vbias.n805 VGND 0.27871f
C12398 Vbias.n806 VGND 0.07848f
C12399 Vbias.n807 VGND 0.16575f
C12400 Vbias.t138 VGND 0.2822f
C12401 Vbias.n808 VGND 0.27871f
C12402 Vbias.n809 VGND 0.07848f
C12403 Vbias.n810 VGND 0.16575f
C12404 Vbias.t163 VGND 0.2822f
C12405 Vbias.n811 VGND 0.27871f
C12406 Vbias.n812 VGND 0.07848f
C12407 Vbias.n813 VGND 0.16575f
C12408 Vbias.t236 VGND 0.2822f
C12409 Vbias.n814 VGND 0.27871f
C12410 Vbias.n815 VGND 0.07848f
C12411 Vbias.n816 VGND 0.16575f
C12412 Vbias.t65 VGND 0.2822f
C12413 Vbias.n817 VGND 0.27871f
C12414 Vbias.n818 VGND 0.07848f
C12415 Vbias.n819 VGND 0.16575f
C12416 Vbias.t90 VGND 0.2822f
C12417 Vbias.n820 VGND 0.27871f
C12418 Vbias.n821 VGND 0.07848f
C12419 Vbias.n822 VGND 0.16575f
C12420 Vbias.t243 VGND 0.2822f
C12421 Vbias.n823 VGND 0.27871f
C12422 Vbias.n824 VGND 0.07848f
C12423 Vbias.n825 VGND 0.16575f
C12424 Vbias.t7 VGND 0.2822f
C12425 Vbias.n826 VGND 0.27871f
C12426 Vbias.n827 VGND 0.07848f
C12427 Vbias.n828 VGND 0.16575f
C12428 Vbias.n829 VGND 0.16575f
C12429 Vbias.n830 VGND 0.07848f
C12430 Vbias.n831 VGND 0.29662f
C12431 Vbias.n832 VGND 0.29662f
C12432 Vbias.n833 VGND 0.07848f
C12433 Vbias.n834 VGND 0.16575f
C12434 Vbias.n835 VGND 0.16575f
C12435 Vbias.n836 VGND 0.07848f
C12436 Vbias.n837 VGND 0.29662f
C12437 Vbias.n838 VGND 0.29662f
C12438 Vbias.n839 VGND 0.07848f
C12439 Vbias.n840 VGND 0.16575f
C12440 Vbias.n841 VGND 0.16575f
C12441 Vbias.n842 VGND 0.07848f
C12442 Vbias.n843 VGND 0.29662f
C12443 Vbias.n844 VGND 0.29662f
C12444 Vbias.n845 VGND 0.07848f
C12445 Vbias.n846 VGND 0.16575f
C12446 Vbias.n847 VGND 0.16575f
C12447 Vbias.n848 VGND 0.07848f
C12448 Vbias.n849 VGND 0.29662f
C12449 Vbias.n850 VGND 0.29662f
C12450 Vbias.n851 VGND 0.07848f
C12451 Vbias.n852 VGND 0.16575f
C12452 Vbias.n853 VGND 0.16575f
C12453 Vbias.n854 VGND 0.07848f
C12454 Vbias.n855 VGND 0.29662f
C12455 Vbias.n856 VGND 0.29662f
C12456 Vbias.n857 VGND 0.07848f
C12457 Vbias.n858 VGND 0.16575f
C12458 Vbias.n859 VGND 0.16575f
C12459 Vbias.n860 VGND 0.07848f
C12460 Vbias.n861 VGND 0.29662f
C12461 Vbias.n862 VGND 0.29662f
C12462 Vbias.n863 VGND 0.07848f
C12463 Vbias.n864 VGND 0.16575f
C12464 Vbias.n865 VGND 0.16575f
C12465 Vbias.n866 VGND 0.07848f
C12466 Vbias.n867 VGND 0.29662f
C12467 Vbias.n868 VGND 0.29662f
C12468 Vbias.n869 VGND 0.07848f
C12469 Vbias.n870 VGND 0.16575f
C12470 Vbias.n871 VGND 0.16575f
C12471 Vbias.n872 VGND 0.07848f
C12472 Vbias.n873 VGND 0.29662f
C12473 Vbias.n874 VGND 0.29662f
C12474 Vbias.n875 VGND 0.07848f
C12475 Vbias.n876 VGND 0.16575f
C12476 Vbias.n877 VGND 0.16575f
C12477 Vbias.n878 VGND 0.07848f
C12478 Vbias.n879 VGND 0.29662f
C12479 Vbias.n880 VGND 0.29662f
C12480 Vbias.n881 VGND 0.07848f
C12481 Vbias.n882 VGND 0.16575f
C12482 Vbias.n883 VGND 0.16575f
C12483 Vbias.n884 VGND 0.07848f
C12484 Vbias.n885 VGND 0.29662f
C12485 Vbias.n886 VGND 0.29662f
C12486 Vbias.n887 VGND 0.07848f
C12487 Vbias.n888 VGND 0.16575f
C12488 Vbias.n889 VGND 0.16575f
C12489 Vbias.n890 VGND 0.07848f
C12490 Vbias.n891 VGND 0.29662f
C12491 Vbias.n892 VGND 0.29662f
C12492 Vbias.n893 VGND 0.07848f
C12493 Vbias.n894 VGND 0.16575f
C12494 Vbias.n895 VGND 0.16575f
C12495 Vbias.n896 VGND 0.07848f
C12496 Vbias.n897 VGND 0.29662f
C12497 Vbias.n898 VGND 0.29662f
C12498 Vbias.n899 VGND 0.07848f
C12499 Vbias.n900 VGND 0.16575f
C12500 Vbias.n901 VGND 0.16575f
C12501 Vbias.n902 VGND 0.07848f
C12502 Vbias.n903 VGND 0.29662f
C12503 Vbias.n904 VGND 0.29662f
C12504 Vbias.n905 VGND 0.07848f
C12505 Vbias.n906 VGND 0.16575f
C12506 Vbias.t198 VGND 0.2822f
C12507 Vbias.n907 VGND 0.27871f
C12508 Vbias.n908 VGND 0.07618f
C12509 Vbias.n909 VGND 0.16575f
C12510 Vbias.n910 VGND 0.07848f
C12511 Vbias.n911 VGND 0.29662f
C12512 Vbias.n912 VGND 0.29662f
C12513 Vbias.n913 VGND 0.07848f
C12514 Vbias.n914 VGND 0.16575f
C12515 Vbias.n915 VGND 0.07618f
C12516 Vbias.n916 VGND 0.29662f
C12517 Vbias.n917 VGND 0.29662f
C12518 Vbias.n918 VGND 0.29418f
C12519 Vbias.n919 VGND 0.07618f
C12520 Vbias.n920 VGND 0.16575f
C12521 Vbias.n921 VGND 0.07848f
C12522 Vbias.n922 VGND 0.29418f
C12523 Vbias.n923 VGND 0.03974f
C12524 Vbias.n924 VGND 0.16575f
C12525 Vbias.n925 VGND 0.16575f
C12526 Vbias.n926 VGND 0.03974f
C12527 Vbias.n927 VGND 0.29418f
C12528 Vbias.n928 VGND 0.07848f
C12529 Vbias.n929 VGND 0.16575f
C12530 Vbias.n930 VGND 0.16575f
C12531 Vbias.n931 VGND 0.07848f
C12532 Vbias.n932 VGND 0.29418f
C12533 Vbias.n933 VGND 0.03974f
C12534 Vbias.n934 VGND 0.16575f
C12535 Vbias.n935 VGND 0.16575f
C12536 Vbias.n936 VGND 0.03974f
C12537 Vbias.n937 VGND 0.29418f
C12538 Vbias.n938 VGND 0.07848f
C12539 Vbias.n939 VGND 0.16575f
C12540 Vbias.n940 VGND 0.16575f
C12541 Vbias.n941 VGND 0.07848f
C12542 Vbias.n942 VGND 0.29418f
C12543 Vbias.n943 VGND 0.03974f
C12544 Vbias.n944 VGND 0.16575f
C12545 Vbias.n945 VGND 0.16575f
C12546 Vbias.n946 VGND 0.03974f
C12547 Vbias.n947 VGND 0.29418f
C12548 Vbias.n948 VGND 0.07848f
C12549 Vbias.n949 VGND 0.16575f
C12550 Vbias.n950 VGND 0.16575f
C12551 Vbias.n951 VGND 0.07848f
C12552 Vbias.n952 VGND 0.29418f
C12553 Vbias.n953 VGND 0.03974f
C12554 Vbias.n954 VGND 0.16575f
C12555 Vbias.n955 VGND 0.16575f
C12556 Vbias.n956 VGND 0.03974f
C12557 Vbias.n957 VGND 0.29418f
C12558 Vbias.n958 VGND 0.07848f
C12559 Vbias.n959 VGND 0.16575f
C12560 Vbias.n960 VGND 0.16575f
C12561 Vbias.n961 VGND 0.07848f
C12562 Vbias.n962 VGND 0.29418f
C12563 Vbias.n963 VGND 0.03974f
C12564 Vbias.n964 VGND 0.16575f
C12565 Vbias.n965 VGND 0.16575f
C12566 Vbias.n966 VGND 0.03974f
C12567 Vbias.n967 VGND 0.29418f
C12568 Vbias.n968 VGND 0.07848f
C12569 Vbias.n969 VGND 0.16575f
C12570 Vbias.n970 VGND 0.16575f
C12571 Vbias.n971 VGND 0.07848f
C12572 Vbias.n972 VGND 0.29418f
C12573 Vbias.n973 VGND 0.03974f
C12574 Vbias.n974 VGND 0.16575f
C12575 Vbias.n975 VGND 0.16575f
C12576 Vbias.n976 VGND 0.03974f
C12577 Vbias.n977 VGND 0.29418f
C12578 Vbias.n978 VGND 0.07848f
C12579 Vbias.n979 VGND 0.16575f
C12580 Vbias.n980 VGND 0.16575f
C12581 Vbias.n981 VGND 0.07848f
C12582 Vbias.n982 VGND 0.29418f
C12583 Vbias.n983 VGND 0.03974f
C12584 Vbias.n984 VGND 0.16575f
C12585 Vbias.n985 VGND 0.16575f
C12586 Vbias.n986 VGND 0.03974f
C12587 Vbias.n987 VGND 0.29418f
C12588 Vbias.n988 VGND 0.29662f
C12589 Vbias.n989 VGND 0.07848f
C12590 Vbias.n990 VGND 0.16575f
C12591 Vbias.n991 VGND 0.16575f
C12592 Vbias.n992 VGND 0.07848f
C12593 Vbias.n993 VGND 0.29662f
C12594 Vbias.n994 VGND 0.29418f
C12595 Vbias.n995 VGND 0.03974f
C12596 Vbias.n996 VGND 0.16575f
C12597 Vbias.n997 VGND 0.80999f
C12598 Vbias.n998 VGND 1.83432f
C12599 XThC.Tn[2].t7 VGND 0.018f
C12600 XThC.Tn[2].t6 VGND 0.018f
C12601 XThC.Tn[2].n0 VGND 0.03633f
C12602 XThC.Tn[2].t5 VGND 0.018f
C12603 XThC.Tn[2].t4 VGND 0.018f
C12604 XThC.Tn[2].n1 VGND 0.04251f
C12605 XThC.Tn[2].n2 VGND 0.119f
C12606 XThC.Tn[2].t11 VGND 0.0117f
C12607 XThC.Tn[2].t10 VGND 0.0117f
C12608 XThC.Tn[2].n3 VGND 0.02664f
C12609 XThC.Tn[2].t9 VGND 0.0117f
C12610 XThC.Tn[2].t8 VGND 0.0117f
C12611 XThC.Tn[2].n4 VGND 0.02664f
C12612 XThC.Tn[2].t1 VGND 0.0117f
C12613 XThC.Tn[2].t2 VGND 0.0117f
C12614 XThC.Tn[2].n5 VGND 0.02664f
C12615 XThC.Tn[2].t0 VGND 0.0117f
C12616 XThC.Tn[2].t3 VGND 0.0117f
C12617 XThC.Tn[2].n6 VGND 0.04439f
C12618 XThC.Tn[2].n7 VGND 0.12687f
C12619 XThC.Tn[2].n8 VGND 0.07843f
C12620 XThC.Tn[2].n9 VGND 0.08852f
C12621 XThC.Tn[2].t20 VGND 0.01427f
C12622 XThC.Tn[2].t18 VGND 0.01558f
C12623 XThC.Tn[2].n10 VGND 0.03478f
C12624 XThC.Tn[2].n11 VGND 0.02383f
C12625 XThC.Tn[2].n12 VGND 0.07822f
C12626 XThC.Tn[2].t38 VGND 0.01427f
C12627 XThC.Tn[2].t35 VGND 0.01558f
C12628 XThC.Tn[2].n13 VGND 0.03478f
C12629 XThC.Tn[2].n14 VGND 0.02383f
C12630 XThC.Tn[2].n15 VGND 0.07844f
C12631 XThC.Tn[2].n16 VGND 0.12927f
C12632 XThC.Tn[2].t43 VGND 0.01427f
C12633 XThC.Tn[2].t37 VGND 0.01558f
C12634 XThC.Tn[2].n17 VGND 0.03478f
C12635 XThC.Tn[2].n18 VGND 0.02383f
C12636 XThC.Tn[2].n19 VGND 0.07844f
C12637 XThC.Tn[2].n20 VGND 0.12927f
C12638 XThC.Tn[2].t12 VGND 0.01427f
C12639 XThC.Tn[2].t39 VGND 0.01558f
C12640 XThC.Tn[2].n21 VGND 0.03478f
C12641 XThC.Tn[2].n22 VGND 0.02383f
C12642 XThC.Tn[2].n23 VGND 0.07844f
C12643 XThC.Tn[2].n24 VGND 0.12927f
C12644 XThC.Tn[2].t31 VGND 0.01427f
C12645 XThC.Tn[2].t28 VGND 0.01558f
C12646 XThC.Tn[2].n25 VGND 0.03478f
C12647 XThC.Tn[2].n26 VGND 0.02383f
C12648 XThC.Tn[2].n27 VGND 0.07844f
C12649 XThC.Tn[2].n28 VGND 0.12927f
C12650 XThC.Tn[2].t32 VGND 0.01427f
C12651 XThC.Tn[2].t29 VGND 0.01558f
C12652 XThC.Tn[2].n29 VGND 0.03478f
C12653 XThC.Tn[2].n30 VGND 0.02383f
C12654 XThC.Tn[2].n31 VGND 0.07844f
C12655 XThC.Tn[2].n32 VGND 0.12927f
C12656 XThC.Tn[2].t16 VGND 0.01427f
C12657 XThC.Tn[2].t42 VGND 0.01558f
C12658 XThC.Tn[2].n33 VGND 0.03478f
C12659 XThC.Tn[2].n34 VGND 0.02383f
C12660 XThC.Tn[2].n35 VGND 0.07844f
C12661 XThC.Tn[2].n36 VGND 0.12927f
C12662 XThC.Tn[2].t23 VGND 0.01427f
C12663 XThC.Tn[2].t19 VGND 0.01558f
C12664 XThC.Tn[2].n37 VGND 0.03478f
C12665 XThC.Tn[2].n38 VGND 0.02383f
C12666 XThC.Tn[2].n39 VGND 0.07844f
C12667 XThC.Tn[2].n40 VGND 0.12927f
C12668 XThC.Tn[2].t25 VGND 0.01427f
C12669 XThC.Tn[2].t21 VGND 0.01558f
C12670 XThC.Tn[2].n41 VGND 0.03478f
C12671 XThC.Tn[2].n42 VGND 0.02383f
C12672 XThC.Tn[2].n43 VGND 0.07844f
C12673 XThC.Tn[2].n44 VGND 0.12927f
C12674 XThC.Tn[2].t13 VGND 0.01427f
C12675 XThC.Tn[2].t40 VGND 0.01558f
C12676 XThC.Tn[2].n45 VGND 0.03478f
C12677 XThC.Tn[2].n46 VGND 0.02383f
C12678 XThC.Tn[2].n47 VGND 0.07844f
C12679 XThC.Tn[2].n48 VGND 0.12927f
C12680 XThC.Tn[2].t15 VGND 0.01427f
C12681 XThC.Tn[2].t41 VGND 0.01558f
C12682 XThC.Tn[2].n49 VGND 0.03478f
C12683 XThC.Tn[2].n50 VGND 0.02383f
C12684 XThC.Tn[2].n51 VGND 0.07844f
C12685 XThC.Tn[2].n52 VGND 0.12927f
C12686 XThC.Tn[2].t26 VGND 0.01427f
C12687 XThC.Tn[2].t22 VGND 0.01558f
C12688 XThC.Tn[2].n53 VGND 0.03478f
C12689 XThC.Tn[2].n54 VGND 0.02383f
C12690 XThC.Tn[2].n55 VGND 0.07844f
C12691 XThC.Tn[2].n56 VGND 0.12927f
C12692 XThC.Tn[2].t34 VGND 0.01427f
C12693 XThC.Tn[2].t30 VGND 0.01558f
C12694 XThC.Tn[2].n57 VGND 0.03478f
C12695 XThC.Tn[2].n58 VGND 0.02383f
C12696 XThC.Tn[2].n59 VGND 0.07844f
C12697 XThC.Tn[2].n60 VGND 0.12927f
C12698 XThC.Tn[2].t36 VGND 0.01427f
C12699 XThC.Tn[2].t33 VGND 0.01558f
C12700 XThC.Tn[2].n61 VGND 0.03478f
C12701 XThC.Tn[2].n62 VGND 0.02383f
C12702 XThC.Tn[2].n63 VGND 0.07844f
C12703 XThC.Tn[2].n64 VGND 0.12927f
C12704 XThC.Tn[2].t17 VGND 0.01427f
C12705 XThC.Tn[2].t14 VGND 0.01558f
C12706 XThC.Tn[2].n65 VGND 0.03478f
C12707 XThC.Tn[2].n66 VGND 0.02383f
C12708 XThC.Tn[2].n67 VGND 0.07844f
C12709 XThC.Tn[2].n68 VGND 0.12927f
C12710 XThC.Tn[2].t27 VGND 0.01427f
C12711 XThC.Tn[2].t24 VGND 0.01558f
C12712 XThC.Tn[2].n69 VGND 0.03478f
C12713 XThC.Tn[2].n70 VGND 0.02383f
C12714 XThC.Tn[2].n71 VGND 0.07844f
C12715 XThC.Tn[2].n72 VGND 0.12927f
C12716 XThC.Tn[2].n73 VGND 0.50031f
C12717 XThC.Tn[2].n74 VGND 0.1061f
C12718 XThC.Tn[2].n75 VGND 0.03766f
C12719 XThC.Tn[4].t8 VGND 0.01183f
C12720 XThC.Tn[4].t11 VGND 0.01183f
C12721 XThC.Tn[4].n0 VGND 0.0449f
C12722 XThC.Tn[4].t10 VGND 0.01183f
C12723 XThC.Tn[4].t9 VGND 0.01183f
C12724 XThC.Tn[4].n1 VGND 0.02695f
C12725 XThC.Tn[4].n2 VGND 0.12834f
C12726 XThC.Tn[4].t7 VGND 0.01183f
C12727 XThC.Tn[4].t6 VGND 0.01183f
C12728 XThC.Tn[4].n3 VGND 0.02695f
C12729 XThC.Tn[4].n4 VGND 0.07934f
C12730 XThC.Tn[4].t5 VGND 0.01183f
C12731 XThC.Tn[4].t4 VGND 0.01183f
C12732 XThC.Tn[4].n5 VGND 0.02695f
C12733 XThC.Tn[4].n6 VGND 0.08954f
C12734 XThC.Tn[4].t28 VGND 0.01443f
C12735 XThC.Tn[4].t26 VGND 0.01576f
C12736 XThC.Tn[4].n7 VGND 0.03519f
C12737 XThC.Tn[4].n8 VGND 0.02411f
C12738 XThC.Tn[4].n9 VGND 0.07913f
C12739 XThC.Tn[4].t14 VGND 0.01443f
C12740 XThC.Tn[4].t43 VGND 0.01576f
C12741 XThC.Tn[4].n10 VGND 0.03519f
C12742 XThC.Tn[4].n11 VGND 0.02411f
C12743 XThC.Tn[4].n12 VGND 0.07935f
C12744 XThC.Tn[4].n13 VGND 0.13077f
C12745 XThC.Tn[4].t19 VGND 0.01443f
C12746 XThC.Tn[4].t13 VGND 0.01576f
C12747 XThC.Tn[4].n14 VGND 0.03519f
C12748 XThC.Tn[4].n15 VGND 0.02411f
C12749 XThC.Tn[4].n16 VGND 0.07935f
C12750 XThC.Tn[4].n17 VGND 0.13077f
C12751 XThC.Tn[4].t20 VGND 0.01443f
C12752 XThC.Tn[4].t15 VGND 0.01576f
C12753 XThC.Tn[4].n18 VGND 0.03519f
C12754 XThC.Tn[4].n19 VGND 0.02411f
C12755 XThC.Tn[4].n20 VGND 0.07935f
C12756 XThC.Tn[4].n21 VGND 0.13077f
C12757 XThC.Tn[4].t39 VGND 0.01443f
C12758 XThC.Tn[4].t36 VGND 0.01576f
C12759 XThC.Tn[4].n22 VGND 0.03519f
C12760 XThC.Tn[4].n23 VGND 0.02411f
C12761 XThC.Tn[4].n24 VGND 0.07935f
C12762 XThC.Tn[4].n25 VGND 0.13077f
C12763 XThC.Tn[4].t40 VGND 0.01443f
C12764 XThC.Tn[4].t37 VGND 0.01576f
C12765 XThC.Tn[4].n26 VGND 0.03519f
C12766 XThC.Tn[4].n27 VGND 0.02411f
C12767 XThC.Tn[4].n28 VGND 0.07935f
C12768 XThC.Tn[4].n29 VGND 0.13077f
C12769 XThC.Tn[4].t24 VGND 0.01443f
C12770 XThC.Tn[4].t18 VGND 0.01576f
C12771 XThC.Tn[4].n30 VGND 0.03519f
C12772 XThC.Tn[4].n31 VGND 0.02411f
C12773 XThC.Tn[4].n32 VGND 0.07935f
C12774 XThC.Tn[4].n33 VGND 0.13077f
C12775 XThC.Tn[4].t31 VGND 0.01443f
C12776 XThC.Tn[4].t27 VGND 0.01576f
C12777 XThC.Tn[4].n34 VGND 0.03519f
C12778 XThC.Tn[4].n35 VGND 0.02411f
C12779 XThC.Tn[4].n36 VGND 0.07935f
C12780 XThC.Tn[4].n37 VGND 0.13077f
C12781 XThC.Tn[4].t33 VGND 0.01443f
C12782 XThC.Tn[4].t29 VGND 0.01576f
C12783 XThC.Tn[4].n38 VGND 0.03519f
C12784 XThC.Tn[4].n39 VGND 0.02411f
C12785 XThC.Tn[4].n40 VGND 0.07935f
C12786 XThC.Tn[4].n41 VGND 0.13077f
C12787 XThC.Tn[4].t21 VGND 0.01443f
C12788 XThC.Tn[4].t16 VGND 0.01576f
C12789 XThC.Tn[4].n42 VGND 0.03519f
C12790 XThC.Tn[4].n43 VGND 0.02411f
C12791 XThC.Tn[4].n44 VGND 0.07935f
C12792 XThC.Tn[4].n45 VGND 0.13077f
C12793 XThC.Tn[4].t23 VGND 0.01443f
C12794 XThC.Tn[4].t17 VGND 0.01576f
C12795 XThC.Tn[4].n46 VGND 0.03519f
C12796 XThC.Tn[4].n47 VGND 0.02411f
C12797 XThC.Tn[4].n48 VGND 0.07935f
C12798 XThC.Tn[4].n49 VGND 0.13077f
C12799 XThC.Tn[4].t34 VGND 0.01443f
C12800 XThC.Tn[4].t30 VGND 0.01576f
C12801 XThC.Tn[4].n50 VGND 0.03519f
C12802 XThC.Tn[4].n51 VGND 0.02411f
C12803 XThC.Tn[4].n52 VGND 0.07935f
C12804 XThC.Tn[4].n53 VGND 0.13077f
C12805 XThC.Tn[4].t42 VGND 0.01443f
C12806 XThC.Tn[4].t38 VGND 0.01576f
C12807 XThC.Tn[4].n54 VGND 0.03519f
C12808 XThC.Tn[4].n55 VGND 0.02411f
C12809 XThC.Tn[4].n56 VGND 0.07935f
C12810 XThC.Tn[4].n57 VGND 0.13077f
C12811 XThC.Tn[4].t12 VGND 0.01443f
C12812 XThC.Tn[4].t41 VGND 0.01576f
C12813 XThC.Tn[4].n58 VGND 0.03519f
C12814 XThC.Tn[4].n59 VGND 0.02411f
C12815 XThC.Tn[4].n60 VGND 0.07935f
C12816 XThC.Tn[4].n61 VGND 0.13077f
C12817 XThC.Tn[4].t25 VGND 0.01443f
C12818 XThC.Tn[4].t22 VGND 0.01576f
C12819 XThC.Tn[4].n62 VGND 0.03519f
C12820 XThC.Tn[4].n63 VGND 0.02411f
C12821 XThC.Tn[4].n64 VGND 0.07935f
C12822 XThC.Tn[4].n65 VGND 0.13077f
C12823 XThC.Tn[4].t35 VGND 0.01443f
C12824 XThC.Tn[4].t32 VGND 0.01576f
C12825 XThC.Tn[4].n66 VGND 0.03519f
C12826 XThC.Tn[4].n67 VGND 0.02411f
C12827 XThC.Tn[4].n68 VGND 0.07935f
C12828 XThC.Tn[4].n69 VGND 0.13077f
C12829 XThC.Tn[4].n70 VGND 0.16028f
C12830 XThC.Tn[4].t1 VGND 0.01821f
C12831 XThC.Tn[4].t0 VGND 0.01821f
C12832 XThC.Tn[4].n71 VGND 0.03675f
C12833 XThC.Tn[4].t3 VGND 0.01821f
C12834 XThC.Tn[4].t2 VGND 0.01821f
C12835 XThC.Tn[4].n72 VGND 0.043f
C12836 XThC.Tn[4].n73 VGND 0.12038f
C12837 XThC.Tn[4].n74 VGND 0.0381f
C12838 XThR.Tn[5].t6 VGND 0.02327f
C12839 XThR.Tn[5].t7 VGND 0.02327f
C12840 XThR.Tn[5].n0 VGND 0.04698f
C12841 XThR.Tn[5].t5 VGND 0.02327f
C12842 XThR.Tn[5].t4 VGND 0.02327f
C12843 XThR.Tn[5].n1 VGND 0.05497f
C12844 XThR.Tn[5].n2 VGND 0.15388f
C12845 XThR.Tn[5].t11 VGND 0.01513f
C12846 XThR.Tn[5].t8 VGND 0.01513f
C12847 XThR.Tn[5].n3 VGND 0.03445f
C12848 XThR.Tn[5].t10 VGND 0.01513f
C12849 XThR.Tn[5].t9 VGND 0.01513f
C12850 XThR.Tn[5].n4 VGND 0.03445f
C12851 XThR.Tn[5].t0 VGND 0.01513f
C12852 XThR.Tn[5].t1 VGND 0.01513f
C12853 XThR.Tn[5].n5 VGND 0.0574f
C12854 XThR.Tn[5].t3 VGND 0.01513f
C12855 XThR.Tn[5].t2 VGND 0.01513f
C12856 XThR.Tn[5].n6 VGND 0.03445f
C12857 XThR.Tn[5].n7 VGND 0.16407f
C12858 XThR.Tn[5].n8 VGND 0.10142f
C12859 XThR.Tn[5].n9 VGND 0.11446f
C12860 XThR.Tn[5].t17 VGND 0.01819f
C12861 XThR.Tn[5].t72 VGND 0.01992f
C12862 XThR.Tn[5].n10 VGND 0.04864f
C12863 XThR.Tn[5].n11 VGND 0.09344f
C12864 XThR.Tn[5].t39 VGND 0.01819f
C12865 XThR.Tn[5].t26 VGND 0.01992f
C12866 XThR.Tn[5].n12 VGND 0.04864f
C12867 XThR.Tn[5].t13 VGND 0.01813f
C12868 XThR.Tn[5].t23 VGND 0.01985f
C12869 XThR.Tn[5].n13 VGND 0.05061f
C12870 XThR.Tn[5].n14 VGND 0.03555f
C12871 XThR.Tn[5].n15 VGND 0.0065f
C12872 XThR.Tn[5].n16 VGND 0.11409f
C12873 XThR.Tn[5].t73 VGND 0.01819f
C12874 XThR.Tn[5].t66 VGND 0.01992f
C12875 XThR.Tn[5].n17 VGND 0.04864f
C12876 XThR.Tn[5].t48 VGND 0.01813f
C12877 XThR.Tn[5].t61 VGND 0.01985f
C12878 XThR.Tn[5].n18 VGND 0.05061f
C12879 XThR.Tn[5].n19 VGND 0.03555f
C12880 XThR.Tn[5].n20 VGND 0.0065f
C12881 XThR.Tn[5].n21 VGND 0.11409f
C12882 XThR.Tn[5].t28 VGND 0.01819f
C12883 XThR.Tn[5].t21 VGND 0.01992f
C12884 XThR.Tn[5].n22 VGND 0.04864f
C12885 XThR.Tn[5].t65 VGND 0.01813f
C12886 XThR.Tn[5].t18 VGND 0.01985f
C12887 XThR.Tn[5].n23 VGND 0.05061f
C12888 XThR.Tn[5].n24 VGND 0.03555f
C12889 XThR.Tn[5].n25 VGND 0.0065f
C12890 XThR.Tn[5].n26 VGND 0.11409f
C12891 XThR.Tn[5].t55 VGND 0.01819f
C12892 XThR.Tn[5].t51 VGND 0.01992f
C12893 XThR.Tn[5].n27 VGND 0.04864f
C12894 XThR.Tn[5].t33 VGND 0.01813f
C12895 XThR.Tn[5].t46 VGND 0.01985f
C12896 XThR.Tn[5].n28 VGND 0.05061f
C12897 XThR.Tn[5].n29 VGND 0.03555f
C12898 XThR.Tn[5].n30 VGND 0.0065f
C12899 XThR.Tn[5].n31 VGND 0.11409f
C12900 XThR.Tn[5].t30 VGND 0.01819f
C12901 XThR.Tn[5].t22 VGND 0.01992f
C12902 XThR.Tn[5].n32 VGND 0.04864f
C12903 XThR.Tn[5].t67 VGND 0.01813f
C12904 XThR.Tn[5].t19 VGND 0.01985f
C12905 XThR.Tn[5].n33 VGND 0.05061f
C12906 XThR.Tn[5].n34 VGND 0.03555f
C12907 XThR.Tn[5].n35 VGND 0.0065f
C12908 XThR.Tn[5].n36 VGND 0.11409f
C12909 XThR.Tn[5].t69 VGND 0.01819f
C12910 XThR.Tn[5].t40 VGND 0.01992f
C12911 XThR.Tn[5].n37 VGND 0.04864f
C12912 XThR.Tn[5].t43 VGND 0.01813f
C12913 XThR.Tn[5].t37 VGND 0.01985f
C12914 XThR.Tn[5].n38 VGND 0.05061f
C12915 XThR.Tn[5].n39 VGND 0.03555f
C12916 XThR.Tn[5].n40 VGND 0.0065f
C12917 XThR.Tn[5].n41 VGND 0.11409f
C12918 XThR.Tn[5].t38 VGND 0.01819f
C12919 XThR.Tn[5].t32 VGND 0.01992f
C12920 XThR.Tn[5].n42 VGND 0.04864f
C12921 XThR.Tn[5].t14 VGND 0.01813f
C12922 XThR.Tn[5].t29 VGND 0.01985f
C12923 XThR.Tn[5].n43 VGND 0.05061f
C12924 XThR.Tn[5].n44 VGND 0.03555f
C12925 XThR.Tn[5].n45 VGND 0.0065f
C12926 XThR.Tn[5].n46 VGND 0.11409f
C12927 XThR.Tn[5].t42 VGND 0.01819f
C12928 XThR.Tn[5].t49 VGND 0.01992f
C12929 XThR.Tn[5].n47 VGND 0.04864f
C12930 XThR.Tn[5].t16 VGND 0.01813f
C12931 XThR.Tn[5].t45 VGND 0.01985f
C12932 XThR.Tn[5].n48 VGND 0.05061f
C12933 XThR.Tn[5].n49 VGND 0.03555f
C12934 XThR.Tn[5].n50 VGND 0.0065f
C12935 XThR.Tn[5].n51 VGND 0.11409f
C12936 XThR.Tn[5].t58 VGND 0.01819f
C12937 XThR.Tn[5].t68 VGND 0.01992f
C12938 XThR.Tn[5].n52 VGND 0.04864f
C12939 XThR.Tn[5].t36 VGND 0.01813f
C12940 XThR.Tn[5].t63 VGND 0.01985f
C12941 XThR.Tn[5].n53 VGND 0.05061f
C12942 XThR.Tn[5].n54 VGND 0.03555f
C12943 XThR.Tn[5].n55 VGND 0.0065f
C12944 XThR.Tn[5].n56 VGND 0.11409f
C12945 XThR.Tn[5].t53 VGND 0.01819f
C12946 XThR.Tn[5].t24 VGND 0.01992f
C12947 XThR.Tn[5].n57 VGND 0.04864f
C12948 XThR.Tn[5].t25 VGND 0.01813f
C12949 XThR.Tn[5].t20 VGND 0.01985f
C12950 XThR.Tn[5].n58 VGND 0.05061f
C12951 XThR.Tn[5].n59 VGND 0.03555f
C12952 XThR.Tn[5].n60 VGND 0.0065f
C12953 XThR.Tn[5].n61 VGND 0.11409f
C12954 XThR.Tn[5].t71 VGND 0.01819f
C12955 XThR.Tn[5].t60 VGND 0.01992f
C12956 XThR.Tn[5].n62 VGND 0.04864f
C12957 XThR.Tn[5].t44 VGND 0.01813f
C12958 XThR.Tn[5].t57 VGND 0.01985f
C12959 XThR.Tn[5].n63 VGND 0.05061f
C12960 XThR.Tn[5].n64 VGND 0.03555f
C12961 XThR.Tn[5].n65 VGND 0.0065f
C12962 XThR.Tn[5].n66 VGND 0.11409f
C12963 XThR.Tn[5].t41 VGND 0.01819f
C12964 XThR.Tn[5].t35 VGND 0.01992f
C12965 XThR.Tn[5].n67 VGND 0.04864f
C12966 XThR.Tn[5].t15 VGND 0.01813f
C12967 XThR.Tn[5].t31 VGND 0.01985f
C12968 XThR.Tn[5].n68 VGND 0.05061f
C12969 XThR.Tn[5].n69 VGND 0.03555f
C12970 XThR.Tn[5].n70 VGND 0.0065f
C12971 XThR.Tn[5].n71 VGND 0.11409f
C12972 XThR.Tn[5].t56 VGND 0.01819f
C12973 XThR.Tn[5].t52 VGND 0.01992f
C12974 XThR.Tn[5].n72 VGND 0.04864f
C12975 XThR.Tn[5].t34 VGND 0.01813f
C12976 XThR.Tn[5].t47 VGND 0.01985f
C12977 XThR.Tn[5].n73 VGND 0.05061f
C12978 XThR.Tn[5].n74 VGND 0.03555f
C12979 XThR.Tn[5].n75 VGND 0.0065f
C12980 XThR.Tn[5].n76 VGND 0.11409f
C12981 XThR.Tn[5].t12 VGND 0.01819f
C12982 XThR.Tn[5].t70 VGND 0.01992f
C12983 XThR.Tn[5].n77 VGND 0.04864f
C12984 XThR.Tn[5].t50 VGND 0.01813f
C12985 XThR.Tn[5].t64 VGND 0.01985f
C12986 XThR.Tn[5].n78 VGND 0.05061f
C12987 XThR.Tn[5].n79 VGND 0.03555f
C12988 XThR.Tn[5].n80 VGND 0.0065f
C12989 XThR.Tn[5].n81 VGND 0.11409f
C12990 XThR.Tn[5].t54 VGND 0.01819f
C12991 XThR.Tn[5].t62 VGND 0.01992f
C12992 XThR.Tn[5].n82 VGND 0.04864f
C12993 XThR.Tn[5].t27 VGND 0.01813f
C12994 XThR.Tn[5].t59 VGND 0.01985f
C12995 XThR.Tn[5].n83 VGND 0.05061f
C12996 XThR.Tn[5].n84 VGND 0.03555f
C12997 XThR.Tn[5].n85 VGND 0.0065f
C12998 XThR.Tn[5].n86 VGND 0.11409f
C12999 XThR.Tn[5].n87 VGND 0.10368f
C13000 XThR.Tn[5].n88 VGND 0.20081f
C13001 XThR.Tn[5].n89 VGND 0.0487f
C13002 XThR.Tn[3].t5 VGND 0.02315f
C13003 XThR.Tn[3].t6 VGND 0.02315f
C13004 XThR.Tn[3].n0 VGND 0.04673f
C13005 XThR.Tn[3].t4 VGND 0.02315f
C13006 XThR.Tn[3].t7 VGND 0.02315f
C13007 XThR.Tn[3].n1 VGND 0.05468f
C13008 XThR.Tn[3].n2 VGND 0.15307f
C13009 XThR.Tn[3].t11 VGND 0.01505f
C13010 XThR.Tn[3].t8 VGND 0.01505f
C13011 XThR.Tn[3].n3 VGND 0.03427f
C13012 XThR.Tn[3].t10 VGND 0.01505f
C13013 XThR.Tn[3].t9 VGND 0.01505f
C13014 XThR.Tn[3].n4 VGND 0.03427f
C13015 XThR.Tn[3].t0 VGND 0.01505f
C13016 XThR.Tn[3].t1 VGND 0.01505f
C13017 XThR.Tn[3].n5 VGND 0.0571f
C13018 XThR.Tn[3].t3 VGND 0.01505f
C13019 XThR.Tn[3].t2 VGND 0.01505f
C13020 XThR.Tn[3].n6 VGND 0.03427f
C13021 XThR.Tn[3].n7 VGND 0.16319f
C13022 XThR.Tn[3].n8 VGND 0.10088f
C13023 XThR.Tn[3].n9 VGND 0.11385f
C13024 XThR.Tn[3].t64 VGND 0.01809f
C13025 XThR.Tn[3].t57 VGND 0.01981f
C13026 XThR.Tn[3].n10 VGND 0.04838f
C13027 XThR.Tn[3].n11 VGND 0.09294f
C13028 XThR.Tn[3].t18 VGND 0.01809f
C13029 XThR.Tn[3].t70 VGND 0.01981f
C13030 XThR.Tn[3].n12 VGND 0.04838f
C13031 XThR.Tn[3].t24 VGND 0.01803f
C13032 XThR.Tn[3].t55 VGND 0.01975f
C13033 XThR.Tn[3].n13 VGND 0.05034f
C13034 XThR.Tn[3].n14 VGND 0.03536f
C13035 XThR.Tn[3].n15 VGND 0.00647f
C13036 XThR.Tn[3].n16 VGND 0.11349f
C13037 XThR.Tn[3].t59 VGND 0.01809f
C13038 XThR.Tn[3].t49 VGND 0.01981f
C13039 XThR.Tn[3].n17 VGND 0.04838f
C13040 XThR.Tn[3].t62 VGND 0.01803f
C13041 XThR.Tn[3].t29 VGND 0.01975f
C13042 XThR.Tn[3].n18 VGND 0.05034f
C13043 XThR.Tn[3].n19 VGND 0.03536f
C13044 XThR.Tn[3].n20 VGND 0.00647f
C13045 XThR.Tn[3].n21 VGND 0.11349f
C13046 XThR.Tn[3].t71 VGND 0.01809f
C13047 XThR.Tn[3].t67 VGND 0.01981f
C13048 XThR.Tn[3].n22 VGND 0.04838f
C13049 XThR.Tn[3].t12 VGND 0.01803f
C13050 XThR.Tn[3].t47 VGND 0.01975f
C13051 XThR.Tn[3].n23 VGND 0.05034f
C13052 XThR.Tn[3].n24 VGND 0.03536f
C13053 XThR.Tn[3].n25 VGND 0.00647f
C13054 XThR.Tn[3].n26 VGND 0.11349f
C13055 XThR.Tn[3].t39 VGND 0.01809f
C13056 XThR.Tn[3].t33 VGND 0.01981f
C13057 XThR.Tn[3].n27 VGND 0.04838f
C13058 XThR.Tn[3].t42 VGND 0.01803f
C13059 XThR.Tn[3].t13 VGND 0.01975f
C13060 XThR.Tn[3].n28 VGND 0.05034f
C13061 XThR.Tn[3].n29 VGND 0.03536f
C13062 XThR.Tn[3].n30 VGND 0.00647f
C13063 XThR.Tn[3].n31 VGND 0.11349f
C13064 XThR.Tn[3].t72 VGND 0.01809f
C13065 XThR.Tn[3].t68 VGND 0.01981f
C13066 XThR.Tn[3].n32 VGND 0.04838f
C13067 XThR.Tn[3].t16 VGND 0.01803f
C13068 XThR.Tn[3].t48 VGND 0.01975f
C13069 XThR.Tn[3].n33 VGND 0.05034f
C13070 XThR.Tn[3].n34 VGND 0.03536f
C13071 XThR.Tn[3].n35 VGND 0.00647f
C13072 XThR.Tn[3].n36 VGND 0.11349f
C13073 XThR.Tn[3].t52 VGND 0.01809f
C13074 XThR.Tn[3].t20 VGND 0.01981f
C13075 XThR.Tn[3].n37 VGND 0.04838f
C13076 XThR.Tn[3].t56 VGND 0.01803f
C13077 XThR.Tn[3].t66 VGND 0.01975f
C13078 XThR.Tn[3].n38 VGND 0.05034f
C13079 XThR.Tn[3].n39 VGND 0.03536f
C13080 XThR.Tn[3].n40 VGND 0.00647f
C13081 XThR.Tn[3].n41 VGND 0.11349f
C13082 XThR.Tn[3].t19 VGND 0.01809f
C13083 XThR.Tn[3].t14 VGND 0.01981f
C13084 XThR.Tn[3].n42 VGND 0.04838f
C13085 XThR.Tn[3].t23 VGND 0.01803f
C13086 XThR.Tn[3].t61 VGND 0.01975f
C13087 XThR.Tn[3].n43 VGND 0.05034f
C13088 XThR.Tn[3].n44 VGND 0.03536f
C13089 XThR.Tn[3].n45 VGND 0.00647f
C13090 XThR.Tn[3].n46 VGND 0.11349f
C13091 XThR.Tn[3].t22 VGND 0.01809f
C13092 XThR.Tn[3].t31 VGND 0.01981f
C13093 XThR.Tn[3].n47 VGND 0.04838f
C13094 XThR.Tn[3].t28 VGND 0.01803f
C13095 XThR.Tn[3].t73 VGND 0.01975f
C13096 XThR.Tn[3].n48 VGND 0.05034f
C13097 XThR.Tn[3].n49 VGND 0.03536f
C13098 XThR.Tn[3].n50 VGND 0.00647f
C13099 XThR.Tn[3].n51 VGND 0.11349f
C13100 XThR.Tn[3].t41 VGND 0.01809f
C13101 XThR.Tn[3].t51 VGND 0.01981f
C13102 XThR.Tn[3].n52 VGND 0.04838f
C13103 XThR.Tn[3].t45 VGND 0.01803f
C13104 XThR.Tn[3].t30 VGND 0.01975f
C13105 XThR.Tn[3].n53 VGND 0.05034f
C13106 XThR.Tn[3].n54 VGND 0.03536f
C13107 XThR.Tn[3].n55 VGND 0.00647f
C13108 XThR.Tn[3].n56 VGND 0.11349f
C13109 XThR.Tn[3].t35 VGND 0.01809f
C13110 XThR.Tn[3].t69 VGND 0.01981f
C13111 XThR.Tn[3].n57 VGND 0.04838f
C13112 XThR.Tn[3].t37 VGND 0.01803f
C13113 XThR.Tn[3].t50 VGND 0.01975f
C13114 XThR.Tn[3].n58 VGND 0.05034f
C13115 XThR.Tn[3].n59 VGND 0.03536f
C13116 XThR.Tn[3].n60 VGND 0.00647f
C13117 XThR.Tn[3].n61 VGND 0.11349f
C13118 XThR.Tn[3].t54 VGND 0.01809f
C13119 XThR.Tn[3].t44 VGND 0.01981f
C13120 XThR.Tn[3].n62 VGND 0.04838f
C13121 XThR.Tn[3].t58 VGND 0.01803f
C13122 XThR.Tn[3].t25 VGND 0.01975f
C13123 XThR.Tn[3].n63 VGND 0.05034f
C13124 XThR.Tn[3].n64 VGND 0.03536f
C13125 XThR.Tn[3].n65 VGND 0.00647f
C13126 XThR.Tn[3].n66 VGND 0.11349f
C13127 XThR.Tn[3].t21 VGND 0.01809f
C13128 XThR.Tn[3].t17 VGND 0.01981f
C13129 XThR.Tn[3].n67 VGND 0.04838f
C13130 XThR.Tn[3].t26 VGND 0.01803f
C13131 XThR.Tn[3].t63 VGND 0.01975f
C13132 XThR.Tn[3].n68 VGND 0.05034f
C13133 XThR.Tn[3].n69 VGND 0.03536f
C13134 XThR.Tn[3].n70 VGND 0.00647f
C13135 XThR.Tn[3].n71 VGND 0.11349f
C13136 XThR.Tn[3].t40 VGND 0.01809f
C13137 XThR.Tn[3].t34 VGND 0.01981f
C13138 XThR.Tn[3].n72 VGND 0.04838f
C13139 XThR.Tn[3].t43 VGND 0.01803f
C13140 XThR.Tn[3].t15 VGND 0.01975f
C13141 XThR.Tn[3].n73 VGND 0.05034f
C13142 XThR.Tn[3].n74 VGND 0.03536f
C13143 XThR.Tn[3].n75 VGND 0.00647f
C13144 XThR.Tn[3].n76 VGND 0.11349f
C13145 XThR.Tn[3].t60 VGND 0.01809f
C13146 XThR.Tn[3].t53 VGND 0.01981f
C13147 XThR.Tn[3].n77 VGND 0.04838f
C13148 XThR.Tn[3].t65 VGND 0.01803f
C13149 XThR.Tn[3].t32 VGND 0.01975f
C13150 XThR.Tn[3].n78 VGND 0.05034f
C13151 XThR.Tn[3].n79 VGND 0.03536f
C13152 XThR.Tn[3].n80 VGND 0.00647f
C13153 XThR.Tn[3].n81 VGND 0.11349f
C13154 XThR.Tn[3].t36 VGND 0.01809f
C13155 XThR.Tn[3].t46 VGND 0.01981f
C13156 XThR.Tn[3].n82 VGND 0.04838f
C13157 XThR.Tn[3].t38 VGND 0.01803f
C13158 XThR.Tn[3].t27 VGND 0.01975f
C13159 XThR.Tn[3].n83 VGND 0.05034f
C13160 XThR.Tn[3].n84 VGND 0.03536f
C13161 XThR.Tn[3].n85 VGND 0.00647f
C13162 XThR.Tn[3].n86 VGND 0.11349f
C13163 XThR.Tn[3].n87 VGND 0.10313f
C13164 XThR.Tn[3].n88 VGND 0.22842f
C13165 XThR.Tn[3].n89 VGND 0.04845f
C13166 XThC.TB4.t1 VGND 0.12238f
C13167 XThC.TB4.n0 VGND 0.16166f
C13168 XThC.TB4.t4 VGND 0.02956f
C13169 XThC.TB4.t13 VGND 0.05016f
C13170 XThC.TB4.n1 VGND 0.05972f
C13171 XThC.TB4.t7 VGND 0.02956f
C13172 XThC.TB4.t17 VGND 0.05016f
C13173 XThC.TB4.n2 VGND 0.03074f
C13174 XThC.TB4.t10 VGND 0.02956f
C13175 XThC.TB4.t2 VGND 0.05016f
C13176 XThC.TB4.n3 VGND 0.06603f
C13177 XThC.TB4.t14 VGND 0.02956f
C13178 XThC.TB4.t3 VGND 0.05016f
C13179 XThC.TB4.n4 VGND 0.0613f
C13180 XThC.TB4.n5 VGND 0.03729f
C13181 XThC.TB4.n6 VGND 0.06174f
C13182 XThC.TB4.n7 VGND 0.02389f
C13183 XThC.TB4.n8 VGND 0.02916f
C13184 XThC.TB4.n9 VGND 0.06603f
C13185 XThC.TB4.n10 VGND 0.0331f
C13186 XThC.TB4.n11 VGND 0.06459f
C13187 XThC.TB4.t5 VGND 0.02956f
C13188 XThC.TB4.t16 VGND 0.05016f
C13189 XThC.TB4.n12 VGND 0.06761f
C13190 XThC.TB4.t9 VGND 0.02956f
C13191 XThC.TB4.t6 VGND 0.05016f
C13192 XThC.TB4.t15 VGND 0.02956f
C13193 XThC.TB4.t12 VGND 0.05016f
C13194 XThC.TB4.t11 VGND 0.02956f
C13195 XThC.TB4.t8 VGND 0.05016f
C13196 XThC.TB4.n13 VGND 0.08416f
C13197 XThC.TB4.n14 VGND 0.08889f
C13198 XThC.TB4.n15 VGND 0.03426f
C13199 XThC.TB4.n16 VGND 0.07234f
C13200 XThC.TB4.n17 VGND 0.0331f
C13201 XThC.TB4.n18 VGND 0.02701f
C13202 XThC.TB4.n19 VGND 0.48759f
C13203 XThC.TB4.n20 VGND 0.34501f
C13204 XThC.TB4.n21 VGND 0.08408f
C13205 XThC.TB4.t0 VGND 0.06491f
C13206 XThC.TB4.n22 VGND 0.04329f
C13207 XThC.Tn[0].t2 VGND 0.01209f
C13208 XThC.Tn[0].t1 VGND 0.01209f
C13209 XThC.Tn[0].n0 VGND 0.0244f
C13210 XThC.Tn[0].t4 VGND 0.01209f
C13211 XThC.Tn[0].t3 VGND 0.01209f
C13212 XThC.Tn[0].n1 VGND 0.02855f
C13213 XThC.Tn[0].n2 VGND 0.07993f
C13214 XThC.Tn[0].t6 VGND 0.00786f
C13215 XThC.Tn[0].t5 VGND 0.00786f
C13216 XThC.Tn[0].n3 VGND 0.01789f
C13217 XThC.Tn[0].t8 VGND 0.00786f
C13218 XThC.Tn[0].t7 VGND 0.00786f
C13219 XThC.Tn[0].n4 VGND 0.01789f
C13220 XThC.Tn[0].t10 VGND 0.00786f
C13221 XThC.Tn[0].t11 VGND 0.00786f
C13222 XThC.Tn[0].n5 VGND 0.01789f
C13223 XThC.Tn[0].t0 VGND 0.00786f
C13224 XThC.Tn[0].t9 VGND 0.00786f
C13225 XThC.Tn[0].n6 VGND 0.02982f
C13226 XThC.Tn[0].n7 VGND 0.08522f
C13227 XThC.Tn[0].n8 VGND 0.05268f
C13228 XThC.Tn[0].n9 VGND 0.05945f
C13229 XThC.Tn[0].t18 VGND 0.00958f
C13230 XThC.Tn[0].t22 VGND 0.01047f
C13231 XThC.Tn[0].n10 VGND 0.02336f
C13232 XThC.Tn[0].n11 VGND 0.01601f
C13233 XThC.Tn[0].n12 VGND 0.05254f
C13234 XThC.Tn[0].t35 VGND 0.00958f
C13235 XThC.Tn[0].t41 VGND 0.01047f
C13236 XThC.Tn[0].n13 VGND 0.02336f
C13237 XThC.Tn[0].n14 VGND 0.01601f
C13238 XThC.Tn[0].n15 VGND 0.05268f
C13239 XThC.Tn[0].n16 VGND 0.08683f
C13240 XThC.Tn[0].t37 VGND 0.00958f
C13241 XThC.Tn[0].t12 VGND 0.01047f
C13242 XThC.Tn[0].n17 VGND 0.02336f
C13243 XThC.Tn[0].n18 VGND 0.01601f
C13244 XThC.Tn[0].n19 VGND 0.05268f
C13245 XThC.Tn[0].n20 VGND 0.08683f
C13246 XThC.Tn[0].t39 VGND 0.00958f
C13247 XThC.Tn[0].t13 VGND 0.01047f
C13248 XThC.Tn[0].n21 VGND 0.02336f
C13249 XThC.Tn[0].n22 VGND 0.01601f
C13250 XThC.Tn[0].n23 VGND 0.05268f
C13251 XThC.Tn[0].n24 VGND 0.08683f
C13252 XThC.Tn[0].t28 VGND 0.00958f
C13253 XThC.Tn[0].t32 VGND 0.01047f
C13254 XThC.Tn[0].n25 VGND 0.02336f
C13255 XThC.Tn[0].n26 VGND 0.01601f
C13256 XThC.Tn[0].n27 VGND 0.05268f
C13257 XThC.Tn[0].n28 VGND 0.08683f
C13258 XThC.Tn[0].t30 VGND 0.00958f
C13259 XThC.Tn[0].t34 VGND 0.01047f
C13260 XThC.Tn[0].n29 VGND 0.02336f
C13261 XThC.Tn[0].n30 VGND 0.01601f
C13262 XThC.Tn[0].n31 VGND 0.05268f
C13263 XThC.Tn[0].n32 VGND 0.08683f
C13264 XThC.Tn[0].t43 VGND 0.00958f
C13265 XThC.Tn[0].t17 VGND 0.01047f
C13266 XThC.Tn[0].n33 VGND 0.02336f
C13267 XThC.Tn[0].n34 VGND 0.01601f
C13268 XThC.Tn[0].n35 VGND 0.05268f
C13269 XThC.Tn[0].n36 VGND 0.08683f
C13270 XThC.Tn[0].t20 VGND 0.00958f
C13271 XThC.Tn[0].t25 VGND 0.01047f
C13272 XThC.Tn[0].n37 VGND 0.02336f
C13273 XThC.Tn[0].n38 VGND 0.01601f
C13274 XThC.Tn[0].n39 VGND 0.05268f
C13275 XThC.Tn[0].n40 VGND 0.08683f
C13276 XThC.Tn[0].t21 VGND 0.00958f
C13277 XThC.Tn[0].t26 VGND 0.01047f
C13278 XThC.Tn[0].n41 VGND 0.02336f
C13279 XThC.Tn[0].n42 VGND 0.01601f
C13280 XThC.Tn[0].n43 VGND 0.05268f
C13281 XThC.Tn[0].n44 VGND 0.08683f
C13282 XThC.Tn[0].t40 VGND 0.00958f
C13283 XThC.Tn[0].t15 VGND 0.01047f
C13284 XThC.Tn[0].n45 VGND 0.02336f
C13285 XThC.Tn[0].n46 VGND 0.01601f
C13286 XThC.Tn[0].n47 VGND 0.05268f
C13287 XThC.Tn[0].n48 VGND 0.08683f
C13288 XThC.Tn[0].t42 VGND 0.00958f
C13289 XThC.Tn[0].t16 VGND 0.01047f
C13290 XThC.Tn[0].n49 VGND 0.02336f
C13291 XThC.Tn[0].n50 VGND 0.01601f
C13292 XThC.Tn[0].n51 VGND 0.05268f
C13293 XThC.Tn[0].n52 VGND 0.08683f
C13294 XThC.Tn[0].t23 VGND 0.00958f
C13295 XThC.Tn[0].t27 VGND 0.01047f
C13296 XThC.Tn[0].n53 VGND 0.02336f
C13297 XThC.Tn[0].n54 VGND 0.01601f
C13298 XThC.Tn[0].n55 VGND 0.05268f
C13299 XThC.Tn[0].n56 VGND 0.08683f
C13300 XThC.Tn[0].t31 VGND 0.00958f
C13301 XThC.Tn[0].t36 VGND 0.01047f
C13302 XThC.Tn[0].n57 VGND 0.02336f
C13303 XThC.Tn[0].n58 VGND 0.01601f
C13304 XThC.Tn[0].n59 VGND 0.05268f
C13305 XThC.Tn[0].n60 VGND 0.08683f
C13306 XThC.Tn[0].t33 VGND 0.00958f
C13307 XThC.Tn[0].t38 VGND 0.01047f
C13308 XThC.Tn[0].n61 VGND 0.02336f
C13309 XThC.Tn[0].n62 VGND 0.01601f
C13310 XThC.Tn[0].n63 VGND 0.05268f
C13311 XThC.Tn[0].n64 VGND 0.08683f
C13312 XThC.Tn[0].t14 VGND 0.00958f
C13313 XThC.Tn[0].t19 VGND 0.01047f
C13314 XThC.Tn[0].n65 VGND 0.02336f
C13315 XThC.Tn[0].n66 VGND 0.01601f
C13316 XThC.Tn[0].n67 VGND 0.05268f
C13317 XThC.Tn[0].n68 VGND 0.08683f
C13318 XThC.Tn[0].t24 VGND 0.00958f
C13319 XThC.Tn[0].t29 VGND 0.01047f
C13320 XThC.Tn[0].n69 VGND 0.02336f
C13321 XThC.Tn[0].n70 VGND 0.01601f
C13322 XThC.Tn[0].n71 VGND 0.05268f
C13323 XThC.Tn[0].n72 VGND 0.08683f
C13324 XThC.Tn[0].n73 VGND 0.53669f
C13325 XThC.Tn[0].n74 VGND 0.06506f
C13326 XThC.Tn[0].n75 VGND 0.0253f
C13327 XThC.Tn[13].t6 VGND 0.0195f
C13328 XThC.Tn[13].t5 VGND 0.0195f
C13329 XThC.Tn[13].n0 VGND 0.04213f
C13330 XThC.Tn[13].t4 VGND 0.0195f
C13331 XThC.Tn[13].t7 VGND 0.0195f
C13332 XThC.Tn[13].n1 VGND 0.06641f
C13333 XThC.Tn[13].n2 VGND 0.17588f
C13334 XThC.Tn[13].t9 VGND 0.0195f
C13335 XThC.Tn[13].t8 VGND 0.0195f
C13336 XThC.Tn[13].n3 VGND 0.05921f
C13337 XThC.Tn[13].t11 VGND 0.0195f
C13338 XThC.Tn[13].t10 VGND 0.0195f
C13339 XThC.Tn[13].n4 VGND 0.04335f
C13340 XThC.Tn[13].n5 VGND 0.19292f
C13341 XThC.Tn[13].n6 VGND 0.01295f
C13342 XThC.Tn[13].t29 VGND 0.01546f
C13343 XThC.Tn[13].t27 VGND 0.01688f
C13344 XThC.Tn[13].n7 VGND 0.03768f
C13345 XThC.Tn[13].n8 VGND 0.02582f
C13346 XThC.Tn[13].n9 VGND 0.08475f
C13347 XThC.Tn[13].t15 VGND 0.01546f
C13348 XThC.Tn[13].t12 VGND 0.01688f
C13349 XThC.Tn[13].n10 VGND 0.03768f
C13350 XThC.Tn[13].n11 VGND 0.02582f
C13351 XThC.Tn[13].n12 VGND 0.08498f
C13352 XThC.Tn[13].n13 VGND 0.14005f
C13353 XThC.Tn[13].t20 VGND 0.01546f
C13354 XThC.Tn[13].t14 VGND 0.01688f
C13355 XThC.Tn[13].n14 VGND 0.03768f
C13356 XThC.Tn[13].n15 VGND 0.02582f
C13357 XThC.Tn[13].n16 VGND 0.08498f
C13358 XThC.Tn[13].n17 VGND 0.14005f
C13359 XThC.Tn[13].t21 VGND 0.01546f
C13360 XThC.Tn[13].t16 VGND 0.01688f
C13361 XThC.Tn[13].n18 VGND 0.03768f
C13362 XThC.Tn[13].n19 VGND 0.02582f
C13363 XThC.Tn[13].n20 VGND 0.08498f
C13364 XThC.Tn[13].n21 VGND 0.14005f
C13365 XThC.Tn[13].t40 VGND 0.01546f
C13366 XThC.Tn[13].t37 VGND 0.01688f
C13367 XThC.Tn[13].n22 VGND 0.03768f
C13368 XThC.Tn[13].n23 VGND 0.02582f
C13369 XThC.Tn[13].n24 VGND 0.08498f
C13370 XThC.Tn[13].n25 VGND 0.14005f
C13371 XThC.Tn[13].t41 VGND 0.01546f
C13372 XThC.Tn[13].t38 VGND 0.01688f
C13373 XThC.Tn[13].n26 VGND 0.03768f
C13374 XThC.Tn[13].n27 VGND 0.02582f
C13375 XThC.Tn[13].n28 VGND 0.08498f
C13376 XThC.Tn[13].n29 VGND 0.14005f
C13377 XThC.Tn[13].t25 VGND 0.01546f
C13378 XThC.Tn[13].t19 VGND 0.01688f
C13379 XThC.Tn[13].n30 VGND 0.03768f
C13380 XThC.Tn[13].n31 VGND 0.02582f
C13381 XThC.Tn[13].n32 VGND 0.08498f
C13382 XThC.Tn[13].n33 VGND 0.14005f
C13383 XThC.Tn[13].t32 VGND 0.01546f
C13384 XThC.Tn[13].t28 VGND 0.01688f
C13385 XThC.Tn[13].n34 VGND 0.03768f
C13386 XThC.Tn[13].n35 VGND 0.02582f
C13387 XThC.Tn[13].n36 VGND 0.08498f
C13388 XThC.Tn[13].n37 VGND 0.14005f
C13389 XThC.Tn[13].t34 VGND 0.01546f
C13390 XThC.Tn[13].t30 VGND 0.01688f
C13391 XThC.Tn[13].n38 VGND 0.03768f
C13392 XThC.Tn[13].n39 VGND 0.02582f
C13393 XThC.Tn[13].n40 VGND 0.08498f
C13394 XThC.Tn[13].n41 VGND 0.14005f
C13395 XThC.Tn[13].t22 VGND 0.01546f
C13396 XThC.Tn[13].t17 VGND 0.01688f
C13397 XThC.Tn[13].n42 VGND 0.03768f
C13398 XThC.Tn[13].n43 VGND 0.02582f
C13399 XThC.Tn[13].n44 VGND 0.08498f
C13400 XThC.Tn[13].n45 VGND 0.14005f
C13401 XThC.Tn[13].t24 VGND 0.01546f
C13402 XThC.Tn[13].t18 VGND 0.01688f
C13403 XThC.Tn[13].n46 VGND 0.03768f
C13404 XThC.Tn[13].n47 VGND 0.02582f
C13405 XThC.Tn[13].n48 VGND 0.08498f
C13406 XThC.Tn[13].n49 VGND 0.14005f
C13407 XThC.Tn[13].t35 VGND 0.01546f
C13408 XThC.Tn[13].t31 VGND 0.01688f
C13409 XThC.Tn[13].n50 VGND 0.03768f
C13410 XThC.Tn[13].n51 VGND 0.02582f
C13411 XThC.Tn[13].n52 VGND 0.08498f
C13412 XThC.Tn[13].n53 VGND 0.14005f
C13413 XThC.Tn[13].t43 VGND 0.01546f
C13414 XThC.Tn[13].t39 VGND 0.01688f
C13415 XThC.Tn[13].n54 VGND 0.03768f
C13416 XThC.Tn[13].n55 VGND 0.02582f
C13417 XThC.Tn[13].n56 VGND 0.08498f
C13418 XThC.Tn[13].n57 VGND 0.14005f
C13419 XThC.Tn[13].t13 VGND 0.01546f
C13420 XThC.Tn[13].t42 VGND 0.01688f
C13421 XThC.Tn[13].n58 VGND 0.03768f
C13422 XThC.Tn[13].n59 VGND 0.02582f
C13423 XThC.Tn[13].n60 VGND 0.08498f
C13424 XThC.Tn[13].n61 VGND 0.14005f
C13425 XThC.Tn[13].t26 VGND 0.01546f
C13426 XThC.Tn[13].t23 VGND 0.01688f
C13427 XThC.Tn[13].n62 VGND 0.03768f
C13428 XThC.Tn[13].n63 VGND 0.02582f
C13429 XThC.Tn[13].n64 VGND 0.08498f
C13430 XThC.Tn[13].n65 VGND 0.14005f
C13431 XThC.Tn[13].t36 VGND 0.01546f
C13432 XThC.Tn[13].t33 VGND 0.01688f
C13433 XThC.Tn[13].n66 VGND 0.03768f
C13434 XThC.Tn[13].n67 VGND 0.02582f
C13435 XThC.Tn[13].n68 VGND 0.08498f
C13436 XThC.Tn[13].n69 VGND 0.14005f
C13437 XThC.Tn[13].n70 VGND 0.72631f
C13438 XThC.Tn[13].n71 VGND 0.25541f
C13439 XThC.Tn[13].t0 VGND 0.01267f
C13440 XThC.Tn[13].t2 VGND 0.01267f
C13441 XThC.Tn[13].n72 VGND 0.02535f
C13442 XThC.Tn[13].t3 VGND 0.01267f
C13443 XThC.Tn[13].t1 VGND 0.01267f
C13444 XThC.Tn[13].n73 VGND 0.03161f
C13445 XThC.Tn[13].n74 VGND 0.05845f
C13446 XThC.Tn[12].t7 VGND 0.01298f
C13447 XThC.Tn[12].t6 VGND 0.01298f
C13448 XThC.Tn[12].n0 VGND 0.03236f
C13449 XThC.Tn[12].t5 VGND 0.01298f
C13450 XThC.Tn[12].t4 VGND 0.01298f
C13451 XThC.Tn[12].n1 VGND 0.02595f
C13452 XThC.Tn[12].n2 VGND 0.06529f
C13453 XThC.Tn[12].t37 VGND 0.01582f
C13454 XThC.Tn[12].t35 VGND 0.01728f
C13455 XThC.Tn[12].n3 VGND 0.03858f
C13456 XThC.Tn[12].n4 VGND 0.02643f
C13457 XThC.Tn[12].n5 VGND 0.08676f
C13458 XThC.Tn[12].t23 VGND 0.01582f
C13459 XThC.Tn[12].t20 VGND 0.01728f
C13460 XThC.Tn[12].n6 VGND 0.03858f
C13461 XThC.Tn[12].n7 VGND 0.02643f
C13462 XThC.Tn[12].n8 VGND 0.087f
C13463 XThC.Tn[12].n9 VGND 0.14339f
C13464 XThC.Tn[12].t28 VGND 0.01582f
C13465 XThC.Tn[12].t22 VGND 0.01728f
C13466 XThC.Tn[12].n10 VGND 0.03858f
C13467 XThC.Tn[12].n11 VGND 0.02643f
C13468 XThC.Tn[12].n12 VGND 0.087f
C13469 XThC.Tn[12].n13 VGND 0.14339f
C13470 XThC.Tn[12].t29 VGND 0.01582f
C13471 XThC.Tn[12].t24 VGND 0.01728f
C13472 XThC.Tn[12].n14 VGND 0.03858f
C13473 XThC.Tn[12].n15 VGND 0.02643f
C13474 XThC.Tn[12].n16 VGND 0.087f
C13475 XThC.Tn[12].n17 VGND 0.14339f
C13476 XThC.Tn[12].t16 VGND 0.01582f
C13477 XThC.Tn[12].t13 VGND 0.01728f
C13478 XThC.Tn[12].n18 VGND 0.03858f
C13479 XThC.Tn[12].n19 VGND 0.02643f
C13480 XThC.Tn[12].n20 VGND 0.087f
C13481 XThC.Tn[12].n21 VGND 0.14339f
C13482 XThC.Tn[12].t17 VGND 0.01582f
C13483 XThC.Tn[12].t14 VGND 0.01728f
C13484 XThC.Tn[12].n22 VGND 0.03858f
C13485 XThC.Tn[12].n23 VGND 0.02643f
C13486 XThC.Tn[12].n24 VGND 0.087f
C13487 XThC.Tn[12].n25 VGND 0.14339f
C13488 XThC.Tn[12].t33 VGND 0.01582f
C13489 XThC.Tn[12].t27 VGND 0.01728f
C13490 XThC.Tn[12].n26 VGND 0.03858f
C13491 XThC.Tn[12].n27 VGND 0.02643f
C13492 XThC.Tn[12].n28 VGND 0.087f
C13493 XThC.Tn[12].n29 VGND 0.14339f
C13494 XThC.Tn[12].t40 VGND 0.01582f
C13495 XThC.Tn[12].t36 VGND 0.01728f
C13496 XThC.Tn[12].n30 VGND 0.03858f
C13497 XThC.Tn[12].n31 VGND 0.02643f
C13498 XThC.Tn[12].n32 VGND 0.087f
C13499 XThC.Tn[12].n33 VGND 0.14339f
C13500 XThC.Tn[12].t42 VGND 0.01582f
C13501 XThC.Tn[12].t38 VGND 0.01728f
C13502 XThC.Tn[12].n34 VGND 0.03858f
C13503 XThC.Tn[12].n35 VGND 0.02643f
C13504 XThC.Tn[12].n36 VGND 0.087f
C13505 XThC.Tn[12].n37 VGND 0.14339f
C13506 XThC.Tn[12].t30 VGND 0.01582f
C13507 XThC.Tn[12].t25 VGND 0.01728f
C13508 XThC.Tn[12].n38 VGND 0.03858f
C13509 XThC.Tn[12].n39 VGND 0.02643f
C13510 XThC.Tn[12].n40 VGND 0.087f
C13511 XThC.Tn[12].n41 VGND 0.14339f
C13512 XThC.Tn[12].t32 VGND 0.01582f
C13513 XThC.Tn[12].t26 VGND 0.01728f
C13514 XThC.Tn[12].n42 VGND 0.03858f
C13515 XThC.Tn[12].n43 VGND 0.02643f
C13516 XThC.Tn[12].n44 VGND 0.087f
C13517 XThC.Tn[12].n45 VGND 0.14339f
C13518 XThC.Tn[12].t43 VGND 0.01582f
C13519 XThC.Tn[12].t39 VGND 0.01728f
C13520 XThC.Tn[12].n46 VGND 0.03858f
C13521 XThC.Tn[12].n47 VGND 0.02643f
C13522 XThC.Tn[12].n48 VGND 0.087f
C13523 XThC.Tn[12].n49 VGND 0.14339f
C13524 XThC.Tn[12].t19 VGND 0.01582f
C13525 XThC.Tn[12].t15 VGND 0.01728f
C13526 XThC.Tn[12].n50 VGND 0.03858f
C13527 XThC.Tn[12].n51 VGND 0.02643f
C13528 XThC.Tn[12].n52 VGND 0.087f
C13529 XThC.Tn[12].n53 VGND 0.14339f
C13530 XThC.Tn[12].t21 VGND 0.01582f
C13531 XThC.Tn[12].t18 VGND 0.01728f
C13532 XThC.Tn[12].n54 VGND 0.03858f
C13533 XThC.Tn[12].n55 VGND 0.02643f
C13534 XThC.Tn[12].n56 VGND 0.087f
C13535 XThC.Tn[12].n57 VGND 0.14339f
C13536 XThC.Tn[12].t34 VGND 0.01582f
C13537 XThC.Tn[12].t31 VGND 0.01728f
C13538 XThC.Tn[12].n58 VGND 0.03858f
C13539 XThC.Tn[12].n59 VGND 0.02643f
C13540 XThC.Tn[12].n60 VGND 0.087f
C13541 XThC.Tn[12].n61 VGND 0.14339f
C13542 XThC.Tn[12].t12 VGND 0.01582f
C13543 XThC.Tn[12].t41 VGND 0.01728f
C13544 XThC.Tn[12].n62 VGND 0.03858f
C13545 XThC.Tn[12].n63 VGND 0.02643f
C13546 XThC.Tn[12].n64 VGND 0.087f
C13547 XThC.Tn[12].n65 VGND 0.14339f
C13548 XThC.Tn[12].n66 VGND 0.68185f
C13549 XThC.Tn[12].n67 VGND 0.24221f
C13550 XThC.Tn[12].t9 VGND 0.01996f
C13551 XThC.Tn[12].t10 VGND 0.01996f
C13552 XThC.Tn[12].n68 VGND 0.04313f
C13553 XThC.Tn[12].t8 VGND 0.01996f
C13554 XThC.Tn[12].t11 VGND 0.01996f
C13555 XThC.Tn[12].n69 VGND 0.06565f
C13556 XThC.Tn[12].n70 VGND 0.18241f
C13557 XThC.Tn[12].n71 VGND 0.02868f
C13558 XThC.Tn[12].t1 VGND 0.01996f
C13559 XThC.Tn[12].t0 VGND 0.01996f
C13560 XThC.Tn[12].n72 VGND 0.06062f
C13561 XThC.Tn[12].t3 VGND 0.01996f
C13562 XThC.Tn[12].t2 VGND 0.01996f
C13563 XThC.Tn[12].n73 VGND 0.04438f
C13564 XThC.Tn[12].n74 VGND 0.19752f
C13565 XThC.Tn[11].t11 VGND 0.01319f
C13566 XThC.Tn[11].t2 VGND 0.01319f
C13567 XThC.Tn[11].n0 VGND 0.0329f
C13568 XThC.Tn[11].t5 VGND 0.01319f
C13569 XThC.Tn[11].t3 VGND 0.01319f
C13570 XThC.Tn[11].n1 VGND 0.02638f
C13571 XThC.Tn[11].n2 VGND 0.06083f
C13572 XThC.Tn[11].t20 VGND 0.01608f
C13573 XThC.Tn[11].t18 VGND 0.01757f
C13574 XThC.Tn[11].n3 VGND 0.03922f
C13575 XThC.Tn[11].n4 VGND 0.02687f
C13576 XThC.Tn[11].n5 VGND 0.08819f
C13577 XThC.Tn[11].t38 VGND 0.01608f
C13578 XThC.Tn[11].t35 VGND 0.01757f
C13579 XThC.Tn[11].n6 VGND 0.03922f
C13580 XThC.Tn[11].n7 VGND 0.02687f
C13581 XThC.Tn[11].n8 VGND 0.08843f
C13582 XThC.Tn[11].n9 VGND 0.14574f
C13583 XThC.Tn[11].t43 VGND 0.01608f
C13584 XThC.Tn[11].t37 VGND 0.01757f
C13585 XThC.Tn[11].n10 VGND 0.03922f
C13586 XThC.Tn[11].n11 VGND 0.02687f
C13587 XThC.Tn[11].n12 VGND 0.08843f
C13588 XThC.Tn[11].n13 VGND 0.14574f
C13589 XThC.Tn[11].t12 VGND 0.01608f
C13590 XThC.Tn[11].t39 VGND 0.01757f
C13591 XThC.Tn[11].n14 VGND 0.03922f
C13592 XThC.Tn[11].n15 VGND 0.02687f
C13593 XThC.Tn[11].n16 VGND 0.08843f
C13594 XThC.Tn[11].n17 VGND 0.14574f
C13595 XThC.Tn[11].t31 VGND 0.01608f
C13596 XThC.Tn[11].t28 VGND 0.01757f
C13597 XThC.Tn[11].n18 VGND 0.03922f
C13598 XThC.Tn[11].n19 VGND 0.02687f
C13599 XThC.Tn[11].n20 VGND 0.08843f
C13600 XThC.Tn[11].n21 VGND 0.14574f
C13601 XThC.Tn[11].t32 VGND 0.01608f
C13602 XThC.Tn[11].t29 VGND 0.01757f
C13603 XThC.Tn[11].n22 VGND 0.03922f
C13604 XThC.Tn[11].n23 VGND 0.02687f
C13605 XThC.Tn[11].n24 VGND 0.08843f
C13606 XThC.Tn[11].n25 VGND 0.14574f
C13607 XThC.Tn[11].t16 VGND 0.01608f
C13608 XThC.Tn[11].t42 VGND 0.01757f
C13609 XThC.Tn[11].n26 VGND 0.03922f
C13610 XThC.Tn[11].n27 VGND 0.02687f
C13611 XThC.Tn[11].n28 VGND 0.08843f
C13612 XThC.Tn[11].n29 VGND 0.14574f
C13613 XThC.Tn[11].t23 VGND 0.01608f
C13614 XThC.Tn[11].t19 VGND 0.01757f
C13615 XThC.Tn[11].n30 VGND 0.03922f
C13616 XThC.Tn[11].n31 VGND 0.02687f
C13617 XThC.Tn[11].n32 VGND 0.08843f
C13618 XThC.Tn[11].n33 VGND 0.14574f
C13619 XThC.Tn[11].t25 VGND 0.01608f
C13620 XThC.Tn[11].t21 VGND 0.01757f
C13621 XThC.Tn[11].n34 VGND 0.03922f
C13622 XThC.Tn[11].n35 VGND 0.02687f
C13623 XThC.Tn[11].n36 VGND 0.08843f
C13624 XThC.Tn[11].n37 VGND 0.14574f
C13625 XThC.Tn[11].t13 VGND 0.01608f
C13626 XThC.Tn[11].t40 VGND 0.01757f
C13627 XThC.Tn[11].n38 VGND 0.03922f
C13628 XThC.Tn[11].n39 VGND 0.02687f
C13629 XThC.Tn[11].n40 VGND 0.08843f
C13630 XThC.Tn[11].n41 VGND 0.14574f
C13631 XThC.Tn[11].t15 VGND 0.01608f
C13632 XThC.Tn[11].t41 VGND 0.01757f
C13633 XThC.Tn[11].n42 VGND 0.03922f
C13634 XThC.Tn[11].n43 VGND 0.02687f
C13635 XThC.Tn[11].n44 VGND 0.08843f
C13636 XThC.Tn[11].n45 VGND 0.14574f
C13637 XThC.Tn[11].t26 VGND 0.01608f
C13638 XThC.Tn[11].t22 VGND 0.01757f
C13639 XThC.Tn[11].n46 VGND 0.03922f
C13640 XThC.Tn[11].n47 VGND 0.02687f
C13641 XThC.Tn[11].n48 VGND 0.08843f
C13642 XThC.Tn[11].n49 VGND 0.14574f
C13643 XThC.Tn[11].t34 VGND 0.01608f
C13644 XThC.Tn[11].t30 VGND 0.01757f
C13645 XThC.Tn[11].n50 VGND 0.03922f
C13646 XThC.Tn[11].n51 VGND 0.02687f
C13647 XThC.Tn[11].n52 VGND 0.08843f
C13648 XThC.Tn[11].n53 VGND 0.14574f
C13649 XThC.Tn[11].t36 VGND 0.01608f
C13650 XThC.Tn[11].t33 VGND 0.01757f
C13651 XThC.Tn[11].n54 VGND 0.03922f
C13652 XThC.Tn[11].n55 VGND 0.02687f
C13653 XThC.Tn[11].n56 VGND 0.08843f
C13654 XThC.Tn[11].n57 VGND 0.14574f
C13655 XThC.Tn[11].t17 VGND 0.01608f
C13656 XThC.Tn[11].t14 VGND 0.01757f
C13657 XThC.Tn[11].n58 VGND 0.03922f
C13658 XThC.Tn[11].n59 VGND 0.02687f
C13659 XThC.Tn[11].n60 VGND 0.08843f
C13660 XThC.Tn[11].n61 VGND 0.14574f
C13661 XThC.Tn[11].t27 VGND 0.01608f
C13662 XThC.Tn[11].t24 VGND 0.01757f
C13663 XThC.Tn[11].n62 VGND 0.03922f
C13664 XThC.Tn[11].n63 VGND 0.02687f
C13665 XThC.Tn[11].n64 VGND 0.08843f
C13666 XThC.Tn[11].n65 VGND 0.14574f
C13667 XThC.Tn[11].n66 VGND 0.6764f
C13668 XThC.Tn[11].n67 VGND 0.26496f
C13669 XThC.Tn[11].t4 VGND 0.02029f
C13670 XThC.Tn[11].t1 VGND 0.02029f
C13671 XThC.Tn[11].n68 VGND 0.04384f
C13672 XThC.Tn[11].t6 VGND 0.02029f
C13673 XThC.Tn[11].t0 VGND 0.02029f
C13674 XThC.Tn[11].n69 VGND 0.06911f
C13675 XThC.Tn[11].n70 VGND 0.18303f
C13676 XThC.Tn[11].n71 VGND 0.01348f
C13677 XThC.Tn[11].t7 VGND 0.02029f
C13678 XThC.Tn[11].t10 VGND 0.02029f
C13679 XThC.Tn[11].n72 VGND 0.06161f
C13680 XThC.Tn[11].t9 VGND 0.02029f
C13681 XThC.Tn[11].t8 VGND 0.02029f
C13682 XThC.Tn[11].n73 VGND 0.04511f
C13683 XThC.Tn[11].n74 VGND 0.20076f
C13684 XThC.Tn[9].t4 VGND 0.02f
C13685 XThC.Tn[9].t7 VGND 0.02f
C13686 XThC.Tn[9].n0 VGND 0.04321f
C13687 XThC.Tn[9].t6 VGND 0.02f
C13688 XThC.Tn[9].t5 VGND 0.02f
C13689 XThC.Tn[9].n1 VGND 0.06812f
C13690 XThC.Tn[9].n2 VGND 0.1804f
C13691 XThC.Tn[9].t9 VGND 0.02f
C13692 XThC.Tn[9].t8 VGND 0.02f
C13693 XThC.Tn[9].n3 VGND 0.06073f
C13694 XThC.Tn[9].t11 VGND 0.02f
C13695 XThC.Tn[9].t10 VGND 0.02f
C13696 XThC.Tn[9].n4 VGND 0.04446f
C13697 XThC.Tn[9].n5 VGND 0.19787f
C13698 XThC.Tn[9].n6 VGND 0.01328f
C13699 XThC.Tn[9].t26 VGND 0.01585f
C13700 XThC.Tn[9].t12 VGND 0.01732f
C13701 XThC.Tn[9].n7 VGND 0.03865f
C13702 XThC.Tn[9].n8 VGND 0.02648f
C13703 XThC.Tn[9].n9 VGND 0.08692f
C13704 XThC.Tn[9].t13 VGND 0.01585f
C13705 XThC.Tn[9].t30 VGND 0.01732f
C13706 XThC.Tn[9].n10 VGND 0.03865f
C13707 XThC.Tn[9].n11 VGND 0.02648f
C13708 XThC.Tn[9].n12 VGND 0.08716f
C13709 XThC.Tn[9].n13 VGND 0.14365f
C13710 XThC.Tn[9].t15 VGND 0.01585f
C13711 XThC.Tn[9].t34 VGND 0.01732f
C13712 XThC.Tn[9].n14 VGND 0.03865f
C13713 XThC.Tn[9].n15 VGND 0.02648f
C13714 XThC.Tn[9].n16 VGND 0.08716f
C13715 XThC.Tn[9].n17 VGND 0.14365f
C13716 XThC.Tn[9].t17 VGND 0.01585f
C13717 XThC.Tn[9].t35 VGND 0.01732f
C13718 XThC.Tn[9].n18 VGND 0.03865f
C13719 XThC.Tn[9].n19 VGND 0.02648f
C13720 XThC.Tn[9].n20 VGND 0.08716f
C13721 XThC.Tn[9].n21 VGND 0.14365f
C13722 XThC.Tn[9].t39 VGND 0.01585f
C13723 XThC.Tn[9].t24 VGND 0.01732f
C13724 XThC.Tn[9].n22 VGND 0.03865f
C13725 XThC.Tn[9].n23 VGND 0.02648f
C13726 XThC.Tn[9].n24 VGND 0.08716f
C13727 XThC.Tn[9].n25 VGND 0.14365f
C13728 XThC.Tn[9].t40 VGND 0.01585f
C13729 XThC.Tn[9].t25 VGND 0.01732f
C13730 XThC.Tn[9].n26 VGND 0.03865f
C13731 XThC.Tn[9].n27 VGND 0.02648f
C13732 XThC.Tn[9].n28 VGND 0.08716f
C13733 XThC.Tn[9].n29 VGND 0.14365f
C13734 XThC.Tn[9].t22 VGND 0.01585f
C13735 XThC.Tn[9].t38 VGND 0.01732f
C13736 XThC.Tn[9].n30 VGND 0.03865f
C13737 XThC.Tn[9].n31 VGND 0.02648f
C13738 XThC.Tn[9].n32 VGND 0.08716f
C13739 XThC.Tn[9].n33 VGND 0.14365f
C13740 XThC.Tn[9].t28 VGND 0.01585f
C13741 XThC.Tn[9].t14 VGND 0.01732f
C13742 XThC.Tn[9].n34 VGND 0.03865f
C13743 XThC.Tn[9].n35 VGND 0.02648f
C13744 XThC.Tn[9].n36 VGND 0.08716f
C13745 XThC.Tn[9].n37 VGND 0.14365f
C13746 XThC.Tn[9].t31 VGND 0.01585f
C13747 XThC.Tn[9].t16 VGND 0.01732f
C13748 XThC.Tn[9].n38 VGND 0.03865f
C13749 XThC.Tn[9].n39 VGND 0.02648f
C13750 XThC.Tn[9].n40 VGND 0.08716f
C13751 XThC.Tn[9].n41 VGND 0.14365f
C13752 XThC.Tn[9].t19 VGND 0.01585f
C13753 XThC.Tn[9].t36 VGND 0.01732f
C13754 XThC.Tn[9].n42 VGND 0.03865f
C13755 XThC.Tn[9].n43 VGND 0.02648f
C13756 XThC.Tn[9].n44 VGND 0.08716f
C13757 XThC.Tn[9].n45 VGND 0.14365f
C13758 XThC.Tn[9].t21 VGND 0.01585f
C13759 XThC.Tn[9].t37 VGND 0.01732f
C13760 XThC.Tn[9].n46 VGND 0.03865f
C13761 XThC.Tn[9].n47 VGND 0.02648f
C13762 XThC.Tn[9].n48 VGND 0.08716f
C13763 XThC.Tn[9].n49 VGND 0.14365f
C13764 XThC.Tn[9].t32 VGND 0.01585f
C13765 XThC.Tn[9].t18 VGND 0.01732f
C13766 XThC.Tn[9].n50 VGND 0.03865f
C13767 XThC.Tn[9].n51 VGND 0.02648f
C13768 XThC.Tn[9].n52 VGND 0.08716f
C13769 XThC.Tn[9].n53 VGND 0.14365f
C13770 XThC.Tn[9].t42 VGND 0.01585f
C13771 XThC.Tn[9].t27 VGND 0.01732f
C13772 XThC.Tn[9].n54 VGND 0.03865f
C13773 XThC.Tn[9].n55 VGND 0.02648f
C13774 XThC.Tn[9].n56 VGND 0.08716f
C13775 XThC.Tn[9].n57 VGND 0.14365f
C13776 XThC.Tn[9].t43 VGND 0.01585f
C13777 XThC.Tn[9].t29 VGND 0.01732f
C13778 XThC.Tn[9].n58 VGND 0.03865f
C13779 XThC.Tn[9].n59 VGND 0.02648f
C13780 XThC.Tn[9].n60 VGND 0.08716f
C13781 XThC.Tn[9].n61 VGND 0.14365f
C13782 XThC.Tn[9].t23 VGND 0.01585f
C13783 XThC.Tn[9].t41 VGND 0.01732f
C13784 XThC.Tn[9].n62 VGND 0.03865f
C13785 XThC.Tn[9].n63 VGND 0.02648f
C13786 XThC.Tn[9].n64 VGND 0.08716f
C13787 XThC.Tn[9].n65 VGND 0.14365f
C13788 XThC.Tn[9].t33 VGND 0.01585f
C13789 XThC.Tn[9].t20 VGND 0.01732f
C13790 XThC.Tn[9].n66 VGND 0.03865f
C13791 XThC.Tn[9].n67 VGND 0.02648f
C13792 XThC.Tn[9].n68 VGND 0.08716f
C13793 XThC.Tn[9].n69 VGND 0.14365f
C13794 XThC.Tn[9].n70 VGND 0.61747f
C13795 XThC.Tn[9].n71 VGND 0.26115f
C13796 XThC.Tn[9].t1 VGND 0.013f
C13797 XThC.Tn[9].t0 VGND 0.013f
C13798 XThC.Tn[9].n72 VGND 0.03242f
C13799 XThC.Tn[9].t2 VGND 0.013f
C13800 XThC.Tn[9].t3 VGND 0.013f
C13801 XThC.Tn[9].n73 VGND 0.026f
C13802 XThC.Tn[9].n74 VGND 0.05995f
C13803 XThC.Tn[5].t7 VGND 0.01807f
C13804 XThC.Tn[5].t6 VGND 0.01807f
C13805 XThC.Tn[5].n0 VGND 0.03647f
C13806 XThC.Tn[5].t5 VGND 0.01807f
C13807 XThC.Tn[5].t4 VGND 0.01807f
C13808 XThC.Tn[5].n1 VGND 0.04267f
C13809 XThC.Tn[5].n2 VGND 0.12799f
C13810 XThC.Tn[5].t9 VGND 0.01174f
C13811 XThC.Tn[5].t8 VGND 0.01174f
C13812 XThC.Tn[5].n3 VGND 0.02674f
C13813 XThC.Tn[5].t11 VGND 0.01174f
C13814 XThC.Tn[5].t10 VGND 0.01174f
C13815 XThC.Tn[5].n4 VGND 0.02674f
C13816 XThC.Tn[5].t2 VGND 0.01174f
C13817 XThC.Tn[5].t1 VGND 0.01174f
C13818 XThC.Tn[5].n5 VGND 0.02674f
C13819 XThC.Tn[5].t0 VGND 0.01174f
C13820 XThC.Tn[5].t3 VGND 0.01174f
C13821 XThC.Tn[5].n6 VGND 0.04456f
C13822 XThC.Tn[5].n7 VGND 0.12735f
C13823 XThC.Tn[5].n8 VGND 0.07873f
C13824 XThC.Tn[5].n9 VGND 0.08885f
C13825 XThC.Tn[5].t15 VGND 0.01432f
C13826 XThC.Tn[5].t33 VGND 0.01564f
C13827 XThC.Tn[5].n10 VGND 0.03492f
C13828 XThC.Tn[5].n11 VGND 0.02392f
C13829 XThC.Tn[5].n12 VGND 0.07852f
C13830 XThC.Tn[5].t34 VGND 0.01432f
C13831 XThC.Tn[5].t19 VGND 0.01564f
C13832 XThC.Tn[5].n13 VGND 0.03492f
C13833 XThC.Tn[5].n14 VGND 0.02392f
C13834 XThC.Tn[5].n15 VGND 0.07873f
C13835 XThC.Tn[5].n16 VGND 0.12976f
C13836 XThC.Tn[5].t36 VGND 0.01432f
C13837 XThC.Tn[5].t23 VGND 0.01564f
C13838 XThC.Tn[5].n17 VGND 0.03492f
C13839 XThC.Tn[5].n18 VGND 0.02392f
C13840 XThC.Tn[5].n19 VGND 0.07873f
C13841 XThC.Tn[5].n20 VGND 0.12976f
C13842 XThC.Tn[5].t38 VGND 0.01432f
C13843 XThC.Tn[5].t24 VGND 0.01564f
C13844 XThC.Tn[5].n21 VGND 0.03492f
C13845 XThC.Tn[5].n22 VGND 0.02392f
C13846 XThC.Tn[5].n23 VGND 0.07873f
C13847 XThC.Tn[5].n24 VGND 0.12976f
C13848 XThC.Tn[5].t28 VGND 0.01432f
C13849 XThC.Tn[5].t13 VGND 0.01564f
C13850 XThC.Tn[5].n25 VGND 0.03492f
C13851 XThC.Tn[5].n26 VGND 0.02392f
C13852 XThC.Tn[5].n27 VGND 0.07873f
C13853 XThC.Tn[5].n28 VGND 0.12976f
C13854 XThC.Tn[5].t29 VGND 0.01432f
C13855 XThC.Tn[5].t14 VGND 0.01564f
C13856 XThC.Tn[5].n29 VGND 0.03492f
C13857 XThC.Tn[5].n30 VGND 0.02392f
C13858 XThC.Tn[5].n31 VGND 0.07873f
C13859 XThC.Tn[5].n32 VGND 0.12976f
C13860 XThC.Tn[5].t43 VGND 0.01432f
C13861 XThC.Tn[5].t27 VGND 0.01564f
C13862 XThC.Tn[5].n33 VGND 0.03492f
C13863 XThC.Tn[5].n34 VGND 0.02392f
C13864 XThC.Tn[5].n35 VGND 0.07873f
C13865 XThC.Tn[5].n36 VGND 0.12976f
C13866 XThC.Tn[5].t17 VGND 0.01432f
C13867 XThC.Tn[5].t35 VGND 0.01564f
C13868 XThC.Tn[5].n37 VGND 0.03492f
C13869 XThC.Tn[5].n38 VGND 0.02392f
C13870 XThC.Tn[5].n39 VGND 0.07873f
C13871 XThC.Tn[5].n40 VGND 0.12976f
C13872 XThC.Tn[5].t20 VGND 0.01432f
C13873 XThC.Tn[5].t37 VGND 0.01564f
C13874 XThC.Tn[5].n41 VGND 0.03492f
C13875 XThC.Tn[5].n42 VGND 0.02392f
C13876 XThC.Tn[5].n43 VGND 0.07873f
C13877 XThC.Tn[5].n44 VGND 0.12976f
C13878 XThC.Tn[5].t40 VGND 0.01432f
C13879 XThC.Tn[5].t25 VGND 0.01564f
C13880 XThC.Tn[5].n45 VGND 0.03492f
C13881 XThC.Tn[5].n46 VGND 0.02392f
C13882 XThC.Tn[5].n47 VGND 0.07873f
C13883 XThC.Tn[5].n48 VGND 0.12976f
C13884 XThC.Tn[5].t42 VGND 0.01432f
C13885 XThC.Tn[5].t26 VGND 0.01564f
C13886 XThC.Tn[5].n49 VGND 0.03492f
C13887 XThC.Tn[5].n50 VGND 0.02392f
C13888 XThC.Tn[5].n51 VGND 0.07873f
C13889 XThC.Tn[5].n52 VGND 0.12976f
C13890 XThC.Tn[5].t21 VGND 0.01432f
C13891 XThC.Tn[5].t39 VGND 0.01564f
C13892 XThC.Tn[5].n53 VGND 0.03492f
C13893 XThC.Tn[5].n54 VGND 0.02392f
C13894 XThC.Tn[5].n55 VGND 0.07873f
C13895 XThC.Tn[5].n56 VGND 0.12976f
C13896 XThC.Tn[5].t31 VGND 0.01432f
C13897 XThC.Tn[5].t16 VGND 0.01564f
C13898 XThC.Tn[5].n57 VGND 0.03492f
C13899 XThC.Tn[5].n58 VGND 0.02392f
C13900 XThC.Tn[5].n59 VGND 0.07873f
C13901 XThC.Tn[5].n60 VGND 0.12976f
C13902 XThC.Tn[5].t32 VGND 0.01432f
C13903 XThC.Tn[5].t18 VGND 0.01564f
C13904 XThC.Tn[5].n61 VGND 0.03492f
C13905 XThC.Tn[5].n62 VGND 0.02392f
C13906 XThC.Tn[5].n63 VGND 0.07873f
C13907 XThC.Tn[5].n64 VGND 0.12976f
C13908 XThC.Tn[5].t12 VGND 0.01432f
C13909 XThC.Tn[5].t30 VGND 0.01564f
C13910 XThC.Tn[5].n65 VGND 0.03492f
C13911 XThC.Tn[5].n66 VGND 0.02392f
C13912 XThC.Tn[5].n67 VGND 0.07873f
C13913 XThC.Tn[5].n68 VGND 0.12976f
C13914 XThC.Tn[5].t22 VGND 0.01432f
C13915 XThC.Tn[5].t41 VGND 0.01564f
C13916 XThC.Tn[5].n69 VGND 0.03492f
C13917 XThC.Tn[5].n70 VGND 0.02392f
C13918 XThC.Tn[5].n71 VGND 0.07873f
C13919 XThC.Tn[5].n72 VGND 0.12976f
C13920 XThC.Tn[5].n73 VGND 0.14766f
C13921 XThR.Tn[9].t2 VGND 0.02425f
C13922 XThR.Tn[9].t0 VGND 0.02425f
C13923 XThR.Tn[9].n0 VGND 0.07362f
C13924 XThR.Tn[9].t3 VGND 0.02425f
C13925 XThR.Tn[9].t1 VGND 0.02425f
C13926 XThR.Tn[9].n1 VGND 0.0539f
C13927 XThR.Tn[9].n2 VGND 0.24507f
C13928 XThR.Tn[9].t5 VGND 0.01576f
C13929 XThR.Tn[9].t7 VGND 0.01576f
C13930 XThR.Tn[9].n3 VGND 0.03931f
C13931 XThR.Tn[9].t4 VGND 0.01576f
C13932 XThR.Tn[9].t6 VGND 0.01576f
C13933 XThR.Tn[9].n4 VGND 0.03152f
C13934 XThR.Tn[9].n5 VGND 0.07929f
C13935 XThR.Tn[9].t17 VGND 0.01895f
C13936 XThR.Tn[9].t71 VGND 0.02075f
C13937 XThR.Tn[9].n6 VGND 0.05067f
C13938 XThR.Tn[9].n7 VGND 0.09733f
C13939 XThR.Tn[9].t35 VGND 0.01895f
C13940 XThR.Tn[9].t28 VGND 0.02075f
C13941 XThR.Tn[9].n8 VGND 0.05067f
C13942 XThR.Tn[9].t50 VGND 0.01889f
C13943 XThR.Tn[9].t19 VGND 0.02068f
C13944 XThR.Tn[9].n9 VGND 0.05272f
C13945 XThR.Tn[9].n10 VGND 0.03704f
C13946 XThR.Tn[9].n11 VGND 0.00677f
C13947 XThR.Tn[9].n12 VGND 0.11885f
C13948 XThR.Tn[9].t72 VGND 0.01895f
C13949 XThR.Tn[9].t64 VGND 0.02075f
C13950 XThR.Tn[9].n13 VGND 0.05067f
C13951 XThR.Tn[9].t26 VGND 0.01889f
C13952 XThR.Tn[9].t59 VGND 0.02068f
C13953 XThR.Tn[9].n14 VGND 0.05272f
C13954 XThR.Tn[9].n15 VGND 0.03704f
C13955 XThR.Tn[9].n16 VGND 0.00677f
C13956 XThR.Tn[9].n17 VGND 0.11885f
C13957 XThR.Tn[9].t29 VGND 0.01895f
C13958 XThR.Tn[9].t21 VGND 0.02075f
C13959 XThR.Tn[9].n18 VGND 0.05067f
C13960 XThR.Tn[9].t41 VGND 0.01889f
C13961 XThR.Tn[9].t15 VGND 0.02068f
C13962 XThR.Tn[9].n19 VGND 0.05272f
C13963 XThR.Tn[9].n20 VGND 0.03704f
C13964 XThR.Tn[9].n21 VGND 0.00677f
C13965 XThR.Tn[9].n22 VGND 0.11885f
C13966 XThR.Tn[9].t56 VGND 0.01895f
C13967 XThR.Tn[9].t46 VGND 0.02075f
C13968 XThR.Tn[9].n23 VGND 0.05067f
C13969 XThR.Tn[9].t73 VGND 0.01889f
C13970 XThR.Tn[9].t42 VGND 0.02068f
C13971 XThR.Tn[9].n24 VGND 0.05272f
C13972 XThR.Tn[9].n25 VGND 0.03704f
C13973 XThR.Tn[9].n26 VGND 0.00677f
C13974 XThR.Tn[9].n27 VGND 0.11885f
C13975 XThR.Tn[9].t31 VGND 0.01895f
C13976 XThR.Tn[9].t23 VGND 0.02075f
C13977 XThR.Tn[9].n28 VGND 0.05067f
C13978 XThR.Tn[9].t44 VGND 0.01889f
C13979 XThR.Tn[9].t16 VGND 0.02068f
C13980 XThR.Tn[9].n29 VGND 0.05272f
C13981 XThR.Tn[9].n30 VGND 0.03704f
C13982 XThR.Tn[9].n31 VGND 0.00677f
C13983 XThR.Tn[9].n32 VGND 0.11885f
C13984 XThR.Tn[9].t67 VGND 0.01895f
C13985 XThR.Tn[9].t37 VGND 0.02075f
C13986 XThR.Tn[9].n33 VGND 0.05067f
C13987 XThR.Tn[9].t20 VGND 0.01889f
C13988 XThR.Tn[9].t33 VGND 0.02068f
C13989 XThR.Tn[9].n34 VGND 0.05272f
C13990 XThR.Tn[9].n35 VGND 0.03704f
C13991 XThR.Tn[9].n36 VGND 0.00677f
C13992 XThR.Tn[9].n37 VGND 0.11885f
C13993 XThR.Tn[9].t36 VGND 0.01895f
C13994 XThR.Tn[9].t32 VGND 0.02075f
C13995 XThR.Tn[9].n38 VGND 0.05067f
C13996 XThR.Tn[9].t51 VGND 0.01889f
C13997 XThR.Tn[9].t25 VGND 0.02068f
C13998 XThR.Tn[9].n39 VGND 0.05272f
C13999 XThR.Tn[9].n40 VGND 0.03704f
C14000 XThR.Tn[9].n41 VGND 0.00677f
C14001 XThR.Tn[9].n42 VGND 0.11885f
C14002 XThR.Tn[9].t39 VGND 0.01895f
C14003 XThR.Tn[9].t45 VGND 0.02075f
C14004 XThR.Tn[9].n43 VGND 0.05067f
C14005 XThR.Tn[9].t55 VGND 0.01889f
C14006 XThR.Tn[9].t40 VGND 0.02068f
C14007 XThR.Tn[9].n44 VGND 0.05272f
C14008 XThR.Tn[9].n45 VGND 0.03704f
C14009 XThR.Tn[9].n46 VGND 0.00677f
C14010 XThR.Tn[9].n47 VGND 0.11885f
C14011 XThR.Tn[9].t58 VGND 0.01895f
C14012 XThR.Tn[9].t66 VGND 0.02075f
C14013 XThR.Tn[9].n48 VGND 0.05067f
C14014 XThR.Tn[9].t13 VGND 0.01889f
C14015 XThR.Tn[9].t60 VGND 0.02068f
C14016 XThR.Tn[9].n49 VGND 0.05272f
C14017 XThR.Tn[9].n50 VGND 0.03704f
C14018 XThR.Tn[9].n51 VGND 0.00677f
C14019 XThR.Tn[9].n52 VGND 0.11885f
C14020 XThR.Tn[9].t48 VGND 0.01895f
C14021 XThR.Tn[9].t24 VGND 0.02075f
C14022 XThR.Tn[9].n53 VGND 0.05067f
C14023 XThR.Tn[9].t65 VGND 0.01889f
C14024 XThR.Tn[9].t18 VGND 0.02068f
C14025 XThR.Tn[9].n54 VGND 0.05272f
C14026 XThR.Tn[9].n55 VGND 0.03704f
C14027 XThR.Tn[9].n56 VGND 0.00677f
C14028 XThR.Tn[9].n57 VGND 0.11885f
C14029 XThR.Tn[9].t70 VGND 0.01895f
C14030 XThR.Tn[9].t62 VGND 0.02075f
C14031 XThR.Tn[9].n58 VGND 0.05067f
C14032 XThR.Tn[9].t22 VGND 0.01889f
C14033 XThR.Tn[9].t52 VGND 0.02068f
C14034 XThR.Tn[9].n59 VGND 0.05272f
C14035 XThR.Tn[9].n60 VGND 0.03704f
C14036 XThR.Tn[9].n61 VGND 0.00677f
C14037 XThR.Tn[9].n62 VGND 0.11885f
C14038 XThR.Tn[9].t38 VGND 0.01895f
C14039 XThR.Tn[9].t34 VGND 0.02075f
C14040 XThR.Tn[9].n63 VGND 0.05067f
C14041 XThR.Tn[9].t53 VGND 0.01889f
C14042 XThR.Tn[9].t27 VGND 0.02068f
C14043 XThR.Tn[9].n64 VGND 0.05272f
C14044 XThR.Tn[9].n65 VGND 0.03704f
C14045 XThR.Tn[9].n66 VGND 0.00677f
C14046 XThR.Tn[9].n67 VGND 0.11885f
C14047 XThR.Tn[9].t57 VGND 0.01895f
C14048 XThR.Tn[9].t47 VGND 0.02075f
C14049 XThR.Tn[9].n68 VGND 0.05067f
C14050 XThR.Tn[9].t12 VGND 0.01889f
C14051 XThR.Tn[9].t43 VGND 0.02068f
C14052 XThR.Tn[9].n69 VGND 0.05272f
C14053 XThR.Tn[9].n70 VGND 0.03704f
C14054 XThR.Tn[9].n71 VGND 0.00677f
C14055 XThR.Tn[9].n72 VGND 0.11885f
C14056 XThR.Tn[9].t14 VGND 0.01895f
C14057 XThR.Tn[9].t69 VGND 0.02075f
C14058 XThR.Tn[9].n73 VGND 0.05067f
C14059 XThR.Tn[9].t30 VGND 0.01889f
C14060 XThR.Tn[9].t61 VGND 0.02068f
C14061 XThR.Tn[9].n74 VGND 0.05272f
C14062 XThR.Tn[9].n75 VGND 0.03704f
C14063 XThR.Tn[9].n76 VGND 0.00677f
C14064 XThR.Tn[9].n77 VGND 0.11885f
C14065 XThR.Tn[9].t49 VGND 0.01895f
C14066 XThR.Tn[9].t63 VGND 0.02075f
C14067 XThR.Tn[9].n78 VGND 0.05067f
C14068 XThR.Tn[9].t68 VGND 0.01889f
C14069 XThR.Tn[9].t54 VGND 0.02068f
C14070 XThR.Tn[9].n79 VGND 0.05272f
C14071 XThR.Tn[9].n80 VGND 0.03704f
C14072 XThR.Tn[9].n81 VGND 0.00677f
C14073 XThR.Tn[9].n82 VGND 0.11885f
C14074 XThR.Tn[9].n83 VGND 0.10801f
C14075 XThR.Tn[9].n84 VGND 0.35039f
C14076 XThR.Tn[9].t10 VGND 0.02425f
C14077 XThR.Tn[9].t8 VGND 0.02425f
C14078 XThR.Tn[9].n85 VGND 0.05239f
C14079 XThR.Tn[9].t11 VGND 0.02425f
C14080 XThR.Tn[9].t9 VGND 0.02425f
C14081 XThR.Tn[9].n86 VGND 0.07973f
C14082 XThR.Tn[9].n87 VGND 0.22139f
C14083 XThR.Tn[9].n88 VGND 0.02964f
C14084 XThC.Tn[6].t7 VGND 0.0182f
C14085 XThC.Tn[6].t6 VGND 0.0182f
C14086 XThC.Tn[6].n0 VGND 0.03674f
C14087 XThC.Tn[6].t5 VGND 0.0182f
C14088 XThC.Tn[6].t4 VGND 0.0182f
C14089 XThC.Tn[6].n1 VGND 0.04298f
C14090 XThC.Tn[6].n2 VGND 0.12033f
C14091 XThC.Tn[6].t8 VGND 0.01183f
C14092 XThC.Tn[6].t11 VGND 0.01183f
C14093 XThC.Tn[6].n3 VGND 0.02694f
C14094 XThC.Tn[6].t10 VGND 0.01183f
C14095 XThC.Tn[6].t9 VGND 0.01183f
C14096 XThC.Tn[6].n4 VGND 0.02694f
C14097 XThC.Tn[6].t1 VGND 0.01183f
C14098 XThC.Tn[6].t0 VGND 0.01183f
C14099 XThC.Tn[6].n5 VGND 0.02694f
C14100 XThC.Tn[6].t3 VGND 0.01183f
C14101 XThC.Tn[6].t2 VGND 0.01183f
C14102 XThC.Tn[6].n6 VGND 0.04489f
C14103 XThC.Tn[6].n7 VGND 0.12829f
C14104 XThC.Tn[6].n8 VGND 0.07931f
C14105 XThC.Tn[6].n9 VGND 0.0895f
C14106 XThC.Tn[6].t23 VGND 0.01443f
C14107 XThC.Tn[6].t26 VGND 0.01576f
C14108 XThC.Tn[6].n10 VGND 0.03517f
C14109 XThC.Tn[6].n11 VGND 0.0241f
C14110 XThC.Tn[6].n12 VGND 0.0791f
C14111 XThC.Tn[6].t40 VGND 0.01443f
C14112 XThC.Tn[6].t13 VGND 0.01576f
C14113 XThC.Tn[6].n13 VGND 0.03517f
C14114 XThC.Tn[6].n14 VGND 0.0241f
C14115 XThC.Tn[6].n15 VGND 0.07932f
C14116 XThC.Tn[6].n16 VGND 0.13072f
C14117 XThC.Tn[6].t42 VGND 0.01443f
C14118 XThC.Tn[6].t17 VGND 0.01576f
C14119 XThC.Tn[6].n17 VGND 0.03517f
C14120 XThC.Tn[6].n18 VGND 0.0241f
C14121 XThC.Tn[6].n19 VGND 0.07932f
C14122 XThC.Tn[6].n20 VGND 0.13072f
C14123 XThC.Tn[6].t12 VGND 0.01443f
C14124 XThC.Tn[6].t18 VGND 0.01576f
C14125 XThC.Tn[6].n21 VGND 0.03517f
C14126 XThC.Tn[6].n22 VGND 0.0241f
C14127 XThC.Tn[6].n23 VGND 0.07932f
C14128 XThC.Tn[6].n24 VGND 0.13072f
C14129 XThC.Tn[6].t33 VGND 0.01443f
C14130 XThC.Tn[6].t37 VGND 0.01576f
C14131 XThC.Tn[6].n25 VGND 0.03517f
C14132 XThC.Tn[6].n26 VGND 0.0241f
C14133 XThC.Tn[6].n27 VGND 0.07932f
C14134 XThC.Tn[6].n28 VGND 0.13072f
C14135 XThC.Tn[6].t35 VGND 0.01443f
C14136 XThC.Tn[6].t38 VGND 0.01576f
C14137 XThC.Tn[6].n29 VGND 0.03517f
C14138 XThC.Tn[6].n30 VGND 0.0241f
C14139 XThC.Tn[6].n31 VGND 0.07932f
C14140 XThC.Tn[6].n32 VGND 0.13072f
C14141 XThC.Tn[6].t16 VGND 0.01443f
C14142 XThC.Tn[6].t22 VGND 0.01576f
C14143 XThC.Tn[6].n33 VGND 0.03517f
C14144 XThC.Tn[6].n34 VGND 0.0241f
C14145 XThC.Tn[6].n35 VGND 0.07932f
C14146 XThC.Tn[6].n36 VGND 0.13072f
C14147 XThC.Tn[6].t25 VGND 0.01443f
C14148 XThC.Tn[6].t29 VGND 0.01576f
C14149 XThC.Tn[6].n37 VGND 0.03517f
C14150 XThC.Tn[6].n38 VGND 0.0241f
C14151 XThC.Tn[6].n39 VGND 0.07932f
C14152 XThC.Tn[6].n40 VGND 0.13072f
C14153 XThC.Tn[6].t27 VGND 0.01443f
C14154 XThC.Tn[6].t31 VGND 0.01576f
C14155 XThC.Tn[6].n41 VGND 0.03517f
C14156 XThC.Tn[6].n42 VGND 0.0241f
C14157 XThC.Tn[6].n43 VGND 0.07932f
C14158 XThC.Tn[6].n44 VGND 0.13072f
C14159 XThC.Tn[6].t14 VGND 0.01443f
C14160 XThC.Tn[6].t19 VGND 0.01576f
C14161 XThC.Tn[6].n45 VGND 0.03517f
C14162 XThC.Tn[6].n46 VGND 0.0241f
C14163 XThC.Tn[6].n47 VGND 0.07932f
C14164 XThC.Tn[6].n48 VGND 0.13072f
C14165 XThC.Tn[6].t15 VGND 0.01443f
C14166 XThC.Tn[6].t21 VGND 0.01576f
C14167 XThC.Tn[6].n49 VGND 0.03517f
C14168 XThC.Tn[6].n50 VGND 0.0241f
C14169 XThC.Tn[6].n51 VGND 0.07932f
C14170 XThC.Tn[6].n52 VGND 0.13072f
C14171 XThC.Tn[6].t28 VGND 0.01443f
C14172 XThC.Tn[6].t32 VGND 0.01576f
C14173 XThC.Tn[6].n53 VGND 0.03517f
C14174 XThC.Tn[6].n54 VGND 0.0241f
C14175 XThC.Tn[6].n55 VGND 0.07932f
C14176 XThC.Tn[6].n56 VGND 0.13072f
C14177 XThC.Tn[6].t36 VGND 0.01443f
C14178 XThC.Tn[6].t41 VGND 0.01576f
C14179 XThC.Tn[6].n57 VGND 0.03517f
C14180 XThC.Tn[6].n58 VGND 0.0241f
C14181 XThC.Tn[6].n59 VGND 0.07932f
C14182 XThC.Tn[6].n60 VGND 0.13072f
C14183 XThC.Tn[6].t39 VGND 0.01443f
C14184 XThC.Tn[6].t43 VGND 0.01576f
C14185 XThC.Tn[6].n61 VGND 0.03517f
C14186 XThC.Tn[6].n62 VGND 0.0241f
C14187 XThC.Tn[6].n63 VGND 0.07932f
C14188 XThC.Tn[6].n64 VGND 0.13072f
C14189 XThC.Tn[6].t20 VGND 0.01443f
C14190 XThC.Tn[6].t24 VGND 0.01576f
C14191 XThC.Tn[6].n65 VGND 0.03517f
C14192 XThC.Tn[6].n66 VGND 0.0241f
C14193 XThC.Tn[6].n67 VGND 0.07932f
C14194 XThC.Tn[6].n68 VGND 0.13072f
C14195 XThC.Tn[6].t30 VGND 0.01443f
C14196 XThC.Tn[6].t34 VGND 0.01576f
C14197 XThC.Tn[6].n69 VGND 0.03517f
C14198 XThC.Tn[6].n70 VGND 0.0241f
C14199 XThC.Tn[6].n71 VGND 0.07932f
C14200 XThC.Tn[6].n72 VGND 0.13072f
C14201 XThC.Tn[6].n73 VGND 0.14537f
C14202 XThC.Tn[6].n74 VGND 0.03808f
C14203 XThC.TBN.n0 VGND 0.01531f
C14204 XThC.TBN.t50 VGND 0.01024f
C14205 XThC.TBN.t118 VGND 0.00603f
C14206 XThC.TBN.t18 VGND 0.01024f
C14207 XThC.TBN.t83 VGND 0.00603f
C14208 XThC.TBN.n1 VGND 0.01477f
C14209 XThC.TBN.n2 VGND 0.00524f
C14210 XThC.TBN.t120 VGND 0.01024f
C14211 XThC.TBN.t71 VGND 0.00603f
C14212 XThC.TBN.t114 VGND 0.01024f
C14213 XThC.TBN.t62 VGND 0.00603f
C14214 XThC.TBN.n3 VGND 0.0138f
C14215 XThC.TBN.n4 VGND 0.00676f
C14216 XThC.TBN.n5 VGND 0.01477f
C14217 XThC.TBN.n6 VGND 0.00676f
C14218 XThC.TBN.n7 VGND 0.00548f
C14219 XThC.TBN.n8 VGND 0.00561f
C14220 XThC.TBN.n9 VGND 0.00676f
C14221 XThC.TBN.n10 VGND 0.02164f
C14222 XThC.TBN.n11 VGND 0.00584f
C14223 XThC.TBN.n12 VGND 0.00877f
C14224 XThC.TBN.t121 VGND 0.00603f
C14225 XThC.TBN.t79 VGND 0.01024f
C14226 XThC.TBN.t84 VGND 0.00603f
C14227 XThC.TBN.t36 VGND 0.01024f
C14228 XThC.TBN.n13 VGND 0.01477f
C14229 XThC.TBN.n14 VGND 0.00524f
C14230 XThC.TBN.t73 VGND 0.00603f
C14231 XThC.TBN.t26 VGND 0.01024f
C14232 XThC.TBN.t64 VGND 0.00603f
C14233 XThC.TBN.t21 VGND 0.01024f
C14234 XThC.TBN.n15 VGND 0.0138f
C14235 XThC.TBN.n16 VGND 0.00676f
C14236 XThC.TBN.n17 VGND 0.01477f
C14237 XThC.TBN.n18 VGND 0.00676f
C14238 XThC.TBN.n19 VGND 0.00548f
C14239 XThC.TBN.n20 VGND 0.00561f
C14240 XThC.TBN.n21 VGND 0.00676f
C14241 XThC.TBN.n22 VGND 0.02164f
C14242 XThC.TBN.n23 VGND 0.00584f
C14243 XThC.TBN.n24 VGND 0.00417f
C14244 XThC.TBN.n25 VGND 0.11789f
C14245 XThC.TBN.t106 VGND 0.01024f
C14246 XThC.TBN.t89 VGND 0.00603f
C14247 XThC.TBN.t70 VGND 0.01024f
C14248 XThC.TBN.t41 VGND 0.00603f
C14249 XThC.TBN.n26 VGND 0.01477f
C14250 XThC.TBN.n27 VGND 0.00524f
C14251 XThC.TBN.t56 VGND 0.01024f
C14252 XThC.TBN.t35 VGND 0.00603f
C14253 XThC.TBN.t48 VGND 0.01024f
C14254 XThC.TBN.t32 VGND 0.00603f
C14255 XThC.TBN.n28 VGND 0.0138f
C14256 XThC.TBN.n29 VGND 0.00676f
C14257 XThC.TBN.n30 VGND 0.01477f
C14258 XThC.TBN.n31 VGND 0.00676f
C14259 XThC.TBN.n32 VGND 0.00548f
C14260 XThC.TBN.n33 VGND 0.00561f
C14261 XThC.TBN.n34 VGND 0.00676f
C14262 XThC.TBN.n35 VGND 0.02164f
C14263 XThC.TBN.n36 VGND 0.00584f
C14264 XThC.TBN.n37 VGND 0.00417f
C14265 XThC.TBN.n38 VGND 0.07443f
C14266 XThC.TBN.t43 VGND 0.00603f
C14267 XThC.TBN.t39 VGND 0.01024f
C14268 XThC.TBN.t10 VGND 0.00603f
C14269 XThC.TBN.t122 VGND 0.01024f
C14270 XThC.TBN.n39 VGND 0.01477f
C14271 XThC.TBN.n40 VGND 0.00524f
C14272 XThC.TBN.t112 VGND 0.00603f
C14273 XThC.TBN.t109 VGND 0.01024f
C14274 XThC.TBN.t108 VGND 0.00603f
C14275 XThC.TBN.t102 VGND 0.01024f
C14276 XThC.TBN.n41 VGND 0.0138f
C14277 XThC.TBN.n42 VGND 0.00676f
C14278 XThC.TBN.n43 VGND 0.01477f
C14279 XThC.TBN.n44 VGND 0.00676f
C14280 XThC.TBN.n45 VGND 0.00548f
C14281 XThC.TBN.n46 VGND 0.00561f
C14282 XThC.TBN.n47 VGND 0.00676f
C14283 XThC.TBN.n48 VGND 0.02164f
C14284 XThC.TBN.n49 VGND 0.00584f
C14285 XThC.TBN.n50 VGND 0.00417f
C14286 XThC.TBN.n51 VGND 0.07443f
C14287 XThC.TBN.t47 VGND 0.01024f
C14288 XThC.TBN.t31 VGND 0.00603f
C14289 XThC.TBN.t17 VGND 0.01024f
C14290 XThC.TBN.t104 VGND 0.00603f
C14291 XThC.TBN.n52 VGND 0.01477f
C14292 XThC.TBN.n53 VGND 0.00524f
C14293 XThC.TBN.t116 VGND 0.01024f
C14294 XThC.TBN.t94 VGND 0.00603f
C14295 XThC.TBN.t111 VGND 0.01024f
C14296 XThC.TBN.t92 VGND 0.00603f
C14297 XThC.TBN.n54 VGND 0.0138f
C14298 XThC.TBN.n55 VGND 0.00676f
C14299 XThC.TBN.n56 VGND 0.01477f
C14300 XThC.TBN.n57 VGND 0.00676f
C14301 XThC.TBN.n58 VGND 0.00548f
C14302 XThC.TBN.n59 VGND 0.00561f
C14303 XThC.TBN.n60 VGND 0.00676f
C14304 XThC.TBN.n61 VGND 0.02164f
C14305 XThC.TBN.n62 VGND 0.00584f
C14306 XThC.TBN.n63 VGND 0.00417f
C14307 XThC.TBN.n64 VGND 0.07443f
C14308 XThC.TBN.t107 VGND 0.00603f
C14309 XThC.TBN.t101 VGND 0.01024f
C14310 XThC.TBN.t72 VGND 0.00603f
C14311 XThC.TBN.t63 VGND 0.01024f
C14312 XThC.TBN.n65 VGND 0.01477f
C14313 XThC.TBN.n66 VGND 0.00524f
C14314 XThC.TBN.t57 VGND 0.00603f
C14315 XThC.TBN.t52 VGND 0.01024f
C14316 XThC.TBN.t49 VGND 0.00603f
C14317 XThC.TBN.t44 VGND 0.01024f
C14318 XThC.TBN.n67 VGND 0.0138f
C14319 XThC.TBN.n68 VGND 0.00676f
C14320 XThC.TBN.n69 VGND 0.01477f
C14321 XThC.TBN.n70 VGND 0.00676f
C14322 XThC.TBN.n71 VGND 0.00548f
C14323 XThC.TBN.n72 VGND 0.00561f
C14324 XThC.TBN.n73 VGND 0.00676f
C14325 XThC.TBN.n74 VGND 0.02164f
C14326 XThC.TBN.n75 VGND 0.00584f
C14327 XThC.TBN.n76 VGND 0.00417f
C14328 XThC.TBN.n77 VGND 0.07443f
C14329 XThC.TBN.t25 VGND 0.01024f
C14330 XThC.TBN.t123 VGND 0.00603f
C14331 XThC.TBN.t100 VGND 0.01024f
C14332 XThC.TBN.t85 VGND 0.00603f
C14333 XThC.TBN.n78 VGND 0.01477f
C14334 XThC.TBN.n79 VGND 0.00524f
C14335 XThC.TBN.t93 VGND 0.01024f
C14336 XThC.TBN.t74 VGND 0.00603f
C14337 XThC.TBN.t90 VGND 0.01024f
C14338 XThC.TBN.t65 VGND 0.00603f
C14339 XThC.TBN.n80 VGND 0.0138f
C14340 XThC.TBN.n81 VGND 0.00676f
C14341 XThC.TBN.n82 VGND 0.01477f
C14342 XThC.TBN.n83 VGND 0.00676f
C14343 XThC.TBN.n84 VGND 0.00548f
C14344 XThC.TBN.n85 VGND 0.00561f
C14345 XThC.TBN.n86 VGND 0.00676f
C14346 XThC.TBN.n87 VGND 0.02164f
C14347 XThC.TBN.n88 VGND 0.00584f
C14348 XThC.TBN.n89 VGND 0.00417f
C14349 XThC.TBN.n90 VGND 0.06238f
C14350 XThC.TBN.n91 VGND 0.03511f
C14351 XThC.TBN.t46 VGND 0.01024f
C14352 XThC.TBN.t67 VGND 0.00603f
C14353 XThC.TBN.n92 VGND 0.00619f
C14354 XThC.TBN.t6 VGND 0.01024f
C14355 XThC.TBN.t24 VGND 0.00603f
C14356 XThC.TBN.n93 VGND 0.01243f
C14357 XThC.TBN.t12 VGND 0.01024f
C14358 XThC.TBN.t29 VGND 0.00603f
C14359 XThC.TBN.n94 VGND 0.01348f
C14360 XThC.TBN.n95 VGND 0.0076f
C14361 XThC.TBN.n96 VGND 0.01252f
C14362 XThC.TBN.n97 VGND 0.00434f
C14363 XThC.TBN.n98 VGND 0.00603f
C14364 XThC.TBN.n99 VGND 0.01348f
C14365 XThC.TBN.t54 VGND 0.01024f
C14366 XThC.TBN.t76 VGND 0.00603f
C14367 XThC.TBN.n100 VGND 0.01227f
C14368 XThC.TBN.n101 VGND 0.00676f
C14369 XThC.TBN.n102 VGND 0.01009f
C14370 XThC.TBN.t55 VGND 0.00603f
C14371 XThC.TBN.t38 VGND 0.01024f
C14372 XThC.TBN.n103 VGND 0.00619f
C14373 XThC.TBN.t16 VGND 0.00603f
C14374 XThC.TBN.t113 VGND 0.01024f
C14375 XThC.TBN.n104 VGND 0.01243f
C14376 XThC.TBN.t19 VGND 0.00603f
C14377 XThC.TBN.t119 VGND 0.01024f
C14378 XThC.TBN.n105 VGND 0.01348f
C14379 XThC.TBN.n106 VGND 0.0076f
C14380 XThC.TBN.n107 VGND 0.01252f
C14381 XThC.TBN.n108 VGND 0.00434f
C14382 XThC.TBN.n109 VGND 0.00603f
C14383 XThC.TBN.n110 VGND 0.01348f
C14384 XThC.TBN.t59 VGND 0.00603f
C14385 XThC.TBN.t42 VGND 0.01024f
C14386 XThC.TBN.n111 VGND 0.01227f
C14387 XThC.TBN.n112 VGND 0.00676f
C14388 XThC.TBN.n113 VGND 0.00747f
C14389 XThC.TBN.n114 VGND 0.11256f
C14390 XThC.TBN.t30 VGND 0.01024f
C14391 XThC.TBN.t8 VGND 0.00603f
C14392 XThC.TBN.n115 VGND 0.00619f
C14393 XThC.TBN.t98 VGND 0.01024f
C14394 XThC.TBN.t82 VGND 0.00603f
C14395 XThC.TBN.n116 VGND 0.01243f
C14396 XThC.TBN.t103 VGND 0.01024f
C14397 XThC.TBN.t87 VGND 0.00603f
C14398 XThC.TBN.n117 VGND 0.01348f
C14399 XThC.TBN.n118 VGND 0.0076f
C14400 XThC.TBN.n119 VGND 0.01252f
C14401 XThC.TBN.n120 VGND 0.00434f
C14402 XThC.TBN.n121 VGND 0.00603f
C14403 XThC.TBN.n122 VGND 0.01348f
C14404 XThC.TBN.t34 VGND 0.01024f
C14405 XThC.TBN.t15 VGND 0.00603f
C14406 XThC.TBN.n123 VGND 0.01227f
C14407 XThC.TBN.n124 VGND 0.00676f
C14408 XThC.TBN.n125 VGND 0.00747f
C14409 XThC.TBN.n126 VGND 0.07521f
C14410 XThC.TBN.t110 VGND 0.00603f
C14411 XThC.TBN.t96 VGND 0.01024f
C14412 XThC.TBN.n127 VGND 0.00619f
C14413 XThC.TBN.t68 VGND 0.00603f
C14414 XThC.TBN.t51 VGND 0.01024f
C14415 XThC.TBN.n128 VGND 0.01243f
C14416 XThC.TBN.t77 VGND 0.00603f
C14417 XThC.TBN.t58 VGND 0.01024f
C14418 XThC.TBN.n129 VGND 0.01348f
C14419 XThC.TBN.n130 VGND 0.0076f
C14420 XThC.TBN.n131 VGND 0.01252f
C14421 XThC.TBN.n132 VGND 0.00434f
C14422 XThC.TBN.n133 VGND 0.00603f
C14423 XThC.TBN.n134 VGND 0.01348f
C14424 XThC.TBN.t115 VGND 0.00603f
C14425 XThC.TBN.t99 VGND 0.01024f
C14426 XThC.TBN.n135 VGND 0.01227f
C14427 XThC.TBN.n136 VGND 0.00676f
C14428 XThC.TBN.n137 VGND 0.00747f
C14429 XThC.TBN.n138 VGND 0.07521f
C14430 XThC.TBN.t88 VGND 0.01024f
C14431 XThC.TBN.t60 VGND 0.00603f
C14432 XThC.TBN.n139 VGND 0.00619f
C14433 XThC.TBN.t37 VGND 0.01024f
C14434 XThC.TBN.t20 VGND 0.00603f
C14435 XThC.TBN.n140 VGND 0.01243f
C14436 XThC.TBN.t40 VGND 0.01024f
C14437 XThC.TBN.t22 VGND 0.00603f
C14438 XThC.TBN.n141 VGND 0.01348f
C14439 XThC.TBN.n142 VGND 0.0076f
C14440 XThC.TBN.n143 VGND 0.01252f
C14441 XThC.TBN.n144 VGND 0.00434f
C14442 XThC.TBN.n145 VGND 0.00603f
C14443 XThC.TBN.n146 VGND 0.01348f
C14444 XThC.TBN.t91 VGND 0.01024f
C14445 XThC.TBN.t66 VGND 0.00603f
C14446 XThC.TBN.n147 VGND 0.01227f
C14447 XThC.TBN.n148 VGND 0.00676f
C14448 XThC.TBN.n149 VGND 0.00747f
C14449 XThC.TBN.n150 VGND 0.07534f
C14450 XThC.TBN.t45 VGND 0.00603f
C14451 XThC.TBN.t7 VGND 0.01024f
C14452 XThC.TBN.n151 VGND 0.00619f
C14453 XThC.TBN.t5 VGND 0.00603f
C14454 XThC.TBN.t81 VGND 0.01024f
C14455 XThC.TBN.n152 VGND 0.01243f
C14456 XThC.TBN.t11 VGND 0.00603f
C14457 XThC.TBN.t86 VGND 0.01024f
C14458 XThC.TBN.n153 VGND 0.01348f
C14459 XThC.TBN.n154 VGND 0.0076f
C14460 XThC.TBN.n155 VGND 0.01252f
C14461 XThC.TBN.n156 VGND 0.00434f
C14462 XThC.TBN.n157 VGND 0.00603f
C14463 XThC.TBN.n158 VGND 0.01348f
C14464 XThC.TBN.t53 VGND 0.00603f
C14465 XThC.TBN.t13 VGND 0.01024f
C14466 XThC.TBN.n159 VGND 0.01227f
C14467 XThC.TBN.n160 VGND 0.00676f
C14468 XThC.TBN.n161 VGND 0.00747f
C14469 XThC.TBN.n162 VGND 0.07521f
C14470 XThC.TBN.t23 VGND 0.01024f
C14471 XThC.TBN.t117 VGND 0.00603f
C14472 XThC.TBN.n163 VGND 0.00619f
C14473 XThC.TBN.t95 VGND 0.01024f
C14474 XThC.TBN.t78 VGND 0.00603f
C14475 XThC.TBN.n164 VGND 0.01243f
C14476 XThC.TBN.t97 VGND 0.01024f
C14477 XThC.TBN.t80 VGND 0.00603f
C14478 XThC.TBN.n165 VGND 0.01348f
C14479 XThC.TBN.n166 VGND 0.0076f
C14480 XThC.TBN.n167 VGND 0.01252f
C14481 XThC.TBN.n168 VGND 0.00434f
C14482 XThC.TBN.n169 VGND 0.00603f
C14483 XThC.TBN.n170 VGND 0.01348f
C14484 XThC.TBN.t28 VGND 0.01024f
C14485 XThC.TBN.t4 VGND 0.00603f
C14486 XThC.TBN.n171 VGND 0.01227f
C14487 XThC.TBN.n172 VGND 0.00676f
C14488 XThC.TBN.n173 VGND 0.00747f
C14489 XThC.TBN.n174 VGND 0.08751f
C14490 XThC.TBN.n175 VGND 0.0808f
C14491 XThC.TBN.t105 VGND 0.00603f
C14492 XThC.TBN.t75 VGND 0.01024f
C14493 XThC.TBN.t69 VGND 0.00603f
C14494 XThC.TBN.t33 VGND 0.01024f
C14495 XThC.TBN.n176 VGND 0.01477f
C14496 XThC.TBN.t61 VGND 0.00603f
C14497 XThC.TBN.t27 VGND 0.01024f
C14498 XThC.TBN.n177 VGND 0.02293f
C14499 XThC.TBN.n178 VGND 0.00676f
C14500 XThC.TBN.n179 VGND 0.00561f
C14501 XThC.TBN.n180 VGND 0.00561f
C14502 XThC.TBN.n181 VGND 0.00676f
C14503 XThC.TBN.n182 VGND 0.01477f
C14504 XThC.TBN.t14 VGND 0.00603f
C14505 XThC.TBN.t9 VGND 0.01024f
C14506 XThC.TBN.n183 VGND 0.0138f
C14507 XThC.TBN.n184 VGND 0.00676f
C14508 XThC.TBN.n185 VGND 0.00372f
C14509 XThC.TBN.n186 VGND 0.00408f
C14510 XThC.TBN.n187 VGND 0.11129f
C14511 XThC.TBN.n188 VGND 0.02169f
C14512 XThC.TBN.t2 VGND 0.00658f
C14513 XThC.TBN.t3 VGND 0.00658f
C14514 XThC.TBN.n189 VGND 0.01513f
C14515 XThC.TBN.n190 VGND 0.0307f
C14516 XThC.TBN.n191 VGND 0.00526f
C14517 XThC.TBN.n192 VGND 0.00607f
C14518 XThC.TBN.t1 VGND 0.00428f
C14519 XThC.TBN.t0 VGND 0.00428f
C14520 XThC.TBN.n193 VGND 0.0094f
C14521 XThR.Tn[12].t11 VGND 0.02425f
C14522 XThR.Tn[12].t9 VGND 0.02425f
C14523 XThR.Tn[12].n0 VGND 0.07362f
C14524 XThR.Tn[12].t8 VGND 0.02425f
C14525 XThR.Tn[12].t10 VGND 0.02425f
C14526 XThR.Tn[12].n1 VGND 0.0539f
C14527 XThR.Tn[12].n2 VGND 0.24508f
C14528 XThR.Tn[12].t6 VGND 0.02425f
C14529 XThR.Tn[12].t4 VGND 0.02425f
C14530 XThR.Tn[12].n3 VGND 0.05239f
C14531 XThR.Tn[12].t7 VGND 0.02425f
C14532 XThR.Tn[12].t5 VGND 0.02425f
C14533 XThR.Tn[12].n4 VGND 0.07973f
C14534 XThR.Tn[12].n5 VGND 0.2214f
C14535 XThR.Tn[12].n6 VGND 0.01091f
C14536 XThR.Tn[12].t36 VGND 0.01895f
C14537 XThR.Tn[12].t28 VGND 0.02075f
C14538 XThR.Tn[12].n7 VGND 0.05067f
C14539 XThR.Tn[12].n8 VGND 0.09734f
C14540 XThR.Tn[12].t53 VGND 0.01895f
C14541 XThR.Tn[12].t43 VGND 0.02075f
C14542 XThR.Tn[12].n9 VGND 0.05067f
C14543 XThR.Tn[12].t71 VGND 0.01889f
C14544 XThR.Tn[12].t21 VGND 0.02068f
C14545 XThR.Tn[12].n10 VGND 0.05272f
C14546 XThR.Tn[12].n11 VGND 0.03704f
C14547 XThR.Tn[12].n12 VGND 0.00677f
C14548 XThR.Tn[12].n13 VGND 0.11886f
C14549 XThR.Tn[12].t30 VGND 0.01895f
C14550 XThR.Tn[12].t20 VGND 0.02075f
C14551 XThR.Tn[12].n14 VGND 0.05067f
C14552 XThR.Tn[12].t49 VGND 0.01889f
C14553 XThR.Tn[12].t60 VGND 0.02068f
C14554 XThR.Tn[12].n15 VGND 0.05272f
C14555 XThR.Tn[12].n16 VGND 0.03704f
C14556 XThR.Tn[12].n17 VGND 0.00677f
C14557 XThR.Tn[12].n18 VGND 0.11886f
C14558 XThR.Tn[12].t45 VGND 0.01895f
C14559 XThR.Tn[12].t38 VGND 0.02075f
C14560 XThR.Tn[12].n19 VGND 0.05067f
C14561 XThR.Tn[12].t63 VGND 0.01889f
C14562 XThR.Tn[12].t15 VGND 0.02068f
C14563 XThR.Tn[12].n20 VGND 0.05272f
C14564 XThR.Tn[12].n21 VGND 0.03704f
C14565 XThR.Tn[12].n22 VGND 0.00677f
C14566 XThR.Tn[12].n23 VGND 0.11886f
C14567 XThR.Tn[12].t70 VGND 0.01895f
C14568 XThR.Tn[12].t66 VGND 0.02075f
C14569 XThR.Tn[12].n24 VGND 0.05067f
C14570 XThR.Tn[12].t33 VGND 0.01889f
C14571 XThR.Tn[12].t46 VGND 0.02068f
C14572 XThR.Tn[12].n25 VGND 0.05272f
C14573 XThR.Tn[12].n26 VGND 0.03704f
C14574 XThR.Tn[12].n27 VGND 0.00677f
C14575 XThR.Tn[12].n28 VGND 0.11886f
C14576 XThR.Tn[12].t48 VGND 0.01895f
C14577 XThR.Tn[12].t39 VGND 0.02075f
C14578 XThR.Tn[12].n29 VGND 0.05067f
C14579 XThR.Tn[12].t64 VGND 0.01889f
C14580 XThR.Tn[12].t17 VGND 0.02068f
C14581 XThR.Tn[12].n30 VGND 0.05272f
C14582 XThR.Tn[12].n31 VGND 0.03704f
C14583 XThR.Tn[12].n32 VGND 0.00677f
C14584 XThR.Tn[12].n33 VGND 0.11886f
C14585 XThR.Tn[12].t23 VGND 0.01895f
C14586 XThR.Tn[12].t56 VGND 0.02075f
C14587 XThR.Tn[12].n34 VGND 0.05067f
C14588 XThR.Tn[12].t41 VGND 0.01889f
C14589 XThR.Tn[12].t37 VGND 0.02068f
C14590 XThR.Tn[12].n35 VGND 0.05272f
C14591 XThR.Tn[12].n36 VGND 0.03704f
C14592 XThR.Tn[12].n37 VGND 0.00677f
C14593 XThR.Tn[12].n38 VGND 0.11886f
C14594 XThR.Tn[12].t54 VGND 0.01895f
C14595 XThR.Tn[12].t51 VGND 0.02075f
C14596 XThR.Tn[12].n39 VGND 0.05067f
C14597 XThR.Tn[12].t72 VGND 0.01889f
C14598 XThR.Tn[12].t29 VGND 0.02068f
C14599 XThR.Tn[12].n40 VGND 0.05272f
C14600 XThR.Tn[12].n41 VGND 0.03704f
C14601 XThR.Tn[12].n42 VGND 0.00677f
C14602 XThR.Tn[12].n43 VGND 0.11886f
C14603 XThR.Tn[12].t59 VGND 0.01895f
C14604 XThR.Tn[12].t65 VGND 0.02075f
C14605 XThR.Tn[12].n44 VGND 0.05067f
C14606 XThR.Tn[12].t14 VGND 0.01889f
C14607 XThR.Tn[12].t44 VGND 0.02068f
C14608 XThR.Tn[12].n45 VGND 0.05272f
C14609 XThR.Tn[12].n46 VGND 0.03704f
C14610 XThR.Tn[12].n47 VGND 0.00677f
C14611 XThR.Tn[12].n48 VGND 0.11886f
C14612 XThR.Tn[12].t12 VGND 0.01895f
C14613 XThR.Tn[12].t22 VGND 0.02075f
C14614 XThR.Tn[12].n49 VGND 0.05067f
C14615 XThR.Tn[12].t35 VGND 0.01889f
C14616 XThR.Tn[12].t61 VGND 0.02068f
C14617 XThR.Tn[12].n50 VGND 0.05272f
C14618 XThR.Tn[12].n51 VGND 0.03704f
C14619 XThR.Tn[12].n52 VGND 0.00677f
C14620 XThR.Tn[12].n53 VGND 0.11886f
C14621 XThR.Tn[12].t68 VGND 0.01895f
C14622 XThR.Tn[12].t40 VGND 0.02075f
C14623 XThR.Tn[12].n54 VGND 0.05067f
C14624 XThR.Tn[12].t26 VGND 0.01889f
C14625 XThR.Tn[12].t19 VGND 0.02068f
C14626 XThR.Tn[12].n55 VGND 0.05272f
C14627 XThR.Tn[12].n56 VGND 0.03704f
C14628 XThR.Tn[12].n57 VGND 0.00677f
C14629 XThR.Tn[12].n58 VGND 0.11886f
C14630 XThR.Tn[12].t25 VGND 0.01895f
C14631 XThR.Tn[12].t16 VGND 0.02075f
C14632 XThR.Tn[12].n59 VGND 0.05067f
C14633 XThR.Tn[12].t42 VGND 0.01889f
C14634 XThR.Tn[12].t55 VGND 0.02068f
C14635 XThR.Tn[12].n60 VGND 0.05272f
C14636 XThR.Tn[12].n61 VGND 0.03704f
C14637 XThR.Tn[12].n62 VGND 0.00677f
C14638 XThR.Tn[12].n63 VGND 0.11886f
C14639 XThR.Tn[12].t57 VGND 0.01895f
C14640 XThR.Tn[12].t52 VGND 0.02075f
C14641 XThR.Tn[12].n64 VGND 0.05067f
C14642 XThR.Tn[12].t13 VGND 0.01889f
C14643 XThR.Tn[12].t31 VGND 0.02068f
C14644 XThR.Tn[12].n65 VGND 0.05272f
C14645 XThR.Tn[12].n66 VGND 0.03704f
C14646 XThR.Tn[12].n67 VGND 0.00677f
C14647 XThR.Tn[12].n68 VGND 0.11886f
C14648 XThR.Tn[12].t73 VGND 0.01895f
C14649 XThR.Tn[12].t67 VGND 0.02075f
C14650 XThR.Tn[12].n69 VGND 0.05067f
C14651 XThR.Tn[12].t34 VGND 0.01889f
C14652 XThR.Tn[12].t47 VGND 0.02068f
C14653 XThR.Tn[12].n70 VGND 0.05272f
C14654 XThR.Tn[12].n71 VGND 0.03704f
C14655 XThR.Tn[12].n72 VGND 0.00677f
C14656 XThR.Tn[12].n73 VGND 0.11886f
C14657 XThR.Tn[12].t32 VGND 0.01895f
C14658 XThR.Tn[12].t24 VGND 0.02075f
C14659 XThR.Tn[12].n74 VGND 0.05067f
C14660 XThR.Tn[12].t50 VGND 0.01889f
C14661 XThR.Tn[12].t62 VGND 0.02068f
C14662 XThR.Tn[12].n75 VGND 0.05272f
C14663 XThR.Tn[12].n76 VGND 0.03704f
C14664 XThR.Tn[12].n77 VGND 0.00677f
C14665 XThR.Tn[12].n78 VGND 0.11886f
C14666 XThR.Tn[12].t69 VGND 0.01895f
C14667 XThR.Tn[12].t18 VGND 0.02075f
C14668 XThR.Tn[12].n79 VGND 0.05067f
C14669 XThR.Tn[12].t27 VGND 0.01889f
C14670 XThR.Tn[12].t58 VGND 0.02068f
C14671 XThR.Tn[12].n80 VGND 0.05272f
C14672 XThR.Tn[12].n81 VGND 0.03704f
C14673 XThR.Tn[12].n82 VGND 0.00677f
C14674 XThR.Tn[12].n83 VGND 0.11886f
C14675 XThR.Tn[12].n84 VGND 0.10802f
C14676 XThR.Tn[12].n85 VGND 0.36839f
C14677 XThR.Tn[12].t2 VGND 0.01576f
C14678 XThR.Tn[12].t0 VGND 0.01576f
C14679 XThR.Tn[12].n86 VGND 0.03152f
C14680 XThR.Tn[12].t3 VGND 0.01576f
C14681 XThR.Tn[12].t1 VGND 0.01576f
C14682 XThR.Tn[12].n87 VGND 0.03931f
C14683 XThR.Tn[12].n88 VGND 0.07268f
C14684 XThR.Tn[14].t8 VGND 0.02436f
C14685 XThR.Tn[14].t9 VGND 0.02436f
C14686 XThR.Tn[14].n0 VGND 0.07395f
C14687 XThR.Tn[14].t10 VGND 0.02436f
C14688 XThR.Tn[14].t11 VGND 0.02436f
C14689 XThR.Tn[14].n1 VGND 0.05414f
C14690 XThR.Tn[14].n2 VGND 0.24618f
C14691 XThR.Tn[14].t6 VGND 0.02436f
C14692 XThR.Tn[14].t7 VGND 0.02436f
C14693 XThR.Tn[14].n3 VGND 0.05262f
C14694 XThR.Tn[14].t4 VGND 0.02436f
C14695 XThR.Tn[14].t5 VGND 0.02436f
C14696 XThR.Tn[14].n4 VGND 0.08009f
C14697 XThR.Tn[14].n5 VGND 0.22239f
C14698 XThR.Tn[14].n6 VGND 0.01096f
C14699 XThR.Tn[14].t69 VGND 0.01904f
C14700 XThR.Tn[14].t62 VGND 0.02084f
C14701 XThR.Tn[14].n7 VGND 0.0509f
C14702 XThR.Tn[14].n8 VGND 0.09778f
C14703 XThR.Tn[14].t24 VGND 0.01904f
C14704 XThR.Tn[14].t13 VGND 0.02084f
C14705 XThR.Tn[14].n9 VGND 0.0509f
C14706 XThR.Tn[14].t28 VGND 0.01897f
C14707 XThR.Tn[14].t60 VGND 0.02078f
C14708 XThR.Tn[14].n10 VGND 0.05296f
C14709 XThR.Tn[14].n11 VGND 0.03721f
C14710 XThR.Tn[14].n12 VGND 0.0068f
C14711 XThR.Tn[14].n13 VGND 0.11939f
C14712 XThR.Tn[14].t64 VGND 0.01904f
C14713 XThR.Tn[14].t54 VGND 0.02084f
C14714 XThR.Tn[14].n14 VGND 0.0509f
C14715 XThR.Tn[14].t67 VGND 0.01897f
C14716 XThR.Tn[14].t34 VGND 0.02078f
C14717 XThR.Tn[14].n15 VGND 0.05296f
C14718 XThR.Tn[14].n16 VGND 0.03721f
C14719 XThR.Tn[14].n17 VGND 0.0068f
C14720 XThR.Tn[14].n18 VGND 0.11939f
C14721 XThR.Tn[14].t14 VGND 0.01904f
C14722 XThR.Tn[14].t72 VGND 0.02084f
C14723 XThR.Tn[14].n19 VGND 0.0509f
C14724 XThR.Tn[14].t17 VGND 0.01897f
C14725 XThR.Tn[14].t52 VGND 0.02078f
C14726 XThR.Tn[14].n20 VGND 0.05296f
C14727 XThR.Tn[14].n21 VGND 0.03721f
C14728 XThR.Tn[14].n22 VGND 0.0068f
C14729 XThR.Tn[14].n23 VGND 0.11939f
C14730 XThR.Tn[14].t44 VGND 0.01904f
C14731 XThR.Tn[14].t38 VGND 0.02084f
C14732 XThR.Tn[14].n24 VGND 0.0509f
C14733 XThR.Tn[14].t47 VGND 0.01897f
C14734 XThR.Tn[14].t18 VGND 0.02078f
C14735 XThR.Tn[14].n25 VGND 0.05296f
C14736 XThR.Tn[14].n26 VGND 0.03721f
C14737 XThR.Tn[14].n27 VGND 0.0068f
C14738 XThR.Tn[14].n28 VGND 0.11939f
C14739 XThR.Tn[14].t15 VGND 0.01904f
C14740 XThR.Tn[14].t73 VGND 0.02084f
C14741 XThR.Tn[14].n29 VGND 0.0509f
C14742 XThR.Tn[14].t21 VGND 0.01897f
C14743 XThR.Tn[14].t53 VGND 0.02078f
C14744 XThR.Tn[14].n30 VGND 0.05296f
C14745 XThR.Tn[14].n31 VGND 0.03721f
C14746 XThR.Tn[14].n32 VGND 0.0068f
C14747 XThR.Tn[14].n33 VGND 0.11939f
C14748 XThR.Tn[14].t57 VGND 0.01904f
C14749 XThR.Tn[14].t25 VGND 0.02084f
C14750 XThR.Tn[14].n34 VGND 0.0509f
C14751 XThR.Tn[14].t61 VGND 0.01897f
C14752 XThR.Tn[14].t71 VGND 0.02078f
C14753 XThR.Tn[14].n35 VGND 0.05296f
C14754 XThR.Tn[14].n36 VGND 0.03721f
C14755 XThR.Tn[14].n37 VGND 0.0068f
C14756 XThR.Tn[14].n38 VGND 0.11939f
C14757 XThR.Tn[14].t23 VGND 0.01904f
C14758 XThR.Tn[14].t19 VGND 0.02084f
C14759 XThR.Tn[14].n39 VGND 0.0509f
C14760 XThR.Tn[14].t29 VGND 0.01897f
C14761 XThR.Tn[14].t66 VGND 0.02078f
C14762 XThR.Tn[14].n40 VGND 0.05296f
C14763 XThR.Tn[14].n41 VGND 0.03721f
C14764 XThR.Tn[14].n42 VGND 0.0068f
C14765 XThR.Tn[14].n43 VGND 0.11939f
C14766 XThR.Tn[14].t27 VGND 0.01904f
C14767 XThR.Tn[14].t36 VGND 0.02084f
C14768 XThR.Tn[14].n44 VGND 0.0509f
C14769 XThR.Tn[14].t33 VGND 0.01897f
C14770 XThR.Tn[14].t16 VGND 0.02078f
C14771 XThR.Tn[14].n45 VGND 0.05296f
C14772 XThR.Tn[14].n46 VGND 0.03721f
C14773 XThR.Tn[14].n47 VGND 0.0068f
C14774 XThR.Tn[14].n48 VGND 0.11939f
C14775 XThR.Tn[14].t46 VGND 0.01904f
C14776 XThR.Tn[14].t56 VGND 0.02084f
C14777 XThR.Tn[14].n49 VGND 0.0509f
C14778 XThR.Tn[14].t50 VGND 0.01897f
C14779 XThR.Tn[14].t35 VGND 0.02078f
C14780 XThR.Tn[14].n50 VGND 0.05296f
C14781 XThR.Tn[14].n51 VGND 0.03721f
C14782 XThR.Tn[14].n52 VGND 0.0068f
C14783 XThR.Tn[14].n53 VGND 0.11939f
C14784 XThR.Tn[14].t40 VGND 0.01904f
C14785 XThR.Tn[14].t12 VGND 0.02084f
C14786 XThR.Tn[14].n54 VGND 0.0509f
C14787 XThR.Tn[14].t42 VGND 0.01897f
C14788 XThR.Tn[14].t55 VGND 0.02078f
C14789 XThR.Tn[14].n55 VGND 0.05296f
C14790 XThR.Tn[14].n56 VGND 0.03721f
C14791 XThR.Tn[14].n57 VGND 0.0068f
C14792 XThR.Tn[14].n58 VGND 0.11939f
C14793 XThR.Tn[14].t59 VGND 0.01904f
C14794 XThR.Tn[14].t49 VGND 0.02084f
C14795 XThR.Tn[14].n59 VGND 0.0509f
C14796 XThR.Tn[14].t63 VGND 0.01897f
C14797 XThR.Tn[14].t30 VGND 0.02078f
C14798 XThR.Tn[14].n60 VGND 0.05296f
C14799 XThR.Tn[14].n61 VGND 0.03721f
C14800 XThR.Tn[14].n62 VGND 0.0068f
C14801 XThR.Tn[14].n63 VGND 0.11939f
C14802 XThR.Tn[14].t26 VGND 0.01904f
C14803 XThR.Tn[14].t22 VGND 0.02084f
C14804 XThR.Tn[14].n64 VGND 0.0509f
C14805 XThR.Tn[14].t31 VGND 0.01897f
C14806 XThR.Tn[14].t68 VGND 0.02078f
C14807 XThR.Tn[14].n65 VGND 0.05296f
C14808 XThR.Tn[14].n66 VGND 0.03721f
C14809 XThR.Tn[14].n67 VGND 0.0068f
C14810 XThR.Tn[14].n68 VGND 0.11939f
C14811 XThR.Tn[14].t45 VGND 0.01904f
C14812 XThR.Tn[14].t39 VGND 0.02084f
C14813 XThR.Tn[14].n69 VGND 0.0509f
C14814 XThR.Tn[14].t48 VGND 0.01897f
C14815 XThR.Tn[14].t20 VGND 0.02078f
C14816 XThR.Tn[14].n70 VGND 0.05296f
C14817 XThR.Tn[14].n71 VGND 0.03721f
C14818 XThR.Tn[14].n72 VGND 0.0068f
C14819 XThR.Tn[14].n73 VGND 0.11939f
C14820 XThR.Tn[14].t65 VGND 0.01904f
C14821 XThR.Tn[14].t58 VGND 0.02084f
C14822 XThR.Tn[14].n74 VGND 0.0509f
C14823 XThR.Tn[14].t70 VGND 0.01897f
C14824 XThR.Tn[14].t37 VGND 0.02078f
C14825 XThR.Tn[14].n75 VGND 0.05296f
C14826 XThR.Tn[14].n76 VGND 0.03721f
C14827 XThR.Tn[14].n77 VGND 0.0068f
C14828 XThR.Tn[14].n78 VGND 0.11939f
C14829 XThR.Tn[14].t41 VGND 0.01904f
C14830 XThR.Tn[14].t51 VGND 0.02084f
C14831 XThR.Tn[14].n79 VGND 0.0509f
C14832 XThR.Tn[14].t43 VGND 0.01897f
C14833 XThR.Tn[14].t32 VGND 0.02078f
C14834 XThR.Tn[14].n80 VGND 0.05296f
C14835 XThR.Tn[14].n81 VGND 0.03721f
C14836 XThR.Tn[14].n82 VGND 0.0068f
C14837 XThR.Tn[14].n83 VGND 0.11939f
C14838 XThR.Tn[14].n84 VGND 0.1085f
C14839 XThR.Tn[14].n85 VGND 0.43585f
C14840 XThR.Tn[14].t0 VGND 0.01583f
C14841 XThR.Tn[14].t1 VGND 0.01583f
C14842 XThR.Tn[14].n86 VGND 0.03166f
C14843 XThR.Tn[14].t2 VGND 0.01583f
C14844 XThR.Tn[14].t3 VGND 0.01583f
C14845 XThR.Tn[14].n87 VGND 0.03948f
C14846 XThR.Tn[14].n88 VGND 0.07301f
C14847 XThR.Tn[6].t7 VGND 0.02335f
C14848 XThR.Tn[6].t4 VGND 0.02335f
C14849 XThR.Tn[6].n0 VGND 0.04712f
C14850 XThR.Tn[6].t6 VGND 0.02335f
C14851 XThR.Tn[6].t5 VGND 0.02335f
C14852 XThR.Tn[6].n1 VGND 0.05514f
C14853 XThR.Tn[6].n2 VGND 0.16538f
C14854 XThR.Tn[6].t8 VGND 0.01517f
C14855 XThR.Tn[6].t9 VGND 0.01517f
C14856 XThR.Tn[6].n3 VGND 0.03456f
C14857 XThR.Tn[6].t11 VGND 0.01517f
C14858 XThR.Tn[6].t10 VGND 0.01517f
C14859 XThR.Tn[6].n4 VGND 0.03456f
C14860 XThR.Tn[6].t0 VGND 0.01517f
C14861 XThR.Tn[6].t1 VGND 0.01517f
C14862 XThR.Tn[6].n5 VGND 0.05758f
C14863 XThR.Tn[6].t3 VGND 0.01517f
C14864 XThR.Tn[6].t2 VGND 0.01517f
C14865 XThR.Tn[6].n6 VGND 0.03456f
C14866 XThR.Tn[6].n7 VGND 0.16456f
C14867 XThR.Tn[6].n8 VGND 0.10173f
C14868 XThR.Tn[6].n9 VGND 0.11481f
C14869 XThR.Tn[6].t62 VGND 0.01825f
C14870 XThR.Tn[6].t56 VGND 0.01998f
C14871 XThR.Tn[6].n10 VGND 0.04879f
C14872 XThR.Tn[6].n11 VGND 0.09372f
C14873 XThR.Tn[6].t20 VGND 0.01825f
C14874 XThR.Tn[6].t72 VGND 0.01998f
C14875 XThR.Tn[6].n12 VGND 0.04879f
C14876 XThR.Tn[6].t36 VGND 0.01819f
C14877 XThR.Tn[6].t68 VGND 0.01991f
C14878 XThR.Tn[6].n13 VGND 0.05076f
C14879 XThR.Tn[6].n14 VGND 0.03566f
C14880 XThR.Tn[6].n15 VGND 0.00652f
C14881 XThR.Tn[6].n16 VGND 0.11444f
C14882 XThR.Tn[6].t57 VGND 0.01825f
C14883 XThR.Tn[6].t49 VGND 0.01998f
C14884 XThR.Tn[6].n17 VGND 0.04879f
C14885 XThR.Tn[6].t14 VGND 0.01819f
C14886 XThR.Tn[6].t45 VGND 0.01991f
C14887 XThR.Tn[6].n18 VGND 0.05076f
C14888 XThR.Tn[6].n19 VGND 0.03566f
C14889 XThR.Tn[6].n20 VGND 0.00652f
C14890 XThR.Tn[6].n21 VGND 0.11444f
C14891 XThR.Tn[6].t73 VGND 0.01825f
C14892 XThR.Tn[6].t66 VGND 0.01998f
C14893 XThR.Tn[6].n22 VGND 0.04879f
C14894 XThR.Tn[6].t26 VGND 0.01819f
C14895 XThR.Tn[6].t63 VGND 0.01991f
C14896 XThR.Tn[6].n23 VGND 0.05076f
C14897 XThR.Tn[6].n24 VGND 0.03566f
C14898 XThR.Tn[6].n25 VGND 0.00652f
C14899 XThR.Tn[6].n26 VGND 0.11444f
C14900 XThR.Tn[6].t35 VGND 0.01825f
C14901 XThR.Tn[6].t31 VGND 0.01998f
C14902 XThR.Tn[6].n27 VGND 0.04879f
C14903 XThR.Tn[6].t59 VGND 0.01819f
C14904 XThR.Tn[6].t27 VGND 0.01991f
C14905 XThR.Tn[6].n28 VGND 0.05076f
C14906 XThR.Tn[6].n29 VGND 0.03566f
C14907 XThR.Tn[6].n30 VGND 0.00652f
C14908 XThR.Tn[6].n31 VGND 0.11444f
C14909 XThR.Tn[6].t13 VGND 0.01825f
C14910 XThR.Tn[6].t67 VGND 0.01998f
C14911 XThR.Tn[6].n32 VGND 0.04879f
C14912 XThR.Tn[6].t29 VGND 0.01819f
C14913 XThR.Tn[6].t64 VGND 0.01991f
C14914 XThR.Tn[6].n33 VGND 0.05076f
C14915 XThR.Tn[6].n34 VGND 0.03566f
C14916 XThR.Tn[6].n35 VGND 0.00652f
C14917 XThR.Tn[6].n36 VGND 0.11444f
C14918 XThR.Tn[6].t51 VGND 0.01825f
C14919 XThR.Tn[6].t22 VGND 0.01998f
C14920 XThR.Tn[6].n37 VGND 0.04879f
C14921 XThR.Tn[6].t70 VGND 0.01819f
C14922 XThR.Tn[6].t19 VGND 0.01991f
C14923 XThR.Tn[6].n38 VGND 0.05076f
C14924 XThR.Tn[6].n39 VGND 0.03566f
C14925 XThR.Tn[6].n40 VGND 0.00652f
C14926 XThR.Tn[6].n41 VGND 0.11444f
C14927 XThR.Tn[6].t21 VGND 0.01825f
C14928 XThR.Tn[6].t17 VGND 0.01998f
C14929 XThR.Tn[6].n42 VGND 0.04879f
C14930 XThR.Tn[6].t37 VGND 0.01819f
C14931 XThR.Tn[6].t12 VGND 0.01991f
C14932 XThR.Tn[6].n43 VGND 0.05076f
C14933 XThR.Tn[6].n44 VGND 0.03566f
C14934 XThR.Tn[6].n45 VGND 0.00652f
C14935 XThR.Tn[6].n46 VGND 0.11444f
C14936 XThR.Tn[6].t24 VGND 0.01825f
C14937 XThR.Tn[6].t30 VGND 0.01998f
C14938 XThR.Tn[6].n47 VGND 0.04879f
C14939 XThR.Tn[6].t43 VGND 0.01819f
C14940 XThR.Tn[6].t25 VGND 0.01991f
C14941 XThR.Tn[6].n48 VGND 0.05076f
C14942 XThR.Tn[6].n49 VGND 0.03566f
C14943 XThR.Tn[6].n50 VGND 0.00652f
C14944 XThR.Tn[6].n51 VGND 0.11444f
C14945 XThR.Tn[6].t40 VGND 0.01825f
C14946 XThR.Tn[6].t50 VGND 0.01998f
C14947 XThR.Tn[6].n52 VGND 0.04879f
C14948 XThR.Tn[6].t61 VGND 0.01819f
C14949 XThR.Tn[6].t47 VGND 0.01991f
C14950 XThR.Tn[6].n53 VGND 0.05076f
C14951 XThR.Tn[6].n54 VGND 0.03566f
C14952 XThR.Tn[6].n55 VGND 0.00652f
C14953 XThR.Tn[6].n56 VGND 0.11444f
C14954 XThR.Tn[6].t33 VGND 0.01825f
C14955 XThR.Tn[6].t69 VGND 0.01998f
C14956 XThR.Tn[6].n57 VGND 0.04879f
C14957 XThR.Tn[6].t54 VGND 0.01819f
C14958 XThR.Tn[6].t65 VGND 0.01991f
C14959 XThR.Tn[6].n58 VGND 0.05076f
C14960 XThR.Tn[6].n59 VGND 0.03566f
C14961 XThR.Tn[6].n60 VGND 0.00652f
C14962 XThR.Tn[6].n61 VGND 0.11444f
C14963 XThR.Tn[6].t53 VGND 0.01825f
C14964 XThR.Tn[6].t44 VGND 0.01998f
C14965 XThR.Tn[6].n62 VGND 0.04879f
C14966 XThR.Tn[6].t71 VGND 0.01819f
C14967 XThR.Tn[6].t39 VGND 0.01991f
C14968 XThR.Tn[6].n63 VGND 0.05076f
C14969 XThR.Tn[6].n64 VGND 0.03566f
C14970 XThR.Tn[6].n65 VGND 0.00652f
C14971 XThR.Tn[6].n66 VGND 0.11444f
C14972 XThR.Tn[6].t23 VGND 0.01825f
C14973 XThR.Tn[6].t18 VGND 0.01998f
C14974 XThR.Tn[6].n67 VGND 0.04879f
C14975 XThR.Tn[6].t41 VGND 0.01819f
C14976 XThR.Tn[6].t15 VGND 0.01991f
C14977 XThR.Tn[6].n68 VGND 0.05076f
C14978 XThR.Tn[6].n69 VGND 0.03566f
C14979 XThR.Tn[6].n70 VGND 0.00652f
C14980 XThR.Tn[6].n71 VGND 0.11444f
C14981 XThR.Tn[6].t38 VGND 0.01825f
C14982 XThR.Tn[6].t32 VGND 0.01998f
C14983 XThR.Tn[6].n72 VGND 0.04879f
C14984 XThR.Tn[6].t60 VGND 0.01819f
C14985 XThR.Tn[6].t28 VGND 0.01991f
C14986 XThR.Tn[6].n73 VGND 0.05076f
C14987 XThR.Tn[6].n74 VGND 0.03566f
C14988 XThR.Tn[6].n75 VGND 0.00652f
C14989 XThR.Tn[6].n76 VGND 0.11444f
C14990 XThR.Tn[6].t58 VGND 0.01825f
C14991 XThR.Tn[6].t52 VGND 0.01998f
C14992 XThR.Tn[6].n77 VGND 0.04879f
C14993 XThR.Tn[6].t16 VGND 0.01819f
C14994 XThR.Tn[6].t48 VGND 0.01991f
C14995 XThR.Tn[6].n78 VGND 0.05076f
C14996 XThR.Tn[6].n79 VGND 0.03566f
C14997 XThR.Tn[6].n80 VGND 0.00652f
C14998 XThR.Tn[6].n81 VGND 0.11444f
C14999 XThR.Tn[6].t34 VGND 0.01825f
C15000 XThR.Tn[6].t46 VGND 0.01998f
C15001 XThR.Tn[6].n82 VGND 0.04879f
C15002 XThR.Tn[6].t55 VGND 0.01819f
C15003 XThR.Tn[6].t42 VGND 0.01991f
C15004 XThR.Tn[6].n83 VGND 0.05076f
C15005 XThR.Tn[6].n84 VGND 0.03566f
C15006 XThR.Tn[6].n85 VGND 0.00652f
C15007 XThR.Tn[6].n86 VGND 0.11444f
C15008 XThR.Tn[6].n87 VGND 0.104f
C15009 XThR.Tn[6].n88 VGND 0.17311f
C15010 XThR.TBN.n0 VGND 0.00433f
C15011 XThR.TBN.t60 VGND 0.01124f
C15012 XThR.TBN.t95 VGND 0.00662f
C15013 XThR.TBN.n1 VGND 0.01347f
C15014 XThR.TBN.t12 VGND 0.01124f
C15015 XThR.TBN.t44 VGND 0.00662f
C15016 XThR.TBN.t81 VGND 0.01124f
C15017 XThR.TBN.t116 VGND 0.00662f
C15018 XThR.TBN.n2 VGND 0.01479f
C15019 XThR.TBN.t121 VGND 0.01124f
C15020 XThR.TBN.t35 VGND 0.00662f
C15021 XThR.TBN.n3 VGND 0.01365f
C15022 XThR.TBN.n4 VGND 0.00834f
C15023 XThR.TBN.n5 VGND 0.01304f
C15024 XThR.TBN.n6 VGND 0.0068f
C15025 XThR.TBN.n7 VGND 0.00662f
C15026 XThR.TBN.n8 VGND 0.01479f
C15027 XThR.TBN.n9 VGND 0.00742f
C15028 XThR.TBN.n10 VGND 0.0122f
C15029 XThR.TBN.n11 VGND 0.00433f
C15030 XThR.TBN.t42 VGND 0.00662f
C15031 XThR.TBN.t115 VGND 0.01124f
C15032 XThR.TBN.n12 VGND 0.01347f
C15033 XThR.TBN.t112 VGND 0.00662f
C15034 XThR.TBN.t65 VGND 0.01124f
C15035 XThR.TBN.t64 VGND 0.00662f
C15036 XThR.TBN.t21 VGND 0.01124f
C15037 XThR.TBN.n13 VGND 0.01479f
C15038 XThR.TBN.t107 VGND 0.00662f
C15039 XThR.TBN.t57 VGND 0.01124f
C15040 XThR.TBN.n14 VGND 0.01365f
C15041 XThR.TBN.n15 VGND 0.00834f
C15042 XThR.TBN.n16 VGND 0.01304f
C15043 XThR.TBN.n17 VGND 0.0068f
C15044 XThR.TBN.n18 VGND 0.00662f
C15045 XThR.TBN.n19 VGND 0.01479f
C15046 XThR.TBN.n20 VGND 0.00742f
C15047 XThR.TBN.n21 VGND 0.00932f
C15048 XThR.TBN.n22 VGND 0.12354f
C15049 XThR.TBN.n23 VGND 0.00433f
C15050 XThR.TBN.t27 VGND 0.01124f
C15051 XThR.TBN.t61 VGND 0.00662f
C15052 XThR.TBN.n24 VGND 0.01347f
C15053 XThR.TBN.t96 VGND 0.01124f
C15054 XThR.TBN.t14 VGND 0.00662f
C15055 XThR.TBN.t46 VGND 0.01124f
C15056 XThR.TBN.t82 VGND 0.00662f
C15057 XThR.TBN.n25 VGND 0.01479f
C15058 XThR.TBN.t89 VGND 0.01124f
C15059 XThR.TBN.t122 VGND 0.00662f
C15060 XThR.TBN.n26 VGND 0.01365f
C15061 XThR.TBN.n27 VGND 0.00834f
C15062 XThR.TBN.n28 VGND 0.01304f
C15063 XThR.TBN.n29 VGND 0.0068f
C15064 XThR.TBN.n30 VGND 0.00662f
C15065 XThR.TBN.n31 VGND 0.01479f
C15066 XThR.TBN.n32 VGND 0.00742f
C15067 XThR.TBN.n33 VGND 0.00932f
C15068 XThR.TBN.n34 VGND 0.08255f
C15069 XThR.TBN.n35 VGND 0.00433f
C15070 XThR.TBN.t11 VGND 0.00662f
C15071 XThR.TBN.t80 VGND 0.01124f
C15072 XThR.TBN.n36 VGND 0.01347f
C15073 XThR.TBN.t79 VGND 0.00662f
C15074 XThR.TBN.t31 VGND 0.01124f
C15075 XThR.TBN.t32 VGND 0.00662f
C15076 XThR.TBN.t102 VGND 0.01124f
C15077 XThR.TBN.n37 VGND 0.01479f
C15078 XThR.TBN.t71 VGND 0.00662f
C15079 XThR.TBN.t25 VGND 0.01124f
C15080 XThR.TBN.n38 VGND 0.01365f
C15081 XThR.TBN.n39 VGND 0.00834f
C15082 XThR.TBN.n40 VGND 0.01304f
C15083 XThR.TBN.n41 VGND 0.0068f
C15084 XThR.TBN.n42 VGND 0.00662f
C15085 XThR.TBN.n43 VGND 0.01479f
C15086 XThR.TBN.n44 VGND 0.00742f
C15087 XThR.TBN.n45 VGND 0.00932f
C15088 XThR.TBN.n46 VGND 0.08255f
C15089 XThR.TBN.n47 VGND 0.00433f
C15090 XThR.TBN.t85 VGND 0.01124f
C15091 XThR.TBN.t29 VGND 0.00662f
C15092 XThR.TBN.n48 VGND 0.01347f
C15093 XThR.TBN.t33 VGND 0.01124f
C15094 XThR.TBN.t98 VGND 0.00662f
C15095 XThR.TBN.t105 VGND 0.01124f
C15096 XThR.TBN.t47 VGND 0.00662f
C15097 XThR.TBN.n49 VGND 0.01479f
C15098 XThR.TBN.t26 VGND 0.01124f
C15099 XThR.TBN.t90 VGND 0.00662f
C15100 XThR.TBN.n50 VGND 0.01365f
C15101 XThR.TBN.n51 VGND 0.00834f
C15102 XThR.TBN.n52 VGND 0.01304f
C15103 XThR.TBN.n53 VGND 0.0068f
C15104 XThR.TBN.n54 VGND 0.00662f
C15105 XThR.TBN.n55 VGND 0.01479f
C15106 XThR.TBN.n56 VGND 0.00742f
C15107 XThR.TBN.n57 VGND 0.00932f
C15108 XThR.TBN.n58 VGND 0.08269f
C15109 XThR.TBN.n59 VGND 0.00433f
C15110 XThR.TBN.t8 VGND 0.00662f
C15111 XThR.TBN.t54 VGND 0.01124f
C15112 XThR.TBN.n60 VGND 0.01347f
C15113 XThR.TBN.t74 VGND 0.00662f
C15114 XThR.TBN.t5 VGND 0.01124f
C15115 XThR.TBN.t28 VGND 0.00662f
C15116 XThR.TBN.t73 VGND 0.01124f
C15117 XThR.TBN.n61 VGND 0.01479f
C15118 XThR.TBN.t67 VGND 0.00662f
C15119 XThR.TBN.t114 VGND 0.01124f
C15120 XThR.TBN.n62 VGND 0.01365f
C15121 XThR.TBN.n63 VGND 0.00834f
C15122 XThR.TBN.n64 VGND 0.01304f
C15123 XThR.TBN.n65 VGND 0.0068f
C15124 XThR.TBN.n66 VGND 0.00662f
C15125 XThR.TBN.n67 VGND 0.01479f
C15126 XThR.TBN.n68 VGND 0.00742f
C15127 XThR.TBN.n69 VGND 0.00932f
C15128 XThR.TBN.n70 VGND 0.08255f
C15129 XThR.TBN.n71 VGND 0.00433f
C15130 XThR.TBN.t49 VGND 0.01124f
C15131 XThR.TBN.t111 VGND 0.00662f
C15132 XThR.TBN.n72 VGND 0.01347f
C15133 XThR.TBN.t119 VGND 0.01124f
C15134 XThR.TBN.t62 VGND 0.00662f
C15135 XThR.TBN.t69 VGND 0.01124f
C15136 XThR.TBN.t18 VGND 0.00662f
C15137 XThR.TBN.n73 VGND 0.01479f
C15138 XThR.TBN.t108 VGND 0.01124f
C15139 XThR.TBN.t53 VGND 0.00662f
C15140 XThR.TBN.n74 VGND 0.01365f
C15141 XThR.TBN.n75 VGND 0.00834f
C15142 XThR.TBN.n76 VGND 0.01304f
C15143 XThR.TBN.n77 VGND 0.0068f
C15144 XThR.TBN.n78 VGND 0.00662f
C15145 XThR.TBN.n79 VGND 0.01479f
C15146 XThR.TBN.n80 VGND 0.00742f
C15147 XThR.TBN.n81 VGND 0.00932f
C15148 XThR.TBN.n82 VGND 0.09424f
C15149 XThR.TBN.t99 VGND 0.01124f
C15150 XThR.TBN.t20 VGND 0.00662f
C15151 XThR.TBN.t87 VGND 0.01124f
C15152 XThR.TBN.t120 VGND 0.00662f
C15153 XThR.TBN.n83 VGND 0.01621f
C15154 XThR.TBN.t77 VGND 0.01124f
C15155 XThR.TBN.t110 VGND 0.00662f
C15156 XThR.TBN.t68 VGND 0.01124f
C15157 XThR.TBN.t103 VGND 0.00662f
C15158 XThR.TBN.n84 VGND 0.01515f
C15159 XThR.TBN.n85 VGND 0.00615f
C15160 XThR.TBN.n86 VGND 0.00742f
C15161 XThR.TBN.n87 VGND 0.01621f
C15162 XThR.TBN.n88 VGND 0.00742f
C15163 XThR.TBN.n89 VGND 0.00615f
C15164 XThR.TBN.n90 VGND 0.00615f
C15165 XThR.TBN.n91 VGND 0.00742f
C15166 XThR.TBN.n92 VGND 0.02375f
C15167 XThR.TBN.n93 VGND 0.01318f
C15168 XThR.TBN.t24 VGND 0.00662f
C15169 XThR.TBN.t66 VGND 0.01124f
C15170 XThR.TBN.t91 VGND 0.00662f
C15171 XThR.TBN.t23 VGND 0.01124f
C15172 XThR.TBN.n94 VGND 0.01621f
C15173 XThR.TBN.t10 VGND 0.00662f
C15174 XThR.TBN.t59 VGND 0.01124f
C15175 XThR.TBN.t48 VGND 0.00662f
C15176 XThR.TBN.t97 VGND 0.01124f
C15177 XThR.TBN.n95 VGND 0.01515f
C15178 XThR.TBN.n96 VGND 0.00615f
C15179 XThR.TBN.n97 VGND 0.00742f
C15180 XThR.TBN.n98 VGND 0.01621f
C15181 XThR.TBN.n99 VGND 0.00742f
C15182 XThR.TBN.n100 VGND 0.00615f
C15183 XThR.TBN.n101 VGND 0.00615f
C15184 XThR.TBN.n102 VGND 0.00742f
C15185 XThR.TBN.n103 VGND 0.02375f
C15186 XThR.TBN.n104 VGND 0.0086f
C15187 XThR.TBN.n105 VGND 0.13142f
C15188 XThR.TBN.t15 VGND 0.01124f
C15189 XThR.TBN.t38 VGND 0.00662f
C15190 XThR.TBN.t83 VGND 0.01124f
C15191 XThR.TBN.t109 VGND 0.00662f
C15192 XThR.TBN.n106 VGND 0.01621f
C15193 XThR.TBN.t123 VGND 0.01124f
C15194 XThR.TBN.t30 VGND 0.00662f
C15195 XThR.TBN.t39 VGND 0.01124f
C15196 XThR.TBN.t70 VGND 0.00662f
C15197 XThR.TBN.n107 VGND 0.01515f
C15198 XThR.TBN.n108 VGND 0.00615f
C15199 XThR.TBN.n109 VGND 0.00742f
C15200 XThR.TBN.n110 VGND 0.01621f
C15201 XThR.TBN.n111 VGND 0.00742f
C15202 XThR.TBN.n112 VGND 0.00615f
C15203 XThR.TBN.n113 VGND 0.00615f
C15204 XThR.TBN.n114 VGND 0.00742f
C15205 XThR.TBN.n115 VGND 0.02375f
C15206 XThR.TBN.n116 VGND 0.0086f
C15207 XThR.TBN.n117 VGND 0.08248f
C15208 XThR.TBN.t51 VGND 0.00662f
C15209 XThR.TBN.t100 VGND 0.01124f
C15210 XThR.TBN.t4 VGND 0.00662f
C15211 XThR.TBN.t50 VGND 0.01124f
C15212 XThR.TBN.n118 VGND 0.01621f
C15213 XThR.TBN.t40 VGND 0.00662f
C15214 XThR.TBN.t92 VGND 0.01124f
C15215 XThR.TBN.t84 VGND 0.00662f
C15216 XThR.TBN.t13 VGND 0.01124f
C15217 XThR.TBN.n119 VGND 0.01515f
C15218 XThR.TBN.n120 VGND 0.00615f
C15219 XThR.TBN.n121 VGND 0.00742f
C15220 XThR.TBN.n122 VGND 0.01621f
C15221 XThR.TBN.n123 VGND 0.00742f
C15222 XThR.TBN.n124 VGND 0.00615f
C15223 XThR.TBN.n125 VGND 0.00615f
C15224 XThR.TBN.n126 VGND 0.00742f
C15225 XThR.TBN.n127 VGND 0.02375f
C15226 XThR.TBN.n128 VGND 0.0086f
C15227 XThR.TBN.n129 VGND 0.08248f
C15228 XThR.TBN.t45 VGND 0.01124f
C15229 XThR.TBN.t104 VGND 0.00662f
C15230 XThR.TBN.t117 VGND 0.01124f
C15231 XThR.TBN.t55 VGND 0.00662f
C15232 XThR.TBN.n130 VGND 0.01621f
C15233 XThR.TBN.t36 VGND 0.01124f
C15234 XThR.TBN.t94 VGND 0.00662f
C15235 XThR.TBN.t75 VGND 0.01124f
C15236 XThR.TBN.t17 VGND 0.00662f
C15237 XThR.TBN.n131 VGND 0.01515f
C15238 XThR.TBN.n132 VGND 0.00615f
C15239 XThR.TBN.n133 VGND 0.00742f
C15240 XThR.TBN.n134 VGND 0.01621f
C15241 XThR.TBN.n135 VGND 0.00742f
C15242 XThR.TBN.n136 VGND 0.00615f
C15243 XThR.TBN.n137 VGND 0.00615f
C15244 XThR.TBN.n138 VGND 0.00742f
C15245 XThR.TBN.n139 VGND 0.02375f
C15246 XThR.TBN.n140 VGND 0.0086f
C15247 XThR.TBN.n141 VGND 0.08248f
C15248 XThR.TBN.t88 VGND 0.00662f
C15249 XThR.TBN.t19 VGND 0.01124f
C15250 XThR.TBN.t37 VGND 0.00662f
C15251 XThR.TBN.t86 VGND 0.01124f
C15252 XThR.TBN.n142 VGND 0.01621f
C15253 XThR.TBN.t76 VGND 0.00662f
C15254 XThR.TBN.t6 VGND 0.01124f
C15255 XThR.TBN.t118 VGND 0.00662f
C15256 XThR.TBN.t43 VGND 0.01124f
C15257 XThR.TBN.n143 VGND 0.01515f
C15258 XThR.TBN.n144 VGND 0.00615f
C15259 XThR.TBN.n145 VGND 0.00742f
C15260 XThR.TBN.n146 VGND 0.01621f
C15261 XThR.TBN.n147 VGND 0.00742f
C15262 XThR.TBN.n148 VGND 0.00615f
C15263 XThR.TBN.n149 VGND 0.00615f
C15264 XThR.TBN.n150 VGND 0.00742f
C15265 XThR.TBN.n151 VGND 0.02375f
C15266 XThR.TBN.n152 VGND 0.0086f
C15267 XThR.TBN.n153 VGND 0.08248f
C15268 XThR.TBN.t41 VGND 0.01124f
C15269 XThR.TBN.t101 VGND 0.00662f
C15270 XThR.TBN.t113 VGND 0.01124f
C15271 XThR.TBN.t52 VGND 0.00662f
C15272 XThR.TBN.n154 VGND 0.01621f
C15273 XThR.TBN.t34 VGND 0.01124f
C15274 XThR.TBN.t93 VGND 0.00662f
C15275 XThR.TBN.t72 VGND 0.01124f
C15276 XThR.TBN.t16 VGND 0.00662f
C15277 XThR.TBN.n155 VGND 0.01515f
C15278 XThR.TBN.n156 VGND 0.00615f
C15279 XThR.TBN.n157 VGND 0.00742f
C15280 XThR.TBN.n158 VGND 0.01621f
C15281 XThR.TBN.n159 VGND 0.00742f
C15282 XThR.TBN.n160 VGND 0.00615f
C15283 XThR.TBN.n161 VGND 0.00615f
C15284 XThR.TBN.n162 VGND 0.00742f
C15285 XThR.TBN.n163 VGND 0.02375f
C15286 XThR.TBN.n164 VGND 0.0086f
C15287 XThR.TBN.n165 VGND 0.07393f
C15288 XThR.TBN.n166 VGND 0.08425f
C15289 XThR.TBN.t58 VGND 0.00662f
C15290 XThR.TBN.t106 VGND 0.01124f
C15291 XThR.TBN.t22 VGND 0.00662f
C15292 XThR.TBN.t63 VGND 0.01124f
C15293 XThR.TBN.n167 VGND 0.01515f
C15294 XThR.TBN.n168 VGND 0.00749f
C15295 XThR.TBN.n169 VGND 0.01621f
C15296 XThR.TBN.t9 VGND 0.00662f
C15297 XThR.TBN.t56 VGND 0.01124f
C15298 XThR.TBN.t78 VGND 0.00662f
C15299 XThR.TBN.t7 VGND 0.01124f
C15300 XThR.TBN.n170 VGND 0.02517f
C15301 XThR.TBN.n171 VGND 0.00814f
C15302 XThR.TBN.n172 VGND 0.00615f
C15303 XThR.TBN.n173 VGND 0.00742f
C15304 XThR.TBN.n174 VGND 0.01621f
C15305 XThR.TBN.n175 VGND 0.00742f
C15306 XThR.TBN.n176 VGND 0.00435f
C15307 XThR.TBN.n177 VGND 0.00502f
C15308 XThR.TBN.n178 VGND 0.12255f
C15309 XThR.TBN.n179 VGND 0.02242f
C15310 XThR.TBN.t3 VGND 0.00722f
C15311 XThR.TBN.t2 VGND 0.00722f
C15312 XThR.TBN.n180 VGND 0.01587f
C15313 XThR.TBN.n181 VGND 0.00684f
C15314 XThR.TBN.n182 VGND 0.00577f
C15315 XThR.TBN.t0 VGND 0.0047f
C15316 XThR.TBN.t1 VGND 0.0047f
C15317 XThR.TBN.n183 VGND 0.0112f
C15318 XThR.TBN.n184 VGND 0.022f
C15319 XThC.Tn[10].t6 VGND 0.01306f
C15320 XThC.Tn[10].t4 VGND 0.01306f
C15321 XThC.Tn[10].n0 VGND 0.03258f
C15322 XThC.Tn[10].t2 VGND 0.01306f
C15323 XThC.Tn[10].t7 VGND 0.01306f
C15324 XThC.Tn[10].n1 VGND 0.02613f
C15325 XThC.Tn[10].n2 VGND 0.06572f
C15326 XThC.Tn[10].n3 VGND 0.02851f
C15327 XThC.Tn[10].t38 VGND 0.01593f
C15328 XThC.Tn[10].t36 VGND 0.0174f
C15329 XThC.Tn[10].n4 VGND 0.03884f
C15330 XThC.Tn[10].n5 VGND 0.02661f
C15331 XThC.Tn[10].n6 VGND 0.08734f
C15332 XThC.Tn[10].t24 VGND 0.01593f
C15333 XThC.Tn[10].t21 VGND 0.0174f
C15334 XThC.Tn[10].n7 VGND 0.03884f
C15335 XThC.Tn[10].n8 VGND 0.02661f
C15336 XThC.Tn[10].n9 VGND 0.08758f
C15337 XThC.Tn[10].n10 VGND 0.14434f
C15338 XThC.Tn[10].t29 VGND 0.01593f
C15339 XThC.Tn[10].t23 VGND 0.0174f
C15340 XThC.Tn[10].n11 VGND 0.03884f
C15341 XThC.Tn[10].n12 VGND 0.02661f
C15342 XThC.Tn[10].n13 VGND 0.08758f
C15343 XThC.Tn[10].n14 VGND 0.14434f
C15344 XThC.Tn[10].t30 VGND 0.01593f
C15345 XThC.Tn[10].t25 VGND 0.0174f
C15346 XThC.Tn[10].n15 VGND 0.03884f
C15347 XThC.Tn[10].n16 VGND 0.02661f
C15348 XThC.Tn[10].n17 VGND 0.08758f
C15349 XThC.Tn[10].n18 VGND 0.14434f
C15350 XThC.Tn[10].t17 VGND 0.01593f
C15351 XThC.Tn[10].t14 VGND 0.0174f
C15352 XThC.Tn[10].n19 VGND 0.03884f
C15353 XThC.Tn[10].n20 VGND 0.02661f
C15354 XThC.Tn[10].n21 VGND 0.08758f
C15355 XThC.Tn[10].n22 VGND 0.14434f
C15356 XThC.Tn[10].t18 VGND 0.01593f
C15357 XThC.Tn[10].t15 VGND 0.0174f
C15358 XThC.Tn[10].n23 VGND 0.03884f
C15359 XThC.Tn[10].n24 VGND 0.02661f
C15360 XThC.Tn[10].n25 VGND 0.08758f
C15361 XThC.Tn[10].n26 VGND 0.14434f
C15362 XThC.Tn[10].t34 VGND 0.01593f
C15363 XThC.Tn[10].t28 VGND 0.0174f
C15364 XThC.Tn[10].n27 VGND 0.03884f
C15365 XThC.Tn[10].n28 VGND 0.02661f
C15366 XThC.Tn[10].n29 VGND 0.08758f
C15367 XThC.Tn[10].n30 VGND 0.14434f
C15368 XThC.Tn[10].t41 VGND 0.01593f
C15369 XThC.Tn[10].t37 VGND 0.0174f
C15370 XThC.Tn[10].n31 VGND 0.03884f
C15371 XThC.Tn[10].n32 VGND 0.02661f
C15372 XThC.Tn[10].n33 VGND 0.08758f
C15373 XThC.Tn[10].n34 VGND 0.14434f
C15374 XThC.Tn[10].t43 VGND 0.01593f
C15375 XThC.Tn[10].t39 VGND 0.0174f
C15376 XThC.Tn[10].n35 VGND 0.03884f
C15377 XThC.Tn[10].n36 VGND 0.02661f
C15378 XThC.Tn[10].n37 VGND 0.08758f
C15379 XThC.Tn[10].n38 VGND 0.14434f
C15380 XThC.Tn[10].t31 VGND 0.01593f
C15381 XThC.Tn[10].t26 VGND 0.0174f
C15382 XThC.Tn[10].n39 VGND 0.03884f
C15383 XThC.Tn[10].n40 VGND 0.02661f
C15384 XThC.Tn[10].n41 VGND 0.08758f
C15385 XThC.Tn[10].n42 VGND 0.14434f
C15386 XThC.Tn[10].t33 VGND 0.01593f
C15387 XThC.Tn[10].t27 VGND 0.0174f
C15388 XThC.Tn[10].n43 VGND 0.03884f
C15389 XThC.Tn[10].n44 VGND 0.02661f
C15390 XThC.Tn[10].n45 VGND 0.08758f
C15391 XThC.Tn[10].n46 VGND 0.14434f
C15392 XThC.Tn[10].t12 VGND 0.01593f
C15393 XThC.Tn[10].t40 VGND 0.0174f
C15394 XThC.Tn[10].n47 VGND 0.03884f
C15395 XThC.Tn[10].n48 VGND 0.02661f
C15396 XThC.Tn[10].n49 VGND 0.08758f
C15397 XThC.Tn[10].n50 VGND 0.14434f
C15398 XThC.Tn[10].t20 VGND 0.01593f
C15399 XThC.Tn[10].t16 VGND 0.0174f
C15400 XThC.Tn[10].n51 VGND 0.03884f
C15401 XThC.Tn[10].n52 VGND 0.02661f
C15402 XThC.Tn[10].n53 VGND 0.08758f
C15403 XThC.Tn[10].n54 VGND 0.14434f
C15404 XThC.Tn[10].t22 VGND 0.01593f
C15405 XThC.Tn[10].t19 VGND 0.0174f
C15406 XThC.Tn[10].n55 VGND 0.03884f
C15407 XThC.Tn[10].n56 VGND 0.02661f
C15408 XThC.Tn[10].n57 VGND 0.08758f
C15409 XThC.Tn[10].n58 VGND 0.14434f
C15410 XThC.Tn[10].t35 VGND 0.01593f
C15411 XThC.Tn[10].t32 VGND 0.0174f
C15412 XThC.Tn[10].n59 VGND 0.03884f
C15413 XThC.Tn[10].n60 VGND 0.02661f
C15414 XThC.Tn[10].n61 VGND 0.08758f
C15415 XThC.Tn[10].n62 VGND 0.14434f
C15416 XThC.Tn[10].t13 VGND 0.01593f
C15417 XThC.Tn[10].t42 VGND 0.0174f
C15418 XThC.Tn[10].n63 VGND 0.03884f
C15419 XThC.Tn[10].n64 VGND 0.02661f
C15420 XThC.Tn[10].n65 VGND 0.08758f
C15421 XThC.Tn[10].n66 VGND 0.14434f
C15422 XThC.Tn[10].n67 VGND 0.61921f
C15423 XThC.Tn[10].n68 VGND 0.2357f
C15424 XThC.Tn[10].t3 VGND 0.0201f
C15425 XThC.Tn[10].t8 VGND 0.0201f
C15426 XThC.Tn[10].n69 VGND 0.04342f
C15427 XThC.Tn[10].t5 VGND 0.0201f
C15428 XThC.Tn[10].t11 VGND 0.0201f
C15429 XThC.Tn[10].n70 VGND 0.06609f
C15430 XThC.Tn[10].n71 VGND 0.18363f
C15431 XThC.Tn[10].n72 VGND 0.02887f
C15432 XThC.Tn[10].t9 VGND 0.0201f
C15433 XThC.Tn[10].t10 VGND 0.0201f
C15434 XThC.Tn[10].n73 VGND 0.06102f
C15435 XThC.Tn[10].t0 VGND 0.0201f
C15436 XThC.Tn[10].t1 VGND 0.0201f
C15437 XThC.Tn[10].n74 VGND 0.04467f
C15438 XThC.Tn[10].n75 VGND 0.19884f
C15439 Iout.n0 VGND 0.23929f
C15440 Iout.n1 VGND 1.25122f
C15441 Iout.n2 VGND 0.23929f
C15442 Iout.n3 VGND 0.23929f
C15443 Iout.t58 VGND 0.02304f
C15444 Iout.n4 VGND 0.05124f
C15445 Iout.n5 VGND 0.20242f
C15446 Iout.n6 VGND 0.23929f
C15447 Iout.n7 VGND 1.25122f
C15448 Iout.n8 VGND 0.23929f
C15449 Iout.t244 VGND 0.02304f
C15450 Iout.n9 VGND 0.05124f
C15451 Iout.n10 VGND 0.20242f
C15452 Iout.n11 VGND 0.23929f
C15453 Iout.n12 VGND 1.25122f
C15454 Iout.n13 VGND 0.23929f
C15455 Iout.t162 VGND 0.02304f
C15456 Iout.n14 VGND 0.05124f
C15457 Iout.n15 VGND 0.20242f
C15458 Iout.n16 VGND 0.23929f
C15459 Iout.n17 VGND 1.25122f
C15460 Iout.n18 VGND 0.23929f
C15461 Iout.t142 VGND 0.02304f
C15462 Iout.n19 VGND 0.05124f
C15463 Iout.n20 VGND 0.20242f
C15464 Iout.n21 VGND 0.49611f
C15465 Iout.t150 VGND 0.02304f
C15466 Iout.n22 VGND 0.05124f
C15467 Iout.n23 VGND 0.29851f
C15468 Iout.n24 VGND 0.23929f
C15469 Iout.n25 VGND 0.23929f
C15470 Iout.n26 VGND 0.23929f
C15471 Iout.n27 VGND 0.23929f
C15472 Iout.n28 VGND 0.23929f
C15473 Iout.n29 VGND 0.23929f
C15474 Iout.n30 VGND 0.23929f
C15475 Iout.n31 VGND 0.23929f
C15476 Iout.n32 VGND 0.23929f
C15477 Iout.n33 VGND 0.23929f
C15478 Iout.n34 VGND 0.23929f
C15479 Iout.n35 VGND 0.23929f
C15480 Iout.n36 VGND 0.23929f
C15481 Iout.n37 VGND 0.23929f
C15482 Iout.t59 VGND 0.02304f
C15483 Iout.n38 VGND 0.05124f
C15484 Iout.n39 VGND 0.02606f
C15485 Iout.n40 VGND 0.23929f
C15486 Iout.n41 VGND 0.04775f
C15487 Iout.t125 VGND 0.02304f
C15488 Iout.n42 VGND 0.05124f
C15489 Iout.n43 VGND 0.02606f
C15490 Iout.t215 VGND 0.02304f
C15491 Iout.n44 VGND 0.05124f
C15492 Iout.n45 VGND 0.02606f
C15493 Iout.n46 VGND 0.23929f
C15494 Iout.t227 VGND 0.02304f
C15495 Iout.n47 VGND 0.05124f
C15496 Iout.n48 VGND 0.02606f
C15497 Iout.n49 VGND 0.23929f
C15498 Iout.t209 VGND 0.02304f
C15499 Iout.n50 VGND 0.05124f
C15500 Iout.n51 VGND 0.02606f
C15501 Iout.n52 VGND 0.23929f
C15502 Iout.t205 VGND 0.02304f
C15503 Iout.n53 VGND 0.05124f
C15504 Iout.n54 VGND 0.02606f
C15505 Iout.n55 VGND 0.23929f
C15506 Iout.t109 VGND 0.02304f
C15507 Iout.n56 VGND 0.05124f
C15508 Iout.n57 VGND 0.02606f
C15509 Iout.n58 VGND 0.23929f
C15510 Iout.t185 VGND 0.02304f
C15511 Iout.n59 VGND 0.05124f
C15512 Iout.n60 VGND 0.02606f
C15513 Iout.n61 VGND 0.23929f
C15514 Iout.t27 VGND 0.02304f
C15515 Iout.n62 VGND 0.05124f
C15516 Iout.n63 VGND 0.02606f
C15517 Iout.n64 VGND 0.23929f
C15518 Iout.t224 VGND 0.02304f
C15519 Iout.n65 VGND 0.05124f
C15520 Iout.n66 VGND 0.02606f
C15521 Iout.n67 VGND 0.23929f
C15522 Iout.t179 VGND 0.02304f
C15523 Iout.n68 VGND 0.05124f
C15524 Iout.n69 VGND 0.02606f
C15525 Iout.n70 VGND 0.23929f
C15526 Iout.t83 VGND 0.02304f
C15527 Iout.n71 VGND 0.05124f
C15528 Iout.n72 VGND 0.02606f
C15529 Iout.n73 VGND 0.23929f
C15530 Iout.t24 VGND 0.02304f
C15531 Iout.n74 VGND 0.05124f
C15532 Iout.n75 VGND 0.02606f
C15533 Iout.n76 VGND 0.23929f
C15534 Iout.t194 VGND 0.02304f
C15535 Iout.n77 VGND 0.05124f
C15536 Iout.n78 VGND 0.02606f
C15537 Iout.n79 VGND 0.23929f
C15538 Iout.n80 VGND 0.23929f
C15539 Iout.t62 VGND 0.02304f
C15540 Iout.n81 VGND 0.05124f
C15541 Iout.n82 VGND 0.02606f
C15542 Iout.n83 VGND 0.23929f
C15543 Iout.n84 VGND 0.04775f
C15544 Iout.t41 VGND 0.02304f
C15545 Iout.n85 VGND 0.05124f
C15546 Iout.n86 VGND 0.02606f
C15547 Iout.t18 VGND 0.02304f
C15548 Iout.n87 VGND 0.05124f
C15549 Iout.n88 VGND 0.02606f
C15550 Iout.n89 VGND 0.23929f
C15551 Iout.t113 VGND 0.02304f
C15552 Iout.n90 VGND 0.05124f
C15553 Iout.n91 VGND 0.02606f
C15554 Iout.n92 VGND 0.23929f
C15555 Iout.t36 VGND 0.02304f
C15556 Iout.n93 VGND 0.05124f
C15557 Iout.n94 VGND 0.02606f
C15558 Iout.n95 VGND 0.23929f
C15559 Iout.t112 VGND 0.02304f
C15560 Iout.n96 VGND 0.05124f
C15561 Iout.n97 VGND 0.02606f
C15562 Iout.n98 VGND 0.23929f
C15563 Iout.t249 VGND 0.02304f
C15564 Iout.n99 VGND 0.05124f
C15565 Iout.n100 VGND 0.02606f
C15566 Iout.n101 VGND 0.23929f
C15567 Iout.t156 VGND 0.02304f
C15568 Iout.n102 VGND 0.05124f
C15569 Iout.n103 VGND 0.02606f
C15570 Iout.n104 VGND 0.23929f
C15571 Iout.t237 VGND 0.02304f
C15572 Iout.n105 VGND 0.05124f
C15573 Iout.n106 VGND 0.02606f
C15574 Iout.n107 VGND 0.23929f
C15575 Iout.t229 VGND 0.02304f
C15576 Iout.n108 VGND 0.05124f
C15577 Iout.n109 VGND 0.02606f
C15578 Iout.n110 VGND 0.23929f
C15579 Iout.t255 VGND 0.02304f
C15580 Iout.n111 VGND 0.05124f
C15581 Iout.n112 VGND 0.02606f
C15582 Iout.n113 VGND 0.23929f
C15583 Iout.t216 VGND 0.02304f
C15584 Iout.n114 VGND 0.05124f
C15585 Iout.n115 VGND 0.02606f
C15586 Iout.n116 VGND 0.23929f
C15587 Iout.t206 VGND 0.02304f
C15588 Iout.n117 VGND 0.05124f
C15589 Iout.n118 VGND 0.02606f
C15590 Iout.n119 VGND 0.23929f
C15591 Iout.t164 VGND 0.02304f
C15592 Iout.n120 VGND 0.05124f
C15593 Iout.n121 VGND 0.02606f
C15594 Iout.n122 VGND 0.04775f
C15595 Iout.t220 VGND 0.02304f
C15596 Iout.n123 VGND 0.05124f
C15597 Iout.n124 VGND 0.02606f
C15598 Iout.n125 VGND 0.23929f
C15599 Iout.n126 VGND 0.23929f
C15600 Iout.t139 VGND 0.02304f
C15601 Iout.n127 VGND 0.05124f
C15602 Iout.n128 VGND 0.02606f
C15603 Iout.n129 VGND 0.04775f
C15604 Iout.t103 VGND 0.02304f
C15605 Iout.n130 VGND 0.05124f
C15606 Iout.n131 VGND 0.02606f
C15607 Iout.n132 VGND 0.23929f
C15608 Iout.t21 VGND 0.02304f
C15609 Iout.n133 VGND 0.05124f
C15610 Iout.n134 VGND 0.02606f
C15611 Iout.n135 VGND 0.04775f
C15612 Iout.t100 VGND 0.02304f
C15613 Iout.n136 VGND 0.05124f
C15614 Iout.n137 VGND 0.02606f
C15615 Iout.n138 VGND 0.23929f
C15616 Iout.n139 VGND 0.23929f
C15617 Iout.t118 VGND 0.02304f
C15618 Iout.n140 VGND 0.05124f
C15619 Iout.n141 VGND 0.02606f
C15620 Iout.n142 VGND 0.04775f
C15621 Iout.t64 VGND 0.02304f
C15622 Iout.n143 VGND 0.05124f
C15623 Iout.n144 VGND 0.02606f
C15624 Iout.n145 VGND 0.14126f
C15625 Iout.t79 VGND 0.02304f
C15626 Iout.n146 VGND 0.05124f
C15627 Iout.n147 VGND 0.02606f
C15628 Iout.n148 VGND 0.04775f
C15629 Iout.t16 VGND 0.02304f
C15630 Iout.n149 VGND 0.05124f
C15631 Iout.n150 VGND 0.02606f
C15632 Iout.n151 VGND 0.23929f
C15633 Iout.n152 VGND 0.14126f
C15634 Iout.n153 VGND 0.23929f
C15635 Iout.n154 VGND 0.23929f
C15636 Iout.n155 VGND 0.23929f
C15637 Iout.t72 VGND 0.02304f
C15638 Iout.n156 VGND 0.05124f
C15639 Iout.n157 VGND 0.02606f
C15640 Iout.n158 VGND 0.23929f
C15641 Iout.n159 VGND 0.23929f
C15642 Iout.n160 VGND 0.23929f
C15643 Iout.n161 VGND 0.23929f
C15644 Iout.n162 VGND 0.23929f
C15645 Iout.n163 VGND 0.23929f
C15646 Iout.n164 VGND 0.23929f
C15647 Iout.n165 VGND 0.23929f
C15648 Iout.n166 VGND 0.23929f
C15649 Iout.n167 VGND 0.23929f
C15650 Iout.t239 VGND 0.02304f
C15651 Iout.n168 VGND 0.05124f
C15652 Iout.n169 VGND 0.02606f
C15653 Iout.n170 VGND 0.23929f
C15654 Iout.n171 VGND 0.04775f
C15655 Iout.t154 VGND 0.02304f
C15656 Iout.n172 VGND 0.05124f
C15657 Iout.n173 VGND 0.02606f
C15658 Iout.t137 VGND 0.02304f
C15659 Iout.n174 VGND 0.05124f
C15660 Iout.n175 VGND 0.02606f
C15661 Iout.n176 VGND 0.23929f
C15662 Iout.t1 VGND 0.02304f
C15663 Iout.n177 VGND 0.05124f
C15664 Iout.n178 VGND 0.02606f
C15665 Iout.n179 VGND 0.23929f
C15666 Iout.t235 VGND 0.02304f
C15667 Iout.n180 VGND 0.05124f
C15668 Iout.n181 VGND 0.02606f
C15669 Iout.n182 VGND 0.23929f
C15670 Iout.t88 VGND 0.02304f
C15671 Iout.n183 VGND 0.05124f
C15672 Iout.n184 VGND 0.02606f
C15673 Iout.n185 VGND 0.23929f
C15674 Iout.t33 VGND 0.02304f
C15675 Iout.n186 VGND 0.05124f
C15676 Iout.n187 VGND 0.02606f
C15677 Iout.n188 VGND 0.23929f
C15678 Iout.t182 VGND 0.02304f
C15679 Iout.n189 VGND 0.05124f
C15680 Iout.n190 VGND 0.02606f
C15681 Iout.n191 VGND 0.14126f
C15682 Iout.t233 VGND 0.02304f
C15683 Iout.n192 VGND 0.05124f
C15684 Iout.n193 VGND 0.02606f
C15685 Iout.n194 VGND 0.04775f
C15686 Iout.t167 VGND 0.02304f
C15687 Iout.n195 VGND 0.05124f
C15688 Iout.n196 VGND 0.02606f
C15689 Iout.n197 VGND 0.14126f
C15690 Iout.n198 VGND 0.04775f
C15691 Iout.t57 VGND 0.02304f
C15692 Iout.n199 VGND 0.05124f
C15693 Iout.n200 VGND 0.02606f
C15694 Iout.n201 VGND 0.04775f
C15695 Iout.t19 VGND 0.02304f
C15696 Iout.n202 VGND 0.05124f
C15697 Iout.n203 VGND 0.02606f
C15698 Iout.n204 VGND 0.14126f
C15699 Iout.n205 VGND 0.04775f
C15700 Iout.t226 VGND 0.02304f
C15701 Iout.n206 VGND 0.05124f
C15702 Iout.n207 VGND 0.02606f
C15703 Iout.n208 VGND 0.14126f
C15704 Iout.n209 VGND 0.04775f
C15705 Iout.t131 VGND 0.02304f
C15706 Iout.n210 VGND 0.05124f
C15707 Iout.n211 VGND 0.02606f
C15708 Iout.n212 VGND 0.14126f
C15709 Iout.n213 VGND 0.04775f
C15710 Iout.t91 VGND 0.02304f
C15711 Iout.n214 VGND 0.05124f
C15712 Iout.n215 VGND 0.02606f
C15713 Iout.n216 VGND 0.14126f
C15714 Iout.n217 VGND 0.04775f
C15715 Iout.t146 VGND 0.02304f
C15716 Iout.n218 VGND 0.05124f
C15717 Iout.n219 VGND 0.02606f
C15718 Iout.n220 VGND 0.14126f
C15719 Iout.n221 VGND 0.04775f
C15720 Iout.t32 VGND 0.02304f
C15721 Iout.n222 VGND 0.05124f
C15722 Iout.n223 VGND 0.02606f
C15723 Iout.n224 VGND 0.14126f
C15724 Iout.n225 VGND 0.04775f
C15725 Iout.t117 VGND 0.02304f
C15726 Iout.n226 VGND 0.05124f
C15727 Iout.n227 VGND 0.02606f
C15728 Iout.n228 VGND 0.04775f
C15729 Iout.n229 VGND 0.14126f
C15730 Iout.n230 VGND 0.23929f
C15731 Iout.n231 VGND 0.04775f
C15732 Iout.t172 VGND 0.02304f
C15733 Iout.n232 VGND 0.05124f
C15734 Iout.n233 VGND 0.02606f
C15735 Iout.n234 VGND 0.04775f
C15736 Iout.t178 VGND 0.02304f
C15737 Iout.n235 VGND 0.05124f
C15738 Iout.n236 VGND 0.02606f
C15739 Iout.n237 VGND 0.04775f
C15740 Iout.t3 VGND 0.02304f
C15741 Iout.n238 VGND 0.05124f
C15742 Iout.n239 VGND 0.02606f
C15743 Iout.n240 VGND 0.04775f
C15744 Iout.t119 VGND 0.02304f
C15745 Iout.n241 VGND 0.05124f
C15746 Iout.n242 VGND 0.02606f
C15747 Iout.n243 VGND 0.04775f
C15748 Iout.t50 VGND 0.02304f
C15749 Iout.n244 VGND 0.05124f
C15750 Iout.n245 VGND 0.02606f
C15751 Iout.n246 VGND 0.04775f
C15752 Iout.t13 VGND 0.02304f
C15753 Iout.n247 VGND 0.05124f
C15754 Iout.n248 VGND 0.02606f
C15755 Iout.n249 VGND 0.04775f
C15756 Iout.t5 VGND 0.02304f
C15757 Iout.n250 VGND 0.05124f
C15758 Iout.n251 VGND 0.02606f
C15759 Iout.t99 VGND 0.02304f
C15760 Iout.n252 VGND 0.05124f
C15761 Iout.n253 VGND 0.02606f
C15762 Iout.n254 VGND 0.04775f
C15763 Iout.t157 VGND 0.02304f
C15764 Iout.n255 VGND 0.05124f
C15765 Iout.n256 VGND 0.02606f
C15766 Iout.n257 VGND 0.04775f
C15767 Iout.n258 VGND 0.23929f
C15768 Iout.t147 VGND 0.02304f
C15769 Iout.n259 VGND 0.05124f
C15770 Iout.n260 VGND 0.02606f
C15771 Iout.n261 VGND 0.04775f
C15772 Iout.n262 VGND 0.23929f
C15773 Iout.n263 VGND 0.23929f
C15774 Iout.n264 VGND 0.04775f
C15775 Iout.t238 VGND 0.02304f
C15776 Iout.n265 VGND 0.05124f
C15777 Iout.n266 VGND 0.02606f
C15778 Iout.n267 VGND 0.04775f
C15779 Iout.n268 VGND 0.23929f
C15780 Iout.n269 VGND 0.23929f
C15781 Iout.n270 VGND 0.04775f
C15782 Iout.t107 VGND 0.02304f
C15783 Iout.n271 VGND 0.05124f
C15784 Iout.n272 VGND 0.02606f
C15785 Iout.n273 VGND 0.04775f
C15786 Iout.n274 VGND 0.23929f
C15787 Iout.n275 VGND 0.23929f
C15788 Iout.n276 VGND 0.04775f
C15789 Iout.t53 VGND 0.02304f
C15790 Iout.n277 VGND 0.05124f
C15791 Iout.n278 VGND 0.02606f
C15792 Iout.n279 VGND 0.04775f
C15793 Iout.n280 VGND 0.23929f
C15794 Iout.n281 VGND 0.23929f
C15795 Iout.n282 VGND 0.04775f
C15796 Iout.t225 VGND 0.02304f
C15797 Iout.n283 VGND 0.05124f
C15798 Iout.n284 VGND 0.02606f
C15799 Iout.n285 VGND 0.04775f
C15800 Iout.n286 VGND 0.23929f
C15801 Iout.n287 VGND 0.23929f
C15802 Iout.n288 VGND 0.04775f
C15803 Iout.t222 VGND 0.02304f
C15804 Iout.n289 VGND 0.05124f
C15805 Iout.n290 VGND 0.02606f
C15806 Iout.n291 VGND 0.04775f
C15807 Iout.n292 VGND 0.23929f
C15808 Iout.n293 VGND 0.23929f
C15809 Iout.n294 VGND 0.04775f
C15810 Iout.t81 VGND 0.02304f
C15811 Iout.n295 VGND 0.05124f
C15812 Iout.n296 VGND 0.02606f
C15813 Iout.n297 VGND 0.04775f
C15814 Iout.n298 VGND 0.23929f
C15815 Iout.n299 VGND 0.23929f
C15816 Iout.n300 VGND 0.04775f
C15817 Iout.t74 VGND 0.02304f
C15818 Iout.n301 VGND 0.05124f
C15819 Iout.n302 VGND 0.02606f
C15820 Iout.n303 VGND 0.04775f
C15821 Iout.n304 VGND 0.23929f
C15822 Iout.t102 VGND 0.02304f
C15823 Iout.n305 VGND 0.05124f
C15824 Iout.n306 VGND 0.02606f
C15825 Iout.n307 VGND 0.04775f
C15826 Iout.t87 VGND 0.02304f
C15827 Iout.n308 VGND 0.05124f
C15828 Iout.n309 VGND 0.02606f
C15829 Iout.n310 VGND 0.04775f
C15830 Iout.t175 VGND 0.02304f
C15831 Iout.n311 VGND 0.05124f
C15832 Iout.n312 VGND 0.02606f
C15833 Iout.n313 VGND 0.04775f
C15834 Iout.t204 VGND 0.02304f
C15835 Iout.n314 VGND 0.05124f
C15836 Iout.n315 VGND 0.02606f
C15837 Iout.n316 VGND 0.04775f
C15838 Iout.t28 VGND 0.02304f
C15839 Iout.n317 VGND 0.05124f
C15840 Iout.n318 VGND 0.02606f
C15841 Iout.n319 VGND 0.04775f
C15842 Iout.t94 VGND 0.02304f
C15843 Iout.n320 VGND 0.05124f
C15844 Iout.n321 VGND 0.02606f
C15845 Iout.n322 VGND 0.04775f
C15846 Iout.t134 VGND 0.02304f
C15847 Iout.n323 VGND 0.05124f
C15848 Iout.n324 VGND 0.02606f
C15849 Iout.n325 VGND 0.04775f
C15850 Iout.t55 VGND 0.02304f
C15851 Iout.n326 VGND 0.05124f
C15852 Iout.n327 VGND 0.02606f
C15853 Iout.n328 VGND 0.04775f
C15854 Iout.t254 VGND 0.02304f
C15855 Iout.n329 VGND 0.05124f
C15856 Iout.n330 VGND 0.02606f
C15857 Iout.n331 VGND 0.04775f
C15858 Iout.n332 VGND 0.23929f
C15859 Iout.t191 VGND 0.02304f
C15860 Iout.n333 VGND 0.05124f
C15861 Iout.n334 VGND 0.02606f
C15862 Iout.n335 VGND 0.04775f
C15863 Iout.t253 VGND 0.02304f
C15864 Iout.n336 VGND 0.05124f
C15865 Iout.n337 VGND 0.02606f
C15866 Iout.n338 VGND 0.04775f
C15867 Iout.t223 VGND 0.02304f
C15868 Iout.n339 VGND 0.05124f
C15869 Iout.n340 VGND 0.02606f
C15870 Iout.n341 VGND 0.04775f
C15871 Iout.t124 VGND 0.02304f
C15872 Iout.n342 VGND 0.05124f
C15873 Iout.n343 VGND 0.02606f
C15874 Iout.n344 VGND 0.04775f
C15875 Iout.t207 VGND 0.02304f
C15876 Iout.n345 VGND 0.05124f
C15877 Iout.n346 VGND 0.02606f
C15878 Iout.n347 VGND 0.04775f
C15879 Iout.t26 VGND 0.02304f
C15880 Iout.n348 VGND 0.05124f
C15881 Iout.n349 VGND 0.02606f
C15882 Iout.n350 VGND 0.04775f
C15883 Iout.t108 VGND 0.02304f
C15884 Iout.n351 VGND 0.05124f
C15885 Iout.n352 VGND 0.02606f
C15886 Iout.n353 VGND 0.04775f
C15887 Iout.t136 VGND 0.02304f
C15888 Iout.n354 VGND 0.05124f
C15889 Iout.n355 VGND 0.02606f
C15890 Iout.n356 VGND 0.04775f
C15891 Iout.t252 VGND 0.02304f
C15892 Iout.n357 VGND 0.05124f
C15893 Iout.n358 VGND 0.02606f
C15894 Iout.n359 VGND 0.04775f
C15895 Iout.t158 VGND 0.02304f
C15896 Iout.n360 VGND 0.05124f
C15897 Iout.n361 VGND 0.02606f
C15898 Iout.n362 VGND 0.04775f
C15899 Iout.t148 VGND 0.02304f
C15900 Iout.n363 VGND 0.05124f
C15901 Iout.n364 VGND 0.02606f
C15902 Iout.n365 VGND 0.04775f
C15903 Iout.t89 VGND 0.02304f
C15904 Iout.n366 VGND 0.05124f
C15905 Iout.n367 VGND 0.02606f
C15906 Iout.n368 VGND 0.04775f
C15907 Iout.n369 VGND 0.23929f
C15908 Iout.t217 VGND 0.02304f
C15909 Iout.n370 VGND 0.05124f
C15910 Iout.n371 VGND 0.02606f
C15911 Iout.n372 VGND 0.04775f
C15912 Iout.n373 VGND 0.23929f
C15913 Iout.n374 VGND 0.23929f
C15914 Iout.n375 VGND 0.04775f
C15915 Iout.t231 VGND 0.02304f
C15916 Iout.n376 VGND 0.05124f
C15917 Iout.n377 VGND 0.02606f
C15918 Iout.t38 VGND 0.02304f
C15919 Iout.n378 VGND 0.05124f
C15920 Iout.n379 VGND 0.02606f
C15921 Iout.n380 VGND 0.04775f
C15922 Iout.n381 VGND 0.23929f
C15923 Iout.n382 VGND 0.23929f
C15924 Iout.n383 VGND 0.04775f
C15925 Iout.t170 VGND 0.02304f
C15926 Iout.n384 VGND 0.05124f
C15927 Iout.n385 VGND 0.02606f
C15928 Iout.t66 VGND 0.02304f
C15929 Iout.n386 VGND 0.05124f
C15930 Iout.n387 VGND 0.02606f
C15931 Iout.n388 VGND 0.04775f
C15932 Iout.n389 VGND 0.23929f
C15933 Iout.n390 VGND 0.23929f
C15934 Iout.n391 VGND 0.04775f
C15935 Iout.t247 VGND 0.02304f
C15936 Iout.n392 VGND 0.05124f
C15937 Iout.n393 VGND 0.02606f
C15938 Iout.t7 VGND 0.02304f
C15939 Iout.n394 VGND 0.05124f
C15940 Iout.n395 VGND 0.02606f
C15941 Iout.n396 VGND 0.04775f
C15942 Iout.n397 VGND 0.23929f
C15943 Iout.n398 VGND 0.23929f
C15944 Iout.n399 VGND 0.04775f
C15945 Iout.t128 VGND 0.02304f
C15946 Iout.n400 VGND 0.05124f
C15947 Iout.n401 VGND 0.02606f
C15948 Iout.t196 VGND 0.02304f
C15949 Iout.n402 VGND 0.05124f
C15950 Iout.n403 VGND 0.02606f
C15951 Iout.n404 VGND 0.04775f
C15952 Iout.n405 VGND 0.23929f
C15953 Iout.n406 VGND 0.23929f
C15954 Iout.n407 VGND 0.04775f
C15955 Iout.t10 VGND 0.02304f
C15956 Iout.n408 VGND 0.05124f
C15957 Iout.n409 VGND 0.02606f
C15958 Iout.t135 VGND 0.02304f
C15959 Iout.n410 VGND 0.05124f
C15960 Iout.n411 VGND 0.02606f
C15961 Iout.n412 VGND 0.04775f
C15962 Iout.n413 VGND 0.23929f
C15963 Iout.n414 VGND 0.23929f
C15964 Iout.n415 VGND 0.04775f
C15965 Iout.t132 VGND 0.02304f
C15966 Iout.n416 VGND 0.05124f
C15967 Iout.n417 VGND 0.02606f
C15968 Iout.t143 VGND 0.02304f
C15969 Iout.n418 VGND 0.05124f
C15970 Iout.n419 VGND 0.02606f
C15971 Iout.n420 VGND 0.04775f
C15972 Iout.n421 VGND 0.23929f
C15973 Iout.n422 VGND 0.23929f
C15974 Iout.n423 VGND 0.04775f
C15975 Iout.t105 VGND 0.02304f
C15976 Iout.n424 VGND 0.05124f
C15977 Iout.n425 VGND 0.02606f
C15978 Iout.t45 VGND 0.02304f
C15979 Iout.n426 VGND 0.05124f
C15980 Iout.n427 VGND 0.02606f
C15981 Iout.n428 VGND 0.04775f
C15982 Iout.n429 VGND 0.23929f
C15983 Iout.n430 VGND 0.23929f
C15984 Iout.n431 VGND 0.04775f
C15985 Iout.t240 VGND 0.02304f
C15986 Iout.n432 VGND 0.05124f
C15987 Iout.n433 VGND 0.02606f
C15988 Iout.t140 VGND 0.02304f
C15989 Iout.n434 VGND 0.05124f
C15990 Iout.n435 VGND 0.02606f
C15991 Iout.n436 VGND 0.23929f
C15992 Iout.n437 VGND 0.04775f
C15993 Iout.t192 VGND 0.02304f
C15994 Iout.n438 VGND 0.05124f
C15995 Iout.n439 VGND 0.02606f
C15996 Iout.n440 VGND 0.04775f
C15997 Iout.t213 VGND 0.02304f
C15998 Iout.n441 VGND 0.05124f
C15999 Iout.n442 VGND 0.02606f
C16000 Iout.n443 VGND 0.04775f
C16001 Iout.n444 VGND 0.23929f
C16002 Iout.n445 VGND 0.23929f
C16003 Iout.n446 VGND 0.04775f
C16004 Iout.t67 VGND 0.02304f
C16005 Iout.n447 VGND 0.05124f
C16006 Iout.n448 VGND 0.02606f
C16007 Iout.t127 VGND 0.02304f
C16008 Iout.n449 VGND 0.05124f
C16009 Iout.n450 VGND 0.02606f
C16010 Iout.n451 VGND 0.04775f
C16011 Iout.t248 VGND 0.02304f
C16012 Iout.n452 VGND 0.05124f
C16013 Iout.n453 VGND 0.02606f
C16014 Iout.n454 VGND 0.04775f
C16015 Iout.n455 VGND 0.23929f
C16016 Iout.n456 VGND 0.23929f
C16017 Iout.n457 VGND 0.04775f
C16018 Iout.t241 VGND 0.02304f
C16019 Iout.n458 VGND 0.05124f
C16020 Iout.n459 VGND 0.02606f
C16021 Iout.t188 VGND 0.02304f
C16022 Iout.n460 VGND 0.05124f
C16023 Iout.n461 VGND 0.02606f
C16024 Iout.n462 VGND 0.04775f
C16025 Iout.t20 VGND 0.02304f
C16026 Iout.n463 VGND 0.05124f
C16027 Iout.n464 VGND 0.02606f
C16028 Iout.n465 VGND 0.04775f
C16029 Iout.n466 VGND 0.23929f
C16030 Iout.n467 VGND 0.23929f
C16031 Iout.n468 VGND 0.04775f
C16032 Iout.t77 VGND 0.02304f
C16033 Iout.n469 VGND 0.05124f
C16034 Iout.n470 VGND 0.02606f
C16035 Iout.n471 VGND 0.04775f
C16036 Iout.t149 VGND 0.02304f
C16037 Iout.n472 VGND 0.05124f
C16038 Iout.n473 VGND 0.02606f
C16039 Iout.n474 VGND 0.04775f
C16040 Iout.n475 VGND 0.23929f
C16041 Iout.n476 VGND 0.23929f
C16042 Iout.n477 VGND 0.04775f
C16043 Iout.t17 VGND 0.02304f
C16044 Iout.n478 VGND 0.05124f
C16045 Iout.n479 VGND 0.02606f
C16046 Iout.t186 VGND 0.02304f
C16047 Iout.n480 VGND 0.05124f
C16048 Iout.n481 VGND 0.02606f
C16049 Iout.n482 VGND 0.04775f
C16050 Iout.t169 VGND 0.02304f
C16051 Iout.n483 VGND 0.05124f
C16052 Iout.n484 VGND 0.02606f
C16053 Iout.n485 VGND 0.04775f
C16054 Iout.n486 VGND 0.23929f
C16055 Iout.n487 VGND 0.23929f
C16056 Iout.n488 VGND 0.04775f
C16057 Iout.t8 VGND 0.02304f
C16058 Iout.n489 VGND 0.05124f
C16059 Iout.n490 VGND 0.02606f
C16060 Iout.t145 VGND 0.02304f
C16061 Iout.n491 VGND 0.05124f
C16062 Iout.n492 VGND 0.02606f
C16063 Iout.n493 VGND 0.04775f
C16064 Iout.t197 VGND 0.02304f
C16065 Iout.n494 VGND 0.05124f
C16066 Iout.n495 VGND 0.02606f
C16067 Iout.n496 VGND 0.04775f
C16068 Iout.n497 VGND 0.23929f
C16069 Iout.n498 VGND 0.14126f
C16070 Iout.n499 VGND 0.04775f
C16071 Iout.t23 VGND 0.02304f
C16072 Iout.n500 VGND 0.05124f
C16073 Iout.n501 VGND 0.02606f
C16074 Iout.n502 VGND 0.14126f
C16075 Iout.n503 VGND 0.04775f
C16076 Iout.t115 VGND 0.02304f
C16077 Iout.n504 VGND 0.05124f
C16078 Iout.n505 VGND 0.02606f
C16079 Iout.n506 VGND 0.04775f
C16080 Iout.t171 VGND 0.02304f
C16081 Iout.n507 VGND 0.05124f
C16082 Iout.n508 VGND 0.02606f
C16083 Iout.t98 VGND 0.02304f
C16084 Iout.n509 VGND 0.05124f
C16085 Iout.n510 VGND 0.02606f
C16086 Iout.n511 VGND 0.14126f
C16087 Iout.n512 VGND 0.04775f
C16088 Iout.t130 VGND 0.02304f
C16089 Iout.n513 VGND 0.05124f
C16090 Iout.n514 VGND 0.02606f
C16091 Iout.n515 VGND 0.04775f
C16092 Iout.n516 VGND 0.14126f
C16093 Iout.n517 VGND 0.23929f
C16094 Iout.n518 VGND 0.04775f
C16095 Iout.t212 VGND 0.02304f
C16096 Iout.n519 VGND 0.05124f
C16097 Iout.n520 VGND 0.02606f
C16098 Iout.n521 VGND 0.04775f
C16099 Iout.n522 VGND 0.23929f
C16100 Iout.n523 VGND 0.23929f
C16101 Iout.n524 VGND 0.04775f
C16102 Iout.t22 VGND 0.02304f
C16103 Iout.n525 VGND 0.05124f
C16104 Iout.n526 VGND 0.02606f
C16105 Iout.n527 VGND 0.04775f
C16106 Iout.n528 VGND 0.23929f
C16107 Iout.n529 VGND 0.23929f
C16108 Iout.n530 VGND 0.04775f
C16109 Iout.t35 VGND 0.02304f
C16110 Iout.n531 VGND 0.05124f
C16111 Iout.n532 VGND 0.02606f
C16112 Iout.n533 VGND 0.04775f
C16113 Iout.t111 VGND 0.02304f
C16114 Iout.n534 VGND 0.05124f
C16115 Iout.n535 VGND 0.02606f
C16116 Iout.t92 VGND 0.02304f
C16117 Iout.n536 VGND 0.05124f
C16118 Iout.n537 VGND 0.02606f
C16119 Iout.n538 VGND 0.04775f
C16120 Iout.n539 VGND 0.23929f
C16121 Iout.n540 VGND 0.23929f
C16122 Iout.n541 VGND 0.04775f
C16123 Iout.t123 VGND 0.02304f
C16124 Iout.n542 VGND 0.05124f
C16125 Iout.n543 VGND 0.02606f
C16126 Iout.n544 VGND 0.04775f
C16127 Iout.n545 VGND 0.23929f
C16128 Iout.n546 VGND 0.23929f
C16129 Iout.n547 VGND 0.04775f
C16130 Iout.t54 VGND 0.02304f
C16131 Iout.n548 VGND 0.05124f
C16132 Iout.n549 VGND 0.02606f
C16133 Iout.n550 VGND 0.04775f
C16134 Iout.n551 VGND 0.23929f
C16135 Iout.n552 VGND 0.23929f
C16136 Iout.n553 VGND 0.04775f
C16137 Iout.t195 VGND 0.02304f
C16138 Iout.n554 VGND 0.05124f
C16139 Iout.n555 VGND 0.02606f
C16140 Iout.n556 VGND 0.04775f
C16141 Iout.t114 VGND 0.02304f
C16142 Iout.n557 VGND 0.05124f
C16143 Iout.n558 VGND 0.02606f
C16144 Iout.t63 VGND 0.02304f
C16145 Iout.n559 VGND 0.05124f
C16146 Iout.n560 VGND 0.02606f
C16147 Iout.n561 VGND 0.04775f
C16148 Iout.n562 VGND 0.23929f
C16149 Iout.t96 VGND 0.02304f
C16150 Iout.n563 VGND 0.05124f
C16151 Iout.n564 VGND 0.02606f
C16152 Iout.n565 VGND 0.04775f
C16153 Iout.n566 VGND 0.23929f
C16154 Iout.n567 VGND 0.23929f
C16155 Iout.n568 VGND 0.04775f
C16156 Iout.t86 VGND 0.02304f
C16157 Iout.n569 VGND 0.05124f
C16158 Iout.n570 VGND 0.02606f
C16159 Iout.n571 VGND 0.04775f
C16160 Iout.n572 VGND 0.23929f
C16161 Iout.t187 VGND 0.02304f
C16162 Iout.n573 VGND 0.05124f
C16163 Iout.n574 VGND 0.02606f
C16164 Iout.n575 VGND 0.04775f
C16165 Iout.t198 VGND 0.02304f
C16166 Iout.n576 VGND 0.05124f
C16167 Iout.n577 VGND 0.02606f
C16168 Iout.n578 VGND 0.04775f
C16169 Iout.n579 VGND 0.23929f
C16170 Iout.n580 VGND 0.23929f
C16171 Iout.n581 VGND 0.04775f
C16172 Iout.t184 VGND 0.02304f
C16173 Iout.n582 VGND 0.05124f
C16174 Iout.n583 VGND 0.02606f
C16175 Iout.n584 VGND 0.04775f
C16176 Iout.n585 VGND 0.23929f
C16177 Iout.n586 VGND 0.23929f
C16178 Iout.n587 VGND 0.04775f
C16179 Iout.t30 VGND 0.02304f
C16180 Iout.n588 VGND 0.05124f
C16181 Iout.n589 VGND 0.02606f
C16182 Iout.n590 VGND 0.04775f
C16183 Iout.n591 VGND 0.23929f
C16184 Iout.n592 VGND 0.23929f
C16185 Iout.n593 VGND 0.04775f
C16186 Iout.t71 VGND 0.02304f
C16187 Iout.n594 VGND 0.05124f
C16188 Iout.n595 VGND 0.02606f
C16189 Iout.n596 VGND 0.04775f
C16190 Iout.n597 VGND 0.23929f
C16191 Iout.n598 VGND 0.23929f
C16192 Iout.n599 VGND 0.04775f
C16193 Iout.t78 VGND 0.02304f
C16194 Iout.n600 VGND 0.05124f
C16195 Iout.n601 VGND 0.02606f
C16196 Iout.n602 VGND 0.04775f
C16197 Iout.n603 VGND 0.23929f
C16198 Iout.n604 VGND 0.23929f
C16199 Iout.n605 VGND 0.04775f
C16200 Iout.t101 VGND 0.02304f
C16201 Iout.n606 VGND 0.05124f
C16202 Iout.n607 VGND 0.02606f
C16203 Iout.n608 VGND 0.04775f
C16204 Iout.n609 VGND 0.23929f
C16205 Iout.n610 VGND 0.23929f
C16206 Iout.n611 VGND 0.04775f
C16207 Iout.t61 VGND 0.02304f
C16208 Iout.n612 VGND 0.05124f
C16209 Iout.n613 VGND 0.02606f
C16210 Iout.n614 VGND 0.04775f
C16211 Iout.n615 VGND 0.23929f
C16212 Iout.n616 VGND 0.23929f
C16213 Iout.n617 VGND 0.04775f
C16214 Iout.t160 VGND 0.02304f
C16215 Iout.n618 VGND 0.05124f
C16216 Iout.n619 VGND 0.02606f
C16217 Iout.n620 VGND 0.04775f
C16218 Iout.n621 VGND 0.23929f
C16219 Iout.n622 VGND 0.23929f
C16220 Iout.n623 VGND 0.04775f
C16221 Iout.t168 VGND 0.02304f
C16222 Iout.n624 VGND 0.05124f
C16223 Iout.n625 VGND 0.02606f
C16224 Iout.n626 VGND 0.04775f
C16225 Iout.n627 VGND 0.23929f
C16226 Iout.n628 VGND 0.23929f
C16227 Iout.n629 VGND 0.04775f
C16228 Iout.t163 VGND 0.02304f
C16229 Iout.n630 VGND 0.05124f
C16230 Iout.n631 VGND 0.02606f
C16231 Iout.n632 VGND 0.04775f
C16232 Iout.n633 VGND 0.23929f
C16233 Iout.n634 VGND 0.23929f
C16234 Iout.n635 VGND 0.04775f
C16235 Iout.t155 VGND 0.02304f
C16236 Iout.n636 VGND 0.05124f
C16237 Iout.n637 VGND 0.02606f
C16238 Iout.n638 VGND 0.04775f
C16239 Iout.n639 VGND 0.23929f
C16240 Iout.n640 VGND 0.23929f
C16241 Iout.n641 VGND 0.04775f
C16242 Iout.t116 VGND 0.02304f
C16243 Iout.n642 VGND 0.05124f
C16244 Iout.n643 VGND 0.02606f
C16245 Iout.n644 VGND 0.04775f
C16246 Iout.n645 VGND 0.23929f
C16247 Iout.n646 VGND 0.23929f
C16248 Iout.n647 VGND 0.04775f
C16249 Iout.t120 VGND 0.02304f
C16250 Iout.n648 VGND 0.05124f
C16251 Iout.n649 VGND 0.02606f
C16252 Iout.n650 VGND 0.04775f
C16253 Iout.n651 VGND 0.23929f
C16254 Iout.n652 VGND 0.23929f
C16255 Iout.n653 VGND 0.04775f
C16256 Iout.t2 VGND 0.02304f
C16257 Iout.n654 VGND 0.05124f
C16258 Iout.n655 VGND 0.02606f
C16259 Iout.n656 VGND 0.04775f
C16260 Iout.t11 VGND 0.02304f
C16261 Iout.n657 VGND 0.05124f
C16262 Iout.n658 VGND 0.02606f
C16263 Iout.n659 VGND 0.04775f
C16264 Iout.t73 VGND 0.02304f
C16265 Iout.n660 VGND 0.05124f
C16266 Iout.n661 VGND 0.02606f
C16267 Iout.n662 VGND 0.04775f
C16268 Iout.t93 VGND 0.02304f
C16269 Iout.n663 VGND 0.05124f
C16270 Iout.n664 VGND 0.02606f
C16271 Iout.n665 VGND 0.04775f
C16272 Iout.t56 VGND 0.02304f
C16273 Iout.n666 VGND 0.05124f
C16274 Iout.n667 VGND 0.02606f
C16275 Iout.n668 VGND 0.04775f
C16276 Iout.t138 VGND 0.02304f
C16277 Iout.n669 VGND 0.05124f
C16278 Iout.n670 VGND 0.02606f
C16279 Iout.n671 VGND 0.04775f
C16280 Iout.t173 VGND 0.02304f
C16281 Iout.n672 VGND 0.05124f
C16282 Iout.n673 VGND 0.02606f
C16283 Iout.n674 VGND 0.04775f
C16284 Iout.t34 VGND 0.02304f
C16285 Iout.n675 VGND 0.05124f
C16286 Iout.n676 VGND 0.02606f
C16287 Iout.n677 VGND 0.04775f
C16288 Iout.t202 VGND 0.02304f
C16289 Iout.n678 VGND 0.05124f
C16290 Iout.n679 VGND 0.02606f
C16291 Iout.n680 VGND 0.04775f
C16292 Iout.t106 VGND 0.02304f
C16293 Iout.n681 VGND 0.05124f
C16294 Iout.n682 VGND 0.02606f
C16295 Iout.n683 VGND 0.04775f
C16296 Iout.t161 VGND 0.02304f
C16297 Iout.n684 VGND 0.05124f
C16298 Iout.n685 VGND 0.02606f
C16299 Iout.n686 VGND 0.04775f
C16300 Iout.t211 VGND 0.02304f
C16301 Iout.n687 VGND 0.05124f
C16302 Iout.n688 VGND 0.02606f
C16303 Iout.n689 VGND 0.04775f
C16304 Iout.t245 VGND 0.02304f
C16305 Iout.n690 VGND 0.05124f
C16306 Iout.n691 VGND 0.02606f
C16307 Iout.t177 VGND 0.02304f
C16308 Iout.n692 VGND 0.05124f
C16309 Iout.n693 VGND 0.02606f
C16310 Iout.n694 VGND 0.04775f
C16311 Iout.t200 VGND 0.02304f
C16312 Iout.n695 VGND 0.05124f
C16313 Iout.n696 VGND 0.02606f
C16314 Iout.n697 VGND 0.04775f
C16315 Iout.n698 VGND 0.23929f
C16316 Iout.t47 VGND 0.02304f
C16317 Iout.n699 VGND 0.05124f
C16318 Iout.n700 VGND 0.02606f
C16319 Iout.n701 VGND 0.04775f
C16320 Iout.n702 VGND 0.23929f
C16321 Iout.n703 VGND 0.23929f
C16322 Iout.n704 VGND 0.04775f
C16323 Iout.t208 VGND 0.02304f
C16324 Iout.n705 VGND 0.05124f
C16325 Iout.n706 VGND 0.02606f
C16326 Iout.n707 VGND 0.04775f
C16327 Iout.n708 VGND 0.23929f
C16328 Iout.n709 VGND 0.23929f
C16329 Iout.n710 VGND 0.04775f
C16330 Iout.t193 VGND 0.02304f
C16331 Iout.n711 VGND 0.05124f
C16332 Iout.n712 VGND 0.02606f
C16333 Iout.n713 VGND 0.04775f
C16334 Iout.n714 VGND 0.23929f
C16335 Iout.n715 VGND 0.23929f
C16336 Iout.n716 VGND 0.04775f
C16337 Iout.t44 VGND 0.02304f
C16338 Iout.n717 VGND 0.05124f
C16339 Iout.n718 VGND 0.02606f
C16340 Iout.n719 VGND 0.04775f
C16341 Iout.n720 VGND 0.23929f
C16342 Iout.n721 VGND 0.23929f
C16343 Iout.n722 VGND 0.04775f
C16344 Iout.t210 VGND 0.02304f
C16345 Iout.n723 VGND 0.05124f
C16346 Iout.n724 VGND 0.02606f
C16347 Iout.n725 VGND 0.04775f
C16348 Iout.n726 VGND 0.23929f
C16349 Iout.n727 VGND 0.23929f
C16350 Iout.n728 VGND 0.04775f
C16351 Iout.t90 VGND 0.02304f
C16352 Iout.n729 VGND 0.05124f
C16353 Iout.n730 VGND 0.02606f
C16354 Iout.n731 VGND 0.04775f
C16355 Iout.n732 VGND 0.23929f
C16356 Iout.n733 VGND 0.23929f
C16357 Iout.n734 VGND 0.04775f
C16358 Iout.t218 VGND 0.02304f
C16359 Iout.n735 VGND 0.05124f
C16360 Iout.n736 VGND 0.02606f
C16361 Iout.n737 VGND 0.04775f
C16362 Iout.n738 VGND 0.23929f
C16363 Iout.n739 VGND 0.23929f
C16364 Iout.n740 VGND 0.04775f
C16365 Iout.t122 VGND 0.02304f
C16366 Iout.n741 VGND 0.05124f
C16367 Iout.n742 VGND 0.02606f
C16368 Iout.n743 VGND 0.04775f
C16369 Iout.n744 VGND 0.23929f
C16370 Iout.n745 VGND 0.23929f
C16371 Iout.n746 VGND 0.04775f
C16372 Iout.t4 VGND 0.02304f
C16373 Iout.n747 VGND 0.05124f
C16374 Iout.n748 VGND 0.02606f
C16375 Iout.n749 VGND 0.04775f
C16376 Iout.n750 VGND 0.23929f
C16377 Iout.n751 VGND 0.23929f
C16378 Iout.n752 VGND 0.04775f
C16379 Iout.t104 VGND 0.02304f
C16380 Iout.n753 VGND 0.05124f
C16381 Iout.n754 VGND 0.02606f
C16382 Iout.n755 VGND 0.04775f
C16383 Iout.n756 VGND 0.23929f
C16384 Iout.n757 VGND 0.23929f
C16385 Iout.n758 VGND 0.04775f
C16386 Iout.t25 VGND 0.02304f
C16387 Iout.n759 VGND 0.05124f
C16388 Iout.n760 VGND 0.02606f
C16389 Iout.n761 VGND 0.04775f
C16390 Iout.n762 VGND 0.23929f
C16391 Iout.n763 VGND 0.23929f
C16392 Iout.n764 VGND 0.04775f
C16393 Iout.t97 VGND 0.02304f
C16394 Iout.n765 VGND 0.05124f
C16395 Iout.n766 VGND 0.02606f
C16396 Iout.n767 VGND 0.04775f
C16397 Iout.n768 VGND 0.23929f
C16398 Iout.n769 VGND 0.23929f
C16399 Iout.n770 VGND 0.04775f
C16400 Iout.t84 VGND 0.02304f
C16401 Iout.n771 VGND 0.05124f
C16402 Iout.n772 VGND 0.02606f
C16403 Iout.n773 VGND 0.04775f
C16404 Iout.n774 VGND 0.23929f
C16405 Iout.n775 VGND 0.23929f
C16406 Iout.n776 VGND 0.04775f
C16407 Iout.t152 VGND 0.02304f
C16408 Iout.n777 VGND 0.05124f
C16409 Iout.n778 VGND 0.02606f
C16410 Iout.n779 VGND 0.04775f
C16411 Iout.n780 VGND 0.23929f
C16412 Iout.t221 VGND 0.02304f
C16413 Iout.n781 VGND 0.05124f
C16414 Iout.n782 VGND 0.02606f
C16415 Iout.n783 VGND 0.04775f
C16416 Iout.t121 VGND 0.02304f
C16417 Iout.n784 VGND 0.05124f
C16418 Iout.n785 VGND 0.02606f
C16419 Iout.n786 VGND 0.04775f
C16420 Iout.t6 VGND 0.02304f
C16421 Iout.n787 VGND 0.05124f
C16422 Iout.n788 VGND 0.02606f
C16423 Iout.n789 VGND 0.04775f
C16424 Iout.t133 VGND 0.02304f
C16425 Iout.n790 VGND 0.05124f
C16426 Iout.n791 VGND 0.02606f
C16427 Iout.n792 VGND 0.04775f
C16428 Iout.t166 VGND 0.02304f
C16429 Iout.n793 VGND 0.05124f
C16430 Iout.n794 VGND 0.02606f
C16431 Iout.n795 VGND 0.04775f
C16432 Iout.t51 VGND 0.02304f
C16433 Iout.n796 VGND 0.05124f
C16434 Iout.n797 VGND 0.02606f
C16435 Iout.n798 VGND 0.04775f
C16436 Iout.t174 VGND 0.02304f
C16437 Iout.n799 VGND 0.05124f
C16438 Iout.n800 VGND 0.02606f
C16439 Iout.n801 VGND 0.04775f
C16440 Iout.t246 VGND 0.02304f
C16441 Iout.n802 VGND 0.05124f
C16442 Iout.n803 VGND 0.02606f
C16443 Iout.n804 VGND 0.04775f
C16444 Iout.t42 VGND 0.02304f
C16445 Iout.n805 VGND 0.05124f
C16446 Iout.n806 VGND 0.02606f
C16447 Iout.n807 VGND 0.04775f
C16448 Iout.t242 VGND 0.02304f
C16449 Iout.n808 VGND 0.05124f
C16450 Iout.n809 VGND 0.02606f
C16451 Iout.n810 VGND 0.04775f
C16452 Iout.t31 VGND 0.02304f
C16453 Iout.n811 VGND 0.05124f
C16454 Iout.n812 VGND 0.02606f
C16455 Iout.n813 VGND 0.04775f
C16456 Iout.t153 VGND 0.02304f
C16457 Iout.n814 VGND 0.05124f
C16458 Iout.n815 VGND 0.02606f
C16459 Iout.n816 VGND 0.04775f
C16460 Iout.t52 VGND 0.02304f
C16461 Iout.n817 VGND 0.05124f
C16462 Iout.n818 VGND 0.02606f
C16463 Iout.n819 VGND 0.04775f
C16464 Iout.t40 VGND 0.02304f
C16465 Iout.n820 VGND 0.05124f
C16466 Iout.n821 VGND 0.02606f
C16467 Iout.n822 VGND 0.04775f
C16468 Iout.t232 VGND 0.02304f
C16469 Iout.n823 VGND 0.05124f
C16470 Iout.n824 VGND 0.02606f
C16471 Iout.n825 VGND 0.04775f
C16472 Iout.n826 VGND 0.23929f
C16473 Iout.t251 VGND 0.02304f
C16474 Iout.n827 VGND 0.05124f
C16475 Iout.n828 VGND 0.02606f
C16476 Iout.n829 VGND 0.08168f
C16477 Iout.n830 VGND 0.49611f
C16478 Iout.n831 VGND 0.04775f
C16479 Iout.t243 VGND 0.02304f
C16480 Iout.n832 VGND 0.05124f
C16481 Iout.n833 VGND 0.02606f
C16482 Iout.t199 VGND 0.02304f
C16483 Iout.n834 VGND 0.05124f
C16484 Iout.n835 VGND 0.02606f
C16485 Iout.n836 VGND 0.04775f
C16486 Iout.n837 VGND 0.49611f
C16487 Iout.n838 VGND 0.08168f
C16488 Iout.t0 VGND 0.02304f
C16489 Iout.n839 VGND 0.05124f
C16490 Iout.n840 VGND 0.02606f
C16491 Iout.t65 VGND 0.02304f
C16492 Iout.n841 VGND 0.05124f
C16493 Iout.n842 VGND 0.02606f
C16494 Iout.n843 VGND 0.08168f
C16495 Iout.n844 VGND 0.49611f
C16496 Iout.n845 VGND 0.04775f
C16497 Iout.t151 VGND 0.02304f
C16498 Iout.n846 VGND 0.05124f
C16499 Iout.n847 VGND 0.02606f
C16500 Iout.t180 VGND 0.02304f
C16501 Iout.n848 VGND 0.05124f
C16502 Iout.n849 VGND 0.02606f
C16503 Iout.n850 VGND 0.04775f
C16504 Iout.n851 VGND 0.49611f
C16505 Iout.n852 VGND 0.08168f
C16506 Iout.t141 VGND 0.02304f
C16507 Iout.n853 VGND 0.05124f
C16508 Iout.n854 VGND 0.02606f
C16509 Iout.t181 VGND 0.02304f
C16510 Iout.n855 VGND 0.05124f
C16511 Iout.n856 VGND 0.02606f
C16512 Iout.n857 VGND 0.08168f
C16513 Iout.n858 VGND 0.49611f
C16514 Iout.n859 VGND 0.04775f
C16515 Iout.t76 VGND 0.02304f
C16516 Iout.n860 VGND 0.05124f
C16517 Iout.n861 VGND 0.02606f
C16518 Iout.t70 VGND 0.02304f
C16519 Iout.n862 VGND 0.05124f
C16520 Iout.n863 VGND 0.02606f
C16521 Iout.n864 VGND 0.04775f
C16522 Iout.n865 VGND 0.49611f
C16523 Iout.n866 VGND 0.08168f
C16524 Iout.t43 VGND 0.02304f
C16525 Iout.n867 VGND 0.05124f
C16526 Iout.n868 VGND 0.02606f
C16527 Iout.t214 VGND 0.02304f
C16528 Iout.n869 VGND 0.05124f
C16529 Iout.n870 VGND 0.02606f
C16530 Iout.n871 VGND 0.08168f
C16531 Iout.n872 VGND 0.49611f
C16532 Iout.n873 VGND 0.04775f
C16533 Iout.t95 VGND 0.02304f
C16534 Iout.n874 VGND 0.05124f
C16535 Iout.n875 VGND 0.02606f
C16536 Iout.t69 VGND 0.02304f
C16537 Iout.n876 VGND 0.05124f
C16538 Iout.n877 VGND 0.02606f
C16539 Iout.n878 VGND 0.04775f
C16540 Iout.n879 VGND 0.49611f
C16541 Iout.n880 VGND 0.08168f
C16542 Iout.t183 VGND 0.02304f
C16543 Iout.n881 VGND 0.05124f
C16544 Iout.n882 VGND 0.02606f
C16545 Iout.t126 VGND 0.02304f
C16546 Iout.n883 VGND 0.05124f
C16547 Iout.n884 VGND 0.02606f
C16548 Iout.n885 VGND 0.08168f
C16549 Iout.n886 VGND 0.49611f
C16550 Iout.n887 VGND 0.04775f
C16551 Iout.t29 VGND 0.02304f
C16552 Iout.n888 VGND 0.05124f
C16553 Iout.n889 VGND 0.02606f
C16554 Iout.t110 VGND 0.02304f
C16555 Iout.n890 VGND 0.05124f
C16556 Iout.n891 VGND 0.02606f
C16557 Iout.n892 VGND 0.04775f
C16558 Iout.n893 VGND 0.49611f
C16559 Iout.n894 VGND 0.08168f
C16560 Iout.t236 VGND 0.02304f
C16561 Iout.n895 VGND 0.05124f
C16562 Iout.n896 VGND 0.02606f
C16563 Iout.t14 VGND 0.02304f
C16564 Iout.n897 VGND 0.05124f
C16565 Iout.n898 VGND 0.02606f
C16566 Iout.n899 VGND 0.08168f
C16567 Iout.n900 VGND 0.49611f
C16568 Iout.n901 VGND 0.04775f
C16569 Iout.t85 VGND 0.02304f
C16570 Iout.n902 VGND 0.05124f
C16571 Iout.n903 VGND 0.02606f
C16572 Iout.t228 VGND 0.02304f
C16573 Iout.n904 VGND 0.05124f
C16574 Iout.n905 VGND 0.02606f
C16575 Iout.n906 VGND 0.04775f
C16576 Iout.n907 VGND 0.49611f
C16577 Iout.n908 VGND 0.08168f
C16578 Iout.t49 VGND 0.02304f
C16579 Iout.n909 VGND 0.05124f
C16580 Iout.n910 VGND 0.02606f
C16581 Iout.t39 VGND 0.02304f
C16582 Iout.n911 VGND 0.05124f
C16583 Iout.n912 VGND 0.02606f
C16584 Iout.n913 VGND 0.08168f
C16585 Iout.n914 VGND 0.49611f
C16586 Iout.n915 VGND 0.04775f
C16587 Iout.t176 VGND 0.02304f
C16588 Iout.n916 VGND 0.05124f
C16589 Iout.n917 VGND 0.02606f
C16590 Iout.t12 VGND 0.02304f
C16591 Iout.n918 VGND 0.05124f
C16592 Iout.n919 VGND 0.02606f
C16593 Iout.n920 VGND 0.04775f
C16594 Iout.n921 VGND 0.49611f
C16595 Iout.n922 VGND 0.08168f
C16596 Iout.t250 VGND 0.02304f
C16597 Iout.n923 VGND 0.05124f
C16598 Iout.n924 VGND 0.02606f
C16599 Iout.n925 VGND 0.08168f
C16600 Iout.t219 VGND 0.02304f
C16601 Iout.n926 VGND 0.05124f
C16602 Iout.n927 VGND 0.02606f
C16603 Iout.n928 VGND 0.08168f
C16604 Iout.n929 VGND 0.49611f
C16605 Iout.n930 VGND 0.04775f
C16606 Iout.t82 VGND 0.02304f
C16607 Iout.n931 VGND 0.05124f
C16608 Iout.n932 VGND 0.02606f
C16609 Iout.n933 VGND 0.04775f
C16610 Iout.t234 VGND 0.02304f
C16611 Iout.n934 VGND 0.05124f
C16612 Iout.n935 VGND 0.20242f
C16613 Iout.n936 VGND 2.65139f
C16614 Iout.n937 VGND 1.25122f
C16615 Iout.t60 VGND 0.02304f
C16616 Iout.n938 VGND 0.05124f
C16617 Iout.n939 VGND 0.20242f
C16618 Iout.n940 VGND 0.04775f
C16619 Iout.n941 VGND 0.23929f
C16620 Iout.n942 VGND 0.23929f
C16621 Iout.n943 VGND 0.04775f
C16622 Iout.t75 VGND 0.02304f
C16623 Iout.n944 VGND 0.05124f
C16624 Iout.n945 VGND 0.02606f
C16625 Iout.n946 VGND 0.04775f
C16626 Iout.n947 VGND 0.23929f
C16627 Iout.n948 VGND 0.23929f
C16628 Iout.n949 VGND 0.04775f
C16629 Iout.t230 VGND 0.02304f
C16630 Iout.n950 VGND 0.05124f
C16631 Iout.n951 VGND 0.02606f
C16632 Iout.n952 VGND 0.04775f
C16633 Iout.t68 VGND 0.02304f
C16634 Iout.n953 VGND 0.05124f
C16635 Iout.n954 VGND 0.20242f
C16636 Iout.n955 VGND 1.25122f
C16637 Iout.n956 VGND 1.25122f
C16638 Iout.t159 VGND 0.02304f
C16639 Iout.n957 VGND 0.05124f
C16640 Iout.n958 VGND 0.20242f
C16641 Iout.n959 VGND 0.04775f
C16642 Iout.n960 VGND 0.23929f
C16643 Iout.n961 VGND 0.23929f
C16644 Iout.n962 VGND 0.04775f
C16645 Iout.t203 VGND 0.02304f
C16646 Iout.n963 VGND 0.05124f
C16647 Iout.n964 VGND 0.02606f
C16648 Iout.n965 VGND 0.04775f
C16649 Iout.n966 VGND 0.23929f
C16650 Iout.n967 VGND 0.23929f
C16651 Iout.n968 VGND 0.04775f
C16652 Iout.t129 VGND 0.02304f
C16653 Iout.n969 VGND 0.05124f
C16654 Iout.n970 VGND 0.02606f
C16655 Iout.n971 VGND 0.04775f
C16656 Iout.t165 VGND 0.02304f
C16657 Iout.n972 VGND 0.05124f
C16658 Iout.n973 VGND 0.20242f
C16659 Iout.n974 VGND 1.25122f
C16660 Iout.n975 VGND 1.25122f
C16661 Iout.t190 VGND 0.02304f
C16662 Iout.n976 VGND 0.05124f
C16663 Iout.n977 VGND 0.20242f
C16664 Iout.n978 VGND 0.04775f
C16665 Iout.n979 VGND 0.23929f
C16666 Iout.n980 VGND 0.23929f
C16667 Iout.n981 VGND 0.04775f
C16668 Iout.t9 VGND 0.02304f
C16669 Iout.n982 VGND 0.05124f
C16670 Iout.n983 VGND 0.02606f
C16671 Iout.n984 VGND 0.04775f
C16672 Iout.n985 VGND 0.23929f
C16673 Iout.n986 VGND 0.23929f
C16674 Iout.n987 VGND 0.04775f
C16675 Iout.t80 VGND 0.02304f
C16676 Iout.n988 VGND 0.05124f
C16677 Iout.n989 VGND 0.02606f
C16678 Iout.n990 VGND 0.04775f
C16679 Iout.t37 VGND 0.02304f
C16680 Iout.n991 VGND 0.05124f
C16681 Iout.n992 VGND 0.20242f
C16682 Iout.n993 VGND 1.25122f
C16683 Iout.n994 VGND 1.25122f
C16684 Iout.t201 VGND 0.02304f
C16685 Iout.n995 VGND 0.05124f
C16686 Iout.n996 VGND 0.20242f
C16687 Iout.n997 VGND 0.04775f
C16688 Iout.n998 VGND 0.23929f
C16689 Iout.n999 VGND 0.23929f
C16690 Iout.n1000 VGND 0.04775f
C16691 Iout.t46 VGND 0.02304f
C16692 Iout.n1001 VGND 0.05124f
C16693 Iout.n1002 VGND 0.02606f
C16694 Iout.n1003 VGND 0.04775f
C16695 Iout.n1004 VGND 0.23929f
C16696 Iout.n1005 VGND 0.23929f
C16697 Iout.n1006 VGND 0.04775f
C16698 Iout.t15 VGND 0.02304f
C16699 Iout.n1007 VGND 0.05124f
C16700 Iout.n1008 VGND 0.02606f
C16701 Iout.n1009 VGND 0.04775f
C16702 Iout.t189 VGND 0.02304f
C16703 Iout.n1010 VGND 0.05124f
C16704 Iout.n1011 VGND 0.20242f
C16705 Iout.n1012 VGND 1.25122f
C16706 Iout.n1013 VGND 1.1235f
C16707 Iout.t48 VGND 0.02304f
C16708 Iout.n1014 VGND 0.05124f
C16709 Iout.n1015 VGND 0.20242f
C16710 Iout.n1016 VGND 0.04775f
C16711 Iout.n1017 VGND 0.23929f
C16712 Iout.n1018 VGND 0.14126f
C16713 Iout.n1019 VGND 0.04775f
C16714 Iout.t144 VGND 0.02304f
C16715 Iout.n1020 VGND 0.05124f
C16716 Iout.n1021 VGND 0.20242f
C16717 Iout.n1022 VGND 0.23244f
C16718 VPWR.n0 VGND 0.04687f
C16719 VPWR.t463 VGND 0.29639f
C16720 VPWR.t557 VGND 0.13116f
C16721 VPWR.t851 VGND 0.37815f
C16722 VPWR.t846 VGND 0.14308f
C16723 VPWR.t831 VGND 0.14308f
C16724 VPWR.t1240 VGND 0.14308f
C16725 VPWR.t1295 VGND 0.14308f
C16726 VPWR.t788 VGND 0.14308f
C16727 VPWR.t784 VGND 0.14308f
C16728 VPWR.t437 VGND 0.1005f
C16729 VPWR.n1 VGND 0.1826f
C16730 VPWR.n2 VGND 0.09661f
C16731 VPWR.t558 VGND 0.05716f
C16732 VPWR.n3 VGND 0.0092f
C16733 VPWR.t438 VGND 0.01433f
C16734 VPWR.t785 VGND 0.01433f
C16735 VPWR.n4 VGND 0.03146f
C16736 VPWR.t789 VGND 0.01433f
C16737 VPWR.t1296 VGND 0.01433f
C16738 VPWR.n5 VGND 0.03141f
C16739 VPWR.n6 VGND 0.0645f
C16740 VPWR.n7 VGND 0.18182f
C16741 VPWR.n8 VGND 0.05756f
C16742 VPWR.n9 VGND 0.04228f
C16743 VPWR.n10 VGND 0.07578f
C16744 VPWR.n11 VGND 0.01119f
C16745 VPWR.n12 VGND 0.0163f
C16746 VPWR.n13 VGND 0.0191f
C16747 VPWR.n14 VGND 0.02802f
C16748 VPWR.n15 VGND 0.08481f
C16749 VPWR.n16 VGND 0.01209f
C16750 VPWR.t464 VGND 0.05714f
C16751 VPWR.n17 VGND 0.0735f
C16752 VPWR.n18 VGND 0.33563f
C16753 VPWR.n19 VGND 0.97868f
C16754 VPWR.n20 VGND 0.31857f
C16755 VPWR.n21 VGND 1.01577f
C16756 VPWR.n22 VGND 0.13887f
C16757 VPWR.t1970 VGND 0.0112f
C16758 VPWR.t1710 VGND 0.01226f
C16759 VPWR.n23 VGND 0.02994f
C16760 VPWR.n24 VGND 0.07953f
C16761 VPWR.t2021 VGND 0.0112f
C16762 VPWR.t1599 VGND 0.01226f
C16763 VPWR.n25 VGND 0.02994f
C16764 VPWR.n26 VGND 0.16006f
C16765 VPWR.t1956 VGND 0.0112f
C16766 VPWR.t1747 VGND 0.01226f
C16767 VPWR.n27 VGND 0.02994f
C16768 VPWR.n28 VGND 0.12753f
C16769 VPWR.t1995 VGND 0.0112f
C16770 VPWR.t1639 VGND 0.01226f
C16771 VPWR.n29 VGND 0.02994f
C16772 VPWR.n30 VGND 0.12753f
C16773 VPWR.t2064 VGND 0.0112f
C16774 VPWR.t1452 VGND 0.01226f
C16775 VPWR.n31 VGND 0.02994f
C16776 VPWR.n32 VGND 0.12753f
C16777 VPWR.t1997 VGND 0.0112f
C16778 VPWR.t1632 VGND 0.01226f
C16779 VPWR.n33 VGND 0.02994f
C16780 VPWR.n34 VGND 0.12753f
C16781 VPWR.t1943 VGND 0.0112f
C16782 VPWR.t1527 VGND 0.01226f
C16783 VPWR.n35 VGND 0.02994f
C16784 VPWR.n36 VGND 0.12753f
C16785 VPWR.t2022 VGND 0.0112f
C16786 VPWR.t1567 VGND 0.01226f
C16787 VPWR.n37 VGND 0.02994f
C16788 VPWR.n38 VGND 0.12753f
C16789 VPWR.t2028 VGND 0.0112f
C16790 VPWR.t1460 VGND 0.01226f
C16791 VPWR.n39 VGND 0.02994f
C16792 VPWR.n40 VGND 0.12753f
C16793 VPWR.t2069 VGND 0.0112f
C16794 VPWR.t1734 VGND 0.01226f
C16795 VPWR.n41 VGND 0.02994f
C16796 VPWR.n42 VGND 0.12753f
C16797 VPWR.t2051 VGND 0.0112f
C16798 VPWR.t1626 VGND 0.01226f
C16799 VPWR.n43 VGND 0.02994f
C16800 VPWR.n44 VGND 0.12753f
C16801 VPWR.t1946 VGND 0.0112f
C16802 VPWR.t1777 VGND 0.01226f
C16803 VPWR.n45 VGND 0.02994f
C16804 VPWR.n46 VGND 0.12753f
C16805 VPWR.t2026 VGND 0.0112f
C16806 VPWR.t1559 VGND 0.01226f
C16807 VPWR.n47 VGND 0.02994f
C16808 VPWR.n48 VGND 0.12753f
C16809 VPWR.t2066 VGND 0.0112f
C16810 VPWR.t1444 VGND 0.01226f
C16811 VPWR.n49 VGND 0.02994f
C16812 VPWR.n50 VGND 0.12753f
C16813 VPWR.t1963 VGND 0.0112f
C16814 VPWR.t1729 VGND 0.01226f
C16815 VPWR.n51 VGND 0.02994f
C16816 VPWR.n52 VGND 0.12753f
C16817 VPWR.t2053 VGND 0.0112f
C16818 VPWR.t1769 VGND 0.01226f
C16819 VPWR.n53 VGND 0.02994f
C16820 VPWR.n54 VGND 0.13808f
C16821 VPWR.n55 VGND 0.11528f
C16822 VPWR.t1558 VGND 0.03331f
C16823 VPWR.t1663 VGND 0.02961f
C16824 VPWR.n56 VGND 0.09152f
C16825 VPWR.t1426 VGND 0.09218f
C16826 VPWR.t1433 VGND 0.03331f
C16827 VPWR.t1427 VGND 0.02961f
C16828 VPWR.n57 VGND 0.09152f
C16829 VPWR.n58 VGND 0.03437f
C16830 VPWR.n59 VGND 0.13913f
C16831 VPWR.n60 VGND 0.13913f
C16832 VPWR.n61 VGND 0.03437f
C16833 VPWR.t1414 VGND 0.03331f
C16834 VPWR.t1787 VGND 0.02961f
C16835 VPWR.n62 VGND 0.09152f
C16836 VPWR.t1653 VGND 0.09218f
C16837 VPWR.t1564 VGND 0.03331f
C16838 VPWR.t1654 VGND 0.02961f
C16839 VPWR.n63 VGND 0.09152f
C16840 VPWR.n64 VGND 0.03437f
C16841 VPWR.n65 VGND 0.13913f
C16842 VPWR.n66 VGND 0.13913f
C16843 VPWR.n67 VGND 0.03437f
C16844 VPWR.t1534 VGND 0.03331f
C16845 VPWR.t1526 VGND 0.02961f
C16846 VPWR.n68 VGND 0.09152f
C16847 VPWR.t1507 VGND 0.09218f
C16848 VPWR.t1790 VGND 0.03331f
C16849 VPWR.t1508 VGND 0.02961f
C16850 VPWR.n69 VGND 0.09152f
C16851 VPWR.n70 VGND 0.03437f
C16852 VPWR.n71 VGND 0.13913f
C16853 VPWR.n72 VGND 0.13913f
C16854 VPWR.n73 VGND 0.03437f
C16855 VPWR.t1660 VGND 0.03331f
C16856 VPWR.t1741 VGND 0.02961f
C16857 VPWR.n74 VGND 0.09152f
C16858 VPWR.t1630 VGND 0.09218f
C16859 VPWR.t1644 VGND 0.03331f
C16860 VPWR.t1631 VGND 0.02961f
C16861 VPWR.n75 VGND 0.09152f
C16862 VPWR.n76 VGND 0.03437f
C16863 VPWR.n77 VGND 0.13913f
C16864 VPWR.n78 VGND 0.13913f
C16865 VPWR.n79 VGND 0.03437f
C16866 VPWR.t1484 VGND 0.03331f
C16867 VPWR.t1503 VGND 0.02961f
C16868 VPWR.n80 VGND 0.09152f
C16869 VPWR.t1467 VGND 0.09218f
C16870 VPWR.t1763 VGND 0.03331f
C16871 VPWR.t1468 VGND 0.02961f
C16872 VPWR.n81 VGND 0.09152f
C16873 VPWR.n82 VGND 0.03437f
C16874 VPWR.n83 VGND 0.13913f
C16875 VPWR.n84 VGND 0.13913f
C16876 VPWR.n85 VGND 0.03437f
C16877 VPWR.t1607 VGND 0.03331f
C16878 VPWR.t1744 VGND 0.02961f
C16879 VPWR.n86 VGND 0.09152f
C16880 VPWR.t1588 VGND 0.09218f
C16881 VPWR.t1595 VGND 0.03331f
C16882 VPWR.t1589 VGND 0.02961f
C16883 VPWR.n87 VGND 0.09152f
C16884 VPWR.n88 VGND 0.03437f
C16885 VPWR.n89 VGND 0.13913f
C16886 VPWR.n90 VGND 0.13913f
C16887 VPWR.n91 VGND 0.03437f
C16888 VPWR.t1487 VGND 0.03331f
C16889 VPWR.t1481 VGND 0.02961f
C16890 VPWR.n92 VGND 0.09152f
C16891 VPWR.t1718 VGND 0.09218f
C16892 VPWR.t1722 VGND 0.03331f
C16893 VPWR.t1719 VGND 0.02961f
C16894 VPWR.n93 VGND 0.09152f
C16895 VPWR.n94 VGND 0.03437f
C16896 VPWR.n95 VGND 0.13913f
C16897 VPWR.n96 VGND 0.13913f
C16898 VPWR.n97 VGND 0.03437f
C16899 VPWR.t1610 VGND 0.03331f
C16900 VPWR.t1701 VGND 0.02961f
C16901 VPWR.n98 VGND 0.09152f
C16902 VPWR.t1464 VGND 0.14512f
C16903 VPWR.t1440 VGND 0.07849f
C16904 VPWR.t1571 VGND 0.09218f
C16905 VPWR.t1465 VGND 0.03331f
C16906 VPWR.t1572 VGND 0.02961f
C16907 VPWR.n99 VGND 0.09152f
C16908 VPWR.t1987 VGND 0.0112f
C16909 VPWR.t1699 VGND 0.01226f
C16910 VPWR.n100 VGND 0.02993f
C16911 VPWR.n101 VGND 0.03284f
C16912 VPWR.n102 VGND 0.00697f
C16913 VPWR.n103 VGND 0.01822f
C16914 VPWR.t2032 VGND 0.0112f
C16915 VPWR.t1570 VGND 0.01226f
C16916 VPWR.n104 VGND 0.02993f
C16917 VPWR.n105 VGND 0.03284f
C16918 VPWR.t1981 VGND 0.01116f
C16919 VPWR.t1463 VGND 0.01222f
C16920 VPWR.n106 VGND 0.03115f
C16921 VPWR.n107 VGND 0.01969f
C16922 VPWR.t1934 VGND 0.01136f
C16923 VPWR.t1439 VGND 0.0124f
C16924 VPWR.n108 VGND 0.02768f
C16925 VPWR.n109 VGND 0.02818f
C16926 VPWR.n110 VGND 0.01776f
C16927 VPWR.n111 VGND 0.00697f
C16928 VPWR.n112 VGND 0.01822f
C16929 VPWR.n113 VGND 0.02654f
C16930 VPWR.t2001 VGND 0.0112f
C16931 VPWR.t1661 VGND 0.01226f
C16932 VPWR.n114 VGND 0.02993f
C16933 VPWR.n115 VGND 0.03284f
C16934 VPWR.t1951 VGND 0.01116f
C16935 VPWR.t1556 VGND 0.01222f
C16936 VPWR.n116 VGND 0.03115f
C16937 VPWR.n117 VGND 0.03694f
C16938 VPWR.n118 VGND 0.00833f
C16939 VPWR.t2048 VGND 0.01136f
C16940 VPWR.t1540 VGND 0.0124f
C16941 VPWR.n119 VGND 0.02768f
C16942 VPWR.n120 VGND 0.02818f
C16943 VPWR.n121 VGND 0.01776f
C16944 VPWR.n122 VGND 0.00697f
C16945 VPWR.n123 VGND 0.01822f
C16946 VPWR.n124 VGND 0.02541f
C16947 VPWR.t1940 VGND 0.0112f
C16948 VPWR.t1425 VGND 0.01226f
C16949 VPWR.n125 VGND 0.02993f
C16950 VPWR.n126 VGND 0.03284f
C16951 VPWR.t1991 VGND 0.01116f
C16952 VPWR.t1431 VGND 0.01222f
C16953 VPWR.n127 VGND 0.03115f
C16954 VPWR.n128 VGND 0.03694f
C16955 VPWR.n129 VGND 0.00833f
C16956 VPWR.t1990 VGND 0.01136f
C16957 VPWR.t1689 VGND 0.0124f
C16958 VPWR.n130 VGND 0.02768f
C16959 VPWR.n131 VGND 0.02818f
C16960 VPWR.n132 VGND 0.01776f
C16961 VPWR.n133 VGND 0.00697f
C16962 VPWR.n134 VGND 0.01822f
C16963 VPWR.n135 VGND 0.02384f
C16964 VPWR.n136 VGND 0.21163f
C16965 VPWR.t1954 VGND 0.0112f
C16966 VPWR.t1785 VGND 0.01226f
C16967 VPWR.n137 VGND 0.02993f
C16968 VPWR.n138 VGND 0.03284f
C16969 VPWR.t2046 VGND 0.01116f
C16970 VPWR.t1412 VGND 0.01222f
C16971 VPWR.n139 VGND 0.03115f
C16972 VPWR.n140 VGND 0.03694f
C16973 VPWR.n141 VGND 0.00833f
C16974 VPWR.t1999 VGND 0.01136f
C16975 VPWR.t1664 VGND 0.0124f
C16976 VPWR.n142 VGND 0.02768f
C16977 VPWR.n143 VGND 0.02818f
C16978 VPWR.n144 VGND 0.01776f
C16979 VPWR.n145 VGND 0.00697f
C16980 VPWR.n146 VGND 0.01822f
C16981 VPWR.n147 VGND 0.02384f
C16982 VPWR.n148 VGND 0.17585f
C16983 VPWR.t2004 VGND 0.0112f
C16984 VPWR.t1652 VGND 0.01226f
C16985 VPWR.n149 VGND 0.02993f
C16986 VPWR.n150 VGND 0.03284f
C16987 VPWR.t1942 VGND 0.01116f
C16988 VPWR.t1562 VGND 0.01222f
C16989 VPWR.n151 VGND 0.03115f
C16990 VPWR.n152 VGND 0.03694f
C16991 VPWR.n153 VGND 0.00833f
C16992 VPWR.t2007 VGND 0.01136f
C16993 VPWR.t1645 VGND 0.0124f
C16994 VPWR.n154 VGND 0.02768f
C16995 VPWR.n155 VGND 0.02818f
C16996 VPWR.n156 VGND 0.01776f
C16997 VPWR.n157 VGND 0.00697f
C16998 VPWR.n158 VGND 0.01822f
C16999 VPWR.n159 VGND 0.02384f
C17000 VPWR.n160 VGND 0.17585f
C17001 VPWR.t2052 VGND 0.0112f
C17002 VPWR.t1524 VGND 0.01226f
C17003 VPWR.n161 VGND 0.02993f
C17004 VPWR.n162 VGND 0.03284f
C17005 VPWR.t1998 VGND 0.01116f
C17006 VPWR.t1532 VGND 0.01222f
C17007 VPWR.n163 VGND 0.03115f
C17008 VPWR.n164 VGND 0.03694f
C17009 VPWR.n165 VGND 0.00833f
C17010 VPWR.t1952 VGND 0.01136f
C17011 VPWR.t1791 VGND 0.0124f
C17012 VPWR.n166 VGND 0.02768f
C17013 VPWR.n167 VGND 0.02818f
C17014 VPWR.n168 VGND 0.01776f
C17015 VPWR.n169 VGND 0.00697f
C17016 VPWR.n170 VGND 0.01822f
C17017 VPWR.n171 VGND 0.02384f
C17018 VPWR.n172 VGND 0.17585f
C17019 VPWR.t2058 VGND 0.0112f
C17020 VPWR.t1506 VGND 0.01226f
C17021 VPWR.n173 VGND 0.02993f
C17022 VPWR.n174 VGND 0.03284f
C17023 VPWR.t2006 VGND 0.01116f
C17024 VPWR.t1788 VGND 0.01222f
C17025 VPWR.n175 VGND 0.03115f
C17026 VPWR.n176 VGND 0.03694f
C17027 VPWR.n177 VGND 0.00833f
C17028 VPWR.t1961 VGND 0.01136f
C17029 VPWR.t1772 VGND 0.0124f
C17030 VPWR.n178 VGND 0.02768f
C17031 VPWR.n179 VGND 0.02818f
C17032 VPWR.n180 VGND 0.01776f
C17033 VPWR.n181 VGND 0.00697f
C17034 VPWR.n182 VGND 0.01822f
C17035 VPWR.n183 VGND 0.02384f
C17036 VPWR.n184 VGND 0.17585f
C17037 VPWR.t1973 VGND 0.0112f
C17038 VPWR.t1739 VGND 0.01226f
C17039 VPWR.n185 VGND 0.02993f
C17040 VPWR.n186 VGND 0.03284f
C17041 VPWR.t2054 VGND 0.01116f
C17042 VPWR.t1658 VGND 0.01222f
C17043 VPWR.n187 VGND 0.03115f
C17044 VPWR.n188 VGND 0.03694f
C17045 VPWR.n189 VGND 0.00833f
C17046 VPWR.t2017 VGND 0.01136f
C17047 VPWR.t1611 VGND 0.0124f
C17048 VPWR.n190 VGND 0.02768f
C17049 VPWR.n191 VGND 0.02818f
C17050 VPWR.n192 VGND 0.01776f
C17051 VPWR.n193 VGND 0.00697f
C17052 VPWR.n194 VGND 0.01822f
C17053 VPWR.n195 VGND 0.02384f
C17054 VPWR.n196 VGND 0.17585f
C17055 VPWR.t2009 VGND 0.0112f
C17056 VPWR.t1629 VGND 0.01226f
C17057 VPWR.n197 VGND 0.02993f
C17058 VPWR.n198 VGND 0.03284f
C17059 VPWR.t1960 VGND 0.01116f
C17060 VPWR.t1642 VGND 0.01222f
C17061 VPWR.n199 VGND 0.03115f
C17062 VPWR.n200 VGND 0.03694f
C17063 VPWR.n201 VGND 0.00833f
C17064 VPWR.t2057 VGND 0.01136f
C17065 VPWR.t1509 VGND 0.0124f
C17066 VPWR.n202 VGND 0.02768f
C17067 VPWR.n203 VGND 0.02818f
C17068 VPWR.n204 VGND 0.01776f
C17069 VPWR.n205 VGND 0.00697f
C17070 VPWR.n206 VGND 0.01822f
C17071 VPWR.n207 VGND 0.02384f
C17072 VPWR.n208 VGND 0.17585f
C17073 VPWR.t2060 VGND 0.0112f
C17074 VPWR.t1501 VGND 0.01226f
C17075 VPWR.n209 VGND 0.02993f
C17076 VPWR.n210 VGND 0.03284f
C17077 VPWR.t1974 VGND 0.01116f
C17078 VPWR.t1482 VGND 0.01222f
C17079 VPWR.n211 VGND 0.03115f
C17080 VPWR.n212 VGND 0.03694f
C17081 VPWR.n213 VGND 0.00833f
C17082 VPWR.t1928 VGND 0.01136f
C17083 VPWR.t1474 VGND 0.0124f
C17084 VPWR.n214 VGND 0.02768f
C17085 VPWR.n215 VGND 0.02818f
C17086 VPWR.n216 VGND 0.01776f
C17087 VPWR.n217 VGND 0.00697f
C17088 VPWR.n218 VGND 0.01822f
C17089 VPWR.n219 VGND 0.02384f
C17090 VPWR.n220 VGND 0.17585f
C17091 VPWR.t1931 VGND 0.0112f
C17092 VPWR.t1466 VGND 0.01226f
C17093 VPWR.n221 VGND 0.02993f
C17094 VPWR.n222 VGND 0.03284f
C17095 VPWR.t2056 VGND 0.01116f
C17096 VPWR.t1761 VGND 0.01222f
C17097 VPWR.n223 VGND 0.03115f
C17098 VPWR.n224 VGND 0.03694f
C17099 VPWR.n225 VGND 0.00833f
C17100 VPWR.t2008 VGND 0.01136f
C17101 VPWR.t1637 VGND 0.0124f
C17102 VPWR.n226 VGND 0.02768f
C17103 VPWR.n227 VGND 0.02818f
C17104 VPWR.n228 VGND 0.01776f
C17105 VPWR.n229 VGND 0.00697f
C17106 VPWR.n230 VGND 0.01822f
C17107 VPWR.n231 VGND 0.02384f
C17108 VPWR.n232 VGND 0.17585f
C17109 VPWR.t1972 VGND 0.0112f
C17110 VPWR.t1742 VGND 0.01226f
C17111 VPWR.n233 VGND 0.02993f
C17112 VPWR.n234 VGND 0.03284f
C17113 VPWR.t1926 VGND 0.01116f
C17114 VPWR.t1605 VGND 0.01222f
C17115 VPWR.n235 VGND 0.03115f
C17116 VPWR.n236 VGND 0.03694f
C17117 VPWR.n237 VGND 0.00833f
C17118 VPWR.t2016 VGND 0.01136f
C17119 VPWR.t1613 VGND 0.0124f
C17120 VPWR.n238 VGND 0.02768f
C17121 VPWR.n239 VGND 0.02818f
C17122 VPWR.n240 VGND 0.01776f
C17123 VPWR.n241 VGND 0.00697f
C17124 VPWR.n242 VGND 0.01822f
C17125 VPWR.n243 VGND 0.02384f
C17126 VPWR.n244 VGND 0.17585f
C17127 VPWR.t2027 VGND 0.0112f
C17128 VPWR.t1587 VGND 0.01226f
C17129 VPWR.n245 VGND 0.02993f
C17130 VPWR.n246 VGND 0.03284f
C17131 VPWR.t1932 VGND 0.01116f
C17132 VPWR.t1593 VGND 0.01222f
C17133 VPWR.n247 VGND 0.03115f
C17134 VPWR.n248 VGND 0.03694f
C17135 VPWR.n249 VGND 0.00833f
C17136 VPWR.t1930 VGND 0.01136f
C17137 VPWR.t1469 VGND 0.0124f
C17138 VPWR.n250 VGND 0.02768f
C17139 VPWR.n251 VGND 0.02818f
C17140 VPWR.n252 VGND 0.01776f
C17141 VPWR.n253 VGND 0.00697f
C17142 VPWR.n254 VGND 0.01822f
C17143 VPWR.n255 VGND 0.02384f
C17144 VPWR.n256 VGND 0.17585f
C17145 VPWR.t2068 VGND 0.0112f
C17146 VPWR.t1479 VGND 0.01226f
C17147 VPWR.n257 VGND 0.02993f
C17148 VPWR.n258 VGND 0.03284f
C17149 VPWR.t2015 VGND 0.01116f
C17150 VPWR.t1485 VGND 0.01222f
C17151 VPWR.n259 VGND 0.03115f
C17152 VPWR.n260 VGND 0.03694f
C17153 VPWR.n261 VGND 0.00833f
C17154 VPWR.t1971 VGND 0.01136f
C17155 VPWR.t1745 VGND 0.0124f
C17156 VPWR.n262 VGND 0.02768f
C17157 VPWR.n263 VGND 0.02818f
C17158 VPWR.n264 VGND 0.01776f
C17159 VPWR.n265 VGND 0.00697f
C17160 VPWR.n266 VGND 0.01822f
C17161 VPWR.n267 VGND 0.02384f
C17162 VPWR.n268 VGND 0.17585f
C17163 VPWR.t1980 VGND 0.0112f
C17164 VPWR.t1717 VGND 0.01226f
C17165 VPWR.n269 VGND 0.02993f
C17166 VPWR.n270 VGND 0.03284f
C17167 VPWR.t2029 VGND 0.01116f
C17168 VPWR.t1720 VGND 0.01222f
C17169 VPWR.n271 VGND 0.03115f
C17170 VPWR.n272 VGND 0.03694f
C17171 VPWR.n273 VGND 0.00833f
C17172 VPWR.t1983 VGND 0.01136f
C17173 VPWR.t1705 VGND 0.0124f
C17174 VPWR.n274 VGND 0.02768f
C17175 VPWR.n275 VGND 0.02818f
C17176 VPWR.n276 VGND 0.01776f
C17177 VPWR.n277 VGND 0.00697f
C17178 VPWR.n278 VGND 0.01822f
C17179 VPWR.n279 VGND 0.02384f
C17180 VPWR.n280 VGND 0.17585f
C17181 VPWR.n281 VGND 0.23724f
C17182 VPWR.n282 VGND 0.02384f
C17183 VPWR.n283 VGND 0.01776f
C17184 VPWR.t2030 VGND 0.01136f
C17185 VPWR.t1575 VGND 0.0124f
C17186 VPWR.n284 VGND 0.02768f
C17187 VPWR.n285 VGND 0.02818f
C17188 VPWR.n286 VGND 0.00833f
C17189 VPWR.t1933 VGND 0.01116f
C17190 VPWR.t1608 VGND 0.01222f
C17191 VPWR.n287 VGND 0.03115f
C17192 VPWR.n288 VGND 0.03694f
C17193 VPWR.n289 VGND 0.03437f
C17194 VPWR.t1083 VGND 0.03331f
C17195 VPWR.t166 VGND 0.02961f
C17196 VPWR.n290 VGND 0.09152f
C17197 VPWR.t1082 VGND 0.14512f
C17198 VPWR.t711 VGND 0.07849f
C17199 VPWR.t165 VGND 0.09218f
C17200 VPWR.t184 VGND 0.03331f
C17201 VPWR.t1771 VGND 0.02961f
C17202 VPWR.n291 VGND 0.09152f
C17203 VPWR.n292 VGND 0.01797f
C17204 VPWR.n293 VGND 0.07618f
C17205 VPWR.t1770 VGND 0.13333f
C17206 VPWR.t1043 VGND 0.07849f
C17207 VPWR.t183 VGND 0.11957f
C17208 VPWR.t436 VGND 0.03331f
C17209 VPWR.t521 VGND 0.02961f
C17210 VPWR.n294 VGND 0.09152f
C17211 VPWR.n295 VGND 0.01797f
C17212 VPWR.n296 VGND 0.00728f
C17213 VPWR.n297 VGND 0.10822f
C17214 VPWR.t520 VGND 0.09218f
C17215 VPWR.t663 VGND 0.07849f
C17216 VPWR.t435 VGND 0.11957f
C17217 VPWR.t97 VGND 0.03331f
C17218 VPWR.t1123 VGND 0.02961f
C17219 VPWR.n298 VGND 0.09152f
C17220 VPWR.n299 VGND 0.01797f
C17221 VPWR.n300 VGND 0.00728f
C17222 VPWR.n301 VGND 0.10822f
C17223 VPWR.t1122 VGND 0.09218f
C17224 VPWR.t1037 VGND 0.07849f
C17225 VPWR.t96 VGND 0.11957f
C17226 VPWR.t856 VGND 0.03331f
C17227 VPWR.t68 VGND 0.02961f
C17228 VPWR.n302 VGND 0.09152f
C17229 VPWR.n303 VGND 0.01797f
C17230 VPWR.n304 VGND 0.00728f
C17231 VPWR.n305 VGND 0.10822f
C17232 VPWR.t67 VGND 0.09218f
C17233 VPWR.t1038 VGND 0.07849f
C17234 VPWR.t855 VGND 0.11957f
C17235 VPWR.t124 VGND 0.03331f
C17236 VPWR.t1847 VGND 0.02961f
C17237 VPWR.n306 VGND 0.09152f
C17238 VPWR.n307 VGND 0.01797f
C17239 VPWR.n308 VGND 0.00728f
C17240 VPWR.n309 VGND 0.10822f
C17241 VPWR.t1846 VGND 0.09218f
C17242 VPWR.t712 VGND 0.07849f
C17243 VPWR.t123 VGND 0.11957f
C17244 VPWR.t1373 VGND 0.03331f
C17245 VPWR.t130 VGND 0.02961f
C17246 VPWR.n310 VGND 0.09152f
C17247 VPWR.n311 VGND 0.01797f
C17248 VPWR.n312 VGND 0.00728f
C17249 VPWR.n313 VGND 0.10822f
C17250 VPWR.t129 VGND 0.09218f
C17251 VPWR.t713 VGND 0.07849f
C17252 VPWR.t1372 VGND 0.11957f
C17253 VPWR.t638 VGND 0.03331f
C17254 VPWR.t1383 VGND 0.02961f
C17255 VPWR.n314 VGND 0.09152f
C17256 VPWR.n315 VGND 0.01797f
C17257 VPWR.n316 VGND 0.00728f
C17258 VPWR.n317 VGND 0.10822f
C17259 VPWR.t1382 VGND 0.09218f
C17260 VPWR.t1041 VGND 0.07849f
C17261 VPWR.t637 VGND 0.11957f
C17262 VPWR.t470 VGND 0.03331f
C17263 VPWR.t644 VGND 0.02961f
C17264 VPWR.n318 VGND 0.09152f
C17265 VPWR.n319 VGND 0.01797f
C17266 VPWR.n320 VGND 0.00728f
C17267 VPWR.n321 VGND 0.10822f
C17268 VPWR.t643 VGND 0.09218f
C17269 VPWR.t708 VGND 0.07849f
C17270 VPWR.t469 VGND 0.11957f
C17271 VPWR.t293 VGND 0.03331f
C17272 VPWR.t582 VGND 0.02961f
C17273 VPWR.n322 VGND 0.09152f
C17274 VPWR.n323 VGND 0.01797f
C17275 VPWR.n324 VGND 0.00728f
C17276 VPWR.n325 VGND 0.10822f
C17277 VPWR.t581 VGND 0.09218f
C17278 VPWR.t709 VGND 0.07849f
C17279 VPWR.t292 VGND 0.11957f
C17280 VPWR.t254 VGND 0.03331f
C17281 VPWR.t299 VGND 0.02961f
C17282 VPWR.n326 VGND 0.09152f
C17283 VPWR.n327 VGND 0.01797f
C17284 VPWR.n328 VGND 0.00728f
C17285 VPWR.n329 VGND 0.10822f
C17286 VPWR.t298 VGND 0.09218f
C17287 VPWR.t1039 VGND 0.07849f
C17288 VPWR.t253 VGND 0.11957f
C17289 VPWR.t170 VGND 0.03331f
C17290 VPWR.t260 VGND 0.02961f
C17291 VPWR.n330 VGND 0.09152f
C17292 VPWR.n331 VGND 0.01797f
C17293 VPWR.n332 VGND 0.00728f
C17294 VPWR.n333 VGND 0.10822f
C17295 VPWR.t259 VGND 0.09218f
C17296 VPWR.t1040 VGND 0.07849f
C17297 VPWR.t169 VGND 0.11957f
C17298 VPWR.t609 VGND 0.03331f
C17299 VPWR.t611 VGND 0.02961f
C17300 VPWR.n334 VGND 0.09152f
C17301 VPWR.n335 VGND 0.01797f
C17302 VPWR.n336 VGND 0.00728f
C17303 VPWR.n337 VGND 0.10822f
C17304 VPWR.t610 VGND 0.09218f
C17305 VPWR.t710 VGND 0.07849f
C17306 VPWR.t608 VGND 0.11957f
C17307 VPWR.t753 VGND 0.03331f
C17308 VPWR.t1010 VGND 0.02961f
C17309 VPWR.n338 VGND 0.09152f
C17310 VPWR.n339 VGND 0.01797f
C17311 VPWR.n340 VGND 0.00728f
C17312 VPWR.n341 VGND 0.10822f
C17313 VPWR.t1009 VGND 0.09218f
C17314 VPWR.t661 VGND 0.07849f
C17315 VPWR.t752 VGND 0.11957f
C17316 VPWR.t506 VGND 0.03331f
C17317 VPWR.t729 VGND 0.02961f
C17318 VPWR.n342 VGND 0.09152f
C17319 VPWR.n343 VGND 0.01797f
C17320 VPWR.n344 VGND 0.00728f
C17321 VPWR.n345 VGND 0.10822f
C17322 VPWR.t728 VGND 0.09218f
C17323 VPWR.t662 VGND 0.07849f
C17324 VPWR.t505 VGND 0.11957f
C17325 VPWR.t178 VGND 0.03331f
C17326 VPWR.t484 VGND 0.02961f
C17327 VPWR.n346 VGND 0.09152f
C17328 VPWR.n347 VGND 0.01797f
C17329 VPWR.n348 VGND 0.00728f
C17330 VPWR.n349 VGND 0.10822f
C17331 VPWR.t483 VGND 0.09218f
C17332 VPWR.t1042 VGND 0.07849f
C17333 VPWR.t177 VGND 0.11957f
C17334 VPWR.n350 VGND 0.10822f
C17335 VPWR.n351 VGND 0.00728f
C17336 VPWR.n352 VGND 0.01797f
C17337 VPWR.n353 VGND 0.13913f
C17338 VPWR.n354 VGND 1.0094f
C17339 VPWR.n355 VGND 0.13913f
C17340 VPWR.t1076 VGND 0.03331f
C17341 VPWR.t1004 VGND 0.02961f
C17342 VPWR.n356 VGND 0.09152f
C17343 VPWR.t1075 VGND 0.14512f
C17344 VPWR.t1356 VGND 0.07849f
C17345 VPWR.t1003 VGND 0.09218f
C17346 VPWR.t487 VGND 0.11957f
C17347 VPWR.t162 VGND 0.03331f
C17348 VPWR.t58 VGND 0.02961f
C17349 VPWR.n357 VGND 0.09152f
C17350 VPWR.n358 VGND 0.13913f
C17351 VPWR.n359 VGND 0.13913f
C17352 VPWR.t488 VGND 0.03331f
C17353 VPWR.t721 VGND 0.02961f
C17354 VPWR.n360 VGND 0.09152f
C17355 VPWR.t816 VGND 0.07849f
C17356 VPWR.t720 VGND 0.09218f
C17357 VPWR.t1172 VGND 0.11957f
C17358 VPWR.t745 VGND 0.03331f
C17359 VPWR.t1054 VGND 0.02961f
C17360 VPWR.n361 VGND 0.09152f
C17361 VPWR.n362 VGND 0.13913f
C17362 VPWR.n363 VGND 0.13913f
C17363 VPWR.t1173 VGND 0.03331f
C17364 VPWR.t621 VGND 0.02961f
C17365 VPWR.n364 VGND 0.09152f
C17366 VPWR.t1355 VGND 0.07849f
C17367 VPWR.t620 VGND 0.09218f
C17368 VPWR.t263 VGND 0.11957f
C17369 VPWR.t615 VGND 0.03331f
C17370 VPWR.t278 VGND 0.02961f
C17371 VPWR.n365 VGND 0.09152f
C17372 VPWR.n366 VGND 0.13913f
C17373 VPWR.n367 VGND 0.13913f
C17374 VPWR.t264 VGND 0.03331f
C17375 VPWR.t309 VGND 0.02961f
C17376 VPWR.n368 VGND 0.09152f
C17377 VPWR.t820 VGND 0.07849f
C17378 VPWR.t308 VGND 0.09218f
C17379 VPWR.t837 VGND 0.11957f
C17380 VPWR.t303 VGND 0.03331f
C17381 VPWR.t592 VGND 0.02961f
C17382 VPWR.n369 VGND 0.09152f
C17383 VPWR.n370 VGND 0.13913f
C17384 VPWR.n371 VGND 0.13913f
C17385 VPWR.t838 VGND 0.03331f
C17386 VPWR.t574 VGND 0.02961f
C17387 VPWR.n372 VGND 0.09152f
C17388 VPWR.t1353 VGND 0.07849f
C17389 VPWR.t573 VGND 0.09218f
C17390 VPWR.t1378 VGND 0.11957f
C17391 VPWR.t568 VGND 0.03331f
C17392 VPWR.t1913 VGND 0.02961f
C17393 VPWR.n373 VGND 0.09152f
C17394 VPWR.n374 VGND 0.13913f
C17395 VPWR.n375 VGND 0.13913f
C17396 VPWR.t1379 VGND 0.03331f
C17397 VPWR.t1362 VGND 0.02961f
C17398 VPWR.n376 VGND 0.09152f
C17399 VPWR.t201 VGND 0.07849f
C17400 VPWR.t1361 VGND 0.09218f
C17401 VPWR.t1102 VGND 0.11957f
C17402 VPWR.t134 VGND 0.03331f
C17403 VPWR.t1853 VGND 0.02961f
C17404 VPWR.n377 VGND 0.09152f
C17405 VPWR.n378 VGND 0.13913f
C17406 VPWR.n379 VGND 0.13913f
C17407 VPWR.t1103 VGND 0.03331f
C17408 VPWR.t1206 VGND 0.02961f
C17409 VPWR.n380 VGND 0.09152f
C17410 VPWR.t819 VGND 0.07849f
C17411 VPWR.t1205 VGND 0.09218f
C17412 VPWR.t411 VGND 0.11957f
C17413 VPWR.t103 VGND 0.03331f
C17414 VPWR.t331 VGND 0.02961f
C17415 VPWR.n381 VGND 0.09152f
C17416 VPWR.n382 VGND 0.13913f
C17417 VPWR.n383 VGND 0.13913f
C17418 VPWR.t412 VGND 0.03331f
C17419 VPWR.t335 VGND 0.02961f
C17420 VPWR.n384 VGND 0.09152f
C17421 VPWR.t817 VGND 0.07849f
C17422 VPWR.t334 VGND 0.09218f
C17423 VPWR.t192 VGND 0.03331f
C17424 VPWR.t1731 VGND 0.02961f
C17425 VPWR.n385 VGND 0.09152f
C17426 VPWR.t321 VGND 0.03331f
C17427 VPWR.t1446 VGND 0.02961f
C17428 VPWR.n386 VGND 0.09152f
C17429 VPWR.t1086 VGND 0.14512f
C17430 VPWR.t678 VGND 0.07849f
C17431 VPWR.t599 VGND 0.09218f
C17432 VPWR.t1087 VGND 0.03331f
C17433 VPWR.t600 VGND 0.02961f
C17434 VPWR.n387 VGND 0.09152f
C17435 VPWR.n388 VGND 0.01797f
C17436 VPWR.n389 VGND 0.00728f
C17437 VPWR.n390 VGND 0.10822f
C17438 VPWR.t149 VGND 0.11957f
C17439 VPWR.t1247 VGND 0.07849f
C17440 VPWR.t491 VGND 0.09218f
C17441 VPWR.t150 VGND 0.03331f
C17442 VPWR.t492 VGND 0.02961f
C17443 VPWR.n391 VGND 0.09152f
C17444 VPWR.n392 VGND 0.01797f
C17445 VPWR.n393 VGND 0.00728f
C17446 VPWR.n394 VGND 0.10822f
C17447 VPWR.t683 VGND 0.11957f
C17448 VPWR.t632 VGND 0.07849f
C17449 VPWR.t738 VGND 0.09218f
C17450 VPWR.t684 VGND 0.03331f
C17451 VPWR.t739 VGND 0.02961f
C17452 VPWR.n395 VGND 0.09152f
C17453 VPWR.n396 VGND 0.01797f
C17454 VPWR.n397 VGND 0.00728f
C17455 VPWR.n398 VGND 0.10822f
C17456 VPWR.t762 VGND 0.11957f
C17457 VPWR.t631 VGND 0.07849f
C17458 VPWR.t1176 VGND 0.09218f
C17459 VPWR.t763 VGND 0.03331f
C17460 VPWR.t1177 VGND 0.02961f
C17461 VPWR.n399 VGND 0.09152f
C17462 VPWR.n400 VGND 0.01797f
C17463 VPWR.n401 VGND 0.00728f
C17464 VPWR.n402 VGND 0.10822f
C17465 VPWR.t1025 VGND 0.11957f
C17466 VPWR.t677 VGND 0.07849f
C17467 VPWR.t1248 VGND 0.09218f
C17468 VPWR.t1026 VGND 0.03331f
C17469 VPWR.t1249 VGND 0.02961f
C17470 VPWR.n403 VGND 0.09152f
C17471 VPWR.n404 VGND 0.01797f
C17472 VPWR.n405 VGND 0.00728f
C17473 VPWR.n406 VGND 0.10822f
C17474 VPWR.t918 VGND 0.11957f
C17475 VPWR.t207 VGND 0.07849f
C17476 VPWR.t271 VGND 0.09218f
C17477 VPWR.t919 VGND 0.03331f
C17478 VPWR.t272 VGND 0.02961f
C17479 VPWR.n407 VGND 0.09152f
C17480 VPWR.n408 VGND 0.01797f
C17481 VPWR.n409 VGND 0.00728f
C17482 VPWR.n410 VGND 0.10822f
C17483 VPWR.t235 VGND 0.11957f
C17484 VPWR.t206 VGND 0.07849f
C17485 VPWR.t1899 VGND 0.09218f
C17486 VPWR.t236 VGND 0.03331f
C17487 VPWR.t1900 VGND 0.02961f
C17488 VPWR.n411 VGND 0.09152f
C17489 VPWR.n412 VGND 0.01797f
C17490 VPWR.n413 VGND 0.00728f
C17491 VPWR.n414 VGND 0.10822f
C17492 VPWR.t1893 VGND 0.11957f
C17493 VPWR.t676 VGND 0.07849f
C17494 VPWR.t843 VGND 0.09218f
C17495 VPWR.t1894 VGND 0.03331f
C17496 VPWR.t844 VGND 0.02961f
C17497 VPWR.n415 VGND 0.09152f
C17498 VPWR.n416 VGND 0.01797f
C17499 VPWR.n417 VGND 0.00728f
C17500 VPWR.n418 VGND 0.10822f
C17501 VPWR.t941 VGND 0.11957f
C17502 VPWR.t675 VGND 0.07849f
C17503 VPWR.t501 VGND 0.09218f
C17504 VPWR.t942 VGND 0.03331f
C17505 VPWR.t502 VGND 0.02961f
C17506 VPWR.n419 VGND 0.09152f
C17507 VPWR.n420 VGND 0.01797f
C17508 VPWR.n421 VGND 0.00728f
C17509 VPWR.n422 VGND 0.10822f
C17510 VPWR.t495 VGND 0.11957f
C17511 VPWR.t208 VGND 0.07849f
C17512 VPWR.t551 VGND 0.09218f
C17513 VPWR.t496 VGND 0.03331f
C17514 VPWR.t552 VGND 0.02961f
C17515 VPWR.n423 VGND 0.09152f
C17516 VPWR.n424 VGND 0.01797f
C17517 VPWR.n425 VGND 0.00728f
C17518 VPWR.n426 VGND 0.10822f
C17519 VPWR.t545 VGND 0.11957f
C17520 VPWR.t630 VGND 0.07849f
C17521 VPWR.t1812 VGND 0.09218f
C17522 VPWR.t546 VGND 0.03331f
C17523 VPWR.t1813 VGND 0.02961f
C17524 VPWR.n427 VGND 0.09152f
C17525 VPWR.n428 VGND 0.01797f
C17526 VPWR.n429 VGND 0.00728f
C17527 VPWR.n430 VGND 0.10822f
C17528 VPWR.t447 VGND 0.11957f
C17529 VPWR.t629 VGND 0.07849f
C17530 VPWR.t865 VGND 0.09218f
C17531 VPWR.t448 VGND 0.03331f
C17532 VPWR.t866 VGND 0.02961f
C17533 VPWR.n431 VGND 0.09152f
C17534 VPWR.n432 VGND 0.01797f
C17535 VPWR.n433 VGND 0.00728f
C17536 VPWR.n434 VGND 0.10822f
C17537 VPWR.t859 VGND 0.11957f
C17538 VPWR.t205 VGND 0.07849f
C17539 VPWR.t108 VGND 0.09218f
C17540 VPWR.t860 VGND 0.03331f
C17541 VPWR.t109 VGND 0.02961f
C17542 VPWR.n435 VGND 0.09152f
C17543 VPWR.n436 VGND 0.01797f
C17544 VPWR.n437 VGND 0.00728f
C17545 VPWR.n438 VGND 0.10822f
C17546 VPWR.t1874 VGND 0.11957f
C17547 VPWR.t204 VGND 0.07849f
C17548 VPWR.t155 VGND 0.09218f
C17549 VPWR.t1875 VGND 0.03331f
C17550 VPWR.t156 VGND 0.02961f
C17551 VPWR.n439 VGND 0.09152f
C17552 VPWR.n440 VGND 0.01797f
C17553 VPWR.n441 VGND 0.00728f
C17554 VPWR.n442 VGND 0.10822f
C17555 VPWR.t1120 VGND 0.11957f
C17556 VPWR.t203 VGND 0.07849f
C17557 VPWR.t195 VGND 0.09218f
C17558 VPWR.t1121 VGND 0.03331f
C17559 VPWR.t196 VGND 0.02961f
C17560 VPWR.n443 VGND 0.09152f
C17561 VPWR.n444 VGND 0.01797f
C17562 VPWR.n445 VGND 0.00728f
C17563 VPWR.n446 VGND 0.10822f
C17564 VPWR.t320 VGND 0.11957f
C17565 VPWR.t674 VGND 0.07849f
C17566 VPWR.t1445 VGND 0.13333f
C17567 VPWR.n447 VGND 0.07618f
C17568 VPWR.n448 VGND 0.01797f
C17569 VPWR.n449 VGND 0.13913f
C17570 VPWR.n450 VGND 1.01577f
C17571 VPWR.n451 VGND 0.13913f
C17572 VPWR.t343 VGND 0.03331f
C17573 VPWR.t1561 VGND 0.02961f
C17574 VPWR.n452 VGND 0.09152f
C17575 VPWR.t322 VGND 0.09218f
C17576 VPWR.t325 VGND 0.03331f
C17577 VPWR.t323 VGND 0.02961f
C17578 VPWR.n453 VGND 0.09152f
C17579 VPWR.n454 VGND 0.13913f
C17580 VPWR.n455 VGND 0.13913f
C17581 VPWR.t1212 VGND 0.03331f
C17582 VPWR.t667 VGND 0.02961f
C17583 VPWR.n456 VGND 0.09152f
C17584 VPWR.t1878 VGND 0.09218f
C17585 VPWR.t1194 VGND 0.03331f
C17586 VPWR.t1879 VGND 0.02961f
C17587 VPWR.n457 VGND 0.09152f
C17588 VPWR.n458 VGND 0.13913f
C17589 VPWR.n459 VGND 0.13913f
C17590 VPWR.t1218 VGND 0.03331f
C17591 VPWR.t1186 VGND 0.02961f
C17592 VPWR.n460 VGND 0.09152f
C17593 VPWR.t1221 VGND 0.09218f
C17594 VPWR.t897 VGND 0.03331f
C17595 VPWR.t1222 VGND 0.02961f
C17596 VPWR.n461 VGND 0.09152f
C17597 VPWR.n462 VGND 0.13913f
C17598 VPWR.n463 VGND 0.13913f
C17599 VPWR.t136 VGND 0.03331f
C17600 VPWR.t905 VGND 0.02961f
C17601 VPWR.n464 VGND 0.09152f
C17602 VPWR.t139 VGND 0.09218f
C17603 VPWR.t286 VGND 0.03331f
C17604 VPWR.t140 VGND 0.02961f
C17605 VPWR.n465 VGND 0.09152f
C17606 VPWR.n466 VGND 0.13913f
C17607 VPWR.n467 VGND 0.13913f
C17608 VPWR.t353 VGND 0.03331f
C17609 VPWR.t556 VGND 0.02961f
C17610 VPWR.n468 VGND 0.09152f
C17611 VPWR.t356 VGND 0.09218f
C17612 VPWR.t793 VGND 0.03331f
C17613 VPWR.t357 VGND 0.02961f
C17614 VPWR.n469 VGND 0.09152f
C17615 VPWR.n470 VGND 0.13913f
C17616 VPWR.n471 VGND 0.13913f
C17617 VPWR.t1389 VGND 0.03331f
C17618 VPWR.t797 VGND 0.02961f
C17619 VPWR.n472 VGND 0.09152f
C17620 VPWR.t1392 VGND 0.09218f
C17621 VPWR.t1062 VGND 0.03331f
C17622 VPWR.t1393 VGND 0.02961f
C17623 VPWR.n473 VGND 0.09152f
C17624 VPWR.n474 VGND 0.13913f
C17625 VPWR.n475 VGND 0.13913f
C17626 VPWR.t779 VGND 0.03331f
C17627 VPWR.t603 VGND 0.02961f
C17628 VPWR.n476 VGND 0.09152f
C17629 VPWR.t756 VGND 0.09218f
C17630 VPWR.t219 VGND 0.03331f
C17631 VPWR.t757 VGND 0.02961f
C17632 VPWR.n477 VGND 0.09152f
C17633 VPWR.n478 VGND 0.13913f
C17634 VPWR.n479 VGND 0.13913f
C17635 VPWR.t1147 VGND 0.03331f
C17636 VPWR.t1288 VGND 0.02961f
C17637 VPWR.n480 VGND 0.09152f
C17638 VPWR.t1094 VGND 0.14512f
C17639 VPWR.t376 VGND 0.07849f
C17640 VPWR.t829 VGND 0.09218f
C17641 VPWR.t1095 VGND 0.03331f
C17642 VPWR.t830 VGND 0.02961f
C17643 VPWR.n481 VGND 0.09152f
C17644 VPWR.t1085 VGND 0.03331f
C17645 VPWR.t164 VGND 0.02961f
C17646 VPWR.n482 VGND 0.09152f
C17647 VPWR.t1084 VGND 0.14512f
C17648 VPWR.t978 VGND 0.07849f
C17649 VPWR.t163 VGND 0.09218f
C17650 VPWR.t182 VGND 0.03331f
C17651 VPWR.t1779 VGND 0.02961f
C17652 VPWR.n483 VGND 0.09152f
C17653 VPWR.n484 VGND 0.01797f
C17654 VPWR.n485 VGND 0.07618f
C17655 VPWR.t1778 VGND 0.13333f
C17656 VPWR.t1366 VGND 0.07849f
C17657 VPWR.t181 VGND 0.11957f
C17658 VPWR.t434 VGND 0.03331f
C17659 VPWR.t519 VGND 0.02961f
C17660 VPWR.n486 VGND 0.09152f
C17661 VPWR.n487 VGND 0.01797f
C17662 VPWR.n488 VGND 0.00728f
C17663 VPWR.n489 VGND 0.10822f
C17664 VPWR.t518 VGND 0.09218f
C17665 VPWR.t950 VGND 0.07849f
C17666 VPWR.t433 VGND 0.11957f
C17667 VPWR.t93 VGND 0.03331f
C17668 VPWR.t414 VGND 0.02961f
C17669 VPWR.n490 VGND 0.09152f
C17670 VPWR.n491 VGND 0.01797f
C17671 VPWR.n492 VGND 0.00728f
C17672 VPWR.n493 VGND 0.10822f
C17673 VPWR.t413 VGND 0.09218f
C17674 VPWR.t973 VGND 0.07849f
C17675 VPWR.t92 VGND 0.11957f
C17676 VPWR.t854 VGND 0.03331f
C17677 VPWR.t64 VGND 0.02961f
C17678 VPWR.n494 VGND 0.09152f
C17679 VPWR.n495 VGND 0.01797f
C17680 VPWR.n496 VGND 0.00728f
C17681 VPWR.n497 VGND 0.10822f
C17682 VPWR.t63 VGND 0.09218f
C17683 VPWR.t974 VGND 0.07849f
C17684 VPWR.t853 VGND 0.11957f
C17685 VPWR.t122 VGND 0.03331f
C17686 VPWR.t1105 VGND 0.02961f
C17687 VPWR.n498 VGND 0.09152f
C17688 VPWR.n499 VGND 0.01797f
C17689 VPWR.n500 VGND 0.00728f
C17690 VPWR.n501 VGND 0.10822f
C17691 VPWR.t1104 VGND 0.09218f
C17692 VPWR.t979 VGND 0.07849f
C17693 VPWR.t121 VGND 0.11957f
C17694 VPWR.t1371 VGND 0.03331f
C17695 VPWR.t126 VGND 0.02961f
C17696 VPWR.n502 VGND 0.09152f
C17697 VPWR.n503 VGND 0.01797f
C17698 VPWR.n504 VGND 0.00728f
C17699 VPWR.n505 VGND 0.10822f
C17700 VPWR.t125 VGND 0.09218f
C17701 VPWR.t980 VGND 0.07849f
C17702 VPWR.t1370 VGND 0.11957f
C17703 VPWR.t512 VGND 0.03331f
C17704 VPWR.t1381 VGND 0.02961f
C17705 VPWR.n506 VGND 0.09152f
C17706 VPWR.n507 VGND 0.01797f
C17707 VPWR.n508 VGND 0.00728f
C17708 VPWR.n509 VGND 0.10822f
C17709 VPWR.t1380 VGND 0.09218f
C17710 VPWR.t977 VGND 0.07849f
C17711 VPWR.t511 VGND 0.11957f
C17712 VPWR.t466 VGND 0.03331f
C17713 VPWR.t640 VGND 0.02961f
C17714 VPWR.n510 VGND 0.09152f
C17715 VPWR.n511 VGND 0.01797f
C17716 VPWR.n512 VGND 0.00728f
C17717 VPWR.n513 VGND 0.10822f
C17718 VPWR.t639 VGND 0.09218f
C17719 VPWR.t1367 VGND 0.07849f
C17720 VPWR.t465 VGND 0.11957f
C17721 VPWR.t291 VGND 0.03331f
C17722 VPWR.t578 VGND 0.02961f
C17723 VPWR.n514 VGND 0.09152f
C17724 VPWR.n515 VGND 0.01797f
C17725 VPWR.n516 VGND 0.00728f
C17726 VPWR.n517 VGND 0.10822f
C17727 VPWR.t577 VGND 0.09218f
C17728 VPWR.t1368 VGND 0.07849f
C17729 VPWR.t290 VGND 0.11957f
C17730 VPWR.t274 VGND 0.03331f
C17731 VPWR.t295 VGND 0.02961f
C17732 VPWR.n518 VGND 0.09152f
C17733 VPWR.n519 VGND 0.01797f
C17734 VPWR.n520 VGND 0.00728f
C17735 VPWR.n521 VGND 0.10822f
C17736 VPWR.t294 VGND 0.09218f
C17737 VPWR.t975 VGND 0.07849f
C17738 VPWR.t273 VGND 0.11957f
C17739 VPWR.t168 VGND 0.03331f
C17740 VPWR.t256 VGND 0.02961f
C17741 VPWR.n522 VGND 0.09152f
C17742 VPWR.n523 VGND 0.01797f
C17743 VPWR.n524 VGND 0.00728f
C17744 VPWR.n525 VGND 0.10822f
C17745 VPWR.t255 VGND 0.09218f
C17746 VPWR.t976 VGND 0.07849f
C17747 VPWR.t167 VGND 0.11957f
C17748 VPWR.t607 VGND 0.03331f
C17749 VPWR.t172 VGND 0.02961f
C17750 VPWR.n526 VGND 0.09152f
C17751 VPWR.n527 VGND 0.01797f
C17752 VPWR.n528 VGND 0.00728f
C17753 VPWR.n529 VGND 0.10822f
C17754 VPWR.t171 VGND 0.09218f
C17755 VPWR.t1369 VGND 0.07849f
C17756 VPWR.t606 VGND 0.11957f
C17757 VPWR.t755 VGND 0.03331f
C17758 VPWR.t1008 VGND 0.02961f
C17759 VPWR.n530 VGND 0.09152f
C17760 VPWR.n531 VGND 0.01797f
C17761 VPWR.n532 VGND 0.00728f
C17762 VPWR.n533 VGND 0.10822f
C17763 VPWR.t1007 VGND 0.09218f
C17764 VPWR.t981 VGND 0.07849f
C17765 VPWR.t754 VGND 0.11957f
C17766 VPWR.t504 VGND 0.03331f
C17767 VPWR.t731 VGND 0.02961f
C17768 VPWR.n534 VGND 0.09152f
C17769 VPWR.n535 VGND 0.01797f
C17770 VPWR.n536 VGND 0.00728f
C17771 VPWR.n537 VGND 0.10822f
C17772 VPWR.t730 VGND 0.09218f
C17773 VPWR.t949 VGND 0.07849f
C17774 VPWR.t503 VGND 0.11957f
C17775 VPWR.t176 VGND 0.03331f
C17776 VPWR.t508 VGND 0.02961f
C17777 VPWR.n538 VGND 0.09152f
C17778 VPWR.n539 VGND 0.01797f
C17779 VPWR.n540 VGND 0.00728f
C17780 VPWR.n541 VGND 0.10822f
C17781 VPWR.t507 VGND 0.09218f
C17782 VPWR.t1365 VGND 0.07849f
C17783 VPWR.t175 VGND 0.11957f
C17784 VPWR.n542 VGND 0.10822f
C17785 VPWR.n543 VGND 0.00728f
C17786 VPWR.n544 VGND 0.01797f
C17787 VPWR.n545 VGND 0.13913f
C17788 VPWR.n546 VGND 1.0094f
C17789 VPWR.n547 VGND 0.13913f
C17790 VPWR.t1070 VGND 0.03331f
C17791 VPWR.t1165 VGND 0.02961f
C17792 VPWR.n548 VGND 0.09152f
C17793 VPWR.t1069 VGND 0.14512f
C17794 VPWR.t1807 VGND 0.07849f
C17795 VPWR.t1164 VGND 0.09218f
C17796 VPWR.t226 VGND 0.11957f
C17797 VPWR.t1157 VGND 0.03331f
C17798 VPWR.t1261 VGND 0.02961f
C17799 VPWR.n549 VGND 0.09152f
C17800 VPWR.n550 VGND 0.13913f
C17801 VPWR.n551 VGND 0.13913f
C17802 VPWR.t227 VGND 0.03331f
C17803 VPWR.t769 VGND 0.02961f
C17804 VPWR.n552 VGND 0.09152f
C17805 VPWR.t1345 VGND 0.07849f
C17806 VPWR.t768 VGND 0.09218f
C17807 VPWR.t1017 VGND 0.11957f
C17808 VPWR.t733 VGND 0.03331f
C17809 VPWR.t1821 VGND 0.02961f
C17810 VPWR.n553 VGND 0.09152f
C17811 VPWR.n554 VGND 0.13913f
C17812 VPWR.n555 VGND 0.13913f
C17813 VPWR.t1018 VGND 0.03331f
C17814 VPWR.t480 VGND 0.02961f
C17815 VPWR.n556 VGND 0.09152f
C17816 VPWR.t1806 VGND 0.07849f
C17817 VPWR.t479 VGND 0.09218f
C17818 VPWR.t241 VGND 0.11957f
C17819 VPWR.t1237 VGND 0.03331f
C17820 VPWR.t250 VGND 0.02961f
C17821 VPWR.n557 VGND 0.09152f
C17822 VPWR.n558 VGND 0.13913f
C17823 VPWR.n559 VGND 0.13913f
C17824 VPWR.t242 VGND 0.03331f
C17825 VPWR.t432 VGND 0.02961f
C17826 VPWR.n560 VGND 0.09152f
C17827 VPWR.t1349 VGND 0.07849f
C17828 VPWR.t431 VGND 0.09218f
C17829 VPWR.t583 VGND 0.11957f
C17830 VPWR.t424 VGND 0.03331f
C17831 VPWR.t993 VGND 0.02961f
C17832 VPWR.n561 VGND 0.09152f
C17833 VPWR.n562 VGND 0.13913f
C17834 VPWR.n563 VGND 0.13913f
C17835 VPWR.t584 VGND 0.03331f
C17836 VPWR.t692 VGND 0.02961f
C17837 VPWR.n564 VGND 0.09152f
C17838 VPWR.t1804 VGND 0.07849f
C17839 VPWR.t691 VGND 0.09218f
C17840 VPWR.t1303 VGND 0.11957f
C17841 VPWR.t1277 VGND 0.03331f
C17842 VPWR.t893 VGND 0.02961f
C17843 VPWR.n565 VGND 0.09152f
C17844 VPWR.n566 VGND 0.13913f
C17845 VPWR.n567 VGND 0.13913f
C17846 VPWR.t1304 VGND 0.03331f
C17847 VPWR.t1319 VGND 0.02961f
C17848 VPWR.n568 VGND 0.09152f
C17849 VPWR.t1343 VGND 0.07849f
C17850 VPWR.t1318 VGND 0.09218f
C17851 VPWR.t1836 VGND 0.11957f
C17852 VPWR.t54 VGND 0.03331f
C17853 VPWR.t1190 VGND 0.02961f
C17854 VPWR.n569 VGND 0.09152f
C17855 VPWR.n570 VGND 0.13913f
C17856 VPWR.n571 VGND 0.13913f
C17857 VPWR.t1837 VGND 0.03331f
C17858 VPWR.t1867 VGND 0.02961f
C17859 VPWR.n572 VGND 0.09152f
C17860 VPWR.t1348 VGND 0.07849f
C17861 VPWR.t1866 VGND 0.09218f
C17862 VPWR.t626 VGND 0.11957f
C17863 VPWR.t70 VGND 0.03331f
C17864 VPWR.t7 VGND 0.02961f
C17865 VPWR.n573 VGND 0.09152f
C17866 VPWR.n574 VGND 0.13913f
C17867 VPWR.n575 VGND 0.13913f
C17868 VPWR.t627 VGND 0.03331f
C17869 VPWR.t311 VGND 0.02961f
C17870 VPWR.n576 VGND 0.09152f
C17871 VPWR.t1346 VGND 0.07849f
C17872 VPWR.t310 VGND 0.09218f
C17873 VPWR.t529 VGND 0.03331f
C17874 VPWR.t1628 VGND 0.02961f
C17875 VPWR.n577 VGND 0.09152f
C17876 VPWR.t188 VGND 0.03331f
C17877 VPWR.t1736 VGND 0.02961f
C17878 VPWR.n578 VGND 0.09152f
C17879 VPWR.t1077 VGND 0.14512f
C17880 VPWR.t944 VGND 0.07849f
C17881 VPWR.t1001 VGND 0.09218f
C17882 VPWR.t1078 VGND 0.03331f
C17883 VPWR.t1002 VGND 0.02961f
C17884 VPWR.n579 VGND 0.09152f
C17885 VPWR.n580 VGND 0.01797f
C17886 VPWR.n581 VGND 0.00728f
C17887 VPWR.n582 VGND 0.10822f
C17888 VPWR.t159 VGND 0.11957f
C17889 VPWR.t1049 VGND 0.07849f
C17890 VPWR.t1285 VGND 0.09218f
C17891 VPWR.t160 VGND 0.03331f
C17892 VPWR.t1286 VGND 0.02961f
C17893 VPWR.n583 VGND 0.09152f
C17894 VPWR.n584 VGND 0.01797f
C17895 VPWR.n585 VGND 0.00728f
C17896 VPWR.n586 VGND 0.10822f
C17897 VPWR.t485 VGND 0.11957f
C17898 VPWR.t948 VGND 0.07849f
C17899 VPWR.t722 VGND 0.09218f
C17900 VPWR.t486 VGND 0.03331f
C17901 VPWR.t723 VGND 0.02961f
C17902 VPWR.n587 VGND 0.09152f
C17903 VPWR.n588 VGND 0.01797f
C17904 VPWR.n589 VGND 0.00728f
C17905 VPWR.n590 VGND 0.10822f
C17906 VPWR.t746 VGND 0.11957f
C17907 VPWR.t947 VGND 0.07849f
C17908 VPWR.t1019 VGND 0.09218f
C17909 VPWR.t747 VGND 0.03331f
C17910 VPWR.t1020 VGND 0.02961f
C17911 VPWR.n591 VGND 0.09152f
C17912 VPWR.n592 VGND 0.01797f
C17913 VPWR.n593 VGND 0.00728f
C17914 VPWR.n594 VGND 0.10822f
C17915 VPWR.t1168 VGND 0.11957f
C17916 VPWR.t943 VGND 0.07849f
C17917 VPWR.t618 VGND 0.09218f
C17918 VPWR.t1169 VGND 0.03331f
C17919 VPWR.t619 VGND 0.02961f
C17920 VPWR.n595 VGND 0.09152f
C17921 VPWR.n596 VGND 0.01797f
C17922 VPWR.n597 VGND 0.00728f
C17923 VPWR.n598 VGND 0.10822f
C17924 VPWR.t612 VGND 0.11957f
C17925 VPWR.t1047 VGND 0.07849f
C17926 VPWR.t275 VGND 0.09218f
C17927 VPWR.t613 VGND 0.03331f
C17928 VPWR.t276 VGND 0.02961f
C17929 VPWR.n599 VGND 0.09152f
C17930 VPWR.n600 VGND 0.01797f
C17931 VPWR.n601 VGND 0.00728f
C17932 VPWR.n602 VGND 0.10822f
C17933 VPWR.t261 VGND 0.11957f
C17934 VPWR.t1046 VGND 0.07849f
C17935 VPWR.t306 VGND 0.09218f
C17936 VPWR.t262 VGND 0.03331f
C17937 VPWR.t307 VGND 0.02961f
C17938 VPWR.n603 VGND 0.09152f
C17939 VPWR.n604 VGND 0.01797f
C17940 VPWR.n605 VGND 0.00728f
C17941 VPWR.n606 VGND 0.10822f
C17942 VPWR.t300 VGND 0.11957f
C17943 VPWR.t1052 VGND 0.07849f
C17944 VPWR.t589 VGND 0.09218f
C17945 VPWR.t301 VGND 0.03331f
C17946 VPWR.t590 VGND 0.02961f
C17947 VPWR.n607 VGND 0.09152f
C17948 VPWR.n608 VGND 0.01797f
C17949 VPWR.n609 VGND 0.00728f
C17950 VPWR.n610 VGND 0.10822f
C17951 VPWR.t473 VGND 0.11957f
C17952 VPWR.t1051 VGND 0.07849f
C17953 VPWR.t571 VGND 0.09218f
C17954 VPWR.t474 VGND 0.03331f
C17955 VPWR.t572 VGND 0.02961f
C17956 VPWR.n611 VGND 0.09152f
C17957 VPWR.n612 VGND 0.01797f
C17958 VPWR.n613 VGND 0.00728f
C17959 VPWR.n614 VGND 0.10822f
C17960 VPWR.t565 VGND 0.11957f
C17961 VPWR.t1048 VGND 0.07849f
C17962 VPWR.t1910 VGND 0.09218f
C17963 VPWR.t566 VGND 0.03331f
C17964 VPWR.t1911 VGND 0.02961f
C17965 VPWR.n615 VGND 0.09152f
C17966 VPWR.n616 VGND 0.01797f
C17967 VPWR.n617 VGND 0.00728f
C17968 VPWR.n618 VGND 0.10822f
C17969 VPWR.t1376 VGND 0.11957f
C17970 VPWR.t946 VGND 0.07849f
C17971 VPWR.t1359 VGND 0.09218f
C17972 VPWR.t1377 VGND 0.03331f
C17973 VPWR.t1360 VGND 0.02961f
C17974 VPWR.n619 VGND 0.09152f
C17975 VPWR.n620 VGND 0.01797f
C17976 VPWR.n621 VGND 0.00728f
C17977 VPWR.n622 VGND 0.10822f
C17978 VPWR.t131 VGND 0.11957f
C17979 VPWR.t945 VGND 0.07849f
C17980 VPWR.t1850 VGND 0.09218f
C17981 VPWR.t132 VGND 0.03331f
C17982 VPWR.t1851 VGND 0.02961f
C17983 VPWR.n623 VGND 0.09152f
C17984 VPWR.n624 VGND 0.01797f
C17985 VPWR.n625 VGND 0.00728f
C17986 VPWR.n626 VGND 0.10822f
C17987 VPWR.t1100 VGND 0.11957f
C17988 VPWR.t1045 VGND 0.07849f
C17989 VPWR.t1203 VGND 0.09218f
C17990 VPWR.t1101 VGND 0.03331f
C17991 VPWR.t1204 VGND 0.02961f
C17992 VPWR.n627 VGND 0.09152f
C17993 VPWR.n628 VGND 0.01797f
C17994 VPWR.n629 VGND 0.00728f
C17995 VPWR.n630 VGND 0.10822f
C17996 VPWR.t100 VGND 0.11957f
C17997 VPWR.t1044 VGND 0.07849f
C17998 VPWR.t1126 VGND 0.09218f
C17999 VPWR.t101 VGND 0.03331f
C18000 VPWR.t1127 VGND 0.02961f
C18001 VPWR.n631 VGND 0.09152f
C18002 VPWR.n632 VGND 0.01797f
C18003 VPWR.n633 VGND 0.00728f
C18004 VPWR.n634 VGND 0.10822f
C18005 VPWR.t409 VGND 0.11957f
C18006 VPWR.t513 VGND 0.07849f
C18007 VPWR.t530 VGND 0.09218f
C18008 VPWR.t410 VGND 0.03331f
C18009 VPWR.t531 VGND 0.02961f
C18010 VPWR.n635 VGND 0.09152f
C18011 VPWR.n636 VGND 0.01797f
C18012 VPWR.n637 VGND 0.00728f
C18013 VPWR.n638 VGND 0.10822f
C18014 VPWR.t187 VGND 0.11957f
C18015 VPWR.t1050 VGND 0.07849f
C18016 VPWR.t1735 VGND 0.13333f
C18017 VPWR.n639 VGND 0.07618f
C18018 VPWR.n640 VGND 0.01797f
C18019 VPWR.n641 VGND 0.13913f
C18020 VPWR.n642 VGND 1.01577f
C18021 VPWR.n643 VGND 0.13913f
C18022 VPWR.t315 VGND 0.03331f
C18023 VPWR.t1462 VGND 0.02961f
C18024 VPWR.n644 VGND 0.09152f
C18025 VPWR.t189 VGND 0.09218f
C18026 VPWR.t1117 VGND 0.03331f
C18027 VPWR.t190 VGND 0.02961f
C18028 VPWR.n645 VGND 0.09152f
C18029 VPWR.n646 VGND 0.13913f
C18030 VPWR.n647 VGND 0.13913f
C18031 VPWR.t1871 VGND 0.03331f
C18032 VPWR.t152 VGND 0.02961f
C18033 VPWR.n648 VGND 0.09152f
C18034 VPWR.t104 VGND 0.09218f
C18035 VPWR.t956 VGND 0.03331f
C18036 VPWR.t105 VGND 0.02961f
C18037 VPWR.n649 VGND 0.09152f
C18038 VPWR.n650 VGND 0.13913f
C18039 VPWR.n651 VGND 0.13913f
C18040 VPWR.t444 VGND 0.03331f
C18041 VPWR.t862 VGND 0.02961f
C18042 VPWR.n652 VGND 0.09152f
C18043 VPWR.t1808 VGND 0.09218f
C18044 VPWR.t542 VGND 0.03331f
C18045 VPWR.t1809 VGND 0.02961f
C18046 VPWR.n653 VGND 0.09152f
C18047 VPWR.n654 VGND 0.13913f
C18048 VPWR.n655 VGND 0.13913f
C18049 VPWR.t371 VGND 0.03331f
C18050 VPWR.t548 VGND 0.02961f
C18051 VPWR.n656 VGND 0.09152f
C18052 VPWR.t497 VGND 0.09218f
C18053 VPWR.t938 VGND 0.03331f
C18054 VPWR.t498 VGND 0.02961f
C18055 VPWR.n657 VGND 0.09152f
C18056 VPWR.n658 VGND 0.13913f
C18057 VPWR.n659 VGND 0.13913f
C18058 VPWR.t1890 VGND 0.03331f
C18059 VPWR.t840 VGND 0.02961f
C18060 VPWR.n660 VGND 0.09152f
C18061 VPWR.t1895 VGND 0.09218f
C18062 VPWR.t232 VGND 0.03331f
C18063 VPWR.t1896 VGND 0.02961f
C18064 VPWR.n661 VGND 0.09152f
C18065 VPWR.n662 VGND 0.13913f
C18066 VPWR.n663 VGND 0.13913f
C18067 VPWR.t1228 VGND 0.03331f
C18068 VPWR.t268 VGND 0.02961f
C18069 VPWR.n664 VGND 0.09152f
C18070 VPWR.t209 VGND 0.09218f
C18071 VPWR.t1825 VGND 0.03331f
C18072 VPWR.t210 VGND 0.02961f
C18073 VPWR.n665 VGND 0.09152f
C18074 VPWR.n666 VGND 0.13913f
C18075 VPWR.n667 VGND 0.13913f
C18076 VPWR.t767 VGND 0.03331f
C18077 VPWR.t1171 VGND 0.02961f
C18078 VPWR.n668 VGND 0.09152f
C18079 VPWR.t742 VGND 0.09218f
C18080 VPWR.t680 VGND 0.03331f
C18081 VPWR.t743 VGND 0.02961f
C18082 VPWR.n669 VGND 0.09152f
C18083 VPWR.n670 VGND 0.13913f
C18084 VPWR.n671 VGND 0.13913f
C18085 VPWR.t146 VGND 0.03331f
C18086 VPWR.t686 VGND 0.02961f
C18087 VPWR.n672 VGND 0.09152f
C18088 VPWR.t1090 VGND 0.14512f
C18089 VPWR.t199 VGND 0.07849f
C18090 VPWR.t595 VGND 0.09218f
C18091 VPWR.t1091 VGND 0.03331f
C18092 VPWR.t596 VGND 0.02961f
C18093 VPWR.n673 VGND 0.09152f
C18094 VPWR.t1097 VGND 0.03331f
C18095 VPWR.t826 VGND 0.02961f
C18096 VPWR.n674 VGND 0.09152f
C18097 VPWR.t1096 VGND 0.14512f
C18098 VPWR.t705 VGND 0.07849f
C18099 VPWR.t825 VGND 0.09218f
C18100 VPWR.t341 VGND 0.03331f
C18101 VPWR.t1569 VGND 0.02961f
C18102 VPWR.n675 VGND 0.09152f
C18103 VPWR.n676 VGND 0.01797f
C18104 VPWR.n677 VGND 0.07618f
C18105 VPWR.t1568 VGND 0.13333f
C18106 VPWR.t47 VGND 0.07849f
C18107 VPWR.t340 VGND 0.11957f
C18108 VPWR.t9 VGND 0.03331f
C18109 VPWR.t319 VGND 0.02961f
C18110 VPWR.n678 VGND 0.09152f
C18111 VPWR.n679 VGND 0.01797f
C18112 VPWR.n680 VGND 0.00728f
C18113 VPWR.n681 VGND 0.10822f
C18114 VPWR.t318 VGND 0.09218f
C18115 VPWR.t908 VGND 0.07849f
C18116 VPWR.t8 VGND 0.11957f
C18117 VPWR.t1210 VGND 0.03331f
C18118 VPWR.t329 VGND 0.02961f
C18119 VPWR.n682 VGND 0.09152f
C18120 VPWR.n683 VGND 0.01797f
C18121 VPWR.n684 VGND 0.00728f
C18122 VPWR.n685 VGND 0.10822f
C18123 VPWR.t328 VGND 0.09218f
C18124 VPWR.t909 VGND 0.07849f
C18125 VPWR.t1209 VGND 0.11957f
C18126 VPWR.t1192 VGND 0.03331f
C18127 VPWR.t1877 VGND 0.02961f
C18128 VPWR.n686 VGND 0.09152f
C18129 VPWR.n687 VGND 0.01797f
C18130 VPWR.n688 VGND 0.00728f
C18131 VPWR.n689 VGND 0.10822f
C18132 VPWR.t1876 VGND 0.09218f
C18133 VPWR.t1197 VGND 0.07849f
C18134 VPWR.t1191 VGND 0.11957f
C18135 VPWR.t1323 VGND 0.03331f
C18136 VPWR.t1182 VGND 0.02961f
C18137 VPWR.n690 VGND 0.09152f
C18138 VPWR.n691 VGND 0.01797f
C18139 VPWR.n692 VGND 0.00728f
C18140 VPWR.n693 VGND 0.10822f
C18141 VPWR.t1181 VGND 0.09218f
C18142 VPWR.t706 VGND 0.07849f
C18143 VPWR.t1322 VGND 0.11957f
C18144 VPWR.t895 VGND 0.03331f
C18145 VPWR.t1220 VGND 0.02961f
C18146 VPWR.n694 VGND 0.09152f
C18147 VPWR.n695 VGND 0.01797f
C18148 VPWR.n696 VGND 0.00728f
C18149 VPWR.n697 VGND 0.10822f
C18150 VPWR.t1219 VGND 0.09218f
C18151 VPWR.t707 VGND 0.07849f
C18152 VPWR.t894 VGND 0.11957f
C18153 VPWR.t696 VGND 0.03331f
C18154 VPWR.t901 VGND 0.02961f
C18155 VPWR.n698 VGND 0.09152f
C18156 VPWR.n699 VGND 0.01797f
C18157 VPWR.n700 VGND 0.00728f
C18158 VPWR.n701 VGND 0.10822f
C18159 VPWR.t900 VGND 0.09218f
C18160 VPWR.t1200 VGND 0.07849f
C18161 VPWR.t695 VGND 0.11957f
C18162 VPWR.t284 VGND 0.03331f
C18163 VPWR.t138 VGND 0.02961f
C18164 VPWR.n702 VGND 0.09152f
C18165 VPWR.n703 VGND 0.01797f
C18166 VPWR.n704 VGND 0.00728f
C18167 VPWR.n705 VGND 0.10822f
C18168 VPWR.t137 VGND 0.09218f
C18169 VPWR.t48 VGND 0.07849f
C18170 VPWR.t283 VGND 0.11957f
C18171 VPWR.t351 VGND 0.03331f
C18172 VPWR.t554 VGND 0.02961f
C18173 VPWR.n706 VGND 0.09152f
C18174 VPWR.n707 VGND 0.01797f
C18175 VPWR.n708 VGND 0.00728f
C18176 VPWR.n709 VGND 0.10822f
C18177 VPWR.t553 VGND 0.09218f
C18178 VPWR.t289 VGND 0.07849f
C18179 VPWR.t350 VGND 0.11957f
C18180 VPWR.t791 VGND 0.03331f
C18181 VPWR.t355 VGND 0.02961f
C18182 VPWR.n710 VGND 0.09152f
C18183 VPWR.n711 VGND 0.01797f
C18184 VPWR.n712 VGND 0.00728f
C18185 VPWR.n713 VGND 0.10822f
C18186 VPWR.t354 VGND 0.09218f
C18187 VPWR.t1198 VGND 0.07849f
C18188 VPWR.t790 VGND 0.11957f
C18189 VPWR.t1387 VGND 0.03331f
C18190 VPWR.t795 VGND 0.02961f
C18191 VPWR.n714 VGND 0.09152f
C18192 VPWR.n715 VGND 0.01797f
C18193 VPWR.n716 VGND 0.00728f
C18194 VPWR.n717 VGND 0.10822f
C18195 VPWR.t794 VGND 0.09218f
C18196 VPWR.t1199 VGND 0.07849f
C18197 VPWR.t1386 VGND 0.11957f
C18198 VPWR.t1060 VGND 0.03331f
C18199 VPWR.t1391 VGND 0.02961f
C18200 VPWR.n718 VGND 0.09152f
C18201 VPWR.n719 VGND 0.01797f
C18202 VPWR.n720 VGND 0.00728f
C18203 VPWR.n721 VGND 0.10822f
C18204 VPWR.t1390 VGND 0.09218f
C18205 VPWR.t704 VGND 0.07849f
C18206 VPWR.t1059 VGND 0.11957f
C18207 VPWR.t781 VGND 0.03331f
C18208 VPWR.t1024 VGND 0.02961f
C18209 VPWR.n722 VGND 0.09152f
C18210 VPWR.n723 VGND 0.01797f
C18211 VPWR.n724 VGND 0.00728f
C18212 VPWR.n725 VGND 0.10822f
C18213 VPWR.t1023 VGND 0.09218f
C18214 VPWR.t906 VGND 0.07849f
C18215 VPWR.t780 VGND 0.11957f
C18216 VPWR.t217 VGND 0.03331f
C18217 VPWR.t759 VGND 0.02961f
C18218 VPWR.n726 VGND 0.09152f
C18219 VPWR.n727 VGND 0.01797f
C18220 VPWR.n728 VGND 0.00728f
C18221 VPWR.n729 VGND 0.10822f
C18222 VPWR.t758 VGND 0.09218f
C18223 VPWR.t907 VGND 0.07849f
C18224 VPWR.t216 VGND 0.11957f
C18225 VPWR.t1145 VGND 0.03331f
C18226 VPWR.t221 VGND 0.02961f
C18227 VPWR.n730 VGND 0.09152f
C18228 VPWR.n731 VGND 0.01797f
C18229 VPWR.n732 VGND 0.00728f
C18230 VPWR.n733 VGND 0.10822f
C18231 VPWR.t220 VGND 0.09218f
C18232 VPWR.t46 VGND 0.07849f
C18233 VPWR.t1144 VGND 0.11957f
C18234 VPWR.n734 VGND 0.10822f
C18235 VPWR.n735 VGND 0.00728f
C18236 VPWR.n736 VGND 0.01797f
C18237 VPWR.n737 VGND 0.13913f
C18238 VPWR.n738 VGND 1.0094f
C18239 VPWR.n739 VGND 0.13913f
C18240 VPWR.t1093 VGND 0.03331f
C18241 VPWR.t144 VGND 0.02961f
C18242 VPWR.n740 VGND 0.09152f
C18243 VPWR.t1092 VGND 0.14512f
C18244 VPWR.t1883 VGND 0.07849f
C18245 VPWR.t143 VGND 0.09218f
C18246 VPWR.t1289 VGND 0.11957f
C18247 VPWR.t828 VGND 0.03331f
C18248 VPWR.t1292 VGND 0.02961f
C18249 VPWR.n741 VGND 0.09152f
C18250 VPWR.n742 VGND 0.13913f
C18251 VPWR.n743 VGND 0.13913f
C18252 VPWR.t1290 VGND 0.03331f
C18253 VPWR.t751 VGND 0.02961f
C18254 VPWR.n744 VGND 0.09152f
C18255 VPWR.t379 VGND 0.07849f
C18256 VPWR.t750 VGND 0.09218f
C18257 VPWR.t1814 VGND 0.11957f
C18258 VPWR.t775 VGND 0.03331f
C18259 VPWR.t605 VGND 0.02961f
C18260 VPWR.n745 VGND 0.09152f
C18261 VPWR.n746 VGND 0.13913f
C18262 VPWR.n747 VGND 0.13913f
C18263 VPWR.t1815 VGND 0.03331f
C18264 VPWR.t1226 VGND 0.02961f
C18265 VPWR.n748 VGND 0.09152f
C18266 VPWR.t1882 VGND 0.07849f
C18267 VPWR.t1225 VGND 0.09218f
C18268 VPWR.t798 VGND 0.11957f
C18269 VPWR.t1224 VGND 0.03331f
C18270 VPWR.t230 VGND 0.02961f
C18271 VPWR.n749 VGND 0.09152f
C18272 VPWR.n750 VGND 0.13913f
C18273 VPWR.n751 VGND 0.13913f
C18274 VPWR.t799 VGND 0.03331f
C18275 VPWR.t1888 VGND 0.02961f
C18276 VPWR.n752 VGND 0.09152f
C18277 VPWR.t383 VGND 0.07849f
C18278 VPWR.t1887 VGND 0.09218f
C18279 VPWR.t986 VGND 0.11957f
C18280 VPWR.t359 VGND 0.03331f
C18281 VPWR.t468 VGND 0.02961f
C18282 VPWR.n753 VGND 0.09152f
C18283 VPWR.n754 VGND 0.13913f
C18284 VPWR.n755 VGND 0.13913f
C18285 VPWR.t987 VGND 0.03331f
C18286 VPWR.t369 VGND 0.02961f
C18287 VPWR.n756 VGND 0.09152f
C18288 VPWR.t1880 VGND 0.07849f
C18289 VPWR.t368 VGND 0.09218f
C18290 VPWR.t902 VGND 0.11957f
C18291 VPWR.t142 VGND 0.03331f
C18292 VPWR.t540 VGND 0.02961f
C18293 VPWR.n757 VGND 0.09152f
C18294 VPWR.n758 VGND 0.13913f
C18295 VPWR.n759 VGND 0.13913f
C18296 VPWR.t903 VGND 0.03331f
C18297 VPWR.t442 VGND 0.02961f
C18298 VPWR.n760 VGND 0.09152f
C18299 VPWR.t1885 VGND 0.07849f
C18300 VPWR.t441 VGND 0.09218f
C18301 VPWR.t1183 VGND 0.11957f
C18302 VPWR.t1115 VGND 0.03331f
C18303 VPWR.t954 VGND 0.02961f
C18304 VPWR.n761 VGND 0.09152f
C18305 VPWR.n762 VGND 0.13913f
C18306 VPWR.n763 VGND 0.13913f
C18307 VPWR.t1184 VGND 0.03331f
C18308 VPWR.t95 VGND 0.02961f
C18309 VPWR.n764 VGND 0.09152f
C18310 VPWR.t382 VGND 0.07849f
C18311 VPWR.t94 VGND 0.09218f
C18312 VPWR.t664 VGND 0.11957f
C18313 VPWR.t1214 VGND 0.03331f
C18314 VPWR.t669 VGND 0.02961f
C18315 VPWR.n765 VGND 0.09152f
C18316 VPWR.n766 VGND 0.13913f
C18317 VPWR.n767 VGND 0.13913f
C18318 VPWR.t665 VGND 0.03331f
C18319 VPWR.t180 VGND 0.02961f
C18320 VPWR.n768 VGND 0.09152f
C18321 VPWR.t380 VGND 0.07849f
C18322 VPWR.t179 VGND 0.09218f
C18323 VPWR.t345 VGND 0.03331f
C18324 VPWR.t1529 VGND 0.02961f
C18325 VPWR.n769 VGND 0.09152f
C18326 VPWR.t525 VGND 0.03331f
C18327 VPWR.t1634 VGND 0.02961f
C18328 VPWR.n770 VGND 0.09152f
C18329 VPWR.t1071 VGND 0.14512f
C18330 VPWR.t1339 VGND 0.07849f
C18331 VPWR.t1162 VGND 0.09218f
C18332 VPWR.t1072 VGND 0.03331f
C18333 VPWR.t1163 VGND 0.02961f
C18334 VPWR.n771 VGND 0.09152f
C18335 VPWR.n772 VGND 0.01797f
C18336 VPWR.n773 VGND 0.00728f
C18337 VPWR.n774 VGND 0.10822f
C18338 VPWR.t458 VGND 0.11957f
C18339 VPWR.t1334 VGND 0.07849f
C18340 VPWR.t1256 VGND 0.09218f
C18341 VPWR.t459 VGND 0.03331f
C18342 VPWR.t1257 VGND 0.02961f
C18343 VPWR.n775 VGND 0.09152f
C18344 VPWR.n776 VGND 0.01797f
C18345 VPWR.n777 VGND 0.00728f
C18346 VPWR.n778 VGND 0.10822f
C18347 VPWR.t224 VGND 0.11957f
C18348 VPWR.t1030 VGND 0.07849f
C18349 VPWR.t770 VGND 0.09218f
C18350 VPWR.t225 VGND 0.03331f
C18351 VPWR.t771 VGND 0.02961f
C18352 VPWR.n779 VGND 0.09152f
C18353 VPWR.n780 VGND 0.01797f
C18354 VPWR.n781 VGND 0.00728f
C18355 VPWR.n782 VGND 0.10822f
C18356 VPWR.t734 VGND 0.11957f
C18357 VPWR.t1029 VGND 0.07849f
C18358 VPWR.t1818 VGND 0.09218f
C18359 VPWR.t735 VGND 0.03331f
C18360 VPWR.t1819 VGND 0.02961f
C18361 VPWR.n783 VGND 0.09152f
C18362 VPWR.n784 VGND 0.01797f
C18363 VPWR.n785 VGND 0.00728f
C18364 VPWR.n786 VGND 0.10822f
C18365 VPWR.t1013 VGND 0.11957f
C18366 VPWR.t1338 VGND 0.07849f
C18367 VPWR.t475 VGND 0.09218f
C18368 VPWR.t1014 VGND 0.03331f
C18369 VPWR.t476 VGND 0.02961f
C18370 VPWR.n787 VGND 0.09152f
C18371 VPWR.n788 VGND 0.01797f
C18372 VPWR.n789 VGND 0.00728f
C18373 VPWR.n790 VGND 0.10822f
C18374 VPWR.t1234 VGND 0.11957f
C18375 VPWR.t1035 VGND 0.07849f
C18376 VPWR.t245 VGND 0.09218f
C18377 VPWR.t1235 VGND 0.03331f
C18378 VPWR.t246 VGND 0.02961f
C18379 VPWR.n791 VGND 0.09152f
C18380 VPWR.n792 VGND 0.01797f
C18381 VPWR.n793 VGND 0.00728f
C18382 VPWR.n794 VGND 0.10822f
C18383 VPWR.t239 VGND 0.11957f
C18384 VPWR.t1034 VGND 0.07849f
C18385 VPWR.t427 VGND 0.09218f
C18386 VPWR.t240 VGND 0.03331f
C18387 VPWR.t428 VGND 0.02961f
C18388 VPWR.n795 VGND 0.09152f
C18389 VPWR.n796 VGND 0.01797f
C18390 VPWR.n797 VGND 0.00728f
C18391 VPWR.n798 VGND 0.10822f
C18392 VPWR.t421 VGND 0.11957f
C18393 VPWR.t1337 VGND 0.07849f
C18394 VPWR.t990 VGND 0.09218f
C18395 VPWR.t422 VGND 0.03331f
C18396 VPWR.t991 VGND 0.02961f
C18397 VPWR.n799 VGND 0.09152f
C18398 VPWR.n800 VGND 0.01797f
C18399 VPWR.n801 VGND 0.00728f
C18400 VPWR.n802 VGND 0.10822f
C18401 VPWR.t579 VGND 0.11957f
C18402 VPWR.t1336 VGND 0.07849f
C18403 VPWR.t1280 VGND 0.09218f
C18404 VPWR.t580 VGND 0.03331f
C18405 VPWR.t1281 VGND 0.02961f
C18406 VPWR.n803 VGND 0.09152f
C18407 VPWR.n804 VGND 0.01797f
C18408 VPWR.n805 VGND 0.00728f
C18409 VPWR.n806 VGND 0.10822f
C18410 VPWR.t1274 VGND 0.11957f
C18411 VPWR.t1036 VGND 0.07849f
C18412 VPWR.t890 VGND 0.09218f
C18413 VPWR.t1275 VGND 0.03331f
C18414 VPWR.t891 VGND 0.02961f
C18415 VPWR.n807 VGND 0.09152f
C18416 VPWR.n808 VGND 0.01797f
C18417 VPWR.n809 VGND 0.00728f
C18418 VPWR.n810 VGND 0.10822f
C18419 VPWR.t1301 VGND 0.11957f
C18420 VPWR.t1028 VGND 0.07849f
C18421 VPWR.t1314 VGND 0.09218f
C18422 VPWR.t1302 VGND 0.03331f
C18423 VPWR.t1315 VGND 0.02961f
C18424 VPWR.n811 VGND 0.09152f
C18425 VPWR.n812 VGND 0.01797f
C18426 VPWR.n813 VGND 0.00728f
C18427 VPWR.n814 VGND 0.10822f
C18428 VPWR.t51 VGND 0.11957f
C18429 VPWR.t1027 VGND 0.07849f
C18430 VPWR.t1187 VGND 0.09218f
C18431 VPWR.t52 VGND 0.03331f
C18432 VPWR.t1188 VGND 0.02961f
C18433 VPWR.n815 VGND 0.09152f
C18434 VPWR.n816 VGND 0.01797f
C18435 VPWR.n817 VGND 0.00728f
C18436 VPWR.n818 VGND 0.10822f
C18437 VPWR.t1834 VGND 0.11957f
C18438 VPWR.t1033 VGND 0.07849f
C18439 VPWR.t1864 VGND 0.09218f
C18440 VPWR.t1835 VGND 0.03331f
C18441 VPWR.t1865 VGND 0.02961f
C18442 VPWR.n819 VGND 0.09152f
C18443 VPWR.n820 VGND 0.01797f
C18444 VPWR.n821 VGND 0.00728f
C18445 VPWR.n822 VGND 0.10822f
C18446 VPWR.t65 VGND 0.11957f
C18447 VPWR.t1032 VGND 0.07849f
C18448 VPWR.t4 VGND 0.09218f
C18449 VPWR.t66 VGND 0.03331f
C18450 VPWR.t5 VGND 0.02961f
C18451 VPWR.n823 VGND 0.09152f
C18452 VPWR.n824 VGND 0.01797f
C18453 VPWR.n825 VGND 0.00728f
C18454 VPWR.n826 VGND 0.10822f
C18455 VPWR.t624 VGND 0.11957f
C18456 VPWR.t1031 VGND 0.07849f
C18457 VPWR.t348 VGND 0.09218f
C18458 VPWR.t625 VGND 0.03331f
C18459 VPWR.t349 VGND 0.02961f
C18460 VPWR.n827 VGND 0.09152f
C18461 VPWR.n828 VGND 0.01797f
C18462 VPWR.n829 VGND 0.00728f
C18463 VPWR.n830 VGND 0.10822f
C18464 VPWR.t524 VGND 0.11957f
C18465 VPWR.t1335 VGND 0.07849f
C18466 VPWR.t1633 VGND 0.13333f
C18467 VPWR.n831 VGND 0.07618f
C18468 VPWR.n832 VGND 0.01797f
C18469 VPWR.n833 VGND 0.13913f
C18470 VPWR.n834 VGND 1.01577f
C18471 VPWR.n835 VGND 0.13913f
C18472 VPWR.t317 VGND 0.03331f
C18473 VPWR.t1454 VGND 0.02961f
C18474 VPWR.n836 VGND 0.09152f
C18475 VPWR.t193 VGND 0.09218f
C18476 VPWR.t1119 VGND 0.03331f
C18477 VPWR.t194 VGND 0.02961f
C18478 VPWR.n837 VGND 0.09152f
C18479 VPWR.n838 VGND 0.13913f
C18480 VPWR.n839 VGND 0.13913f
C18481 VPWR.t1873 VGND 0.03331f
C18482 VPWR.t154 VGND 0.02961f
C18483 VPWR.n840 VGND 0.09152f
C18484 VPWR.t106 VGND 0.09218f
C18485 VPWR.t858 VGND 0.03331f
C18486 VPWR.t107 VGND 0.02961f
C18487 VPWR.n841 VGND 0.09152f
C18488 VPWR.n842 VGND 0.13913f
C18489 VPWR.n843 VGND 0.13913f
C18490 VPWR.t446 VGND 0.03331f
C18491 VPWR.t864 VGND 0.02961f
C18492 VPWR.n844 VGND 0.09152f
C18493 VPWR.t1810 VGND 0.09218f
C18494 VPWR.t544 VGND 0.03331f
C18495 VPWR.t1811 VGND 0.02961f
C18496 VPWR.n845 VGND 0.09152f
C18497 VPWR.n846 VGND 0.13913f
C18498 VPWR.n847 VGND 0.13913f
C18499 VPWR.t494 VGND 0.03331f
C18500 VPWR.t550 VGND 0.02961f
C18501 VPWR.n848 VGND 0.09152f
C18502 VPWR.t499 VGND 0.09218f
C18503 VPWR.t940 VGND 0.03331f
C18504 VPWR.t500 VGND 0.02961f
C18505 VPWR.n849 VGND 0.09152f
C18506 VPWR.n850 VGND 0.13913f
C18507 VPWR.n851 VGND 0.13913f
C18508 VPWR.t1892 VGND 0.03331f
C18509 VPWR.t842 VGND 0.02961f
C18510 VPWR.n852 VGND 0.09152f
C18511 VPWR.t1897 VGND 0.09218f
C18512 VPWR.t234 VGND 0.03331f
C18513 VPWR.t1898 VGND 0.02961f
C18514 VPWR.n853 VGND 0.09152f
C18515 VPWR.n854 VGND 0.13913f
C18516 VPWR.n855 VGND 0.13913f
C18517 VPWR.t917 VGND 0.03331f
C18518 VPWR.t270 VGND 0.02961f
C18519 VPWR.n856 VGND 0.09152f
C18520 VPWR.t211 VGND 0.09218f
C18521 VPWR.t1022 VGND 0.03331f
C18522 VPWR.t212 VGND 0.02961f
C18523 VPWR.n857 VGND 0.09152f
C18524 VPWR.n858 VGND 0.13913f
C18525 VPWR.n859 VGND 0.13913f
C18526 VPWR.t765 VGND 0.03331f
C18527 VPWR.t1175 VGND 0.02961f
C18528 VPWR.n860 VGND 0.09152f
C18529 VPWR.t740 VGND 0.09218f
C18530 VPWR.t682 VGND 0.03331f
C18531 VPWR.t741 VGND 0.02961f
C18532 VPWR.n861 VGND 0.09152f
C18533 VPWR.n862 VGND 0.13913f
C18534 VPWR.n863 VGND 0.13913f
C18535 VPWR.t148 VGND 0.03331f
C18536 VPWR.t688 VGND 0.02961f
C18537 VPWR.n864 VGND 0.09152f
C18538 VPWR.t1088 VGND 0.14512f
C18539 VPWR.t363 VGND 0.07849f
C18540 VPWR.t597 VGND 0.09218f
C18541 VPWR.t1089 VGND 0.03331f
C18542 VPWR.t598 VGND 0.02961f
C18543 VPWR.n865 VGND 0.09152f
C18544 VPWR.t1074 VGND 0.03331f
C18545 VPWR.t1161 VGND 0.02961f
C18546 VPWR.n866 VGND 0.09152f
C18547 VPWR.t1073 VGND 0.14512f
C18548 VPWR.t120 VGND 0.07849f
C18549 VPWR.t1160 VGND 0.09218f
C18550 VPWR.t523 VGND 0.03331f
C18551 VPWR.t1641 VGND 0.02961f
C18552 VPWR.n867 VGND 0.09152f
C18553 VPWR.n868 VGND 0.01797f
C18554 VPWR.n869 VGND 0.07618f
C18555 VPWR.t1640 VGND 0.13333f
C18556 VPWR.t116 VGND 0.07849f
C18557 VPWR.t522 VGND 0.11957f
C18558 VPWR.t623 VGND 0.03331f
C18559 VPWR.t347 VGND 0.02961f
C18560 VPWR.n870 VGND 0.09152f
C18561 VPWR.n871 VGND 0.01797f
C18562 VPWR.n872 VGND 0.00728f
C18563 VPWR.n873 VGND 0.10822f
C18564 VPWR.t346 VGND 0.09218f
C18565 VPWR.t872 VGND 0.07849f
C18566 VPWR.t622 VGND 0.11957f
C18567 VPWR.t62 VGND 0.03331f
C18568 VPWR.t3 VGND 0.02961f
C18569 VPWR.n874 VGND 0.09152f
C18570 VPWR.n875 VGND 0.01797f
C18571 VPWR.n876 VGND 0.00728f
C18572 VPWR.n877 VGND 0.10822f
C18573 VPWR.t2 VGND 0.09218f
C18574 VPWR.t873 VGND 0.07849f
C18575 VPWR.t61 VGND 0.11957f
C18576 VPWR.t1833 VGND 0.03331f
C18577 VPWR.t1863 VGND 0.02961f
C18578 VPWR.n878 VGND 0.09152f
C18579 VPWR.n879 VGND 0.01797f
C18580 VPWR.n880 VGND 0.00728f
C18581 VPWR.n881 VGND 0.10822f
C18582 VPWR.t1862 VGND 0.09218f
C18583 VPWR.t874 VGND 0.07849f
C18584 VPWR.t1832 VGND 0.11957f
C18585 VPWR.t50 VGND 0.03331f
C18586 VPWR.t1841 VGND 0.02961f
C18587 VPWR.n882 VGND 0.09152f
C18588 VPWR.n883 VGND 0.01797f
C18589 VPWR.n884 VGND 0.00728f
C18590 VPWR.n885 VGND 0.10822f
C18591 VPWR.t1840 VGND 0.09218f
C18592 VPWR.t1229 VGND 0.07849f
C18593 VPWR.t49 VGND 0.11957f
C18594 VPWR.t1300 VGND 0.03331f
C18595 VPWR.t56 VGND 0.02961f
C18596 VPWR.n886 VGND 0.09152f
C18597 VPWR.n887 VGND 0.01797f
C18598 VPWR.n888 VGND 0.00728f
C18599 VPWR.n889 VGND 0.10822f
C18600 VPWR.t55 VGND 0.09218f
C18601 VPWR.t1230 VGND 0.07849f
C18602 VPWR.t1299 VGND 0.11957f
C18603 VPWR.t1273 VGND 0.03331f
C18604 VPWR.t889 VGND 0.02961f
C18605 VPWR.n890 VGND 0.09152f
C18606 VPWR.n891 VGND 0.01797f
C18607 VPWR.n892 VGND 0.00728f
C18608 VPWR.n893 VGND 0.10822f
C18609 VPWR.t888 VGND 0.09218f
C18610 VPWR.t877 VGND 0.07849f
C18611 VPWR.t1272 VGND 0.11957f
C18612 VPWR.t576 VGND 0.03331f
C18613 VPWR.t1279 VGND 0.02961f
C18614 VPWR.n894 VGND 0.09152f
C18615 VPWR.n895 VGND 0.01797f
C18616 VPWR.n896 VGND 0.00728f
C18617 VPWR.n897 VGND 0.10822f
C18618 VPWR.t1278 VGND 0.09218f
C18619 VPWR.t117 VGND 0.07849f
C18620 VPWR.t575 VGND 0.11957f
C18621 VPWR.t420 VGND 0.03331f
C18622 VPWR.t989 VGND 0.02961f
C18623 VPWR.n898 VGND 0.09152f
C18624 VPWR.n899 VGND 0.01797f
C18625 VPWR.n900 VGND 0.00728f
C18626 VPWR.n901 VGND 0.10822f
C18627 VPWR.t988 VGND 0.09218f
C18628 VPWR.t118 VGND 0.07849f
C18629 VPWR.t419 VGND 0.11957f
C18630 VPWR.t238 VGND 0.03331f
C18631 VPWR.t426 VGND 0.02961f
C18632 VPWR.n902 VGND 0.09152f
C18633 VPWR.n903 VGND 0.01797f
C18634 VPWR.n904 VGND 0.00728f
C18635 VPWR.n905 VGND 0.10822f
C18636 VPWR.t425 VGND 0.09218f
C18637 VPWR.t875 VGND 0.07849f
C18638 VPWR.t237 VGND 0.11957f
C18639 VPWR.t1233 VGND 0.03331f
C18640 VPWR.t244 VGND 0.02961f
C18641 VPWR.n906 VGND 0.09152f
C18642 VPWR.n907 VGND 0.01797f
C18643 VPWR.n908 VGND 0.00728f
C18644 VPWR.n909 VGND 0.10822f
C18645 VPWR.t243 VGND 0.09218f
C18646 VPWR.t876 VGND 0.07849f
C18647 VPWR.t1232 VGND 0.11957f
C18648 VPWR.t1012 VGND 0.03331f
C18649 VPWR.t1239 VGND 0.02961f
C18650 VPWR.n910 VGND 0.09152f
C18651 VPWR.n911 VGND 0.01797f
C18652 VPWR.n912 VGND 0.00728f
C18653 VPWR.n913 VGND 0.10822f
C18654 VPWR.t1238 VGND 0.09218f
C18655 VPWR.t119 VGND 0.07849f
C18656 VPWR.t1011 VGND 0.11957f
C18657 VPWR.t737 VGND 0.03331f
C18658 VPWR.t1817 VGND 0.02961f
C18659 VPWR.n914 VGND 0.09152f
C18660 VPWR.n915 VGND 0.01797f
C18661 VPWR.n916 VGND 0.00728f
C18662 VPWR.n917 VGND 0.10822f
C18663 VPWR.t1816 VGND 0.09218f
C18664 VPWR.t1231 VGND 0.07849f
C18665 VPWR.t736 VGND 0.11957f
C18666 VPWR.t223 VGND 0.03331f
C18667 VPWR.t773 VGND 0.02961f
C18668 VPWR.n918 VGND 0.09152f
C18669 VPWR.n919 VGND 0.01797f
C18670 VPWR.n920 VGND 0.00728f
C18671 VPWR.n921 VGND 0.10822f
C18672 VPWR.t772 VGND 0.09218f
C18673 VPWR.t871 VGND 0.07849f
C18674 VPWR.t222 VGND 0.11957f
C18675 VPWR.t457 VGND 0.03331f
C18676 VPWR.t1255 VGND 0.02961f
C18677 VPWR.n922 VGND 0.09152f
C18678 VPWR.n923 VGND 0.01797f
C18679 VPWR.n924 VGND 0.00728f
C18680 VPWR.n925 VGND 0.10822f
C18681 VPWR.t1254 VGND 0.09218f
C18682 VPWR.t115 VGND 0.07849f
C18683 VPWR.t456 VGND 0.11957f
C18684 VPWR.n926 VGND 0.10822f
C18685 VPWR.n927 VGND 0.00728f
C18686 VPWR.n928 VGND 0.01797f
C18687 VPWR.n929 VGND 0.13913f
C18688 VPWR.n930 VGND 1.0094f
C18689 VPWR.n931 VGND 0.13913f
C18690 VPWR.t1080 VGND 0.03331f
C18691 VPWR.t1000 VGND 0.02961f
C18692 VPWR.n932 VGND 0.09152f
C18693 VPWR.t1079 VGND 0.14512f
C18694 VPWR.t21 VGND 0.07849f
C18695 VPWR.t999 VGND 0.09218f
C18696 VPWR.t509 VGND 0.11957f
C18697 VPWR.t158 VGND 0.03331f
C18698 VPWR.t490 VGND 0.02961f
C18699 VPWR.n933 VGND 0.09152f
C18700 VPWR.n934 VGND 0.13913f
C18701 VPWR.n935 VGND 0.13913f
C18702 VPWR.t510 VGND 0.03331f
C18703 VPWR.t725 VGND 0.02961f
C18704 VPWR.n936 VGND 0.09152f
C18705 VPWR.t1333 VGND 0.07849f
C18706 VPWR.t724 VGND 0.09218f
C18707 VPWR.t1166 VGND 0.11957f
C18708 VPWR.t749 VGND 0.03331f
C18709 VPWR.t1016 VGND 0.02961f
C18710 VPWR.n937 VGND 0.09152f
C18711 VPWR.n938 VGND 0.13913f
C18712 VPWR.n939 VGND 0.13913f
C18713 VPWR.t1167 VGND 0.03331f
C18714 VPWR.t617 VGND 0.02961f
C18715 VPWR.n940 VGND 0.09152f
C18716 VPWR.t20 VGND 0.07849f
C18717 VPWR.t616 VGND 0.09218f
C18718 VPWR.t257 VGND 0.11957f
C18719 VPWR.t174 VGND 0.03331f
C18720 VPWR.t266 VGND 0.02961f
C18721 VPWR.n941 VGND 0.09152f
C18722 VPWR.n942 VGND 0.13913f
C18723 VPWR.n943 VGND 0.13913f
C18724 VPWR.t258 VGND 0.03331f
C18725 VPWR.t305 VGND 0.02961f
C18726 VPWR.n944 VGND 0.09152f
C18727 VPWR.t1153 VGND 0.07849f
C18728 VPWR.t304 VGND 0.09218f
C18729 VPWR.t471 VGND 0.11957f
C18730 VPWR.t297 VGND 0.03331f
C18731 VPWR.t586 VGND 0.02961f
C18732 VPWR.n945 VGND 0.09152f
C18733 VPWR.n946 VGND 0.13913f
C18734 VPWR.n947 VGND 0.13913f
C18735 VPWR.t472 VGND 0.03331f
C18736 VPWR.t570 VGND 0.02961f
C18737 VPWR.n948 VGND 0.09152f
C18738 VPWR.t1332 VGND 0.07849f
C18739 VPWR.t569 VGND 0.09218f
C18740 VPWR.t1374 VGND 0.11957f
C18741 VPWR.t642 VGND 0.03331f
C18742 VPWR.t1385 VGND 0.02961f
C18743 VPWR.n949 VGND 0.09152f
C18744 VPWR.n950 VGND 0.13913f
C18745 VPWR.n951 VGND 0.13913f
C18746 VPWR.t1375 VGND 0.03331f
C18747 VPWR.t1358 VGND 0.02961f
C18748 VPWR.n952 VGND 0.09152f
C18749 VPWR.t23 VGND 0.07849f
C18750 VPWR.t1357 VGND 0.09218f
C18751 VPWR.t1098 VGND 0.11957f
C18752 VPWR.t128 VGND 0.03331f
C18753 VPWR.t1849 VGND 0.02961f
C18754 VPWR.n953 VGND 0.09152f
C18755 VPWR.n954 VGND 0.13913f
C18756 VPWR.n955 VGND 0.13913f
C18757 VPWR.t1099 VGND 0.03331f
C18758 VPWR.t72 VGND 0.02961f
C18759 VPWR.n956 VGND 0.09152f
C18760 VPWR.t1152 VGND 0.07849f
C18761 VPWR.t71 VGND 0.09218f
C18762 VPWR.t407 VGND 0.11957f
C18763 VPWR.t99 VGND 0.03331f
C18764 VPWR.t1125 VGND 0.02961f
C18765 VPWR.n957 VGND 0.09152f
C18766 VPWR.n958 VGND 0.13913f
C18767 VPWR.n959 VGND 0.13913f
C18768 VPWR.t408 VGND 0.03331f
C18769 VPWR.t527 VGND 0.02961f
C18770 VPWR.n960 VGND 0.09152f
C18771 VPWR.t1150 VGND 0.07849f
C18772 VPWR.t526 VGND 0.09218f
C18773 VPWR.t186 VGND 0.03331f
C18774 VPWR.t1749 VGND 0.02961f
C18775 VPWR.n961 VGND 0.09152f
C18776 VPWR.t337 VGND 0.03331f
C18777 VPWR.t1601 VGND 0.02961f
C18778 VPWR.n962 VGND 0.09152f
C18779 VPWR.t1067 VGND 0.14512f
C18780 VPWR.t697 VGND 0.07849f
C18781 VPWR.t1148 VGND 0.09218f
C18782 VPWR.t1068 VGND 0.03331f
C18783 VPWR.t1149 VGND 0.02961f
C18784 VPWR.n963 VGND 0.09152f
C18785 VPWR.n964 VGND 0.01797f
C18786 VPWR.n965 VGND 0.00728f
C18787 VPWR.n966 VGND 0.10822f
C18788 VPWR.t1158 VGND 0.11957f
C18789 VPWR.t215 VGND 0.07849f
C18790 VPWR.t1262 VGND 0.09218f
C18791 VPWR.t1159 VGND 0.03331f
C18792 VPWR.t1263 VGND 0.02961f
C18793 VPWR.n967 VGND 0.09152f
C18794 VPWR.n968 VGND 0.01797f
C18795 VPWR.n969 VGND 0.00728f
C18796 VPWR.n970 VGND 0.10822f
C18797 VPWR.t1258 VGND 0.11957f
C18798 VPWR.t701 VGND 0.07849f
C18799 VPWR.t760 VGND 0.09218f
C18800 VPWR.t1259 VGND 0.03331f
C18801 VPWR.t761 VGND 0.02961f
C18802 VPWR.n971 VGND 0.09152f
C18803 VPWR.n972 VGND 0.01797f
C18804 VPWR.n973 VGND 0.00728f
C18805 VPWR.n974 VGND 0.10822f
C18806 VPWR.t726 VGND 0.11957f
C18807 VPWR.t700 VGND 0.07849f
C18808 VPWR.t1822 VGND 0.09218f
C18809 VPWR.t727 VGND 0.03331f
C18810 VPWR.t1823 VGND 0.02961f
C18811 VPWR.n975 VGND 0.09152f
C18812 VPWR.n976 VGND 0.01797f
C18813 VPWR.n977 VGND 0.00728f
C18814 VPWR.n978 VGND 0.10822f
C18815 VPWR.t1055 VGND 0.11957f
C18816 VPWR.t636 VGND 0.07849f
C18817 VPWR.t481 VGND 0.09218f
C18818 VPWR.t1056 VGND 0.03331f
C18819 VPWR.t482 VGND 0.02961f
C18820 VPWR.n979 VGND 0.09152f
C18821 VPWR.n980 VGND 0.01797f
C18822 VPWR.n981 VGND 0.00728f
C18823 VPWR.n982 VGND 0.10822f
C18824 VPWR.t477 VGND 0.11957f
C18825 VPWR.t213 VGND 0.07849f
C18826 VPWR.t251 VGND 0.09218f
C18827 VPWR.t478 VGND 0.03331f
C18828 VPWR.t252 VGND 0.02961f
C18829 VPWR.n983 VGND 0.09152f
C18830 VPWR.n984 VGND 0.01797f
C18831 VPWR.n985 VGND 0.00728f
C18832 VPWR.n986 VGND 0.10822f
C18833 VPWR.t247 VGND 0.11957f
C18834 VPWR.t985 VGND 0.07849f
C18835 VPWR.t1005 VGND 0.09218f
C18836 VPWR.t248 VGND 0.03331f
C18837 VPWR.t1006 VGND 0.02961f
C18838 VPWR.n987 VGND 0.09152f
C18839 VPWR.n988 VGND 0.01797f
C18840 VPWR.n989 VGND 0.00728f
C18841 VPWR.n990 VGND 0.10822f
C18842 VPWR.t429 VGND 0.11957f
C18843 VPWR.t635 VGND 0.07849f
C18844 VPWR.t935 VGND 0.09218f
C18845 VPWR.t430 VGND 0.03331f
C18846 VPWR.t936 VGND 0.02961f
C18847 VPWR.n991 VGND 0.09152f
C18848 VPWR.n992 VGND 0.01797f
C18849 VPWR.n993 VGND 0.00728f
C18850 VPWR.n994 VGND 0.10822f
C18851 VPWR.t587 VGND 0.11957f
C18852 VPWR.t634 VGND 0.07849f
C18853 VPWR.t693 VGND 0.09218f
C18854 VPWR.t588 VGND 0.03331f
C18855 VPWR.t694 VGND 0.02961f
C18856 VPWR.n995 VGND 0.09152f
C18857 VPWR.n996 VGND 0.01797f
C18858 VPWR.n997 VGND 0.00728f
C18859 VPWR.n998 VGND 0.10822f
C18860 VPWR.t689 VGND 0.11957f
C18861 VPWR.t214 VGND 0.07849f
C18862 VPWR.t898 VGND 0.09218f
C18863 VPWR.t690 VGND 0.03331f
C18864 VPWR.t899 VGND 0.02961f
C18865 VPWR.n999 VGND 0.09152f
C18866 VPWR.n1000 VGND 0.01797f
C18867 VPWR.n1001 VGND 0.00728f
C18868 VPWR.n1002 VGND 0.10822f
C18869 VPWR.t1305 VGND 0.11957f
C18870 VPWR.t699 VGND 0.07849f
C18871 VPWR.t1320 VGND 0.09218f
C18872 VPWR.t1306 VGND 0.03331f
C18873 VPWR.t1321 VGND 0.02961f
C18874 VPWR.n1003 VGND 0.09152f
C18875 VPWR.n1004 VGND 0.01797f
C18876 VPWR.n1005 VGND 0.00728f
C18877 VPWR.n1006 VGND 0.10822f
C18878 VPWR.t1316 VGND 0.11957f
C18879 VPWR.t698 VGND 0.07849f
C18880 VPWR.t1195 VGND 0.09218f
C18881 VPWR.t1317 VGND 0.03331f
C18882 VPWR.t1196 VGND 0.02961f
C18883 VPWR.n1007 VGND 0.09152f
C18884 VPWR.n1008 VGND 0.01797f
C18885 VPWR.n1009 VGND 0.00728f
C18886 VPWR.n1010 VGND 0.10822f
C18887 VPWR.t1838 VGND 0.11957f
C18888 VPWR.t984 VGND 0.07849f
C18889 VPWR.t1868 VGND 0.09218f
C18890 VPWR.t1839 VGND 0.03331f
C18891 VPWR.t1869 VGND 0.02961f
C18892 VPWR.n1011 VGND 0.09152f
C18893 VPWR.n1012 VGND 0.01797f
C18894 VPWR.n1013 VGND 0.00728f
C18895 VPWR.n1014 VGND 0.10822f
C18896 VPWR.t1201 VGND 0.11957f
C18897 VPWR.t983 VGND 0.07849f
C18898 VPWR.t326 VGND 0.09218f
C18899 VPWR.t1202 VGND 0.03331f
C18900 VPWR.t327 VGND 0.02961f
C18901 VPWR.n1015 VGND 0.09152f
C18902 VPWR.n1016 VGND 0.01797f
C18903 VPWR.n1017 VGND 0.00728f
C18904 VPWR.n1018 VGND 0.10822f
C18905 VPWR.t0 VGND 0.11957f
C18906 VPWR.t982 VGND 0.07849f
C18907 VPWR.t312 VGND 0.09218f
C18908 VPWR.t1 VGND 0.03331f
C18909 VPWR.t313 VGND 0.02961f
C18910 VPWR.n1019 VGND 0.09152f
C18911 VPWR.n1020 VGND 0.01797f
C18912 VPWR.n1021 VGND 0.00728f
C18913 VPWR.n1022 VGND 0.10822f
C18914 VPWR.t336 VGND 0.11957f
C18915 VPWR.t633 VGND 0.07849f
C18916 VPWR.t1600 VGND 0.13333f
C18917 VPWR.n1023 VGND 0.07618f
C18918 VPWR.n1024 VGND 0.01797f
C18919 VPWR.n1025 VGND 0.13913f
C18920 VPWR.n1026 VGND 6.02311f
C18921 VPWR.n1027 VGND 0.06567f
C18922 VPWR.n1028 VGND -0.01866f
C18923 VPWR.t2061 VGND 0.01116f
C18924 VPWR.t1602 VGND 0.01222f
C18925 VPWR.n1029 VGND 0.03042f
C18926 VPWR.n1030 VGND 0.00581f
C18927 VPWR.t1604 VGND 0.02679f
C18928 VPWR.n1031 VGND 0.05724f
C18929 VPWR.t1712 VGND 0.02961f
C18930 VPWR.n1032 VGND 0.04692f
C18931 VPWR.t338 VGND 0.09218f
C18932 VPWR.t1957 VGND 0.01116f
C18933 VPWR.t1494 VGND 0.01222f
C18934 VPWR.n1033 VGND 0.03042f
C18935 VPWR.n1034 VGND 0.00581f
C18936 VPWR.t1496 VGND 0.02679f
C18937 VPWR.n1035 VGND 0.05724f
C18938 VPWR.t339 VGND 0.02961f
C18939 VPWR.n1036 VGND 0.04692f
C18940 VPWR.n1037 VGND -0.01866f
C18941 VPWR.n1038 VGND 0.06567f
C18942 VPWR.t2065 VGND 0.01136f
C18943 VPWR.t1450 VGND 0.0124f
C18944 VPWR.n1039 VGND 0.02769f
C18945 VPWR.n1040 VGND 0.01897f
C18946 VPWR.n1041 VGND 0.06244f
C18947 VPWR.n1042 VGND 0.09746f
C18948 VPWR.n1043 VGND 0.0544f
C18949 VPWR.n1044 VGND 0.06567f
C18950 VPWR.n1045 VGND -0.01866f
C18951 VPWR.t1967 VGND 0.01116f
C18952 VPWR.t1580 VGND 0.01222f
C18953 VPWR.n1046 VGND 0.03042f
C18954 VPWR.n1047 VGND 0.00581f
C18955 VPWR.t1582 VGND 0.02679f
C18956 VPWR.n1048 VGND 0.05724f
C18957 VPWR.t114 VGND 0.02961f
C18958 VPWR.n1049 VGND 0.04692f
C18959 VPWR.t113 VGND 0.09218f
C18960 VPWR.t1458 VGND 0.11957f
C18961 VPWR.t2055 VGND 0.01116f
C18962 VPWR.t1621 VGND 0.01222f
C18963 VPWR.n1050 VGND 0.03042f
C18964 VPWR.n1051 VGND 0.00581f
C18965 VPWR.t1623 VGND 0.02679f
C18966 VPWR.n1052 VGND 0.05724f
C18967 VPWR.t1208 VGND 0.02961f
C18968 VPWR.n1053 VGND 0.04692f
C18969 VPWR.n1054 VGND 0.00805f
C18970 VPWR.n1055 VGND 0.19371f
C18971 VPWR.n1056 VGND 0.08351f
C18972 VPWR.n1057 VGND 0.03437f
C18973 VPWR.t1676 VGND 0.03331f
C18974 VPWR.t1668 VGND 0.02961f
C18975 VPWR.n1058 VGND 0.09152f
C18976 VPWR.t1667 VGND 0.09218f
C18977 VPWR.t1423 VGND 0.11957f
C18978 VPWR.t1704 VGND 0.03331f
C18979 VPWR.t1696 VGND 0.02961f
C18980 VPWR.n1059 VGND 0.09152f
C18981 VPWR.n1060 VGND 0.00805f
C18982 VPWR.t1424 VGND 0.03331f
C18983 VPWR.t1547 VGND 0.02961f
C18984 VPWR.n1061 VGND 0.09152f
C18985 VPWR.t1419 VGND 0.07849f
C18986 VPWR.t1546 VGND 0.13333f
C18987 VPWR.n1062 VGND 0.07615f
C18988 VPWR.n1063 VGND 0.01698f
C18989 VPWR.t2034 VGND 0.0112f
C18990 VPWR.t1545 VGND 0.01226f
C18991 VPWR.n1064 VGND 0.02993f
C18992 VPWR.n1065 VGND 0.03284f
C18993 VPWR.n1066 VGND 0.00697f
C18994 VPWR.n1067 VGND 0.01822f
C18995 VPWR.n1068 VGND 0.17585f
C18996 VPWR.t1989 VGND 0.0112f
C18997 VPWR.t1666 VGND 0.01226f
C18998 VPWR.n1069 VGND 0.02993f
C18999 VPWR.n1070 VGND 0.03284f
C19000 VPWR.n1071 VGND 0.01714f
C19001 VPWR.n1072 VGND 0.00697f
C19002 VPWR.n1073 VGND 0.00805f
C19003 VPWR.n1074 VGND 0.01714f
C19004 VPWR.n1075 VGND 0.00697f
C19005 VPWR.t1988 VGND 0.01136f
C19006 VPWR.t1672 VGND 0.0124f
C19007 VPWR.n1076 VGND 0.02768f
C19008 VPWR.n1077 VGND 0.02818f
C19009 VPWR.n1078 VGND 0.01822f
C19010 VPWR.n1079 VGND 0.17585f
C19011 VPWR.t1947 VGND 0.0112f
C19012 VPWR.t1774 VGND 0.01226f
C19013 VPWR.n1080 VGND 0.02993f
C19014 VPWR.n1081 VGND 0.03284f
C19015 VPWR.n1082 VGND 0.01714f
C19016 VPWR.n1083 VGND 0.00697f
C19017 VPWR.n1084 VGND 0.01714f
C19018 VPWR.n1085 VGND 0.00697f
C19019 VPWR.t1945 VGND 0.01136f
C19020 VPWR.t1780 VGND 0.0124f
C19021 VPWR.n1086 VGND 0.02768f
C19022 VPWR.n1087 VGND 0.02818f
C19023 VPWR.n1088 VGND 0.01822f
C19024 VPWR.n1089 VGND 0.17585f
C19025 VPWR.t1949 VGND 0.0112f
C19026 VPWR.t1766 VGND 0.01226f
C19027 VPWR.n1090 VGND 0.02993f
C19028 VPWR.n1091 VGND 0.03284f
C19029 VPWR.n1092 VGND 0.01714f
C19030 VPWR.n1093 VGND 0.00697f
C19031 VPWR.n1094 VGND 0.01714f
C19032 VPWR.n1095 VGND 0.00697f
C19033 VPWR.t2049 VGND 0.01136f
C19034 VPWR.t1499 VGND 0.0124f
C19035 VPWR.n1096 VGND 0.02768f
C19036 VPWR.n1097 VGND 0.02818f
C19037 VPWR.n1098 VGND 0.01822f
C19038 VPWR.n1099 VGND 0.17585f
C19039 VPWR.t2059 VGND 0.0112f
C19040 VPWR.t1471 VGND 0.01226f
C19041 VPWR.n1100 VGND 0.02993f
C19042 VPWR.n1101 VGND 0.03284f
C19043 VPWR.n1102 VGND 0.01714f
C19044 VPWR.n1103 VGND 0.00697f
C19045 VPWR.n1104 VGND 0.01714f
C19046 VPWR.n1105 VGND 0.00697f
C19047 VPWR.t2014 VGND 0.01136f
C19048 VPWR.t1583 VGND 0.0124f
C19049 VPWR.n1106 VGND 0.02768f
C19050 VPWR.n1107 VGND 0.02818f
C19051 VPWR.n1108 VGND 0.01822f
C19052 VPWR.n1109 VGND 0.02654f
C19053 VPWR.t2018 VGND 0.0112f
C19054 VPWR.t1577 VGND 0.01226f
C19055 VPWR.n1110 VGND 0.02993f
C19056 VPWR.n1111 VGND 0.03284f
C19057 VPWR.n1112 VGND 0.01822f
C19058 VPWR.n1113 VGND 0.00697f
C19059 VPWR.t2012 VGND 0.01116f
C19060 VPWR.t1723 VGND 0.01222f
C19061 VPWR.n1114 VGND 0.03115f
C19062 VPWR.n1115 VGND 0.01969f
C19063 VPWR.t1969 VGND 0.01136f
C19064 VPWR.t1713 VGND 0.0124f
C19065 VPWR.n1116 VGND 0.02768f
C19066 VPWR.n1117 VGND 0.02818f
C19067 VPWR.n1118 VGND 0.01776f
C19068 VPWR.t2067 VGND 0.0112f
C19069 VPWR.t1441 VGND 0.01226f
C19070 VPWR.n1119 VGND 0.02993f
C19071 VPWR.n1120 VGND 0.03284f
C19072 VPWR.n1121 VGND 0.00805f
C19073 VPWR.t1725 VGND 0.03331f
C19074 VPWR.t1443 VGND 0.02961f
C19075 VPWR.n1122 VGND 0.09152f
C19076 VPWR.t1724 VGND 0.14512f
C19077 VPWR.t1714 VGND 0.07849f
C19078 VPWR.t1442 VGND 0.09218f
C19079 VPWR.t1597 VGND 0.11957f
C19080 VPWR.t1493 VGND 0.03331f
C19081 VPWR.t1579 VGND 0.02961f
C19082 VPWR.n1123 VGND 0.09152f
C19083 VPWR.n1124 VGND 0.00833f
C19084 VPWR.t2062 VGND 0.01116f
C19085 VPWR.t1596 VGND 0.01222f
C19086 VPWR.n1125 VGND 0.03115f
C19087 VPWR.n1126 VGND 0.03694f
C19088 VPWR.n1127 VGND 0.03437f
C19089 VPWR.n1128 VGND 0.13913f
C19090 VPWR.n1129 VGND 0.00805f
C19091 VPWR.n1130 VGND 0.01797f
C19092 VPWR.n1131 VGND 0.06567f
C19093 VPWR.n1132 VGND 0.0544f
C19094 VPWR.t1950 VGND 0.01136f
C19095 VPWR.t1764 VGND 0.0124f
C19096 VPWR.n1133 VGND 0.02769f
C19097 VPWR.n1134 VGND 0.01897f
C19098 VPWR.n1135 VGND 0.06244f
C19099 VPWR.n1136 VGND 0.09746f
C19100 VPWR.n1137 VGND 0.06567f
C19101 VPWR.n1138 VGND 0.06567f
C19102 VPWR.n1139 VGND 0.06567f
C19103 VPWR.n1140 VGND 0.06567f
C19104 VPWR.n1141 VGND 0.06567f
C19105 VPWR.n1142 VGND 0.06567f
C19106 VPWR.n1143 VGND 0.0544f
C19107 VPWR.n1144 VGND 0.00805f
C19108 VPWR.n1145 VGND -0.01866f
C19109 VPWR.t2020 VGND 0.01116f
C19110 VPWR.t1707 VGND 0.01222f
C19111 VPWR.n1146 VGND 0.03042f
C19112 VPWR.n1147 VGND 0.00581f
C19113 VPWR.t1709 VGND 0.02679f
C19114 VPWR.n1148 VGND 0.05724f
C19115 VPWR.t1915 VGND 0.02961f
C19116 VPWR.n1149 VGND 0.04692f
C19117 VPWR.t1914 VGND 0.09218f
C19118 VPWR.t1451 VGND 0.07849f
C19119 VPWR.t1581 VGND 0.11957f
C19120 VPWR.t1975 VGND 0.01116f
C19121 VPWR.t1447 VGND 0.01222f
C19122 VPWR.n1150 VGND 0.03042f
C19123 VPWR.n1151 VGND 0.00581f
C19124 VPWR.t1449 VGND 0.02679f
C19125 VPWR.n1152 VGND 0.05724f
C19126 VPWR.t1364 VGND 0.02961f
C19127 VPWR.n1153 VGND 0.04692f
C19128 VPWR.n1154 VGND 0.00805f
C19129 VPWR.n1155 VGND 0.00805f
C19130 VPWR.t1927 VGND 0.01116f
C19131 VPWR.t1691 VGND 0.01222f
C19132 VPWR.n1156 VGND 0.03042f
C19133 VPWR.n1157 VGND 0.00581f
C19134 VPWR.t1693 VGND 0.02679f
C19135 VPWR.n1158 VGND 0.05724f
C19136 VPWR.t824 VGND 0.02961f
C19137 VPWR.n1159 VGND 0.04692f
C19138 VPWR.t281 VGND 0.09218f
C19139 VPWR.t1938 VGND 0.01116f
C19140 VPWR.t1550 VGND 0.01222f
C19141 VPWR.n1160 VGND 0.03042f
C19142 VPWR.n1161 VGND 0.00581f
C19143 VPWR.t1552 VGND 0.02679f
C19144 VPWR.n1162 VGND 0.05724f
C19145 VPWR.t282 VGND 0.02961f
C19146 VPWR.n1163 VGND 0.04692f
C19147 VPWR.n1164 VGND 0.00805f
C19148 VPWR.n1165 VGND 0.00805f
C19149 VPWR.t2023 VGND 0.01116f
C19150 VPWR.t1428 VGND 0.01222f
C19151 VPWR.n1166 VGND 0.03042f
C19152 VPWR.n1167 VGND 0.00581f
C19153 VPWR.t1430 VGND 0.02679f
C19154 VPWR.n1168 VGND 0.05724f
C19155 VPWR.t418 VGND 0.02961f
C19156 VPWR.n1169 VGND 0.04692f
C19157 VPWR.t279 VGND 0.09218f
C19158 VPWR.t2035 VGND 0.01116f
C19159 VPWR.t1677 VGND 0.01222f
C19160 VPWR.n1170 VGND 0.03042f
C19161 VPWR.n1171 VGND 0.00581f
C19162 VPWR.t1679 VGND 0.02679f
C19163 VPWR.n1172 VGND 0.05724f
C19164 VPWR.t280 VGND 0.02961f
C19165 VPWR.n1173 VGND 0.04692f
C19166 VPWR.n1174 VGND 0.00805f
C19167 VPWR.n1175 VGND 0.00833f
C19168 VPWR.t1958 VGND 0.01116f
C19169 VPWR.t1488 VGND 0.01222f
C19170 VPWR.n1176 VGND 0.03115f
C19171 VPWR.n1177 VGND 0.03694f
C19172 VPWR.n1178 VGND 0.03437f
C19173 VPWR.t1478 VGND 0.03331f
C19174 VPWR.t1473 VGND 0.02961f
C19175 VPWR.n1179 VGND 0.09152f
C19176 VPWR.t1584 VGND 0.07849f
C19177 VPWR.t1591 VGND 0.09218f
C19178 VPWR.t1598 VGND 0.03331f
C19179 VPWR.t1592 VGND 0.02961f
C19180 VPWR.n1180 VGND 0.09152f
C19181 VPWR.n1181 VGND 0.00725f
C19182 VPWR.n1182 VGND 0.10822f
C19183 VPWR.t1759 VGND 0.11957f
C19184 VPWR.t1625 VGND 0.07849f
C19185 VPWR.t1751 VGND 0.09218f
C19186 VPWR.t1760 VGND 0.03331f
C19187 VPWR.t1752 VGND 0.02961f
C19188 VPWR.n1183 VGND 0.09152f
C19189 VPWR.n1184 VGND 0.00725f
C19190 VPWR.n1185 VGND 0.10822f
C19191 VPWR.t1477 VGND 0.11957f
C19192 VPWR.t1733 VGND 0.07849f
C19193 VPWR.t1472 VGND 0.09218f
C19194 VPWR.t1549 VGND 0.07849f
C19195 VPWR.t1675 VGND 0.11957f
C19196 VPWR.t1438 VGND 0.03331f
C19197 VPWR.t1539 VGND 0.02961f
C19198 VPWR.n1186 VGND 0.09152f
C19199 VPWR.n1187 VGND 0.00725f
C19200 VPWR.n1188 VGND 0.10822f
C19201 VPWR.t1538 VGND 0.09218f
C19202 VPWR.t1523 VGND 0.07849f
C19203 VPWR.t1437 VGND 0.11957f
C19204 VPWR.t1417 VGND 0.03331f
C19205 VPWR.t1795 VGND 0.02961f
C19206 VPWR.n1189 VGND 0.09152f
C19207 VPWR.n1190 VGND 0.00725f
C19208 VPWR.n1191 VGND 0.10822f
C19209 VPWR.t1794 VGND 0.09218f
C19210 VPWR.t1673 VGND 0.07849f
C19211 VPWR.t1416 VGND 0.11957f
C19212 VPWR.t1671 VGND 0.03331f
C19213 VPWR.t1776 VGND 0.02961f
C19214 VPWR.n1192 VGND 0.09152f
C19215 VPWR.n1193 VGND 0.00833f
C19216 VPWR.t2031 VGND 0.01116f
C19217 VPWR.t1415 VGND 0.01222f
C19218 VPWR.n1194 VGND 0.03115f
C19219 VPWR.n1195 VGND 0.03694f
C19220 VPWR.n1196 VGND 0.03437f
C19221 VPWR.n1197 VGND 0.01714f
C19222 VPWR.n1198 VGND 0.00725f
C19223 VPWR.n1199 VGND 0.10822f
C19224 VPWR.t1775 VGND 0.09218f
C19225 VPWR.t1651 VGND 0.07849f
C19226 VPWR.t1670 VGND 0.11957f
C19227 VPWR.t1544 VGND 0.03331f
C19228 VPWR.t1617 VGND 0.02961f
C19229 VPWR.n1200 VGND 0.09152f
C19230 VPWR.n1201 VGND 0.00725f
C19231 VPWR.n1202 VGND 0.10822f
C19232 VPWR.t1616 VGND 0.09218f
C19233 VPWR.t1498 VGND 0.07849f
C19234 VPWR.t1543 VGND 0.11957f
C19235 VPWR.t1518 VGND 0.03331f
C19236 VPWR.t1513 VGND 0.02961f
C19237 VPWR.n1203 VGND 0.09152f
C19238 VPWR.n1204 VGND 0.00725f
C19239 VPWR.n1205 VGND 0.10822f
C19240 VPWR.t1512 VGND 0.09218f
C19241 VPWR.t1781 VGND 0.07849f
C19242 VPWR.t1517 VGND 0.11957f
C19243 VPWR.t1757 VGND 0.03331f
C19244 VPWR.t1768 VGND 0.02961f
C19245 VPWR.n1206 VGND 0.09152f
C19246 VPWR.n1207 VGND 0.00833f
C19247 VPWR.t1992 VGND 0.01116f
C19248 VPWR.t1516 VGND 0.01222f
C19249 VPWR.n1208 VGND 0.03115f
C19250 VPWR.n1209 VGND 0.03694f
C19251 VPWR.n1210 VGND 0.03437f
C19252 VPWR.n1211 VGND 0.01714f
C19253 VPWR.n1212 VGND 0.00725f
C19254 VPWR.n1213 VGND 0.10822f
C19255 VPWR.t1767 VGND 0.09218f
C19256 VPWR.t1738 VGND 0.07849f
C19257 VPWR.t1756 VGND 0.11957f
C19258 VPWR.t1649 VGND 0.03331f
C19259 VPWR.t1728 VGND 0.02961f
C19260 VPWR.n1214 VGND 0.09152f
C19261 VPWR.n1215 VGND 0.00725f
C19262 VPWR.n1216 VGND 0.10822f
C19263 VPWR.t1727 VGND 0.09218f
C19264 VPWR.t1515 VGND 0.07849f
C19265 VPWR.t1648 VGND 0.11957f
C19266 VPWR.t1490 VGND 0.03331f
C19267 VPWR.t1620 VGND 0.02961f
C19268 VPWR.n1217 VGND 0.09152f
C19269 VPWR.n1218 VGND 0.00725f
C19270 VPWR.n1219 VGND 0.10822f
C19271 VPWR.t1619 VGND 0.09218f
C19272 VPWR.t1500 VGND 0.07849f
C19273 VPWR.t1489 VGND 0.11957f
C19274 VPWR.n1220 VGND 0.10822f
C19275 VPWR.n1221 VGND 0.00725f
C19276 VPWR.n1222 VGND 0.01714f
C19277 VPWR.n1223 VGND 0.00805f
C19278 VPWR.t2041 VGND 0.01116f
C19279 VPWR.t1655 VGND 0.01222f
C19280 VPWR.n1224 VGND 0.03042f
C19281 VPWR.n1225 VGND 0.00581f
C19282 VPWR.t1657 VGND 0.02679f
C19283 VPWR.n1226 VGND 0.05724f
C19284 VPWR.t416 VGND 0.02961f
C19285 VPWR.n1227 VGND 0.04692f
C19286 VPWR.t1520 VGND 0.14512f
C19287 VPWR.t1505 VGND 0.07849f
C19288 VPWR.t454 VGND 0.09218f
C19289 VPWR.t1948 VGND 0.01116f
C19290 VPWR.t1519 VGND 0.01222f
C19291 VPWR.n1228 VGND 0.03042f
C19292 VPWR.n1229 VGND 0.00581f
C19293 VPWR.t1521 VGND 0.02679f
C19294 VPWR.n1230 VGND 0.05724f
C19295 VPWR.t455 VGND 0.02961f
C19296 VPWR.n1231 VGND 0.04692f
C19297 VPWR.n1232 VGND -0.01866f
C19298 VPWR.n1233 VGND 0.04687f
C19299 VPWR.t38 VGND 0.97566f
C19300 VPWR.n1234 VGND 0.53213f
C19301 VPWR.t43 VGND 0.97566f
C19302 VPWR.n1235 VGND 0.41384f
C19303 VPWR.n1236 VGND 0.2908f
C19304 VPWR.t560 VGND 0.05716f
C19305 VPWR.n1237 VGND 0.0092f
C19306 VPWR.t702 VGND 0.01433f
C19307 VPWR.t646 VGND 0.01433f
C19308 VPWR.n1238 VGND 0.03146f
C19309 VPWR.t647 VGND 0.01433f
C19310 VPWR.t951 VGND 0.01433f
C19311 VPWR.n1239 VGND 0.03141f
C19312 VPWR.t401 VGND 0.01433f
C19313 VPWR.t400 VGND 0.01433f
C19314 VPWR.n1240 VGND 0.03141f
C19315 VPWR.n1241 VGND 0.1042f
C19316 VPWR.n1242 VGND 0.18182f
C19317 VPWR.n1243 VGND 0.05756f
C19318 VPWR.n1244 VGND 0.04228f
C19319 VPWR.t396 VGND 0.01433f
C19320 VPWR.t402 VGND 0.01433f
C19321 VPWR.n1245 VGND 0.03146f
C19322 VPWR.n1246 VGND 0.12902f
C19323 VPWR.n1247 VGND 0.01119f
C19324 VPWR.n1248 VGND 0.0163f
C19325 VPWR.n1249 VGND 0.0191f
C19326 VPWR.n1250 VGND 0.02802f
C19327 VPWR.t559 VGND 0.05716f
C19328 VPWR.n1251 VGND 0.15059f
C19329 VPWR.n1252 VGND 0.01209f
C19330 VPWR.t1154 VGND 0.05714f
C19331 VPWR.t715 VGND 0.05714f
C19332 VPWR.n1253 VGND 0.13446f
C19333 VPWR.n1254 VGND 0.33563f
C19334 VPWR.n1255 VGND 1.64092f
C19335 VPWR.n1256 VGND 0.04687f
C19336 VPWR.t42 VGND 0.97566f
C19337 VPWR.n1257 VGND 0.53213f
C19338 VPWR.t561 VGND 0.97566f
C19339 VPWR.n1258 VGND 0.41384f
C19340 VPWR.n1259 VGND 0.29342f
C19341 VPWR.n1260 VGND 0.0092f
C19342 VPWR.t1269 VGND 0.01433f
C19343 VPWR.t1267 VGND 0.01433f
C19344 VPWR.n1261 VGND 0.03146f
C19345 VPWR.t1266 VGND 0.01433f
C19346 VPWR.t1264 VGND 0.01433f
C19347 VPWR.n1262 VGND 0.03141f
C19348 VPWR.t1340 VGND 0.01433f
C19349 VPWR.t1341 VGND 0.01433f
C19350 VPWR.n1263 VGND 0.03141f
C19351 VPWR.n1264 VGND 0.1042f
C19352 VPWR.n1265 VGND 0.18182f
C19353 VPWR.n1266 VGND 0.05756f
C19354 VPWR.n1267 VGND 0.04228f
C19355 VPWR.t933 VGND 0.01433f
C19356 VPWR.t1402 VGND 0.01433f
C19357 VPWR.n1268 VGND 0.03146f
C19358 VPWR.n1269 VGND 0.12902f
C19359 VPWR.n1270 VGND 0.01119f
C19360 VPWR.n1271 VGND 0.0163f
C19361 VPWR.n1272 VGND 0.0191f
C19362 VPWR.n1273 VGND 0.02751f
C19363 VPWR.n1274 VGND 0.00767f
C19364 VPWR.t562 VGND 0.05708f
C19365 VPWR.n1275 VGND 0.06101f
C19366 VPWR.n1276 VGND 0.00731f
C19367 VPWR.t462 VGND 0.0572f
C19368 VPWR.n1277 VGND 0.0911f
C19369 VPWR.n1278 VGND 0.33563f
C19370 VPWR.n1279 VGND 1.64092f
C19371 VPWR.n1280 VGND 0.04687f
C19372 VPWR.t37 VGND 0.97566f
C19373 VPWR.n1281 VGND 0.53213f
C19374 VPWR.t387 VGND 0.97566f
C19375 VPWR.n1282 VGND 0.41384f
C19376 VPWR.n1283 VGND 0.29342f
C19377 VPWR.n1284 VGND 0.0092f
C19378 VPWR.t658 VGND 0.01433f
C19379 VPWR.t656 VGND 0.01433f
C19380 VPWR.n1285 VGND 0.03146f
C19381 VPWR.t655 VGND 0.01433f
C19382 VPWR.t654 VGND 0.01433f
C19383 VPWR.n1286 VGND 0.03141f
C19384 VPWR.t388 VGND 0.01433f
C19385 VPWR.t395 VGND 0.01433f
C19386 VPWR.n1287 VGND 0.03141f
C19387 VPWR.n1288 VGND 0.1042f
C19388 VPWR.n1289 VGND 0.18182f
C19389 VPWR.n1290 VGND 0.05756f
C19390 VPWR.n1291 VGND 0.04228f
C19391 VPWR.t392 VGND 0.01433f
C19392 VPWR.t389 VGND 0.01433f
C19393 VPWR.n1292 VGND 0.03146f
C19394 VPWR.n1293 VGND 0.12902f
C19395 VPWR.n1294 VGND 0.01119f
C19396 VPWR.n1295 VGND 0.0163f
C19397 VPWR.n1296 VGND 0.0191f
C19398 VPWR.n1297 VGND 0.02751f
C19399 VPWR.n1298 VGND 0.01398f
C19400 VPWR.n1299 VGND 0.01308f
C19401 VPWR.t1155 VGND 0.0572f
C19402 VPWR.t716 VGND 0.0572f
C19403 VPWR.n1300 VGND 0.16894f
C19404 VPWR.n1301 VGND 0.33563f
C19405 VPWR.n1302 VGND 1.64092f
C19406 VPWR.t1251 VGND 0.05711f
C19407 VPWR.t650 VGND 0.0572f
C19408 VPWR.t1253 VGND 0.05672f
C19409 VPWR.n1303 VGND 0.14706f
C19410 VPWR.t36 VGND 0.05606f
C19411 VPWR.n1304 VGND 0.06775f
C19412 VPWR.n1305 VGND 0.04687f
C19413 VPWR.t440 VGND 0.05397f
C19414 VPWR.n1306 VGND 0.05133f
C19415 VPWR.t1294 VGND 0.01433f
C19416 VPWR.t1308 VGND 0.01433f
C19417 VPWR.n1307 VGND 0.03131f
C19418 VPWR.t1242 VGND 0.05015f
C19419 VPWR.n1308 VGND 0.07521f
C19420 VPWR.n1309 VGND 0.04687f
C19421 VPWR.t836 VGND 0.05714f
C19422 VPWR.n1310 VGND 0.07193f
C19423 VPWR.n1311 VGND 0.02751f
C19424 VPWR.n1312 VGND 0.04687f
C19425 VPWR.n1313 VGND 0.01209f
C19426 VPWR.t1310 VGND 0.01433f
C19427 VPWR.t1312 VGND 0.01433f
C19428 VPWR.n1314 VGND 0.03131f
C19429 VPWR.n1315 VGND 0.04588f
C19430 VPWR.n1316 VGND 0.01209f
C19431 VPWR.n1317 VGND 0.03515f
C19432 VPWR.n1318 VGND 0.03515f
C19433 VPWR.n1319 VGND 0.04687f
C19434 VPWR.n1320 VGND 0.0083f
C19435 VPWR.t787 VGND 0.01433f
C19436 VPWR.t1298 VGND 0.01433f
C19437 VPWR.n1321 VGND 0.03131f
C19438 VPWR.n1322 VGND 0.03605f
C19439 VPWR.t40 VGND 0.01433f
C19440 VPWR.t1799 VGND 0.01433f
C19441 VPWR.n1323 VGND 0.03131f
C19442 VPWR.n1324 VGND 0.03983f
C19443 VPWR.n1325 VGND 0.01055f
C19444 VPWR.n1326 VGND 0.04254f
C19445 VPWR.n1327 VGND 0.01605f
C19446 VPWR.n1328 VGND 0.00631f
C19447 VPWR.t998 VGND 0.04806f
C19448 VPWR.t1250 VGND 0.10812f
C19449 VPWR.t649 VGND 0.12614f
C19450 VPWR.t1252 VGND 0.23427f
C19451 VPWR.t835 VGND 0.12605f
C19452 VPWR.t1311 VGND 0.14308f
C19453 VPWR.t1309 VGND 0.1391f
C19454 VPWR.t1307 VGND 0.22247f
C19455 VPWR.t1293 VGND 0.18922f
C19456 VPWR.t1241 VGND 0.12614f
C19457 VPWR.t1297 VGND 0.12614f
C19458 VPWR.t1798 VGND 0.12614f
C19459 VPWR.t786 VGND 0.12614f
C19460 VPWR.t39 VGND 0.12614f
C19461 VPWR.t439 VGND 0.12614f
C19462 VPWR.t35 VGND 0.12464f
C19463 VPWR.n1329 VGND 0.4287f
C19464 VPWR.n1330 VGND 0.17419f
C19465 VPWR.n1331 VGND 0.0191f
C19466 VPWR.n1332 VGND 0.03515f
C19467 VPWR.n1333 VGND 0.04228f
C19468 VPWR.n1334 VGND 0.01083f
C19469 VPWR.n1335 VGND 0.06357f
C19470 VPWR.n1336 VGND 0.31652f
C19471 VPWR.n1337 VGND 1.64092f
C19472 VPWR.t1909 VGND 0.05619f
C19473 VPWR.t714 VGND 0.05603f
C19474 VPWR.t717 VGND 0.05714f
C19475 VPWR.n1338 VGND 0.07963f
C19476 VPWR.t648 VGND 0.05456f
C19477 VPWR.t403 VGND 0.05456f
C19478 VPWR.n1339 VGND 0.09898f
C19479 VPWR.n1340 VGND 0.04687f
C19480 VPWR.n1341 VGND 0.00911f
C19481 VPWR.n1342 VGND 0.04687f
C19482 VPWR.t703 VGND 0.01433f
C19483 VPWR.t78 VGND 0.01433f
C19484 VPWR.n1343 VGND 0.03131f
C19485 VPWR.t404 VGND 0.01433f
C19486 VPWR.t845 VGND 0.01433f
C19487 VPWR.n1344 VGND 0.03131f
C19488 VPWR.n1345 VGND 0.06379f
C19489 VPWR.t847 VGND 0.05714f
C19490 VPWR.t1313 VGND 0.05714f
C19491 VPWR.n1346 VGND 0.13169f
C19492 VPWR.n1347 VGND 0.02751f
C19493 VPWR.n1348 VGND 0.04687f
C19494 VPWR.n1349 VGND 0.01209f
C19495 VPWR.t110 VGND 0.01433f
C19496 VPWR.t832 VGND 0.01433f
C19497 VPWR.n1350 VGND 0.03131f
C19498 VPWR.t850 VGND 0.01433f
C19499 VPWR.t1796 VGND 0.01433f
C19500 VPWR.n1351 VGND 0.03131f
C19501 VPWR.n1352 VGND 0.07209f
C19502 VPWR.n1353 VGND 0.01209f
C19503 VPWR.n1354 VGND 0.04687f
C19504 VPWR.n1355 VGND 0.04687f
C19505 VPWR.n1356 VGND 0.04687f
C19506 VPWR.n1357 VGND 0.01128f
C19507 VPWR.t952 VGND 0.01433f
C19508 VPWR.t645 VGND 0.01433f
C19509 VPWR.n1358 VGND 0.03131f
C19510 VPWR.t399 VGND 0.01433f
C19511 VPWR.t398 VGND 0.01433f
C19512 VPWR.n1359 VGND 0.03131f
C19513 VPWR.n1360 VGND 0.06379f
C19514 VPWR.n1361 VGND 0.01055f
C19515 VPWR.n1362 VGND 0.00983f
C19516 VPWR.n1363 VGND 0.04687f
C19517 VPWR.n1364 VGND 0.03515f
C19518 VPWR.n1365 VGND 0.00794f
C19519 VPWR.t77 VGND 0.97566f
C19520 VPWR.n1366 VGND 0.53213f
C19521 VPWR.t397 VGND 0.97566f
C19522 VPWR.n1367 VGND 0.41384f
C19523 VPWR.n1368 VGND 0.2908f
C19524 VPWR.n1369 VGND 0.0191f
C19525 VPWR.n1370 VGND 0.03515f
C19526 VPWR.n1371 VGND 0.04254f
C19527 VPWR.n1372 VGND 0.01064f
C19528 VPWR.n1373 VGND 0.05827f
C19529 VPWR.n1374 VGND 0.07893f
C19530 VPWR.n1375 VGND 0.31627f
C19531 VPWR.n1376 VGND 1.64092f
C19532 VPWR.t367 VGND 0.05708f
C19533 VPWR.t1284 VGND 0.05708f
C19534 VPWR.n1377 VGND 0.01398f
C19535 VPWR.t1265 VGND 0.05456f
C19536 VPWR.t934 VGND 0.05456f
C19537 VPWR.n1378 VGND 0.09898f
C19538 VPWR.n1379 VGND 0.04687f
C19539 VPWR.n1380 VGND 0.00911f
C19540 VPWR.n1381 VGND 0.04687f
C19541 VPWR.t1270 VGND 0.01433f
C19542 VPWR.t848 VGND 0.01433f
C19543 VPWR.n1382 VGND 0.03131f
C19544 VPWR.t288 VGND 0.01433f
C19545 VPWR.t73 VGND 0.01433f
C19546 VPWR.n1383 VGND 0.03131f
C19547 VPWR.n1384 VGND 0.06379f
C19548 VPWR.t75 VGND 0.05714f
C19549 VPWR.t45 VGND 0.05714f
C19550 VPWR.n1385 VGND 0.13169f
C19551 VPWR.n1386 VGND 0.02751f
C19552 VPWR.n1387 VGND 0.04687f
C19553 VPWR.n1388 VGND 0.01209f
C19554 VPWR.t852 VGND 0.01433f
C19555 VPWR.t1797 VGND 0.01433f
C19556 VPWR.n1389 VGND 0.03131f
C19557 VPWR.t76 VGND 0.01433f
C19558 VPWR.t112 VGND 0.01433f
C19559 VPWR.n1390 VGND 0.03131f
C19560 VPWR.n1391 VGND 0.07209f
C19561 VPWR.n1392 VGND 0.01209f
C19562 VPWR.n1393 VGND 0.04687f
C19563 VPWR.n1394 VGND 0.04687f
C19564 VPWR.n1395 VGND 0.04687f
C19565 VPWR.n1396 VGND 0.01128f
C19566 VPWR.t1271 VGND 0.01433f
C19567 VPWR.t1268 VGND 0.01433f
C19568 VPWR.n1397 VGND 0.03131f
C19569 VPWR.t287 VGND 0.01433f
C19570 VPWR.t932 VGND 0.01433f
C19571 VPWR.n1398 VGND 0.03131f
C19572 VPWR.n1399 VGND 0.06379f
C19573 VPWR.n1400 VGND 0.01055f
C19574 VPWR.n1401 VGND 0.00983f
C19575 VPWR.n1402 VGND 0.04687f
C19576 VPWR.n1403 VGND 0.03515f
C19577 VPWR.n1404 VGND 0.00794f
C19578 VPWR.t74 VGND 0.97566f
C19579 VPWR.n1405 VGND 0.53213f
C19580 VPWR.t44 VGND 0.97566f
C19581 VPWR.n1406 VGND 0.41384f
C19582 VPWR.n1407 VGND 0.29342f
C19583 VPWR.n1408 VGND 0.0191f
C19584 VPWR.n1409 VGND 0.03515f
C19585 VPWR.n1410 VGND 0.04254f
C19586 VPWR.n1411 VGND 0.01083f
C19587 VPWR.n1412 VGND 0.11537f
C19588 VPWR.n1413 VGND 0.32137f
C19589 VPWR.n1414 VGND 1.64092f
C19590 VPWR.t657 VGND 0.05456f
C19591 VPWR.t390 VGND 0.05456f
C19592 VPWR.n1415 VGND 0.09898f
C19593 VPWR.n1416 VGND 0.04687f
C19594 VPWR.n1417 VGND 0.00911f
C19595 VPWR.n1418 VGND 0.04687f
C19596 VPWR.t652 VGND 0.01433f
C19597 VPWR.t80 VGND 0.01433f
C19598 VPWR.n1419 VGND 0.03131f
C19599 VPWR.t391 VGND 0.01433f
C19600 VPWR.t834 VGND 0.01433f
C19601 VPWR.n1420 VGND 0.03131f
C19602 VPWR.n1421 VGND 0.06379f
C19603 VPWR.t849 VGND 0.05714f
C19604 VPWR.t601 VGND 0.05714f
C19605 VPWR.n1422 VGND 0.13169f
C19606 VPWR.n1423 VGND 0.02751f
C19607 VPWR.n1424 VGND 0.04687f
C19608 VPWR.n1425 VGND 0.01209f
C19609 VPWR.t111 VGND 0.01433f
C19610 VPWR.t833 VGND 0.01433f
C19611 VPWR.n1426 VGND 0.03131f
C19612 VPWR.t34 VGND 0.01433f
C19613 VPWR.t41 VGND 0.01433f
C19614 VPWR.n1427 VGND 0.03131f
C19615 VPWR.n1428 VGND 0.07209f
C19616 VPWR.n1429 VGND 0.01209f
C19617 VPWR.n1430 VGND 0.04687f
C19618 VPWR.n1431 VGND 0.04687f
C19619 VPWR.n1432 VGND 0.04687f
C19620 VPWR.n1433 VGND 0.01128f
C19621 VPWR.t653 VGND 0.01433f
C19622 VPWR.t651 VGND 0.01433f
C19623 VPWR.n1434 VGND 0.03131f
C19624 VPWR.t394 VGND 0.01433f
C19625 VPWR.t393 VGND 0.01433f
C19626 VPWR.n1435 VGND 0.03131f
C19627 VPWR.n1436 VGND 0.06379f
C19628 VPWR.n1437 VGND 0.01055f
C19629 VPWR.n1438 VGND 0.00983f
C19630 VPWR.n1439 VGND 0.04687f
C19631 VPWR.n1440 VGND 0.03515f
C19632 VPWR.n1441 VGND 0.00794f
C19633 VPWR.t79 VGND 0.74843f
C19634 VPWR.n1442 VGND 0.4282f
C19635 VPWR.t33 VGND 0.74843f
C19636 VPWR.n1443 VGND 0.33553f
C19637 VPWR.n1444 VGND 0.28129f
C19638 VPWR.n1445 VGND 0.43003f
C19639 VPWR.n1446 VGND 6.17638f
C19640 VPWR.n1447 VGND 9.5664f
C19641 VPWR.n1448 VGND 0.08351f
C19642 VPWR.n1449 VGND 1.09982f
C19643 VPWR.n1450 VGND 1.0094f
C19644 VPWR.n1451 VGND 0.06482f
C19645 VPWR.n1452 VGND 0.0544f
C19646 VPWR.t2045 VGND 0.01136f
C19647 VPWR.t1504 VGND 0.0124f
C19648 VPWR.n1453 VGND 0.02769f
C19649 VPWR.n1454 VGND 0.01897f
C19650 VPWR.n1455 VGND 0.06244f
C19651 VPWR.n1456 VGND 0.07762f
C19652 VPWR.n1457 VGND 0.09174f
C19653 VPWR.t1996 VGND 0.01136f
C19654 VPWR.t1635 VGND 0.0124f
C19655 VPWR.n1458 VGND 0.02769f
C19656 VPWR.n1459 VGND 0.01897f
C19657 VPWR.n1460 VGND 0.06244f
C19658 VPWR.n1461 VGND 0.09746f
C19659 VPWR.n1462 VGND 0.09174f
C19660 VPWR.n1463 VGND 0.06567f
C19661 VPWR.n1464 VGND 0.0544f
C19662 VPWR.n1465 VGND 0.13913f
C19663 VPWR.n1466 VGND 0.01797f
C19664 VPWR.n1467 VGND 0.00728f
C19665 VPWR.n1468 VGND 0.10822f
C19666 VPWR.t1681 VGND 0.11957f
C19667 VPWR.t1636 VGND 0.07849f
C19668 VPWR.t59 VGND 0.09218f
C19669 VPWR.t2044 VGND 0.01116f
C19670 VPWR.t1680 VGND 0.01222f
C19671 VPWR.n1469 VGND 0.03042f
C19672 VPWR.n1470 VGND 0.00581f
C19673 VPWR.t1682 VGND 0.02679f
C19674 VPWR.n1471 VGND 0.05724f
C19675 VPWR.t60 VGND 0.02961f
C19676 VPWR.n1472 VGND 0.04692f
C19677 VPWR.n1473 VGND 0.01797f
C19678 VPWR.n1474 VGND 0.00728f
C19679 VPWR.n1475 VGND 0.10822f
C19680 VPWR.t1783 VGND 0.11957f
C19681 VPWR.t1765 VGND 0.07849f
C19682 VPWR.t776 VGND 0.09218f
C19683 VPWR.t1994 VGND 0.01116f
C19684 VPWR.t1782 VGND 0.01222f
C19685 VPWR.n1476 VGND 0.03042f
C19686 VPWR.n1477 VGND 0.00581f
C19687 VPWR.t1784 VGND 0.02679f
C19688 VPWR.n1478 VGND 0.05724f
C19689 VPWR.t777 VGND 0.02961f
C19690 VPWR.n1479 VGND 0.04692f
C19691 VPWR.n1480 VGND 0.00728f
C19692 VPWR.n1481 VGND 0.10822f
C19693 VPWR.t1554 VGND 0.11957f
C19694 VPWR.t1421 VGND 0.07849f
C19695 VPWR.t1057 VGND 0.09218f
C19696 VPWR.t1982 VGND 0.01116f
C19697 VPWR.t1553 VGND 0.01222f
C19698 VPWR.n1482 VGND 0.03042f
C19699 VPWR.n1483 VGND 0.00581f
C19700 VPWR.t1555 VGND 0.02679f
C19701 VPWR.n1484 VGND 0.05724f
C19702 VPWR.t1058 VGND 0.02961f
C19703 VPWR.n1485 VGND 0.04692f
C19704 VPWR.n1486 VGND 0.00805f
C19705 VPWR.n1487 VGND 0.08351f
C19706 VPWR.n1488 VGND -0.01866f
C19707 VPWR.n1489 VGND 0.13913f
C19708 VPWR.n1490 VGND 0.01797f
C19709 VPWR.n1491 VGND 0.00728f
C19710 VPWR.n1492 VGND 0.10822f
C19711 VPWR.t1656 VGND 0.11957f
C19712 VPWR.t1531 VGND 0.07849f
C19713 VPWR.t415 VGND 0.09218f
C19714 VPWR.t1686 VGND 0.07849f
C19715 VPWR.t1678 VGND 0.11957f
C19716 VPWR.n1493 VGND 0.10822f
C19717 VPWR.n1494 VGND 0.00728f
C19718 VPWR.n1495 VGND 0.01797f
C19719 VPWR.n1496 VGND 0.0544f
C19720 VPWR.n1497 VGND 0.13913f
C19721 VPWR.n1498 VGND -0.01866f
C19722 VPWR.n1499 VGND 0.08351f
C19723 VPWR.n1500 VGND 0.08351f
C19724 VPWR.n1501 VGND -0.01866f
C19725 VPWR.n1502 VGND 0.0544f
C19726 VPWR.n1503 VGND 0.13913f
C19727 VPWR.n1504 VGND 0.01797f
C19728 VPWR.n1505 VGND 0.00728f
C19729 VPWR.n1506 VGND 0.10822f
C19730 VPWR.t1429 VGND 0.11957f
C19731 VPWR.t1688 VGND 0.07849f
C19732 VPWR.t417 VGND 0.09218f
C19733 VPWR.t1536 VGND 0.07849f
C19734 VPWR.t1551 VGND 0.11957f
C19735 VPWR.n1507 VGND 0.10822f
C19736 VPWR.n1508 VGND 0.00728f
C19737 VPWR.n1509 VGND 0.01797f
C19738 VPWR.n1510 VGND 0.0544f
C19739 VPWR.n1511 VGND 0.13913f
C19740 VPWR.n1512 VGND -0.01866f
C19741 VPWR.n1513 VGND 0.08351f
C19742 VPWR.n1514 VGND 0.08351f
C19743 VPWR.n1515 VGND -0.01866f
C19744 VPWR.n1516 VGND 0.0544f
C19745 VPWR.n1517 VGND 0.13913f
C19746 VPWR.n1518 VGND 0.01797f
C19747 VPWR.n1519 VGND 0.00728f
C19748 VPWR.n1520 VGND 0.10822f
C19749 VPWR.t1692 VGND 0.11957f
C19750 VPWR.t1566 VGND 0.07849f
C19751 VPWR.t823 VGND 0.09218f
C19752 VPWR.t1684 VGND 0.07849f
C19753 VPWR.t1708 VGND 0.11957f
C19754 VPWR.n1521 VGND 0.10822f
C19755 VPWR.n1522 VGND 0.00728f
C19756 VPWR.n1523 VGND 0.01797f
C19757 VPWR.n1524 VGND 0.0544f
C19758 VPWR.n1525 VGND 0.13913f
C19759 VPWR.n1526 VGND -0.01866f
C19760 VPWR.n1527 VGND 0.08351f
C19761 VPWR.n1528 VGND 0.08351f
C19762 VPWR.n1529 VGND 0.08351f
C19763 VPWR.n1530 VGND 0.08351f
C19764 VPWR.n1531 VGND -0.01866f
C19765 VPWR.n1532 VGND 0.13913f
C19766 VPWR.n1533 VGND 0.01797f
C19767 VPWR.n1534 VGND 0.00728f
C19768 VPWR.n1535 VGND 0.10822f
C19769 VPWR.t1363 VGND 0.09218f
C19770 VPWR.t1435 VGND 0.07849f
C19771 VPWR.t1448 VGND 0.11957f
C19772 VPWR.n1536 VGND 0.10822f
C19773 VPWR.n1537 VGND 0.00728f
C19774 VPWR.n1538 VGND 0.01797f
C19775 VPWR.n1539 VGND 0.13913f
C19776 VPWR.n1540 VGND 0.0544f
C19777 VPWR.n1541 VGND 0.06567f
C19778 VPWR.n1542 VGND 0.09174f
C19779 VPWR.t1929 VGND 0.01136f
C19780 VPWR.t1434 VGND 0.0124f
C19781 VPWR.n1543 VGND 0.02769f
C19782 VPWR.n1544 VGND 0.01897f
C19783 VPWR.n1545 VGND 0.06244f
C19784 VPWR.n1546 VGND 0.09746f
C19785 VPWR.n1547 VGND 0.09174f
C19786 VPWR.t1986 VGND 0.01136f
C19787 VPWR.t1683 VGND 0.0124f
C19788 VPWR.n1548 VGND 0.02769f
C19789 VPWR.n1549 VGND 0.01897f
C19790 VPWR.n1550 VGND 0.06244f
C19791 VPWR.n1551 VGND 0.09746f
C19792 VPWR.n1552 VGND 0.09174f
C19793 VPWR.t2025 VGND 0.01136f
C19794 VPWR.t1565 VGND 0.0124f
C19795 VPWR.n1553 VGND 0.02769f
C19796 VPWR.n1554 VGND 0.01897f
C19797 VPWR.n1555 VGND 0.06244f
C19798 VPWR.n1556 VGND 0.09746f
C19799 VPWR.n1557 VGND 0.09174f
C19800 VPWR.t2037 VGND 0.01136f
C19801 VPWR.t1535 VGND 0.0124f
C19802 VPWR.n1558 VGND 0.02769f
C19803 VPWR.n1559 VGND 0.01897f
C19804 VPWR.n1560 VGND 0.06244f
C19805 VPWR.n1561 VGND 0.09746f
C19806 VPWR.n1562 VGND 0.09174f
C19807 VPWR.t1979 VGND 0.01136f
C19808 VPWR.t1687 VGND 0.0124f
C19809 VPWR.n1563 VGND 0.02769f
C19810 VPWR.n1564 VGND 0.01897f
C19811 VPWR.n1565 VGND 0.06244f
C19812 VPWR.n1566 VGND 0.09746f
C19813 VPWR.n1567 VGND 0.09174f
C19814 VPWR.t1985 VGND 0.01136f
C19815 VPWR.t1685 VGND 0.0124f
C19816 VPWR.n1568 VGND 0.02769f
C19817 VPWR.n1569 VGND 0.01897f
C19818 VPWR.n1570 VGND 0.06244f
C19819 VPWR.n1571 VGND 0.09746f
C19820 VPWR.n1572 VGND 0.09174f
C19821 VPWR.t2039 VGND 0.01136f
C19822 VPWR.t1530 VGND 0.0124f
C19823 VPWR.n1573 VGND 0.02769f
C19824 VPWR.n1574 VGND 0.01897f
C19825 VPWR.n1575 VGND 0.06244f
C19826 VPWR.n1576 VGND 0.09746f
C19827 VPWR.n1577 VGND 0.09174f
C19828 VPWR.t1936 VGND 0.01136f
C19829 VPWR.t1420 VGND 0.0124f
C19830 VPWR.n1578 VGND 0.02769f
C19831 VPWR.n1579 VGND 0.01897f
C19832 VPWR.n1580 VGND 0.06244f
C19833 VPWR.n1581 VGND 0.09746f
C19834 VPWR.n1582 VGND 0.09174f
C19835 VPWR.n1583 VGND 0.06567f
C19836 VPWR.n1584 VGND 0.0544f
C19837 VPWR.n1585 VGND 0.13913f
C19838 VPWR.n1586 VGND -0.01866f
C19839 VPWR.n1587 VGND 0.08351f
C19840 VPWR.n1588 VGND 0.08351f
C19841 VPWR.n1589 VGND -0.01866f
C19842 VPWR.n1590 VGND 0.00805f
C19843 VPWR.n1591 VGND 0.01714f
C19844 VPWR.n1592 VGND 0.00725f
C19845 VPWR.n1593 VGND 0.10822f
C19846 VPWR.t1578 VGND 0.09218f
C19847 VPWR.t1456 VGND 0.07849f
C19848 VPWR.t1492 VGND 0.11957f
C19849 VPWR.n1594 VGND 0.10822f
C19850 VPWR.n1595 VGND 0.00725f
C19851 VPWR.n1596 VGND 0.01714f
C19852 VPWR.n1597 VGND 0.03437f
C19853 VPWR.t1966 VGND 0.01116f
C19854 VPWR.t1491 VGND 0.01222f
C19855 VPWR.n1598 VGND 0.03115f
C19856 VPWR.n1599 VGND 0.03694f
C19857 VPWR.n1600 VGND 0.00833f
C19858 VPWR.t2063 VGND 0.01136f
C19859 VPWR.t1455 VGND 0.0124f
C19860 VPWR.n1601 VGND 0.02768f
C19861 VPWR.n1602 VGND 0.02818f
C19862 VPWR.n1603 VGND 0.01776f
C19863 VPWR.n1604 VGND 0.00697f
C19864 VPWR.n1605 VGND 0.01822f
C19865 VPWR.n1606 VGND 0.02384f
C19866 VPWR.n1607 VGND 0.23724f
C19867 VPWR.n1608 VGND 0.17585f
C19868 VPWR.n1609 VGND 0.02384f
C19869 VPWR.n1610 VGND 0.01776f
C19870 VPWR.t2010 VGND 0.0112f
C19871 VPWR.t1590 VGND 0.01226f
C19872 VPWR.n1611 VGND 0.02993f
C19873 VPWR.n1612 VGND 0.03284f
C19874 VPWR.n1613 VGND 0.03437f
C19875 VPWR.t2047 VGND 0.01116f
C19876 VPWR.t1758 VGND 0.01222f
C19877 VPWR.n1614 VGND 0.03115f
C19878 VPWR.n1615 VGND 0.03694f
C19879 VPWR.n1616 VGND 0.00833f
C19880 VPWR.t2000 VGND 0.01136f
C19881 VPWR.t1624 VGND 0.0124f
C19882 VPWR.n1617 VGND 0.02768f
C19883 VPWR.n1618 VGND 0.02818f
C19884 VPWR.n1619 VGND 0.01822f
C19885 VPWR.n1620 VGND 0.02384f
C19886 VPWR.n1621 VGND 0.01776f
C19887 VPWR.t1955 VGND 0.0112f
C19888 VPWR.t1750 VGND 0.01226f
C19889 VPWR.n1622 VGND 0.02993f
C19890 VPWR.n1623 VGND 0.03284f
C19891 VPWR.n1624 VGND 0.03437f
C19892 VPWR.t1965 VGND 0.01116f
C19893 VPWR.t1476 VGND 0.01222f
C19894 VPWR.n1625 VGND 0.03115f
C19895 VPWR.n1626 VGND 0.03694f
C19896 VPWR.n1627 VGND 0.00833f
C19897 VPWR.t1962 VGND 0.01136f
C19898 VPWR.t1732 VGND 0.0124f
C19899 VPWR.n1628 VGND 0.02768f
C19900 VPWR.n1629 VGND 0.02818f
C19901 VPWR.n1630 VGND 0.01776f
C19902 VPWR.n1631 VGND 0.00697f
C19903 VPWR.n1632 VGND 0.01822f
C19904 VPWR.n1633 VGND 0.02384f
C19905 VPWR.n1634 VGND 0.17585f
C19906 VPWR.n1635 VGND 0.17585f
C19907 VPWR.n1636 VGND 0.02384f
C19908 VPWR.n1637 VGND 0.01776f
C19909 VPWR.t2002 VGND 0.0112f
C19910 VPWR.t1618 VGND 0.01226f
C19911 VPWR.n1638 VGND 0.02993f
C19912 VPWR.n1639 VGND 0.03284f
C19913 VPWR.n1640 VGND 0.03437f
C19914 VPWR.t1944 VGND 0.01116f
C19915 VPWR.t1647 VGND 0.01222f
C19916 VPWR.n1641 VGND 0.03115f
C19917 VPWR.n1642 VGND 0.03694f
C19918 VPWR.n1643 VGND 0.00833f
C19919 VPWR.t2042 VGND 0.01136f
C19920 VPWR.t1514 VGND 0.0124f
C19921 VPWR.n1644 VGND 0.02768f
C19922 VPWR.n1645 VGND 0.02818f
C19923 VPWR.n1646 VGND 0.01822f
C19924 VPWR.n1647 VGND 0.02384f
C19925 VPWR.n1648 VGND 0.01776f
C19926 VPWR.t1964 VGND 0.0112f
C19927 VPWR.t1726 VGND 0.01226f
C19928 VPWR.n1649 VGND 0.02993f
C19929 VPWR.n1650 VGND 0.03284f
C19930 VPWR.n1651 VGND 0.03437f
C19931 VPWR.t2005 VGND 0.01116f
C19932 VPWR.t1755 VGND 0.01222f
C19933 VPWR.n1652 VGND 0.03115f
C19934 VPWR.n1653 VGND 0.03694f
C19935 VPWR.n1654 VGND 0.00833f
C19936 VPWR.t1959 VGND 0.01136f
C19937 VPWR.t1737 VGND 0.0124f
C19938 VPWR.n1655 VGND 0.02768f
C19939 VPWR.n1656 VGND 0.02818f
C19940 VPWR.n1657 VGND 0.01776f
C19941 VPWR.n1658 VGND 0.00697f
C19942 VPWR.n1659 VGND 0.01822f
C19943 VPWR.n1660 VGND 0.02384f
C19944 VPWR.n1661 VGND 0.17585f
C19945 VPWR.n1662 VGND 0.17585f
C19946 VPWR.n1663 VGND 0.02384f
C19947 VPWR.n1664 VGND 0.01776f
C19948 VPWR.t2043 VGND 0.0112f
C19949 VPWR.t1511 VGND 0.01226f
C19950 VPWR.n1665 VGND 0.02993f
C19951 VPWR.n1666 VGND 0.03284f
C19952 VPWR.n1667 VGND 0.03437f
C19953 VPWR.t1941 VGND 0.01116f
C19954 VPWR.t1542 VGND 0.01222f
C19955 VPWR.n1668 VGND 0.03115f
C19956 VPWR.n1669 VGND 0.03694f
C19957 VPWR.n1670 VGND 0.00833f
C19958 VPWR.t2050 VGND 0.01136f
C19959 VPWR.t1497 VGND 0.0124f
C19960 VPWR.n1671 VGND 0.02768f
C19961 VPWR.n1672 VGND 0.02818f
C19962 VPWR.n1673 VGND 0.01822f
C19963 VPWR.n1674 VGND 0.02384f
C19964 VPWR.n1675 VGND 0.01776f
C19965 VPWR.t2003 VGND 0.0112f
C19966 VPWR.t1615 VGND 0.01226f
C19967 VPWR.n1676 VGND 0.02993f
C19968 VPWR.n1677 VGND 0.03284f
C19969 VPWR.n1678 VGND 0.03437f
C19970 VPWR.t2038 VGND 0.01116f
C19971 VPWR.t1669 VGND 0.01222f
C19972 VPWR.n1679 VGND 0.03115f
C19973 VPWR.n1680 VGND 0.03694f
C19974 VPWR.n1681 VGND 0.00833f
C19975 VPWR.t1993 VGND 0.01136f
C19976 VPWR.t1650 VGND 0.0124f
C19977 VPWR.n1682 VGND 0.02768f
C19978 VPWR.n1683 VGND 0.02818f
C19979 VPWR.n1684 VGND 0.01776f
C19980 VPWR.n1685 VGND 0.00697f
C19981 VPWR.n1686 VGND 0.01822f
C19982 VPWR.n1687 VGND 0.02384f
C19983 VPWR.n1688 VGND 0.17585f
C19984 VPWR.n1689 VGND 0.17585f
C19985 VPWR.n1690 VGND 0.02384f
C19986 VPWR.n1691 VGND 0.01776f
C19987 VPWR.t1939 VGND 0.0112f
C19988 VPWR.t1793 VGND 0.01226f
C19989 VPWR.n1692 VGND 0.02993f
C19990 VPWR.n1693 VGND 0.03284f
C19991 VPWR.n1694 VGND 0.03437f
C19992 VPWR.t1978 VGND 0.01116f
C19993 VPWR.t1436 VGND 0.01222f
C19994 VPWR.n1695 VGND 0.03115f
C19995 VPWR.n1696 VGND 0.03694f
C19996 VPWR.n1697 VGND 0.00833f
C19997 VPWR.t2040 VGND 0.01136f
C19998 VPWR.t1522 VGND 0.0124f
C19999 VPWR.n1698 VGND 0.02768f
C20000 VPWR.n1699 VGND 0.02818f
C20001 VPWR.n1700 VGND 0.01822f
C20002 VPWR.n1701 VGND 0.02384f
C20003 VPWR.n1702 VGND 0.01776f
C20004 VPWR.t2036 VGND 0.0112f
C20005 VPWR.t1537 VGND 0.01226f
C20006 VPWR.n1703 VGND 0.02993f
C20007 VPWR.n1704 VGND 0.03284f
C20008 VPWR.n1705 VGND 0.03437f
C20009 VPWR.t1935 VGND 0.01116f
C20010 VPWR.t1674 VGND 0.01222f
C20011 VPWR.n1706 VGND 0.03115f
C20012 VPWR.n1707 VGND 0.03694f
C20013 VPWR.n1708 VGND 0.00833f
C20014 VPWR.t2033 VGND 0.01136f
C20015 VPWR.t1548 VGND 0.0124f
C20016 VPWR.n1709 VGND 0.02768f
C20017 VPWR.n1710 VGND 0.02818f
C20018 VPWR.n1711 VGND 0.01776f
C20019 VPWR.n1712 VGND 0.00697f
C20020 VPWR.n1713 VGND 0.01822f
C20021 VPWR.n1714 VGND 0.02384f
C20022 VPWR.n1715 VGND 0.17585f
C20023 VPWR.t1977 VGND 0.0112f
C20024 VPWR.t1694 VGND 0.01226f
C20025 VPWR.n1716 VGND 0.02993f
C20026 VPWR.n1717 VGND 0.03284f
C20027 VPWR.t2024 VGND 0.01116f
C20028 VPWR.t1702 VGND 0.01222f
C20029 VPWR.n1718 VGND 0.03115f
C20030 VPWR.n1719 VGND 0.03694f
C20031 VPWR.n1720 VGND 0.00833f
C20032 VPWR.t2019 VGND 0.01136f
C20033 VPWR.t1573 VGND 0.0124f
C20034 VPWR.n1721 VGND 0.02768f
C20035 VPWR.n1722 VGND 0.02818f
C20036 VPWR.n1723 VGND 0.01776f
C20037 VPWR.n1724 VGND 0.00697f
C20038 VPWR.n1725 VGND 0.01822f
C20039 VPWR.n1726 VGND 0.02384f
C20040 VPWR.n1727 VGND 0.21163f
C20041 VPWR.n1728 VGND 0.02541f
C20042 VPWR.n1729 VGND 0.01776f
C20043 VPWR.t1937 VGND 0.01136f
C20044 VPWR.t1418 VGND 0.0124f
C20045 VPWR.n1730 VGND 0.02768f
C20046 VPWR.n1731 VGND 0.02818f
C20047 VPWR.n1732 VGND 0.00833f
C20048 VPWR.t1984 VGND 0.01116f
C20049 VPWR.t1422 VGND 0.01222f
C20050 VPWR.n1733 VGND 0.03115f
C20051 VPWR.n1734 VGND 0.03694f
C20052 VPWR.n1735 VGND 0.03437f
C20053 VPWR.n1736 VGND 0.00805f
C20054 VPWR.n1737 VGND 0.01714f
C20055 VPWR.n1738 VGND 0.00725f
C20056 VPWR.n1739 VGND 0.10822f
C20057 VPWR.t1695 VGND 0.09218f
C20058 VPWR.t1574 VGND 0.07849f
C20059 VPWR.t1703 VGND 0.11957f
C20060 VPWR.n1740 VGND 0.10822f
C20061 VPWR.n1741 VGND 0.00725f
C20062 VPWR.n1742 VGND 0.01714f
C20063 VPWR.n1743 VGND 0.00805f
C20064 VPWR.n1744 VGND 0.0544f
C20065 VPWR.t2011 VGND 0.01116f
C20066 VPWR.t1457 VGND 0.01222f
C20067 VPWR.n1745 VGND 0.03042f
C20068 VPWR.n1746 VGND 0.00581f
C20069 VPWR.t1459 VGND 0.02679f
C20070 VPWR.n1747 VGND 0.05724f
C20071 VPWR.t333 VGND 0.02961f
C20072 VPWR.n1748 VGND 0.04692f
C20073 VPWR.t1716 VGND 0.07849f
C20074 VPWR.t332 VGND 0.09218f
C20075 VPWR.t1754 VGND 0.07849f
C20076 VPWR.t1495 VGND 0.11957f
C20077 VPWR.n1749 VGND 0.10822f
C20078 VPWR.n1750 VGND 0.00728f
C20079 VPWR.n1751 VGND 0.01797f
C20080 VPWR.n1752 VGND 0.13913f
C20081 VPWR.n1753 VGND -0.01866f
C20082 VPWR.n1754 VGND 0.08351f
C20083 VPWR.n1755 VGND 0.08351f
C20084 VPWR.n1756 VGND -0.01866f
C20085 VPWR.n1757 VGND 0.13913f
C20086 VPWR.n1758 VGND 0.01797f
C20087 VPWR.n1759 VGND 0.00728f
C20088 VPWR.n1760 VGND 0.10822f
C20089 VPWR.t1207 VGND 0.09218f
C20090 VPWR.t1698 VGND 0.07849f
C20091 VPWR.t1622 VGND 0.11957f
C20092 VPWR.n1761 VGND 0.10822f
C20093 VPWR.n1762 VGND 0.00728f
C20094 VPWR.n1763 VGND 0.01797f
C20095 VPWR.n1764 VGND 0.13913f
C20096 VPWR.n1765 VGND 0.0544f
C20097 VPWR.n1766 VGND 0.06567f
C20098 VPWR.n1767 VGND 0.09174f
C20099 VPWR.t1976 VGND 0.01136f
C20100 VPWR.t1697 VGND 0.0124f
C20101 VPWR.n1768 VGND 0.02769f
C20102 VPWR.n1769 VGND 0.01897f
C20103 VPWR.n1770 VGND 0.06244f
C20104 VPWR.n1771 VGND 0.09746f
C20105 VPWR.n1772 VGND 0.09174f
C20106 VPWR.t1968 VGND 0.01136f
C20107 VPWR.t1715 VGND 0.0124f
C20108 VPWR.n1773 VGND 0.02769f
C20109 VPWR.n1774 VGND 0.01897f
C20110 VPWR.n1775 VGND 0.06244f
C20111 VPWR.n1776 VGND 0.09746f
C20112 VPWR.t2013 VGND 0.01136f
C20113 VPWR.t1585 VGND 0.0124f
C20114 VPWR.n1777 VGND 0.02769f
C20115 VPWR.n1778 VGND 0.01897f
C20116 VPWR.n1779 VGND 0.06242f
C20117 VPWR.n1780 VGND 0.05139f
C20118 VPWR.t1953 VGND 0.01136f
C20119 VPWR.t1753 VGND 0.0124f
C20120 VPWR.n1781 VGND 0.02769f
C20121 VPWR.n1782 VGND 0.01897f
C20122 VPWR.n1783 VGND 0.06244f
C20123 VPWR.n1784 VGND 0.09746f
C20124 VPWR.n1785 VGND 0.09174f
C20125 VPWR.n1786 VGND 0.06567f
C20126 VPWR.n1787 VGND 0.0544f
C20127 VPWR.n1788 VGND 0.13913f
C20128 VPWR.n1789 VGND 0.01797f
C20129 VPWR.n1790 VGND 0.00728f
C20130 VPWR.n1791 VGND 0.10822f
C20131 VPWR.t1603 VGND 0.11957f
C20132 VPWR.t1586 VGND 0.07849f
C20133 VPWR.t1711 VGND 0.13333f
C20134 VPWR.n1792 VGND 0.07618f
C20135 VPWR.n1793 VGND 0.01797f
C20136 VPWR.n1794 VGND 0.13913f
C20137 VPWR.n1795 VGND 0.1646f
C20138 VPWR.n1796 VGND 1.01577f
C20139 VPWR.n1797 VGND 0.08351f
C20140 VPWR.n1798 VGND 0.08351f
C20141 VPWR.n1799 VGND 0.08351f
C20142 VPWR.n1800 VGND 0.08351f
C20143 VPWR.n1801 VGND 0.08351f
C20144 VPWR.n1802 VGND 0.08351f
C20145 VPWR.n1803 VGND 0.08351f
C20146 VPWR.n1804 VGND 0.08351f
C20147 VPWR.n1805 VGND 0.08351f
C20148 VPWR.n1806 VGND 0.08351f
C20149 VPWR.n1807 VGND 0.08351f
C20150 VPWR.n1808 VGND 0.08351f
C20151 VPWR.n1809 VGND 0.08351f
C20152 VPWR.n1810 VGND 0.08351f
C20153 VPWR.n1811 VGND 0.08351f
C20154 VPWR.n1812 VGND 0.19371f
C20155 VPWR.n1813 VGND 1.01577f
C20156 VPWR.n1814 VGND 1.01577f
C20157 VPWR.n1815 VGND 0.19371f
C20158 VPWR.n1816 VGND 0.13913f
C20159 VPWR.n1817 VGND 0.01797f
C20160 VPWR.n1818 VGND 0.07618f
C20161 VPWR.t1748 VGND 0.13333f
C20162 VPWR.t1331 VGND 0.07849f
C20163 VPWR.t185 VGND 0.11957f
C20164 VPWR.n1819 VGND 0.10822f
C20165 VPWR.n1820 VGND 0.00728f
C20166 VPWR.n1821 VGND 0.01797f
C20167 VPWR.n1822 VGND 0.13913f
C20168 VPWR.n1823 VGND 0.08351f
C20169 VPWR.n1824 VGND 0.08351f
C20170 VPWR.n1825 VGND 0.13913f
C20171 VPWR.n1826 VGND 0.01797f
C20172 VPWR.n1827 VGND 0.00728f
C20173 VPWR.n1828 VGND 0.10822f
C20174 VPWR.t1124 VGND 0.09218f
C20175 VPWR.t1151 VGND 0.07849f
C20176 VPWR.t98 VGND 0.11957f
C20177 VPWR.n1829 VGND 0.10822f
C20178 VPWR.n1830 VGND 0.00728f
C20179 VPWR.n1831 VGND 0.01797f
C20180 VPWR.n1832 VGND 0.13913f
C20181 VPWR.n1833 VGND 0.08351f
C20182 VPWR.n1834 VGND 0.08351f
C20183 VPWR.n1835 VGND 0.13913f
C20184 VPWR.n1836 VGND 0.01797f
C20185 VPWR.n1837 VGND 0.00728f
C20186 VPWR.n1838 VGND 0.10822f
C20187 VPWR.t1848 VGND 0.09218f
C20188 VPWR.t22 VGND 0.07849f
C20189 VPWR.t127 VGND 0.11957f
C20190 VPWR.n1839 VGND 0.10822f
C20191 VPWR.n1840 VGND 0.00728f
C20192 VPWR.n1841 VGND 0.01797f
C20193 VPWR.n1842 VGND 0.13913f
C20194 VPWR.n1843 VGND 0.08351f
C20195 VPWR.n1844 VGND 0.08351f
C20196 VPWR.n1845 VGND 0.13913f
C20197 VPWR.n1846 VGND 0.01797f
C20198 VPWR.n1847 VGND 0.00728f
C20199 VPWR.n1848 VGND 0.10822f
C20200 VPWR.t1384 VGND 0.09218f
C20201 VPWR.t1329 VGND 0.07849f
C20202 VPWR.t641 VGND 0.11957f
C20203 VPWR.n1849 VGND 0.10822f
C20204 VPWR.n1850 VGND 0.00728f
C20205 VPWR.n1851 VGND 0.01797f
C20206 VPWR.n1852 VGND 0.13913f
C20207 VPWR.n1853 VGND 0.08351f
C20208 VPWR.n1854 VGND 0.08351f
C20209 VPWR.n1855 VGND 0.13913f
C20210 VPWR.n1856 VGND 0.01797f
C20211 VPWR.n1857 VGND 0.00728f
C20212 VPWR.n1858 VGND 0.10822f
C20213 VPWR.t585 VGND 0.09218f
C20214 VPWR.t19 VGND 0.07849f
C20215 VPWR.t296 VGND 0.11957f
C20216 VPWR.n1859 VGND 0.10822f
C20217 VPWR.n1860 VGND 0.00728f
C20218 VPWR.n1861 VGND 0.01797f
C20219 VPWR.n1862 VGND 0.13913f
C20220 VPWR.n1863 VGND 0.08351f
C20221 VPWR.n1864 VGND 0.08351f
C20222 VPWR.n1865 VGND 0.13913f
C20223 VPWR.n1866 VGND 0.01797f
C20224 VPWR.n1867 VGND 0.00728f
C20225 VPWR.n1868 VGND 0.10822f
C20226 VPWR.t265 VGND 0.09218f
C20227 VPWR.t1328 VGND 0.07849f
C20228 VPWR.t173 VGND 0.11957f
C20229 VPWR.n1869 VGND 0.10822f
C20230 VPWR.n1870 VGND 0.00728f
C20231 VPWR.n1871 VGND 0.01797f
C20232 VPWR.n1872 VGND 0.13913f
C20233 VPWR.n1873 VGND 0.08351f
C20234 VPWR.n1874 VGND 0.08351f
C20235 VPWR.n1875 VGND 0.13913f
C20236 VPWR.n1876 VGND 0.01797f
C20237 VPWR.n1877 VGND 0.00728f
C20238 VPWR.n1878 VGND 0.10822f
C20239 VPWR.t1015 VGND 0.09218f
C20240 VPWR.t24 VGND 0.07849f
C20241 VPWR.t748 VGND 0.11957f
C20242 VPWR.n1879 VGND 0.10822f
C20243 VPWR.n1880 VGND 0.00728f
C20244 VPWR.n1881 VGND 0.01797f
C20245 VPWR.n1882 VGND 0.13913f
C20246 VPWR.n1883 VGND 0.08351f
C20247 VPWR.n1884 VGND 0.08351f
C20248 VPWR.n1885 VGND 0.13913f
C20249 VPWR.n1886 VGND 0.01797f
C20250 VPWR.n1887 VGND 0.00728f
C20251 VPWR.n1888 VGND 0.10822f
C20252 VPWR.t489 VGND 0.09218f
C20253 VPWR.t1330 VGND 0.07849f
C20254 VPWR.t157 VGND 0.11957f
C20255 VPWR.n1889 VGND 0.10822f
C20256 VPWR.n1890 VGND 0.00728f
C20257 VPWR.n1891 VGND 0.01797f
C20258 VPWR.n1892 VGND 0.13913f
C20259 VPWR.n1893 VGND 0.08351f
C20260 VPWR.n1894 VGND 1.0094f
C20261 VPWR.n1895 VGND 0.19371f
C20262 VPWR.n1896 VGND 0.08351f
C20263 VPWR.n1897 VGND 0.08351f
C20264 VPWR.n1898 VGND 0.08351f
C20265 VPWR.n1899 VGND 0.08351f
C20266 VPWR.n1900 VGND 0.08351f
C20267 VPWR.n1901 VGND 0.08351f
C20268 VPWR.n1902 VGND 0.08351f
C20269 VPWR.n1903 VGND 0.08351f
C20270 VPWR.n1904 VGND 0.08351f
C20271 VPWR.n1905 VGND 0.08351f
C20272 VPWR.n1906 VGND 0.08351f
C20273 VPWR.n1907 VGND 0.08351f
C20274 VPWR.n1908 VGND 0.08351f
C20275 VPWR.n1909 VGND 0.08351f
C20276 VPWR.n1910 VGND 0.08351f
C20277 VPWR.n1911 VGND 1.0094f
C20278 VPWR.n1912 VGND 1.0094f
C20279 VPWR.n1913 VGND 0.08351f
C20280 VPWR.n1914 VGND 0.13913f
C20281 VPWR.n1915 VGND 0.01797f
C20282 VPWR.n1916 VGND 0.00728f
C20283 VPWR.n1917 VGND 0.10822f
C20284 VPWR.t147 VGND 0.11957f
C20285 VPWR.t1826 VGND 0.07849f
C20286 VPWR.t687 VGND 0.09218f
C20287 VPWR.t532 VGND 0.07849f
C20288 VPWR.t681 VGND 0.11957f
C20289 VPWR.n1918 VGND 0.10822f
C20290 VPWR.n1919 VGND 0.00728f
C20291 VPWR.n1920 VGND 0.01797f
C20292 VPWR.n1921 VGND 0.13913f
C20293 VPWR.n1922 VGND 0.08351f
C20294 VPWR.n1923 VGND 0.08351f
C20295 VPWR.n1924 VGND 0.13913f
C20296 VPWR.n1925 VGND 0.01797f
C20297 VPWR.n1926 VGND 0.00728f
C20298 VPWR.n1927 VGND 0.10822f
C20299 VPWR.t764 VGND 0.11957f
C20300 VPWR.t366 VGND 0.07849f
C20301 VPWR.t1174 VGND 0.09218f
C20302 VPWR.t362 VGND 0.07849f
C20303 VPWR.t1021 VGND 0.11957f
C20304 VPWR.n1928 VGND 0.10822f
C20305 VPWR.n1929 VGND 0.00728f
C20306 VPWR.n1930 VGND 0.01797f
C20307 VPWR.n1931 VGND 0.13913f
C20308 VPWR.n1932 VGND 0.08351f
C20309 VPWR.n1933 VGND 0.08351f
C20310 VPWR.n1934 VGND 0.13913f
C20311 VPWR.n1935 VGND 0.01797f
C20312 VPWR.n1936 VGND 0.00728f
C20313 VPWR.n1937 VGND 0.10822f
C20314 VPWR.t916 VGND 0.11957f
C20315 VPWR.t537 VGND 0.07849f
C20316 VPWR.t269 VGND 0.09218f
C20317 VPWR.t536 VGND 0.07849f
C20318 VPWR.t233 VGND 0.11957f
C20319 VPWR.n1938 VGND 0.10822f
C20320 VPWR.n1939 VGND 0.00728f
C20321 VPWR.n1940 VGND 0.01797f
C20322 VPWR.n1941 VGND 0.13913f
C20323 VPWR.n1942 VGND 0.08351f
C20324 VPWR.n1943 VGND 0.08351f
C20325 VPWR.n1944 VGND 0.13913f
C20326 VPWR.n1945 VGND 0.01797f
C20327 VPWR.n1946 VGND 0.00728f
C20328 VPWR.n1947 VGND 0.10822f
C20329 VPWR.t1891 VGND 0.11957f
C20330 VPWR.t361 VGND 0.07849f
C20331 VPWR.t841 VGND 0.09218f
C20332 VPWR.t360 VGND 0.07849f
C20333 VPWR.t939 VGND 0.11957f
C20334 VPWR.n1948 VGND 0.10822f
C20335 VPWR.n1949 VGND 0.00728f
C20336 VPWR.n1950 VGND 0.01797f
C20337 VPWR.n1951 VGND 0.13913f
C20338 VPWR.n1952 VGND 0.08351f
C20339 VPWR.n1953 VGND 0.08351f
C20340 VPWR.n1954 VGND 0.13913f
C20341 VPWR.n1955 VGND 0.01797f
C20342 VPWR.n1956 VGND 0.00728f
C20343 VPWR.n1957 VGND 0.10822f
C20344 VPWR.t493 VGND 0.11957f
C20345 VPWR.t538 VGND 0.07849f
C20346 VPWR.t549 VGND 0.09218f
C20347 VPWR.t365 VGND 0.07849f
C20348 VPWR.t543 VGND 0.11957f
C20349 VPWR.n1958 VGND 0.10822f
C20350 VPWR.n1959 VGND 0.00728f
C20351 VPWR.n1960 VGND 0.01797f
C20352 VPWR.n1961 VGND 0.13913f
C20353 VPWR.n1962 VGND 0.08351f
C20354 VPWR.n1963 VGND 0.08351f
C20355 VPWR.n1964 VGND 0.13913f
C20356 VPWR.n1965 VGND 0.01797f
C20357 VPWR.n1966 VGND 0.00728f
C20358 VPWR.n1967 VGND 0.10822f
C20359 VPWR.t445 VGND 0.11957f
C20360 VPWR.t364 VGND 0.07849f
C20361 VPWR.t863 VGND 0.09218f
C20362 VPWR.t535 VGND 0.07849f
C20363 VPWR.t857 VGND 0.11957f
C20364 VPWR.n1968 VGND 0.10822f
C20365 VPWR.n1969 VGND 0.00728f
C20366 VPWR.n1970 VGND 0.01797f
C20367 VPWR.n1971 VGND 0.13913f
C20368 VPWR.n1972 VGND 0.08351f
C20369 VPWR.n1973 VGND 0.08351f
C20370 VPWR.n1974 VGND 0.13913f
C20371 VPWR.n1975 VGND 0.01797f
C20372 VPWR.n1976 VGND 0.00728f
C20373 VPWR.n1977 VGND 0.10822f
C20374 VPWR.t1872 VGND 0.11957f
C20375 VPWR.t534 VGND 0.07849f
C20376 VPWR.t153 VGND 0.09218f
C20377 VPWR.t533 VGND 0.07849f
C20378 VPWR.t1118 VGND 0.11957f
C20379 VPWR.n1978 VGND 0.10822f
C20380 VPWR.n1979 VGND 0.00728f
C20381 VPWR.n1980 VGND 0.01797f
C20382 VPWR.n1981 VGND 0.13913f
C20383 VPWR.n1982 VGND 0.08351f
C20384 VPWR.n1983 VGND 0.08351f
C20385 VPWR.n1984 VGND 0.13913f
C20386 VPWR.n1985 VGND 0.01797f
C20387 VPWR.n1986 VGND 0.00728f
C20388 VPWR.n1987 VGND 0.10822f
C20389 VPWR.t316 VGND 0.11957f
C20390 VPWR.t1827 VGND 0.07849f
C20391 VPWR.t1453 VGND 0.13333f
C20392 VPWR.n1988 VGND 0.07618f
C20393 VPWR.n1989 VGND 0.01797f
C20394 VPWR.n1990 VGND 0.13913f
C20395 VPWR.n1991 VGND 0.19371f
C20396 VPWR.n1992 VGND 1.01577f
C20397 VPWR.n1993 VGND 0.08351f
C20398 VPWR.n1994 VGND 0.08351f
C20399 VPWR.n1995 VGND 0.08351f
C20400 VPWR.n1996 VGND 0.08351f
C20401 VPWR.n1997 VGND 0.08351f
C20402 VPWR.n1998 VGND 0.08351f
C20403 VPWR.n1999 VGND 0.08351f
C20404 VPWR.n2000 VGND 0.08351f
C20405 VPWR.n2001 VGND 0.08351f
C20406 VPWR.n2002 VGND 0.08351f
C20407 VPWR.n2003 VGND 0.08351f
C20408 VPWR.n2004 VGND 0.08351f
C20409 VPWR.n2005 VGND 0.08351f
C20410 VPWR.n2006 VGND 0.08351f
C20411 VPWR.n2007 VGND 0.08351f
C20412 VPWR.n2008 VGND 0.19371f
C20413 VPWR.n2009 VGND 1.01577f
C20414 VPWR.n2010 VGND 1.01577f
C20415 VPWR.n2011 VGND 0.19371f
C20416 VPWR.n2012 VGND 0.13913f
C20417 VPWR.n2013 VGND 0.01797f
C20418 VPWR.n2014 VGND 0.07618f
C20419 VPWR.t1528 VGND 0.13333f
C20420 VPWR.t378 VGND 0.07849f
C20421 VPWR.t344 VGND 0.11957f
C20422 VPWR.n2015 VGND 0.10822f
C20423 VPWR.n2016 VGND 0.00728f
C20424 VPWR.n2017 VGND 0.01797f
C20425 VPWR.n2018 VGND 0.13913f
C20426 VPWR.n2019 VGND 0.08351f
C20427 VPWR.n2020 VGND 0.08351f
C20428 VPWR.n2021 VGND 0.13913f
C20429 VPWR.n2022 VGND 0.01797f
C20430 VPWR.n2023 VGND 0.00728f
C20431 VPWR.n2024 VGND 0.10822f
C20432 VPWR.t668 VGND 0.09218f
C20433 VPWR.t381 VGND 0.07849f
C20434 VPWR.t1213 VGND 0.11957f
C20435 VPWR.n2025 VGND 0.10822f
C20436 VPWR.n2026 VGND 0.00728f
C20437 VPWR.n2027 VGND 0.01797f
C20438 VPWR.n2028 VGND 0.13913f
C20439 VPWR.n2029 VGND 0.08351f
C20440 VPWR.n2030 VGND 0.08351f
C20441 VPWR.n2031 VGND 0.13913f
C20442 VPWR.n2032 VGND 0.01797f
C20443 VPWR.n2033 VGND 0.00728f
C20444 VPWR.n2034 VGND 0.10822f
C20445 VPWR.t953 VGND 0.09218f
C20446 VPWR.t1884 VGND 0.07849f
C20447 VPWR.t1114 VGND 0.11957f
C20448 VPWR.n2035 VGND 0.10822f
C20449 VPWR.n2036 VGND 0.00728f
C20450 VPWR.n2037 VGND 0.01797f
C20451 VPWR.n2038 VGND 0.13913f
C20452 VPWR.n2039 VGND 0.08351f
C20453 VPWR.n2040 VGND 0.08351f
C20454 VPWR.n2041 VGND 0.13913f
C20455 VPWR.n2042 VGND 0.01797f
C20456 VPWR.n2043 VGND 0.00728f
C20457 VPWR.n2044 VGND 0.10822f
C20458 VPWR.t539 VGND 0.09218f
C20459 VPWR.t385 VGND 0.07849f
C20460 VPWR.t141 VGND 0.11957f
C20461 VPWR.n2045 VGND 0.10822f
C20462 VPWR.n2046 VGND 0.00728f
C20463 VPWR.n2047 VGND 0.01797f
C20464 VPWR.n2048 VGND 0.13913f
C20465 VPWR.n2049 VGND 0.08351f
C20466 VPWR.n2050 VGND 0.08351f
C20467 VPWR.n2051 VGND 0.13913f
C20468 VPWR.n2052 VGND 0.01797f
C20469 VPWR.n2053 VGND 0.00728f
C20470 VPWR.n2054 VGND 0.10822f
C20471 VPWR.t467 VGND 0.09218f
C20472 VPWR.t1881 VGND 0.07849f
C20473 VPWR.t358 VGND 0.11957f
C20474 VPWR.n2055 VGND 0.10822f
C20475 VPWR.n2056 VGND 0.00728f
C20476 VPWR.n2057 VGND 0.01797f
C20477 VPWR.n2058 VGND 0.13913f
C20478 VPWR.n2059 VGND 0.08351f
C20479 VPWR.n2060 VGND 0.08351f
C20480 VPWR.n2061 VGND 0.13913f
C20481 VPWR.n2062 VGND 0.01797f
C20482 VPWR.n2063 VGND 0.00728f
C20483 VPWR.n2064 VGND 0.10822f
C20484 VPWR.t229 VGND 0.09218f
C20485 VPWR.t384 VGND 0.07849f
C20486 VPWR.t1223 VGND 0.11957f
C20487 VPWR.n2065 VGND 0.10822f
C20488 VPWR.n2066 VGND 0.00728f
C20489 VPWR.n2067 VGND 0.01797f
C20490 VPWR.n2068 VGND 0.13913f
C20491 VPWR.n2069 VGND 0.08351f
C20492 VPWR.n2070 VGND 0.08351f
C20493 VPWR.n2071 VGND 0.13913f
C20494 VPWR.n2072 VGND 0.01797f
C20495 VPWR.n2073 VGND 0.00728f
C20496 VPWR.n2074 VGND 0.10822f
C20497 VPWR.t604 VGND 0.09218f
C20498 VPWR.t1886 VGND 0.07849f
C20499 VPWR.t774 VGND 0.11957f
C20500 VPWR.n2075 VGND 0.10822f
C20501 VPWR.n2076 VGND 0.00728f
C20502 VPWR.n2077 VGND 0.01797f
C20503 VPWR.n2078 VGND 0.13913f
C20504 VPWR.n2079 VGND 0.08351f
C20505 VPWR.n2080 VGND 0.08351f
C20506 VPWR.n2081 VGND 0.13913f
C20507 VPWR.n2082 VGND 0.01797f
C20508 VPWR.n2083 VGND 0.00728f
C20509 VPWR.n2084 VGND 0.10822f
C20510 VPWR.t1291 VGND 0.09218f
C20511 VPWR.t386 VGND 0.07849f
C20512 VPWR.t827 VGND 0.11957f
C20513 VPWR.n2085 VGND 0.10822f
C20514 VPWR.n2086 VGND 0.00728f
C20515 VPWR.n2087 VGND 0.01797f
C20516 VPWR.n2088 VGND 0.13913f
C20517 VPWR.n2089 VGND 0.08351f
C20518 VPWR.n2090 VGND 1.0094f
C20519 VPWR.n2091 VGND 0.19371f
C20520 VPWR.n2092 VGND 0.08351f
C20521 VPWR.n2093 VGND 0.08351f
C20522 VPWR.n2094 VGND 0.08351f
C20523 VPWR.n2095 VGND 0.08351f
C20524 VPWR.n2096 VGND 0.08351f
C20525 VPWR.n2097 VGND 0.08351f
C20526 VPWR.n2098 VGND 0.08351f
C20527 VPWR.n2099 VGND 0.08351f
C20528 VPWR.n2100 VGND 0.08351f
C20529 VPWR.n2101 VGND 0.08351f
C20530 VPWR.n2102 VGND 0.08351f
C20531 VPWR.n2103 VGND 0.08351f
C20532 VPWR.n2104 VGND 0.08351f
C20533 VPWR.n2105 VGND 0.08351f
C20534 VPWR.n2106 VGND 0.08351f
C20535 VPWR.n2107 VGND 1.0094f
C20536 VPWR.n2108 VGND 1.0094f
C20537 VPWR.n2109 VGND 0.08351f
C20538 VPWR.n2110 VGND 0.13913f
C20539 VPWR.n2111 VGND 0.01797f
C20540 VPWR.n2112 VGND 0.00728f
C20541 VPWR.n2113 VGND 0.10822f
C20542 VPWR.t145 VGND 0.11957f
C20543 VPWR.t1178 VGND 0.07849f
C20544 VPWR.t685 VGND 0.09218f
C20545 VPWR.t594 VGND 0.07849f
C20546 VPWR.t679 VGND 0.11957f
C20547 VPWR.n2114 VGND 0.10822f
C20548 VPWR.n2115 VGND 0.00728f
C20549 VPWR.n2116 VGND 0.01797f
C20550 VPWR.n2117 VGND 0.13913f
C20551 VPWR.n2118 VGND 0.08351f
C20552 VPWR.n2119 VGND 0.08351f
C20553 VPWR.n2120 VGND 0.13913f
C20554 VPWR.n2121 VGND 0.01797f
C20555 VPWR.n2122 VGND 0.00728f
C20556 VPWR.n2123 VGND 0.10822f
C20557 VPWR.t766 VGND 0.11957f
C20558 VPWR.t593 VGND 0.07849f
C20559 VPWR.t1170 VGND 0.09218f
C20560 VPWR.t198 VGND 0.07849f
C20561 VPWR.t1824 VGND 0.11957f
C20562 VPWR.n2124 VGND 0.10822f
C20563 VPWR.n2125 VGND 0.00728f
C20564 VPWR.n2126 VGND 0.01797f
C20565 VPWR.n2127 VGND 0.13913f
C20566 VPWR.n2128 VGND 0.08351f
C20567 VPWR.n2129 VGND 0.08351f
C20568 VPWR.n2130 VGND 0.13913f
C20569 VPWR.n2131 VGND 0.01797f
C20570 VPWR.n2132 VGND 0.00728f
C20571 VPWR.n2133 VGND 0.10822f
C20572 VPWR.t1227 VGND 0.11957f
C20573 VPWR.t1245 VGND 0.07849f
C20574 VPWR.t267 VGND 0.09218f
C20575 VPWR.t1244 VGND 0.07849f
C20576 VPWR.t231 VGND 0.11957f
C20577 VPWR.n2134 VGND 0.10822f
C20578 VPWR.n2135 VGND 0.00728f
C20579 VPWR.n2136 VGND 0.01797f
C20580 VPWR.n2137 VGND 0.13913f
C20581 VPWR.n2138 VGND 0.08351f
C20582 VPWR.n2139 VGND 0.08351f
C20583 VPWR.n2140 VGND 0.13913f
C20584 VPWR.n2141 VGND 0.01797f
C20585 VPWR.n2142 VGND 0.00728f
C20586 VPWR.n2143 VGND 0.10822f
C20587 VPWR.t1889 VGND 0.11957f
C20588 VPWR.t197 VGND 0.07849f
C20589 VPWR.t839 VGND 0.09218f
C20590 VPWR.t1180 VGND 0.07849f
C20591 VPWR.t937 VGND 0.11957f
C20592 VPWR.n2144 VGND 0.10822f
C20593 VPWR.n2145 VGND 0.00728f
C20594 VPWR.n2146 VGND 0.01797f
C20595 VPWR.n2147 VGND 0.13913f
C20596 VPWR.n2148 VGND 0.08351f
C20597 VPWR.n2149 VGND 0.08351f
C20598 VPWR.n2150 VGND 0.13913f
C20599 VPWR.n2151 VGND 0.01797f
C20600 VPWR.n2152 VGND 0.00728f
C20601 VPWR.n2153 VGND 0.10822f
C20602 VPWR.t370 VGND 0.11957f
C20603 VPWR.t1246 VGND 0.07849f
C20604 VPWR.t547 VGND 0.09218f
C20605 VPWR.t671 VGND 0.07849f
C20606 VPWR.t541 VGND 0.11957f
C20607 VPWR.n2154 VGND 0.10822f
C20608 VPWR.n2155 VGND 0.00728f
C20609 VPWR.n2156 VGND 0.01797f
C20610 VPWR.n2157 VGND 0.13913f
C20611 VPWR.n2158 VGND 0.08351f
C20612 VPWR.n2159 VGND 0.08351f
C20613 VPWR.n2160 VGND 0.13913f
C20614 VPWR.n2161 VGND 0.01797f
C20615 VPWR.n2162 VGND 0.00728f
C20616 VPWR.n2163 VGND 0.10822f
C20617 VPWR.t443 VGND 0.11957f
C20618 VPWR.t670 VGND 0.07849f
C20619 VPWR.t861 VGND 0.09218f
C20620 VPWR.t1243 VGND 0.07849f
C20621 VPWR.t955 VGND 0.11957f
C20622 VPWR.n2164 VGND 0.10822f
C20623 VPWR.n2165 VGND 0.00728f
C20624 VPWR.n2166 VGND 0.01797f
C20625 VPWR.n2167 VGND 0.13913f
C20626 VPWR.n2168 VGND 0.08351f
C20627 VPWR.n2169 VGND 0.08351f
C20628 VPWR.n2170 VGND 0.13913f
C20629 VPWR.n2171 VGND 0.01797f
C20630 VPWR.n2172 VGND 0.00728f
C20631 VPWR.n2173 VGND 0.10822f
C20632 VPWR.t1870 VGND 0.11957f
C20633 VPWR.t673 VGND 0.07849f
C20634 VPWR.t151 VGND 0.09218f
C20635 VPWR.t672 VGND 0.07849f
C20636 VPWR.t1116 VGND 0.11957f
C20637 VPWR.n2174 VGND 0.10822f
C20638 VPWR.n2175 VGND 0.00728f
C20639 VPWR.n2176 VGND 0.01797f
C20640 VPWR.n2177 VGND 0.13913f
C20641 VPWR.n2178 VGND 0.08351f
C20642 VPWR.n2179 VGND 0.08351f
C20643 VPWR.n2180 VGND 0.13913f
C20644 VPWR.n2181 VGND 0.01797f
C20645 VPWR.n2182 VGND 0.00728f
C20646 VPWR.n2183 VGND 0.10822f
C20647 VPWR.t314 VGND 0.11957f
C20648 VPWR.t1179 VGND 0.07849f
C20649 VPWR.t1461 VGND 0.13333f
C20650 VPWR.n2184 VGND 0.07618f
C20651 VPWR.n2185 VGND 0.01797f
C20652 VPWR.n2186 VGND 0.13913f
C20653 VPWR.n2187 VGND 0.19371f
C20654 VPWR.n2188 VGND 1.01577f
C20655 VPWR.n2189 VGND 0.08351f
C20656 VPWR.n2190 VGND 0.08351f
C20657 VPWR.n2191 VGND 0.08351f
C20658 VPWR.n2192 VGND 0.08351f
C20659 VPWR.n2193 VGND 0.08351f
C20660 VPWR.n2194 VGND 0.08351f
C20661 VPWR.n2195 VGND 0.08351f
C20662 VPWR.n2196 VGND 0.08351f
C20663 VPWR.n2197 VGND 0.08351f
C20664 VPWR.n2198 VGND 0.08351f
C20665 VPWR.n2199 VGND 0.08351f
C20666 VPWR.n2200 VGND 0.08351f
C20667 VPWR.n2201 VGND 0.08351f
C20668 VPWR.n2202 VGND 0.08351f
C20669 VPWR.n2203 VGND 0.08351f
C20670 VPWR.n2204 VGND 0.19371f
C20671 VPWR.n2205 VGND 1.01577f
C20672 VPWR.n2206 VGND 1.01577f
C20673 VPWR.n2207 VGND 0.19371f
C20674 VPWR.n2208 VGND 0.13913f
C20675 VPWR.n2209 VGND 0.01797f
C20676 VPWR.n2210 VGND 0.07618f
C20677 VPWR.t1627 VGND 0.13333f
C20678 VPWR.t1803 VGND 0.07849f
C20679 VPWR.t528 VGND 0.11957f
C20680 VPWR.n2211 VGND 0.10822f
C20681 VPWR.n2212 VGND 0.00728f
C20682 VPWR.n2213 VGND 0.01797f
C20683 VPWR.n2214 VGND 0.13913f
C20684 VPWR.n2215 VGND 0.08351f
C20685 VPWR.n2216 VGND 0.08351f
C20686 VPWR.n2217 VGND 0.13913f
C20687 VPWR.n2218 VGND 0.01797f
C20688 VPWR.n2219 VGND 0.00728f
C20689 VPWR.n2220 VGND 0.10822f
C20690 VPWR.t6 VGND 0.09218f
C20691 VPWR.t1347 VGND 0.07849f
C20692 VPWR.t69 VGND 0.11957f
C20693 VPWR.n2221 VGND 0.10822f
C20694 VPWR.n2222 VGND 0.00728f
C20695 VPWR.n2223 VGND 0.01797f
C20696 VPWR.n2224 VGND 0.13913f
C20697 VPWR.n2225 VGND 0.08351f
C20698 VPWR.n2226 VGND 0.08351f
C20699 VPWR.n2227 VGND 0.13913f
C20700 VPWR.n2228 VGND 0.01797f
C20701 VPWR.n2229 VGND 0.00728f
C20702 VPWR.n2230 VGND 0.10822f
C20703 VPWR.t1189 VGND 0.09218f
C20704 VPWR.t1342 VGND 0.07849f
C20705 VPWR.t53 VGND 0.11957f
C20706 VPWR.n2231 VGND 0.10822f
C20707 VPWR.n2232 VGND 0.00728f
C20708 VPWR.n2233 VGND 0.01797f
C20709 VPWR.n2234 VGND 0.13913f
C20710 VPWR.n2235 VGND 0.08351f
C20711 VPWR.n2236 VGND 0.08351f
C20712 VPWR.n2237 VGND 0.13913f
C20713 VPWR.n2238 VGND 0.01797f
C20714 VPWR.n2239 VGND 0.00728f
C20715 VPWR.n2240 VGND 0.10822f
C20716 VPWR.t892 VGND 0.09218f
C20717 VPWR.t1351 VGND 0.07849f
C20718 VPWR.t1276 VGND 0.11957f
C20719 VPWR.n2241 VGND 0.10822f
C20720 VPWR.n2242 VGND 0.00728f
C20721 VPWR.n2243 VGND 0.01797f
C20722 VPWR.n2244 VGND 0.13913f
C20723 VPWR.n2245 VGND 0.08351f
C20724 VPWR.n2246 VGND 0.08351f
C20725 VPWR.n2247 VGND 0.13913f
C20726 VPWR.n2248 VGND 0.01797f
C20727 VPWR.n2249 VGND 0.00728f
C20728 VPWR.n2250 VGND 0.10822f
C20729 VPWR.t992 VGND 0.09218f
C20730 VPWR.t1805 VGND 0.07849f
C20731 VPWR.t423 VGND 0.11957f
C20732 VPWR.n2251 VGND 0.10822f
C20733 VPWR.n2252 VGND 0.00728f
C20734 VPWR.n2253 VGND 0.01797f
C20735 VPWR.n2254 VGND 0.13913f
C20736 VPWR.n2255 VGND 0.08351f
C20737 VPWR.n2256 VGND 0.08351f
C20738 VPWR.n2257 VGND 0.13913f
C20739 VPWR.n2258 VGND 0.01797f
C20740 VPWR.n2259 VGND 0.00728f
C20741 VPWR.n2260 VGND 0.10822f
C20742 VPWR.t249 VGND 0.09218f
C20743 VPWR.t1350 VGND 0.07849f
C20744 VPWR.t1236 VGND 0.11957f
C20745 VPWR.n2261 VGND 0.10822f
C20746 VPWR.n2262 VGND 0.00728f
C20747 VPWR.n2263 VGND 0.01797f
C20748 VPWR.n2264 VGND 0.13913f
C20749 VPWR.n2265 VGND 0.08351f
C20750 VPWR.n2266 VGND 0.08351f
C20751 VPWR.n2267 VGND 0.13913f
C20752 VPWR.n2268 VGND 0.01797f
C20753 VPWR.n2269 VGND 0.00728f
C20754 VPWR.n2270 VGND 0.10822f
C20755 VPWR.t1820 VGND 0.09218f
C20756 VPWR.t1344 VGND 0.07849f
C20757 VPWR.t732 VGND 0.11957f
C20758 VPWR.n2271 VGND 0.10822f
C20759 VPWR.n2272 VGND 0.00728f
C20760 VPWR.n2273 VGND 0.01797f
C20761 VPWR.n2274 VGND 0.13913f
C20762 VPWR.n2275 VGND 0.08351f
C20763 VPWR.n2276 VGND 0.08351f
C20764 VPWR.n2277 VGND 0.13913f
C20765 VPWR.n2278 VGND 0.01797f
C20766 VPWR.n2279 VGND 0.00728f
C20767 VPWR.n2280 VGND 0.10822f
C20768 VPWR.t1260 VGND 0.09218f
C20769 VPWR.t1802 VGND 0.07849f
C20770 VPWR.t1156 VGND 0.11957f
C20771 VPWR.n2281 VGND 0.10822f
C20772 VPWR.n2282 VGND 0.00728f
C20773 VPWR.n2283 VGND 0.01797f
C20774 VPWR.n2284 VGND 0.13913f
C20775 VPWR.n2285 VGND 0.08351f
C20776 VPWR.n2286 VGND 1.0094f
C20777 VPWR.n2287 VGND 0.19371f
C20778 VPWR.n2288 VGND 0.08351f
C20779 VPWR.n2289 VGND 0.08351f
C20780 VPWR.n2290 VGND 0.08351f
C20781 VPWR.n2291 VGND 0.08351f
C20782 VPWR.n2292 VGND 0.08351f
C20783 VPWR.n2293 VGND 0.08351f
C20784 VPWR.n2294 VGND 0.08351f
C20785 VPWR.n2295 VGND 0.08351f
C20786 VPWR.n2296 VGND 0.08351f
C20787 VPWR.n2297 VGND 0.08351f
C20788 VPWR.n2298 VGND 0.08351f
C20789 VPWR.n2299 VGND 0.08351f
C20790 VPWR.n2300 VGND 0.08351f
C20791 VPWR.n2301 VGND 0.08351f
C20792 VPWR.n2302 VGND 0.08351f
C20793 VPWR.n2303 VGND 1.0094f
C20794 VPWR.n2304 VGND 1.0094f
C20795 VPWR.n2305 VGND 0.08351f
C20796 VPWR.n2306 VGND 0.13913f
C20797 VPWR.n2307 VGND 0.01797f
C20798 VPWR.n2308 VGND 0.00728f
C20799 VPWR.n2309 VGND 0.10822f
C20800 VPWR.t1146 VGND 0.11957f
C20801 VPWR.t453 VGND 0.07849f
C20802 VPWR.t1287 VGND 0.09218f
C20803 VPWR.t1856 VGND 0.07849f
C20804 VPWR.t218 VGND 0.11957f
C20805 VPWR.n2310 VGND 0.10822f
C20806 VPWR.n2311 VGND 0.00728f
C20807 VPWR.n2312 VGND 0.01797f
C20808 VPWR.n2313 VGND 0.13913f
C20809 VPWR.n2314 VGND 0.08351f
C20810 VPWR.n2315 VGND 0.08351f
C20811 VPWR.n2316 VGND 0.13913f
C20812 VPWR.n2317 VGND 0.01797f
C20813 VPWR.n2318 VGND 0.00728f
C20814 VPWR.n2319 VGND 0.10822f
C20815 VPWR.t778 VGND 0.11957f
C20816 VPWR.t1855 VGND 0.07849f
C20817 VPWR.t602 VGND 0.09218f
C20818 VPWR.t375 VGND 0.07849f
C20819 VPWR.t1061 VGND 0.11957f
C20820 VPWR.n2320 VGND 0.10822f
C20821 VPWR.n2321 VGND 0.00728f
C20822 VPWR.n2322 VGND 0.01797f
C20823 VPWR.n2323 VGND 0.13913f
C20824 VPWR.n2324 VGND 0.08351f
C20825 VPWR.n2325 VGND 0.08351f
C20826 VPWR.n2326 VGND 0.13913f
C20827 VPWR.n2327 VGND 0.01797f
C20828 VPWR.n2328 VGND 0.00728f
C20829 VPWR.n2329 VGND 0.10822f
C20830 VPWR.t1388 VGND 0.11957f
C20831 VPWR.t451 VGND 0.07849f
C20832 VPWR.t796 VGND 0.09218f
C20833 VPWR.t450 VGND 0.07849f
C20834 VPWR.t792 VGND 0.11957f
C20835 VPWR.n2330 VGND 0.10822f
C20836 VPWR.n2331 VGND 0.00728f
C20837 VPWR.n2332 VGND 0.01797f
C20838 VPWR.n2333 VGND 0.13913f
C20839 VPWR.n2334 VGND 0.08351f
C20840 VPWR.n2335 VGND 0.08351f
C20841 VPWR.n2336 VGND 0.13913f
C20842 VPWR.n2337 VGND 0.01797f
C20843 VPWR.n2338 VGND 0.00728f
C20844 VPWR.n2339 VGND 0.10822f
C20845 VPWR.t352 VGND 0.11957f
C20846 VPWR.t374 VGND 0.07849f
C20847 VPWR.t555 VGND 0.09218f
C20848 VPWR.t1216 VGND 0.07849f
C20849 VPWR.t285 VGND 0.11957f
C20850 VPWR.n2340 VGND 0.10822f
C20851 VPWR.n2341 VGND 0.00728f
C20852 VPWR.n2342 VGND 0.01797f
C20853 VPWR.n2343 VGND 0.13913f
C20854 VPWR.n2344 VGND 0.08351f
C20855 VPWR.n2345 VGND 0.08351f
C20856 VPWR.n2346 VGND 0.13913f
C20857 VPWR.n2347 VGND 0.01797f
C20858 VPWR.n2348 VGND 0.00728f
C20859 VPWR.n2349 VGND 0.10822f
C20860 VPWR.t135 VGND 0.11957f
C20861 VPWR.t452 VGND 0.07849f
C20862 VPWR.t904 VGND 0.09218f
C20863 VPWR.t1854 VGND 0.07849f
C20864 VPWR.t896 VGND 0.11957f
C20865 VPWR.n2350 VGND 0.10822f
C20866 VPWR.n2351 VGND 0.00728f
C20867 VPWR.n2352 VGND 0.01797f
C20868 VPWR.n2353 VGND 0.13913f
C20869 VPWR.n2354 VGND 0.08351f
C20870 VPWR.n2355 VGND 0.08351f
C20871 VPWR.n2356 VGND 0.13913f
C20872 VPWR.n2357 VGND 0.01797f
C20873 VPWR.n2358 VGND 0.00728f
C20874 VPWR.n2359 VGND 0.10822f
C20875 VPWR.t1217 VGND 0.11957f
C20876 VPWR.t377 VGND 0.07849f
C20877 VPWR.t1185 VGND 0.09218f
C20878 VPWR.t449 VGND 0.07849f
C20879 VPWR.t1193 VGND 0.11957f
C20880 VPWR.n2360 VGND 0.10822f
C20881 VPWR.n2361 VGND 0.00728f
C20882 VPWR.n2362 VGND 0.01797f
C20883 VPWR.n2363 VGND 0.13913f
C20884 VPWR.n2364 VGND 0.08351f
C20885 VPWR.n2365 VGND 0.08351f
C20886 VPWR.n2366 VGND 0.13913f
C20887 VPWR.n2367 VGND 0.01797f
C20888 VPWR.n2368 VGND 0.00728f
C20889 VPWR.n2369 VGND 0.10822f
C20890 VPWR.t1211 VGND 0.11957f
C20891 VPWR.t1858 VGND 0.07849f
C20892 VPWR.t666 VGND 0.09218f
C20893 VPWR.t1857 VGND 0.07849f
C20894 VPWR.t324 VGND 0.11957f
C20895 VPWR.n2370 VGND 0.10822f
C20896 VPWR.n2371 VGND 0.00728f
C20897 VPWR.n2372 VGND 0.01797f
C20898 VPWR.n2373 VGND 0.13913f
C20899 VPWR.n2374 VGND 0.08351f
C20900 VPWR.n2375 VGND 0.08351f
C20901 VPWR.n2376 VGND 0.13913f
C20902 VPWR.n2377 VGND 0.01797f
C20903 VPWR.n2378 VGND 0.00728f
C20904 VPWR.n2379 VGND 0.10822f
C20905 VPWR.t342 VGND 0.11957f
C20906 VPWR.t1215 VGND 0.07849f
C20907 VPWR.t1560 VGND 0.13333f
C20908 VPWR.n2380 VGND 0.07618f
C20909 VPWR.n2381 VGND 0.01797f
C20910 VPWR.n2382 VGND 0.13913f
C20911 VPWR.n2383 VGND 0.19371f
C20912 VPWR.n2384 VGND 1.01577f
C20913 VPWR.n2385 VGND 0.08351f
C20914 VPWR.n2386 VGND 0.08351f
C20915 VPWR.n2387 VGND 0.08351f
C20916 VPWR.n2388 VGND 0.08351f
C20917 VPWR.n2389 VGND 0.08351f
C20918 VPWR.n2390 VGND 0.08351f
C20919 VPWR.n2391 VGND 0.08351f
C20920 VPWR.n2392 VGND 0.08351f
C20921 VPWR.n2393 VGND 0.08351f
C20922 VPWR.n2394 VGND 0.08351f
C20923 VPWR.n2395 VGND 0.08351f
C20924 VPWR.n2396 VGND 0.08351f
C20925 VPWR.n2397 VGND 0.08351f
C20926 VPWR.n2398 VGND 0.08351f
C20927 VPWR.n2399 VGND 0.08351f
C20928 VPWR.n2400 VGND 0.19371f
C20929 VPWR.n2401 VGND 1.01577f
C20930 VPWR.n2402 VGND 1.01577f
C20931 VPWR.n2403 VGND 0.19371f
C20932 VPWR.n2404 VGND 0.13913f
C20933 VPWR.n2405 VGND 0.01797f
C20934 VPWR.n2406 VGND 0.07618f
C20935 VPWR.t1730 VGND 0.13333f
C20936 VPWR.t1352 VGND 0.07849f
C20937 VPWR.t191 VGND 0.11957f
C20938 VPWR.n2407 VGND 0.10822f
C20939 VPWR.n2408 VGND 0.00728f
C20940 VPWR.n2409 VGND 0.01797f
C20941 VPWR.n2410 VGND 0.13913f
C20942 VPWR.n2411 VGND 0.08351f
C20943 VPWR.n2412 VGND 0.08351f
C20944 VPWR.n2413 VGND 0.13913f
C20945 VPWR.n2414 VGND 0.01797f
C20946 VPWR.n2415 VGND 0.00728f
C20947 VPWR.n2416 VGND 0.10822f
C20948 VPWR.t330 VGND 0.09218f
C20949 VPWR.t818 VGND 0.07849f
C20950 VPWR.t102 VGND 0.11957f
C20951 VPWR.n2417 VGND 0.10822f
C20952 VPWR.n2418 VGND 0.00728f
C20953 VPWR.n2419 VGND 0.01797f
C20954 VPWR.n2420 VGND 0.13913f
C20955 VPWR.n2421 VGND 0.08351f
C20956 VPWR.n2422 VGND 0.08351f
C20957 VPWR.n2423 VGND 0.13913f
C20958 VPWR.n2424 VGND 0.01797f
C20959 VPWR.n2425 VGND 0.00728f
C20960 VPWR.n2426 VGND 0.10822f
C20961 VPWR.t1852 VGND 0.09218f
C20962 VPWR.t200 VGND 0.07849f
C20963 VPWR.t133 VGND 0.11957f
C20964 VPWR.n2427 VGND 0.10822f
C20965 VPWR.n2428 VGND 0.00728f
C20966 VPWR.n2429 VGND 0.01797f
C20967 VPWR.n2430 VGND 0.13913f
C20968 VPWR.n2431 VGND 0.08351f
C20969 VPWR.n2432 VGND 0.08351f
C20970 VPWR.n2433 VGND 0.13913f
C20971 VPWR.n2434 VGND 0.01797f
C20972 VPWR.n2435 VGND 0.00728f
C20973 VPWR.n2436 VGND 0.10822f
C20974 VPWR.t1912 VGND 0.09218f
C20975 VPWR.t1860 VGND 0.07849f
C20976 VPWR.t567 VGND 0.11957f
C20977 VPWR.n2437 VGND 0.10822f
C20978 VPWR.n2438 VGND 0.00728f
C20979 VPWR.n2439 VGND 0.01797f
C20980 VPWR.n2440 VGND 0.13913f
C20981 VPWR.n2441 VGND 0.08351f
C20982 VPWR.n2442 VGND 0.08351f
C20983 VPWR.n2443 VGND 0.13913f
C20984 VPWR.n2444 VGND 0.01797f
C20985 VPWR.n2445 VGND 0.00728f
C20986 VPWR.n2446 VGND 0.10822f
C20987 VPWR.t591 VGND 0.09218f
C20988 VPWR.t1354 VGND 0.07849f
C20989 VPWR.t302 VGND 0.11957f
C20990 VPWR.n2447 VGND 0.10822f
C20991 VPWR.n2448 VGND 0.00728f
C20992 VPWR.n2449 VGND 0.01797f
C20993 VPWR.n2450 VGND 0.13913f
C20994 VPWR.n2451 VGND 0.08351f
C20995 VPWR.n2452 VGND 0.08351f
C20996 VPWR.n2453 VGND 0.13913f
C20997 VPWR.n2454 VGND 0.01797f
C20998 VPWR.n2455 VGND 0.00728f
C20999 VPWR.n2456 VGND 0.10822f
C21000 VPWR.t277 VGND 0.09218f
C21001 VPWR.t1859 VGND 0.07849f
C21002 VPWR.t614 VGND 0.11957f
C21003 VPWR.n2457 VGND 0.10822f
C21004 VPWR.n2458 VGND 0.00728f
C21005 VPWR.n2459 VGND 0.01797f
C21006 VPWR.n2460 VGND 0.13913f
C21007 VPWR.n2461 VGND 0.08351f
C21008 VPWR.n2462 VGND 0.08351f
C21009 VPWR.n2463 VGND 0.13913f
C21010 VPWR.n2464 VGND 0.01797f
C21011 VPWR.n2465 VGND 0.00728f
C21012 VPWR.n2466 VGND 0.10822f
C21013 VPWR.t1053 VGND 0.09218f
C21014 VPWR.t202 VGND 0.07849f
C21015 VPWR.t744 VGND 0.11957f
C21016 VPWR.n2467 VGND 0.10822f
C21017 VPWR.n2468 VGND 0.00728f
C21018 VPWR.n2469 VGND 0.01797f
C21019 VPWR.n2470 VGND 0.13913f
C21020 VPWR.n2471 VGND 0.08351f
C21021 VPWR.n2472 VGND 0.08351f
C21022 VPWR.n2473 VGND 0.13913f
C21023 VPWR.n2474 VGND 0.01797f
C21024 VPWR.n2475 VGND 0.00728f
C21025 VPWR.n2476 VGND 0.10822f
C21026 VPWR.t57 VGND 0.09218f
C21027 VPWR.t1861 VGND 0.07849f
C21028 VPWR.t161 VGND 0.11957f
C21029 VPWR.n2477 VGND 0.10822f
C21030 VPWR.n2478 VGND 0.00728f
C21031 VPWR.n2479 VGND 0.01797f
C21032 VPWR.n2480 VGND 0.13913f
C21033 VPWR.n2481 VGND 0.08351f
C21034 VPWR.n2482 VGND 1.0094f
C21035 VPWR.n2483 VGND 0.19371f
C21036 VPWR.n2484 VGND 0.08351f
C21037 VPWR.n2485 VGND 0.08351f
C21038 VPWR.n2486 VGND 0.08351f
C21039 VPWR.n2487 VGND 0.08351f
C21040 VPWR.n2488 VGND 0.08351f
C21041 VPWR.n2489 VGND 0.08351f
C21042 VPWR.n2490 VGND 0.08351f
C21043 VPWR.n2491 VGND 0.08351f
C21044 VPWR.n2492 VGND 0.08351f
C21045 VPWR.n2493 VGND 0.08351f
C21046 VPWR.n2494 VGND 0.08351f
C21047 VPWR.n2495 VGND 0.08351f
C21048 VPWR.n2496 VGND 0.08351f
C21049 VPWR.n2497 VGND 0.08351f
C21050 VPWR.n2498 VGND 0.08351f
C21051 VPWR.n2499 VGND 1.0094f
C21052 VPWR.n2500 VGND 0.5713f
C21053 VPWR.n2501 VGND 0.08351f
C21054 VPWR.n2502 VGND 0.08654f
C21055 VPWR.n2503 VGND 0.00805f
C21056 VPWR.n2504 VGND 0.01714f
C21057 VPWR.n2505 VGND 0.00725f
C21058 VPWR.n2506 VGND 0.10822f
C21059 VPWR.t1609 VGND 0.11957f
C21060 VPWR.t1576 VGND 0.07849f
C21061 VPWR.t1700 VGND 0.09218f
C21062 VPWR.t1706 VGND 0.07849f
C21063 VPWR.t1721 VGND 0.11957f
C21064 VPWR.n2507 VGND 0.10822f
C21065 VPWR.n2508 VGND 0.00725f
C21066 VPWR.n2509 VGND 0.01714f
C21067 VPWR.n2510 VGND 0.00805f
C21068 VPWR.n2511 VGND 0.08654f
C21069 VPWR.n2512 VGND 0.08351f
C21070 VPWR.n2513 VGND 0.08351f
C21071 VPWR.n2514 VGND 0.08654f
C21072 VPWR.n2515 VGND 0.00805f
C21073 VPWR.n2516 VGND 0.01714f
C21074 VPWR.n2517 VGND 0.00725f
C21075 VPWR.n2518 VGND 0.10822f
C21076 VPWR.t1486 VGND 0.11957f
C21077 VPWR.t1746 VGND 0.07849f
C21078 VPWR.t1480 VGND 0.09218f
C21079 VPWR.t1470 VGND 0.07849f
C21080 VPWR.t1594 VGND 0.11957f
C21081 VPWR.n2519 VGND 0.10822f
C21082 VPWR.n2520 VGND 0.00725f
C21083 VPWR.n2521 VGND 0.01714f
C21084 VPWR.n2522 VGND 0.00805f
C21085 VPWR.n2523 VGND 0.08654f
C21086 VPWR.n2524 VGND 0.08351f
C21087 VPWR.n2525 VGND 0.08351f
C21088 VPWR.n2526 VGND 0.08654f
C21089 VPWR.n2527 VGND 0.00805f
C21090 VPWR.n2528 VGND 0.01714f
C21091 VPWR.n2529 VGND 0.00725f
C21092 VPWR.n2530 VGND 0.10822f
C21093 VPWR.t1606 VGND 0.11957f
C21094 VPWR.t1614 VGND 0.07849f
C21095 VPWR.t1743 VGND 0.09218f
C21096 VPWR.t1638 VGND 0.07849f
C21097 VPWR.t1762 VGND 0.11957f
C21098 VPWR.n2531 VGND 0.10822f
C21099 VPWR.n2532 VGND 0.00725f
C21100 VPWR.n2533 VGND 0.01714f
C21101 VPWR.n2534 VGND 0.00805f
C21102 VPWR.n2535 VGND 0.08654f
C21103 VPWR.n2536 VGND 0.08351f
C21104 VPWR.n2537 VGND 0.08351f
C21105 VPWR.n2538 VGND 0.08654f
C21106 VPWR.n2539 VGND 0.00805f
C21107 VPWR.n2540 VGND 0.01714f
C21108 VPWR.n2541 VGND 0.00725f
C21109 VPWR.n2542 VGND 0.10822f
C21110 VPWR.t1483 VGND 0.11957f
C21111 VPWR.t1475 VGND 0.07849f
C21112 VPWR.t1502 VGND 0.09218f
C21113 VPWR.t1510 VGND 0.07849f
C21114 VPWR.t1643 VGND 0.11957f
C21115 VPWR.n2543 VGND 0.10822f
C21116 VPWR.n2544 VGND 0.00725f
C21117 VPWR.n2545 VGND 0.01714f
C21118 VPWR.n2546 VGND 0.00805f
C21119 VPWR.n2547 VGND 0.08654f
C21120 VPWR.n2548 VGND 0.08351f
C21121 VPWR.n2549 VGND 0.08351f
C21122 VPWR.n2550 VGND 0.08654f
C21123 VPWR.n2551 VGND 0.00805f
C21124 VPWR.n2552 VGND 0.01714f
C21125 VPWR.n2553 VGND 0.00725f
C21126 VPWR.n2554 VGND 0.10822f
C21127 VPWR.t1659 VGND 0.11957f
C21128 VPWR.t1612 VGND 0.07849f
C21129 VPWR.t1740 VGND 0.09218f
C21130 VPWR.t1773 VGND 0.07849f
C21131 VPWR.t1789 VGND 0.11957f
C21132 VPWR.n2555 VGND 0.10822f
C21133 VPWR.n2556 VGND 0.00725f
C21134 VPWR.n2557 VGND 0.01714f
C21135 VPWR.n2558 VGND 0.00805f
C21136 VPWR.n2559 VGND 0.08654f
C21137 VPWR.n2560 VGND 0.08351f
C21138 VPWR.n2561 VGND 0.08351f
C21139 VPWR.n2562 VGND 0.08654f
C21140 VPWR.n2563 VGND 0.00805f
C21141 VPWR.n2564 VGND 0.01714f
C21142 VPWR.n2565 VGND 0.00725f
C21143 VPWR.n2566 VGND 0.10822f
C21144 VPWR.t1533 VGND 0.11957f
C21145 VPWR.t1792 VGND 0.07849f
C21146 VPWR.t1525 VGND 0.09218f
C21147 VPWR.t1646 VGND 0.07849f
C21148 VPWR.t1563 VGND 0.11957f
C21149 VPWR.n2567 VGND 0.10822f
C21150 VPWR.n2568 VGND 0.00725f
C21151 VPWR.n2569 VGND 0.01714f
C21152 VPWR.n2570 VGND 0.00805f
C21153 VPWR.n2571 VGND 0.08654f
C21154 VPWR.n2572 VGND 0.08351f
C21155 VPWR.n2573 VGND 0.08351f
C21156 VPWR.n2574 VGND 0.08654f
C21157 VPWR.n2575 VGND 0.00805f
C21158 VPWR.n2576 VGND 0.01714f
C21159 VPWR.n2577 VGND 0.00725f
C21160 VPWR.n2578 VGND 0.10822f
C21161 VPWR.t1413 VGND 0.11957f
C21162 VPWR.t1665 VGND 0.07849f
C21163 VPWR.t1786 VGND 0.09218f
C21164 VPWR.t1690 VGND 0.07849f
C21165 VPWR.t1432 VGND 0.11957f
C21166 VPWR.n2579 VGND 0.10822f
C21167 VPWR.n2580 VGND 0.00725f
C21168 VPWR.n2581 VGND 0.01714f
C21169 VPWR.n2582 VGND 0.00805f
C21170 VPWR.n2583 VGND 0.08654f
C21171 VPWR.n2584 VGND 0.08351f
C21172 VPWR.n2585 VGND 0.08351f
C21173 VPWR.n2586 VGND 0.08654f
C21174 VPWR.n2587 VGND 0.00805f
C21175 VPWR.n2588 VGND 0.01714f
C21176 VPWR.n2589 VGND 0.00725f
C21177 VPWR.n2590 VGND 0.10822f
C21178 VPWR.t1557 VGND 0.11957f
C21179 VPWR.t1541 VGND 0.07849f
C21180 VPWR.t1662 VGND 0.13333f
C21181 VPWR.n2591 VGND 0.07615f
C21182 VPWR.n2592 VGND 0.01698f
C21183 VPWR.n2593 VGND 0.00805f
C21184 VPWR.n2594 VGND 0.10853f
C21185 VPWR.n2595 VGND 0.19371f
C21186 VPWR.n2596 VGND 2.66265f
C21187 VPWR.n2597 VGND 1.08435f
C21188 VPWR.n2598 VGND 0.45434f
C21189 VPWR.t1135 VGND 0.05456f
C21190 VPWR.t805 VGND 0.05456f
C21191 VPWR.n2599 VGND 0.09898f
C21192 VPWR.n2600 VGND 0.04687f
C21193 VPWR.t1134 VGND 0.01433f
C21194 VPWR.t1138 VGND 0.01433f
C21195 VPWR.n2601 VGND 0.03076f
C21196 VPWR.t815 VGND 0.01433f
C21197 VPWR.t803 VGND 0.01433f
C21198 VPWR.n2602 VGND 0.03076f
C21199 VPWR.n2603 VGND 0.01064f
C21200 VPWR.n2604 VGND 0.04687f
C21201 VPWR.t90 VGND 0.01433f
C21202 VPWR.t886 VGND 0.01433f
C21203 VPWR.n2605 VGND 0.03076f
C21204 VPWR.t915 VGND 0.01433f
C21205 VPWR.t910 VGND 0.01433f
C21206 VPWR.n2606 VGND 0.03076f
C21207 VPWR.t924 VGND 0.05714f
C21208 VPWR.t1844 VGND 0.05714f
C21209 VPWR.n2607 VGND 0.13176f
C21210 VPWR.n2608 VGND 0.04228f
C21211 VPWR.n2609 VGND 0.01362f
C21212 VPWR.n2610 VGND 0.06183f
C21213 VPWR.n2611 VGND 0.0092f
C21214 VPWR.t1843 VGND 0.01433f
C21215 VPWR.t1137 VGND 0.01433f
C21216 VPWR.n2612 VGND 0.03076f
C21217 VPWR.t926 VGND 0.01433f
C21218 VPWR.t811 VGND 0.01433f
C21219 VPWR.n2613 VGND 0.03076f
C21220 VPWR.n2614 VGND 0.06183f
C21221 VPWR.n2615 VGND 0.01425f
C21222 VPWR.n2616 VGND 0.04687f
C21223 VPWR.n2617 VGND 0.04687f
C21224 VPWR.n2618 VGND 0.04687f
C21225 VPWR.n2619 VGND 0.01281f
C21226 VPWR.n2620 VGND 0.06183f
C21227 VPWR.n2621 VGND 0.01209f
C21228 VPWR.n2622 VGND 0.00983f
C21229 VPWR.n2623 VGND 0.04687f
C21230 VPWR.n2624 VGND 0.03515f
C21231 VPWR.n2625 VGND 0.00794f
C21232 VPWR.t923 VGND 0.1712f
C21233 VPWR.t89 VGND 0.25229f
C21234 VPWR.t885 VGND 0.25229f
C21235 VPWR.t925 VGND 0.25229f
C21236 VPWR.t810 VGND 0.25229f
C21237 VPWR.t814 VGND 0.25229f
C21238 VPWR.t802 VGND 0.25229f
C21239 VPWR.t804 VGND 0.56168f
C21240 VPWR.n2626 VGND 0.61307f
C21241 VPWR.n2627 VGND 0.01783f
C21242 VPWR.n2628 VGND 1.07531f
C21243 VPWR.n2629 VGND 0.04687f
C21244 VPWR.t84 VGND 0.1712f
C21245 VPWR.t880 VGND 0.25229f
C21246 VPWR.t1326 VGND 0.25229f
C21247 VPWR.t82 VGND 0.25229f
C21248 VPWR.t967 VGND 0.25229f
C21249 VPWR.t959 VGND 0.25229f
C21250 VPWR.t971 VGND 0.25229f
C21251 VPWR.t963 VGND 0.41448f
C21252 VPWR.t514 VGND 0.44001f
C21253 VPWR.n2630 VGND 0.62092f
C21254 VPWR.n2631 VGND 0.17663f
C21255 VPWR.n2632 VGND 0.04687f
C21256 VPWR.t1399 VGND 0.01433f
C21257 VPWR.t1395 VGND 0.01433f
C21258 VPWR.n2633 VGND 0.03076f
C21259 VPWR.t960 VGND 0.01433f
C21260 VPWR.t972 VGND 0.01433f
C21261 VPWR.n2634 VGND 0.03076f
C21262 VPWR.n2635 VGND 0.06183f
C21263 VPWR.n2636 VGND 0.04687f
C21264 VPWR.t83 VGND 0.01433f
C21265 VPWR.t1394 VGND 0.01433f
C21266 VPWR.n2637 VGND 0.03076f
C21267 VPWR.t1922 VGND 0.01433f
C21268 VPWR.t968 VGND 0.01433f
C21269 VPWR.n2638 VGND 0.03076f
C21270 VPWR.n2639 VGND 0.0092f
C21271 VPWR.t1845 VGND 0.05714f
C21272 VPWR.t85 VGND 0.05714f
C21273 VPWR.n2640 VGND 0.13176f
C21274 VPWR.t881 VGND 0.01433f
C21275 VPWR.t1842 VGND 0.01433f
C21276 VPWR.n2641 VGND 0.03076f
C21277 VPWR.t913 VGND 0.01433f
C21278 VPWR.t1327 VGND 0.01433f
C21279 VPWR.n2642 VGND 0.03076f
C21280 VPWR.n2643 VGND 0.06183f
C21281 VPWR.n2644 VGND 0.01362f
C21282 VPWR.n2645 VGND 0.04228f
C21283 VPWR.n2646 VGND 0.04687f
C21284 VPWR.n2647 VGND 0.04687f
C21285 VPWR.n2648 VGND 0.01425f
C21286 VPWR.n2649 VGND 0.06183f
C21287 VPWR.n2650 VGND 0.01064f
C21288 VPWR.n2651 VGND 0.01281f
C21289 VPWR.n2652 VGND 0.04687f
C21290 VPWR.n2653 VGND 0.04687f
C21291 VPWR.n2654 VGND 0.01209f
C21292 VPWR.n2655 VGND 0.00983f
C21293 VPWR.t1400 VGND 0.05456f
C21294 VPWR.t964 VGND 0.05456f
C21295 VPWR.n2656 VGND 0.09898f
C21296 VPWR.n2657 VGND 0.00794f
C21297 VPWR.n2658 VGND 0.03515f
C21298 VPWR.n2659 VGND 0.01783f
C21299 VPWR.n2660 VGND 0.03515f
C21300 VPWR.n2661 VGND 0.01398f
C21301 VPWR.n2662 VGND 0.01083f
C21302 VPWR.t628 VGND 0.05708f
C21303 VPWR.t515 VGND 0.05708f
C21304 VPWR.n2663 VGND 0.11537f
C21305 VPWR.n2664 VGND 0.03261f
C21306 VPWR.n2665 VGND 1.63658f
C21307 VPWR.n2666 VGND 0.04687f
C21308 VPWR.t1283 VGND 0.05603f
C21309 VPWR.t86 VGND 0.1712f
C21310 VPWR.t17 VGND 0.25229f
C21311 VPWR.t1828 VGND 0.25229f
C21312 VPWR.t930 VGND 0.25229f
C21313 VPWR.t1130 VGND 0.25229f
C21314 VPWR.t782 VGND 0.25229f
C21315 VPWR.t372 VGND 0.25229f
C21316 VPWR.t1142 VGND 0.41448f
C21317 VPWR.t460 VGND 0.15918f
C21318 VPWR.t1282 VGND 0.12614f
C21319 VPWR.t563 VGND 0.28082f
C21320 VPWR.n2667 VGND 0.55034f
C21321 VPWR.n2668 VGND 0.17401f
C21322 VPWR.n2669 VGND 0.04687f
C21323 VPWR.t1903 VGND 0.01433f
C21324 VPWR.t1907 VGND 0.01433f
C21325 VPWR.n2670 VGND 0.03076f
C21326 VPWR.t783 VGND 0.01433f
C21327 VPWR.t373 VGND 0.01433f
C21328 VPWR.n2671 VGND 0.03076f
C21329 VPWR.n2672 VGND 0.06183f
C21330 VPWR.n2673 VGND 0.04687f
C21331 VPWR.t1925 VGND 0.01433f
C21332 VPWR.t1906 VGND 0.01433f
C21333 VPWR.n2674 VGND 0.03076f
C21334 VPWR.t931 VGND 0.01433f
C21335 VPWR.t1131 VGND 0.01433f
C21336 VPWR.n2675 VGND 0.03076f
C21337 VPWR.n2676 VGND 0.0092f
C21338 VPWR.t87 VGND 0.05714f
C21339 VPWR.t878 VGND 0.05714f
C21340 VPWR.n2677 VGND 0.13176f
C21341 VPWR.t914 VGND 0.01433f
C21342 VPWR.t1829 VGND 0.01433f
C21343 VPWR.n2678 VGND 0.03076f
C21344 VPWR.t18 VGND 0.01433f
C21345 VPWR.t1921 VGND 0.01433f
C21346 VPWR.n2679 VGND 0.03076f
C21347 VPWR.n2680 VGND 0.06183f
C21348 VPWR.n2681 VGND 0.01362f
C21349 VPWR.n2682 VGND 0.04228f
C21350 VPWR.n2683 VGND 0.04687f
C21351 VPWR.n2684 VGND 0.04687f
C21352 VPWR.n2685 VGND 0.01425f
C21353 VPWR.n2686 VGND 0.06183f
C21354 VPWR.n2687 VGND 0.01064f
C21355 VPWR.n2688 VGND 0.01281f
C21356 VPWR.n2689 VGND 0.04687f
C21357 VPWR.n2690 VGND 0.04687f
C21358 VPWR.n2691 VGND 0.01209f
C21359 VPWR.n2692 VGND 0.00983f
C21360 VPWR.t1904 VGND 0.05456f
C21361 VPWR.t1143 VGND 0.05456f
C21362 VPWR.n2693 VGND 0.09898f
C21363 VPWR.n2694 VGND 0.00794f
C21364 VPWR.n2695 VGND 0.03515f
C21365 VPWR.n2696 VGND 0.01783f
C21366 VPWR.n2697 VGND 0.03515f
C21367 VPWR.t564 VGND 0.05714f
C21368 VPWR.n2698 VGND 0.07963f
C21369 VPWR.n2699 VGND 0.01064f
C21370 VPWR.n2700 VGND 0.05827f
C21371 VPWR.t461 VGND 0.05618f
C21372 VPWR.n2701 VGND 0.07281f
C21373 VPWR.n2702 VGND 0.02776f
C21374 VPWR.n2703 VGND 1.63658f
C21375 VPWR.n2704 VGND 0.04687f
C21376 VPWR.t1923 VGND 0.09709f
C21377 VPWR.t14 VGND 0.14308f
C21378 VPWR.t1919 VGND 0.1391f
C21379 VPWR.t928 VGND 0.22247f
C21380 VPWR.t1108 VGND 0.18922f
C21381 VPWR.t920 VGND 0.12614f
C21382 VPWR.t867 VGND 0.12614f
C21383 VPWR.t11 VGND 0.12614f
C21384 VPWR.t1106 VGND 0.12614f
C21385 VPWR.t882 VGND 0.12614f
C21386 VPWR.t1112 VGND 0.12614f
C21387 VPWR.t1830 VGND 0.1757f
C21388 VPWR.t228 VGND 0.09911f
C21389 VPWR.t994 VGND 0.10812f
C21390 VPWR.t821 VGND 0.12614f
C21391 VPWR.t996 VGND 0.23427f
C21392 VPWR.n2705 VGND 0.37764f
C21393 VPWR.n2706 VGND 0.17419f
C21394 VPWR.t997 VGND 0.05672f
C21395 VPWR.n2707 VGND 0.04687f
C21396 VPWR.t1831 VGND 0.05606f
C21397 VPWR.t1113 VGND 0.05397f
C21398 VPWR.t12 VGND 0.01433f
C21399 VPWR.t883 VGND 0.01433f
C21400 VPWR.n2708 VGND 0.03076f
C21401 VPWR.t868 VGND 0.01433f
C21402 VPWR.t1107 VGND 0.01433f
C21403 VPWR.n2709 VGND 0.03076f
C21404 VPWR.n2710 VGND 0.03507f
C21405 VPWR.n2711 VGND 0.04687f
C21406 VPWR.t929 VGND 0.01433f
C21407 VPWR.t1109 VGND 0.01433f
C21408 VPWR.n2712 VGND 0.03076f
C21409 VPWR.n2713 VGND 0.0092f
C21410 VPWR.t1924 VGND 0.05714f
C21411 VPWR.n2714 VGND 0.072f
C21412 VPWR.t15 VGND 0.01433f
C21413 VPWR.t1920 VGND 0.01433f
C21414 VPWR.n2715 VGND 0.03076f
C21415 VPWR.n2716 VGND 0.03507f
C21416 VPWR.n2717 VGND 0.01362f
C21417 VPWR.n2718 VGND 0.04228f
C21418 VPWR.n2719 VGND 0.04687f
C21419 VPWR.n2720 VGND 0.04687f
C21420 VPWR.n2721 VGND 0.01425f
C21421 VPWR.n2722 VGND 0.03425f
C21422 VPWR.t921 VGND 0.05015f
C21423 VPWR.n2723 VGND 0.03998f
C21424 VPWR.n2724 VGND 0.00983f
C21425 VPWR.n2725 VGND 0.04687f
C21426 VPWR.n2726 VGND 0.04687f
C21427 VPWR.n2727 VGND 0.03885f
C21428 VPWR.n2728 VGND 0.01209f
C21429 VPWR.n2729 VGND 0.05142f
C21430 VPWR.n2730 VGND 0.06775f
C21431 VPWR.n2731 VGND 0.00622f
C21432 VPWR.n2732 VGND 0.02776f
C21433 VPWR.n2733 VGND 0.01783f
C21434 VPWR.n2734 VGND 0.03515f
C21435 VPWR.t822 VGND 0.0572f
C21436 VPWR.n2735 VGND 0.14706f
C21437 VPWR.n2736 VGND 0.01083f
C21438 VPWR.t995 VGND 0.05711f
C21439 VPWR.n2737 VGND 0.06357f
C21440 VPWR.n2738 VGND 0.02751f
C21441 VPWR.n2739 VGND 1.63658f
C21442 VPWR.n2740 VGND 0.04228f
C21443 VPWR.t879 VGND 0.66677f
C21444 VPWR.t1324 VGND 0.25229f
C21445 VPWR.t927 VGND 0.25229f
C21446 VPWR.t13 VGND 0.25229f
C21447 VPWR.t808 VGND 0.25229f
C21448 VPWR.t806 VGND 0.25229f
C21449 VPWR.t812 VGND 0.25229f
C21450 VPWR.t800 VGND 0.22826f
C21451 VPWR.t29 VGND 0.55264f
C21452 VPWR.t1405 VGND 0.15318f
C21453 VPWR.n2741 VGND 0.33109f
C21454 VPWR.n2742 VGND 0.17663f
C21455 VPWR.t1139 VGND 0.01433f
C21456 VPWR.t1136 VGND 0.01433f
C21457 VPWR.n2743 VGND 0.03141f
C21458 VPWR.t809 VGND 0.01433f
C21459 VPWR.t807 VGND 0.01433f
C21460 VPWR.n2744 VGND 0.03141f
C21461 VPWR.n2745 VGND 0.1192f
C21462 VPWR.n2746 VGND 0.09664f
C21463 VPWR.t1140 VGND 0.01433f
C21464 VPWR.t1141 VGND 0.01433f
C21465 VPWR.n2747 VGND 0.03146f
C21466 VPWR.t813 VGND 0.01433f
C21467 VPWR.t801 VGND 0.01433f
C21468 VPWR.n2748 VGND 0.03146f
C21469 VPWR.n2749 VGND 0.13065f
C21470 VPWR.n2750 VGND 0.01119f
C21471 VPWR.n2751 VGND 0.37741f
C21472 VPWR.n2752 VGND 0.01783f
C21473 VPWR.n2753 VGND 0.0163f
C21474 VPWR.n2754 VGND 0.01398f
C21475 VPWR.n2755 VGND 0.01308f
C21476 VPWR.t30 VGND 0.0572f
C21477 VPWR.t1917 VGND 0.0572f
C21478 VPWR.n2756 VGND 0.16894f
C21479 VPWR.n2757 VGND 0.03515f
C21480 VPWR.n2758 VGND 1.63658f
C21481 VPWR.n2759 VGND 0.04228f
C21482 VPWR.t911 VGND 0.66677f
C21483 VPWR.t1918 VGND 0.25229f
C21484 VPWR.t10 VGND 0.25229f
C21485 VPWR.t91 VGND 0.25229f
C21486 VPWR.t957 VGND 0.25229f
C21487 VPWR.t969 VGND 0.25229f
C21488 VPWR.t961 VGND 0.25229f
C21489 VPWR.t965 VGND 0.22826f
C21490 VPWR.t27 VGND 0.49107f
C21491 VPWR.t1407 VGND 0.10812f
C21492 VPWR.t1411 VGND 0.10662f
C21493 VPWR.n2760 VGND 0.32959f
C21494 VPWR.n2761 VGND 0.17663f
C21495 VPWR.t1396 VGND 0.01433f
C21496 VPWR.t1401 VGND 0.01433f
C21497 VPWR.n2762 VGND 0.03141f
C21498 VPWR.t958 VGND 0.01433f
C21499 VPWR.t970 VGND 0.01433f
C21500 VPWR.n2763 VGND 0.03141f
C21501 VPWR.n2764 VGND 0.1192f
C21502 VPWR.n2765 VGND 0.09664f
C21503 VPWR.t1397 VGND 0.01433f
C21504 VPWR.t1398 VGND 0.01433f
C21505 VPWR.n2766 VGND 0.03146f
C21506 VPWR.t962 VGND 0.01433f
C21507 VPWR.t966 VGND 0.01433f
C21508 VPWR.n2767 VGND 0.03146f
C21509 VPWR.n2768 VGND 0.13065f
C21510 VPWR.n2769 VGND 0.01119f
C21511 VPWR.n2770 VGND 0.37741f
C21512 VPWR.n2771 VGND 0.01783f
C21513 VPWR.n2772 VGND 0.01605f
C21514 VPWR.n2773 VGND 0.00767f
C21515 VPWR.t1408 VGND 0.05708f
C21516 VPWR.n2774 VGND 0.06101f
C21517 VPWR.n2775 VGND 0.00731f
C21518 VPWR.t28 VGND 0.0572f
C21519 VPWR.n2776 VGND 0.0911f
C21520 VPWR.n2777 VGND 0.03515f
C21521 VPWR.n2778 VGND 1.63658f
C21522 VPWR.n2779 VGND 0.04279f
C21523 VPWR.t16 VGND 0.66677f
C21524 VPWR.t922 VGND 0.25229f
C21525 VPWR.t88 VGND 0.25229f
C21526 VPWR.t884 VGND 0.25229f
C21527 VPWR.t659 VGND 0.25229f
C21528 VPWR.t405 VGND 0.25229f
C21529 VPWR.t1132 VGND 0.25229f
C21530 VPWR.t1128 VGND 0.22826f
C21531 VPWR.t31 VGND 0.5226f
C21532 VPWR.t1403 VGND 0.18021f
C21533 VPWR.n2780 VGND 0.32809f
C21534 VPWR.n2781 VGND 0.17401f
C21535 VPWR.t1406 VGND 0.05716f
C21536 VPWR.t1908 VGND 0.01433f
C21537 VPWR.t1905 VGND 0.01433f
C21538 VPWR.n2782 VGND 0.03141f
C21539 VPWR.t660 VGND 0.01433f
C21540 VPWR.t406 VGND 0.01433f
C21541 VPWR.n2783 VGND 0.03141f
C21542 VPWR.n2784 VGND 0.1192f
C21543 VPWR.n2785 VGND 0.09664f
C21544 VPWR.t1901 VGND 0.01433f
C21545 VPWR.t1902 VGND 0.01433f
C21546 VPWR.n2786 VGND 0.03146f
C21547 VPWR.t1133 VGND 0.01433f
C21548 VPWR.t1129 VGND 0.01433f
C21549 VPWR.n2787 VGND 0.03146f
C21550 VPWR.n2788 VGND 0.13065f
C21551 VPWR.n2789 VGND 0.01119f
C21552 VPWR.n2790 VGND 0.37741f
C21553 VPWR.n2791 VGND 0.01783f
C21554 VPWR.n2792 VGND 0.01579f
C21555 VPWR.t1404 VGND 0.05716f
C21556 VPWR.n2793 VGND 0.15059f
C21557 VPWR.n2794 VGND 0.01209f
C21558 VPWR.t32 VGND 0.05714f
C21559 VPWR.t1916 VGND 0.05714f
C21560 VPWR.n2795 VGND 0.13446f
C21561 VPWR.n2796 VGND 0.03515f
C21562 VPWR.n2797 VGND 1.63658f
C21563 VPWR.n2798 VGND 0.04279f
C21564 VPWR.t26 VGND 0.05714f
C21565 VPWR.n2799 VGND 0.01579f
C21566 VPWR.t1410 VGND 0.05716f
C21567 VPWR.n2800 VGND 0.01783f
C21568 VPWR.t887 VGND 0.37815f
C21569 VPWR.t81 VGND 0.14308f
C21570 VPWR.t912 VGND 0.14308f
C21571 VPWR.t1325 VGND 0.14308f
C21572 VPWR.t1110 VGND 0.14308f
C21573 VPWR.t869 VGND 0.14308f
C21574 VPWR.t1065 VGND 0.14308f
C21575 VPWR.t1063 VGND 0.12946f
C21576 VPWR.t25 VGND 0.29639f
C21577 VPWR.t1409 VGND 0.1022f
C21578 VPWR.n2801 VGND 0.1826f
C21579 VPWR.t1066 VGND 0.01433f
C21580 VPWR.t1064 VGND 0.01433f
C21581 VPWR.n2802 VGND 0.03146f
C21582 VPWR.n2803 VGND 0.07742f
C21583 VPWR.t1111 VGND 0.01433f
C21584 VPWR.t870 VGND 0.01433f
C21585 VPWR.n2804 VGND 0.03274f
C21586 VPWR.n2805 VGND 0.1748f
C21587 VPWR.n2806 VGND 0.37741f
C21588 VPWR.n2807 VGND 0.01119f
C21589 VPWR.n2808 VGND 0.09661f
C21590 VPWR.n2809 VGND 0.08481f
C21591 VPWR.n2810 VGND 0.01209f
C21592 VPWR.n2811 VGND 0.0735f
C21593 VPWR.n2812 VGND 0.03515f
C21594 VPWR.n2813 VGND 2.3816f
C21595 VPWR.n2814 VGND 1.92879f
C21596 VPWR.t517 VGND 0.02906f
C21597 VPWR.n2815 VGND 0.13023f
C21598 VPWR.n2816 VGND 0.28666f
C21599 VPWR.n2817 VGND 0.0756f
C21600 VPWR.n2818 VGND 0.0359f
C21601 VPWR.n2819 VGND 0.04384f
C21602 VPWR.n2820 VGND 0.08886f
C21603 VPWR.n2821 VGND 0.11583f
C21604 VPWR.n2822 VGND 0.08886f
C21605 VPWR.t718 VGND 2.79496f
C21606 VPWR.t516 VGND 0.88276f
C21607 VPWR.n2823 VGND 0.11674f
C21608 VPWR.n2824 VGND 0.46189f
C21609 VPWR.t719 VGND 0.02904f
C21610 VPWR.n2825 VGND 0.17782f
C21611 VPWR.n2826 VGND 0.01795f
C21612 VPWR.n2827 VGND 0.09797f
C21613 VPWR.n2828 VGND 0.08795f
C21614 VPWR.n2829 VGND 0.11674f
C21615 VPWR.n2830 VGND 0.07352f
C21616 VPWR.t1081 VGND 0.02904f
C21617 VPWR.n2831 VGND 0.17782f
C21618 VPWR.n2832 VGND 0.01795f
C21619 VPWR.n2833 VGND 0.11674f
C21620 VPWR.n2834 VGND 0.0764f
C21621 VPWR.n2835 VGND 0.08713f
C21622 VPWR.n2836 VGND 1.67029f
C21623 VPWR.n2837 VGND 0.08713f
C21624 VPWR.n2838 VGND 0.0764f
C21625 VPWR.n2839 VGND 0.11674f
C21626 VPWR.n2840 VGND 0.09788f
C21627 VPWR.n2841 VGND 0.08096f
C21628 VPWR.n2842 VGND 1.00402f
C21629 VPWR.n2843 VGND 0.06317f
C21630 VPWR.n2844 VGND 0.08837f
C21631 VPWR.n2845 VGND 0.06143f
C21632 VPWR.n2846 VGND 0.01795f
C21633 VPWR.n2847 VGND 0.06317f
C21634 VPWR.n2848 VGND 0.04851f
C21635 VPWR.n2849 VGND 0.17356f
C21636 VPWR.n2850 VGND 0.06838f
C21637 VPWR.n2851 VGND 0.04384f
C21638 VPWR.t1800 VGND 0.34561f
C21639 VPWR.n2852 VGND 0.08096f
C21640 VPWR.n2853 VGND 0.09788f
C21641 VPWR.n2854 VGND 0.0359f
C21642 VPWR.n2855 VGND 2.02287f
C21643 VPWR.n2856 VGND 0.0359f
C21644 VPWR.n2857 VGND 0.0359f
C21645 VPWR.n2858 VGND 0.08922f
C21646 VPWR.n2859 VGND 0.04898f
C21647 VPWR.n2860 VGND 0.37936f
C21648 VPWR.n2861 VGND 0.31214f
C21649 VPWR.t1801 VGND 0.02903f
C21650 VPWR.n2862 VGND 0.21967f
C21651 VPWR.n2863 VGND 3.34958f
C21652 XThR.Tn[2].t11 VGND 0.02313f
C21653 XThR.Tn[2].t10 VGND 0.02313f
C21654 XThR.Tn[2].n0 VGND 0.04668f
C21655 XThR.Tn[2].t4 VGND 0.02313f
C21656 XThR.Tn[2].t7 VGND 0.02313f
C21657 XThR.Tn[2].n1 VGND 0.05462f
C21658 XThR.Tn[2].n2 VGND 0.16384f
C21659 XThR.Tn[2].t8 VGND 0.01503f
C21660 XThR.Tn[2].t1 VGND 0.01503f
C21661 XThR.Tn[2].n3 VGND 0.05704f
C21662 XThR.Tn[2].t3 VGND 0.01503f
C21663 XThR.Tn[2].t2 VGND 0.01503f
C21664 XThR.Tn[2].n4 VGND 0.03423f
C21665 XThR.Tn[2].n5 VGND 0.16303f
C21666 XThR.Tn[2].t6 VGND 0.01503f
C21667 XThR.Tn[2].t9 VGND 0.01503f
C21668 XThR.Tn[2].n6 VGND 0.03423f
C21669 XThR.Tn[2].n7 VGND 0.10078f
C21670 XThR.Tn[2].t5 VGND 0.01503f
C21671 XThR.Tn[2].t0 VGND 0.01503f
C21672 XThR.Tn[2].n8 VGND 0.03423f
C21673 XThR.Tn[2].n9 VGND 0.11374f
C21674 XThR.Tn[2].t21 VGND 0.01808f
C21675 XThR.Tn[2].t14 VGND 0.01979f
C21676 XThR.Tn[2].n10 VGND 0.04833f
C21677 XThR.Tn[2].n11 VGND 0.09285f
C21678 XThR.Tn[2].t40 VGND 0.01808f
C21679 XThR.Tn[2].t31 VGND 0.01979f
C21680 XThR.Tn[2].n12 VGND 0.04833f
C21681 XThR.Tn[2].t55 VGND 0.01802f
C21682 XThR.Tn[2].t66 VGND 0.01973f
C21683 XThR.Tn[2].n13 VGND 0.05029f
C21684 XThR.Tn[2].n14 VGND 0.03533f
C21685 XThR.Tn[2].n15 VGND 0.00646f
C21686 XThR.Tn[2].n16 VGND 0.11337f
C21687 XThR.Tn[2].t15 VGND 0.01808f
C21688 XThR.Tn[2].t67 VGND 0.01979f
C21689 XThR.Tn[2].n17 VGND 0.04833f
C21690 XThR.Tn[2].t30 VGND 0.01802f
C21691 XThR.Tn[2].t43 VGND 0.01973f
C21692 XThR.Tn[2].n18 VGND 0.05029f
C21693 XThR.Tn[2].n19 VGND 0.03533f
C21694 XThR.Tn[2].n20 VGND 0.00646f
C21695 XThR.Tn[2].n21 VGND 0.11337f
C21696 XThR.Tn[2].t32 VGND 0.01808f
C21697 XThR.Tn[2].t23 VGND 0.01979f
C21698 XThR.Tn[2].n22 VGND 0.04833f
C21699 XThR.Tn[2].t47 VGND 0.01802f
C21700 XThR.Tn[2].t60 VGND 0.01973f
C21701 XThR.Tn[2].n23 VGND 0.05029f
C21702 XThR.Tn[2].n24 VGND 0.03533f
C21703 XThR.Tn[2].n25 VGND 0.00646f
C21704 XThR.Tn[2].n26 VGND 0.11337f
C21705 XThR.Tn[2].t58 VGND 0.01808f
C21706 XThR.Tn[2].t50 VGND 0.01979f
C21707 XThR.Tn[2].n27 VGND 0.04833f
C21708 XThR.Tn[2].t16 VGND 0.01802f
C21709 XThR.Tn[2].t28 VGND 0.01973f
C21710 XThR.Tn[2].n28 VGND 0.05029f
C21711 XThR.Tn[2].n29 VGND 0.03533f
C21712 XThR.Tn[2].n30 VGND 0.00646f
C21713 XThR.Tn[2].n31 VGND 0.11337f
C21714 XThR.Tn[2].t34 VGND 0.01808f
C21715 XThR.Tn[2].t25 VGND 0.01979f
C21716 XThR.Tn[2].n32 VGND 0.04833f
C21717 XThR.Tn[2].t48 VGND 0.01802f
C21718 XThR.Tn[2].t62 VGND 0.01973f
C21719 XThR.Tn[2].n33 VGND 0.05029f
C21720 XThR.Tn[2].n34 VGND 0.03533f
C21721 XThR.Tn[2].n35 VGND 0.00646f
C21722 XThR.Tn[2].n36 VGND 0.11337f
C21723 XThR.Tn[2].t70 VGND 0.01808f
C21724 XThR.Tn[2].t41 VGND 0.01979f
C21725 XThR.Tn[2].n37 VGND 0.04833f
C21726 XThR.Tn[2].t22 VGND 0.01802f
C21727 XThR.Tn[2].t20 VGND 0.01973f
C21728 XThR.Tn[2].n38 VGND 0.05029f
C21729 XThR.Tn[2].n39 VGND 0.03533f
C21730 XThR.Tn[2].n40 VGND 0.00646f
C21731 XThR.Tn[2].n41 VGND 0.11337f
C21732 XThR.Tn[2].t39 VGND 0.01808f
C21733 XThR.Tn[2].t35 VGND 0.01979f
C21734 XThR.Tn[2].n42 VGND 0.04833f
C21735 XThR.Tn[2].t54 VGND 0.01802f
C21736 XThR.Tn[2].t12 VGND 0.01973f
C21737 XThR.Tn[2].n43 VGND 0.05029f
C21738 XThR.Tn[2].n44 VGND 0.03533f
C21739 XThR.Tn[2].n45 VGND 0.00646f
C21740 XThR.Tn[2].n46 VGND 0.11337f
C21741 XThR.Tn[2].t44 VGND 0.01808f
C21742 XThR.Tn[2].t49 VGND 0.01979f
C21743 XThR.Tn[2].n47 VGND 0.04833f
C21744 XThR.Tn[2].t57 VGND 0.01802f
C21745 XThR.Tn[2].t27 VGND 0.01973f
C21746 XThR.Tn[2].n48 VGND 0.05029f
C21747 XThR.Tn[2].n49 VGND 0.03533f
C21748 XThR.Tn[2].n50 VGND 0.00646f
C21749 XThR.Tn[2].n51 VGND 0.11337f
C21750 XThR.Tn[2].t61 VGND 0.01808f
C21751 XThR.Tn[2].t69 VGND 0.01979f
C21752 XThR.Tn[2].n52 VGND 0.04833f
C21753 XThR.Tn[2].t18 VGND 0.01802f
C21754 XThR.Tn[2].t45 VGND 0.01973f
C21755 XThR.Tn[2].n53 VGND 0.05029f
C21756 XThR.Tn[2].n54 VGND 0.03533f
C21757 XThR.Tn[2].n55 VGND 0.00646f
C21758 XThR.Tn[2].n56 VGND 0.11337f
C21759 XThR.Tn[2].t52 VGND 0.01808f
C21760 XThR.Tn[2].t26 VGND 0.01979f
C21761 XThR.Tn[2].n57 VGND 0.04833f
C21762 XThR.Tn[2].t68 VGND 0.01802f
C21763 XThR.Tn[2].t63 VGND 0.01973f
C21764 XThR.Tn[2].n58 VGND 0.05029f
C21765 XThR.Tn[2].n59 VGND 0.03533f
C21766 XThR.Tn[2].n60 VGND 0.00646f
C21767 XThR.Tn[2].n61 VGND 0.11337f
C21768 XThR.Tn[2].t73 VGND 0.01808f
C21769 XThR.Tn[2].t64 VGND 0.01979f
C21770 XThR.Tn[2].n62 VGND 0.04833f
C21771 XThR.Tn[2].t24 VGND 0.01802f
C21772 XThR.Tn[2].t37 VGND 0.01973f
C21773 XThR.Tn[2].n63 VGND 0.05029f
C21774 XThR.Tn[2].n64 VGND 0.03533f
C21775 XThR.Tn[2].n65 VGND 0.00646f
C21776 XThR.Tn[2].n66 VGND 0.11337f
C21777 XThR.Tn[2].t42 VGND 0.01808f
C21778 XThR.Tn[2].t36 VGND 0.01979f
C21779 XThR.Tn[2].n67 VGND 0.04833f
C21780 XThR.Tn[2].t56 VGND 0.01802f
C21781 XThR.Tn[2].t13 VGND 0.01973f
C21782 XThR.Tn[2].n68 VGND 0.05029f
C21783 XThR.Tn[2].n69 VGND 0.03533f
C21784 XThR.Tn[2].n70 VGND 0.00646f
C21785 XThR.Tn[2].n71 VGND 0.11337f
C21786 XThR.Tn[2].t59 VGND 0.01808f
C21787 XThR.Tn[2].t51 VGND 0.01979f
C21788 XThR.Tn[2].n72 VGND 0.04833f
C21789 XThR.Tn[2].t17 VGND 0.01802f
C21790 XThR.Tn[2].t29 VGND 0.01973f
C21791 XThR.Tn[2].n73 VGND 0.05029f
C21792 XThR.Tn[2].n74 VGND 0.03533f
C21793 XThR.Tn[2].n75 VGND 0.00646f
C21794 XThR.Tn[2].n76 VGND 0.11337f
C21795 XThR.Tn[2].t19 VGND 0.01808f
C21796 XThR.Tn[2].t72 VGND 0.01979f
C21797 XThR.Tn[2].n77 VGND 0.04833f
C21798 XThR.Tn[2].t33 VGND 0.01802f
C21799 XThR.Tn[2].t46 VGND 0.01973f
C21800 XThR.Tn[2].n78 VGND 0.05029f
C21801 XThR.Tn[2].n79 VGND 0.03533f
C21802 XThR.Tn[2].n80 VGND 0.00646f
C21803 XThR.Tn[2].n81 VGND 0.11337f
C21804 XThR.Tn[2].t53 VGND 0.01808f
C21805 XThR.Tn[2].t65 VGND 0.01979f
C21806 XThR.Tn[2].n82 VGND 0.04833f
C21807 XThR.Tn[2].t71 VGND 0.01802f
C21808 XThR.Tn[2].t38 VGND 0.01973f
C21809 XThR.Tn[2].n83 VGND 0.05029f
C21810 XThR.Tn[2].n84 VGND 0.03533f
C21811 XThR.Tn[2].n85 VGND 0.00646f
C21812 XThR.Tn[2].n86 VGND 0.11337f
C21813 XThR.Tn[2].n87 VGND 0.10303f
C21814 XThR.Tn[2].n88 VGND 0.22327f
.ends

