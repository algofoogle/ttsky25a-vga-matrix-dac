magic
tech sky130A
timestamp 1755581908
<< nwell >>
rect -360 -60 -105 30
<< pwell >>
rect -90 -60 190 185
<< nmos >>
rect -310 120 -295 170
rect -265 120 -250 170
rect -220 120 -205 170
<< pmos >>
rect -310 -40 -295 10
rect -265 -40 -250 10
rect -220 -40 -205 10
<< mvnmos >>
rect 0 75 100 125
rect 0 0 100 50
<< ndiff >>
rect -340 162 -310 170
rect -340 125 -334 162
rect -316 125 -310 162
rect -340 120 -310 125
rect -295 166 -265 170
rect -295 149 -289 166
rect -271 149 -265 166
rect -295 120 -265 149
rect -250 162 -220 170
rect -250 125 -244 162
rect -226 125 -220 162
rect -250 120 -220 125
rect -205 162 -175 170
rect -205 125 -199 162
rect -181 125 -175 162
rect -205 120 -175 125
<< pdiff >>
rect -340 0 -310 10
rect -340 -21 -335 0
rect -317 -21 -310 0
rect -340 -40 -310 -21
rect -295 -40 -265 10
rect -250 6 -220 10
rect -250 -11 -244 6
rect -226 -11 -220 6
rect -250 -40 -220 -11
rect -205 -19 -175 10
rect -205 -36 -199 -19
rect -181 -36 -175 -19
rect -205 -40 -175 -36
<< mvndiff >>
rect 0 155 100 160
rect 0 135 10 155
rect 90 135 100 155
rect 0 125 100 135
rect 0 50 100 75
rect 0 -10 100 0
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< ndiffc >>
rect -334 125 -316 162
rect -289 149 -271 166
rect -244 125 -226 162
rect -199 125 -181 162
<< pdiffc >>
rect -335 -21 -317 0
rect -244 -11 -226 6
rect -199 -36 -181 -19
<< mvndiffc >>
rect 10 135 90 155
rect 10 -30 90 -10
<< nsubdiff >>
rect -145 -5 -125 10
rect -145 -40 -125 -25
<< mvpsubdiff >>
rect -90 175 -40 185
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect -90 145 -40 155
rect 140 155 155 175
rect 175 155 190 175
rect 140 145 190 155
rect -90 -30 -40 -20
rect -90 -50 -75 -30
rect -55 -50 -40 -30
rect 140 -30 190 -20
rect -90 -60 -40 -50
rect 140 -50 155 -30
rect 175 -50 190 -30
rect 140 -60 190 -50
<< nsubdiffcont >>
rect -145 -25 -125 -5
<< mvpsubdiffcont >>
rect -75 155 -55 175
rect 155 155 175 175
rect -75 -50 -55 -30
rect 155 -50 175 -30
<< poly >>
rect -310 170 -295 185
rect -265 170 -250 185
rect -220 170 -205 185
rect -310 90 -295 120
rect -265 90 -250 120
rect -328 80 -295 90
rect -328 63 -320 80
rect -303 63 -295 80
rect -328 53 -295 63
rect -274 80 -241 90
rect -274 63 -266 80
rect -249 63 -241 80
rect -274 53 -241 63
rect -220 62 -205 120
rect -45 115 0 125
rect -45 85 -40 115
rect -20 85 0 115
rect -45 75 0 85
rect 100 115 145 125
rect 100 85 120 115
rect 140 85 145 115
rect 100 75 145 85
rect -220 53 -165 62
rect -310 10 -295 53
rect -265 10 -250 53
rect -220 36 -188 53
rect -171 36 -165 53
rect -220 25 -165 36
rect -45 40 0 50
rect -220 10 -205 25
rect -45 10 -40 40
rect -20 10 0 40
rect -45 0 0 10
rect 100 40 145 50
rect 100 10 120 40
rect 140 10 145 40
rect 100 0 145 10
rect -310 -55 -295 -40
rect -265 -55 -250 -40
rect -220 -55 -205 -40
<< polycont >>
rect -320 63 -303 80
rect -266 63 -249 80
rect -40 85 -20 115
rect 120 85 140 115
rect -188 36 -171 53
rect -40 10 -20 40
rect 120 10 140 40
<< locali >>
rect -334 162 -316 172
rect -289 166 -271 183
rect -90 175 -40 185
rect -289 141 -271 149
rect -244 162 -226 172
rect -334 124 -316 125
rect -244 124 -226 125
rect -334 107 -226 124
rect -199 162 -181 172
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect 140 155 155 175
rect 175 155 190 175
rect -90 145 -40 155
rect 0 135 10 155
rect 90 135 100 155
rect 140 145 190 155
rect -199 115 -181 125
rect -45 115 -15 125
rect -199 90 -40 115
rect -320 80 -303 89
rect -320 54 -303 63
rect -266 80 -249 89
rect -266 54 -249 63
rect -232 85 -40 90
rect -20 85 -15 115
rect -232 75 -15 85
rect 115 115 145 125
rect 115 85 120 115
rect 140 85 145 115
rect 115 75 145 85
rect -232 73 -181 75
rect -232 23 -215 73
rect -197 36 -188 53
rect -171 36 -156 53
rect -45 40 -15 50
rect -335 0 -317 8
rect -244 6 -215 23
rect -45 10 -40 40
rect -20 10 -15 40
rect -155 -5 -125 10
rect -45 0 -15 10
rect 115 40 145 50
rect 115 10 120 40
rect 140 10 145 40
rect 115 0 145 10
rect -244 -19 -226 -11
rect -199 -19 -181 -11
rect -335 -38 -317 -21
rect -199 -38 -181 -36
rect -335 -55 -181 -38
rect -155 -25 -145 -5
rect 0 -20 10 -10
rect -155 -40 -125 -25
rect -90 -30 10 -20
rect 90 -20 100 -10
rect 90 -30 190 -20
rect -90 -50 -75 -30
rect -55 -50 155 -30
rect 175 -50 190 -30
rect -90 -60 190 -50
<< viali >>
rect 10 135 90 155
rect -40 10 -20 40
rect 120 10 140 40
rect 10 -30 90 -10
<< metal1 >>
rect 0 155 100 185
rect 0 135 10 155
rect 90 135 100 155
rect 0 130 100 135
rect -45 40 190 50
rect -45 10 -40 40
rect -20 10 120 40
rect 140 10 190 40
rect -45 0 -15 10
rect 115 0 190 10
rect 0 -10 100 -5
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< labels >>
flabel mvndiff 5 55 95 70 0 FreeSans 80 0 0 0 SM
flabel metal1 150 5 185 45 0 FreeSans 80 0 0 0 Vbias
port 1 nsew
flabel metal1 5 165 95 180 0 FreeSans 80 0 0 0 Iout
port 2 nsew
<< end >>
