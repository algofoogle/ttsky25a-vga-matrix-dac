magic
tech sky130A
magscale 1 2
timestamp 1757695336
<< nwell >>
rect -296 -269 296 269
<< pmos >>
rect -100 -50 100 50
<< pdiff >>
rect -158 38 -100 50
rect -158 -38 -146 38
rect -112 -38 -100 38
rect -158 -50 -100 -38
rect 100 38 158 50
rect 100 -38 112 38
rect 146 -38 158 38
rect 100 -50 158 -38
<< pdiffc >>
rect -146 -38 -112 38
rect 112 -38 146 38
<< nsubdiff >>
rect -260 199 260 233
rect -260 137 -226 199
rect 226 137 260 199
rect -260 -199 -226 -137
rect 226 -199 260 -137
rect -260 -233 -164 -199
rect 164 -233 260 -199
<< nsubdiffcont >>
rect -260 -137 -226 137
rect 226 -137 260 137
rect -164 -233 164 -199
<< poly >>
rect -100 131 100 147
rect -100 97 -84 131
rect 84 97 100 131
rect -100 50 100 97
rect -100 -97 100 -50
rect -100 -131 -84 -97
rect 84 -131 100 -97
rect -100 -147 100 -131
<< polycont >>
rect -84 97 84 131
rect -84 -131 84 -97
<< locali >>
rect -260 199 260 233
rect -260 137 -226 199
rect 226 137 260 199
rect -100 97 -84 131
rect 84 97 100 131
rect -146 38 -112 54
rect -146 -54 -112 -38
rect 112 38 146 54
rect 112 -54 146 -38
rect -100 -131 -84 -97
rect 84 -131 100 -97
rect -260 -199 -226 -137
rect 226 -199 260 -137
rect -260 -233 -164 -199
rect 164 -233 260 -199
<< viali >>
rect -84 97 84 131
rect -146 -38 -112 38
rect 112 -38 146 38
rect -84 -131 84 -97
<< metal1 >>
rect -96 131 96 137
rect -96 97 -84 131
rect 84 97 96 131
rect -96 91 96 97
rect -152 38 -106 50
rect -152 -38 -146 38
rect -112 -38 -106 38
rect -152 -50 -106 -38
rect 106 38 152 50
rect 106 -38 112 38
rect 146 -38 152 38
rect 106 -50 152 -38
rect -96 -97 96 -91
rect -96 -131 -84 -97
rect 84 -131 96 -97
rect -96 -137 96 -131
<< properties >>
string FIXED_BBOX -243 -216 243 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
