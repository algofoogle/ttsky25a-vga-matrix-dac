magic
tech sky130A
timestamp 1757605323
<< nwell >>
rect 0 -27 86 0
<< pwell >>
rect 86 -27 393 0
<< nsubdiff >>
rect 18 -9 68 19
<< metal1 >>
rect 100 212 118 243
rect 89 163 118 212
rect 60 158 118 163
rect 60 127 65 158
rect 94 127 118 158
rect 60 122 118 127
rect 100 77 118 122
rect 0 72 118 77
rect 0 41 5 72
rect 34 63 118 72
rect 34 41 39 63
rect 0 36 39 41
rect 100 0 118 63
rect 173 167 217 243
rect 173 126 178 167
rect 212 126 217 167
rect 324 169 363 174
rect 324 138 329 169
rect 358 138 363 169
rect 324 133 363 138
rect 173 0 217 126
rect 260 43 299 48
rect 260 12 265 43
rect 294 12 299 43
rect 260 7 299 12
<< via1 >>
rect 65 127 94 158
rect 5 41 34 72
rect 178 126 212 167
rect 329 138 358 169
rect 265 12 294 43
<< metal2 >>
rect 173 167 217 172
rect 60 158 100 163
rect 60 127 65 158
rect 94 127 100 158
rect 60 121 100 127
rect 173 126 178 167
rect 212 145 217 167
rect 324 169 363 174
rect 324 145 329 169
rect 212 138 329 145
rect 358 138 363 169
rect 212 130 363 138
rect 212 126 217 130
rect 173 121 217 126
rect 0 72 393 77
rect 0 41 5 72
rect 34 63 393 72
rect 34 41 39 63
rect 0 36 39 41
rect 260 43 299 48
rect 260 12 265 43
rect 294 12 299 43
rect 260 7 299 12
<< via2 >>
rect 65 127 94 158
rect 178 126 212 167
rect 329 138 358 169
rect 5 41 34 72
rect 265 12 294 43
<< metal3 >>
rect 0 77 30 243
rect 69 163 99 243
rect 60 158 99 163
rect 60 127 65 158
rect 94 127 99 158
rect 60 122 99 127
rect 0 72 39 77
rect 0 41 5 72
rect 34 41 39 72
rect 0 36 39 41
rect 0 0 30 36
rect 69 0 99 122
rect 173 167 217 243
rect 173 126 178 167
rect 212 126 217 167
rect 173 0 217 126
rect 260 49 290 202
rect 333 174 363 243
rect 324 169 363 174
rect 324 138 329 169
rect 358 138 363 169
rect 324 133 363 138
rect 260 44 302 49
rect 260 12 265 44
rect 297 12 302 44
rect 260 7 302 12
rect 333 0 363 133
<< via3 >>
rect 178 126 212 167
rect 265 43 297 44
rect 265 12 294 43
rect 294 12 297 43
<< metal4 >>
rect 0 167 393 172
rect 0 126 178 167
rect 212 126 393 167
rect 0 121 393 126
rect 240 44 320 48
rect 240 12 265 44
rect 297 12 320 44
rect 240 7 320 12
use icell  icell
timestamp 1757605323
transform 1 0 0 0 1 0
box 0 0 393 243
<< labels >>
flabel metal3 0 220 30 232 0 FreeSans 40 0 0 0 VPWR
port 1 nsew
flabel metal3 173 220 217 232 0 FreeSans 40 0 0 0 VGND
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 393 232
<< end >>
