magic
tech sky130A
timestamp 1756363220
<< nwell >>
rect 0 -11 86 232
<< pwell >>
rect 86 -11 393 232
<< nmos >>
rect 131 167 182 182
rect 131 122 182 137
rect 131 77 182 92
<< pmos >>
rect 18 167 68 182
rect 18 122 68 137
rect 18 77 68 92
<< mvnmos >>
rect 260 122 310 172
rect 260 47 310 97
<< ndiff >>
rect 131 206 182 210
rect 131 188 139 206
rect 176 188 182 206
rect 131 182 182 188
rect 131 161 182 167
rect 131 143 135 161
rect 152 143 182 161
rect 131 137 182 143
rect 131 116 182 122
rect 131 98 139 116
rect 176 98 182 116
rect 131 92 182 98
rect 131 71 182 77
rect 131 53 141 71
rect 174 53 182 71
rect 131 49 182 53
<< pdiff >>
rect 18 207 68 212
rect 18 189 37 207
rect 58 189 68 207
rect 18 182 68 189
rect 18 137 68 167
rect 18 116 68 122
rect 18 98 47 116
rect 64 98 68 116
rect 18 92 68 98
rect 18 70 68 77
rect 18 53 22 70
rect 39 53 68 70
rect 18 47 68 53
<< mvndiff >>
rect 260 203 310 207
rect 260 182 268 203
rect 302 182 310 203
rect 260 172 310 182
rect 260 97 310 122
rect 260 37 310 47
rect 260 17 268 37
rect 302 17 310 37
rect 260 12 310 17
<< ndiffc >>
rect 139 188 176 206
rect 135 143 152 161
rect 139 98 176 116
rect 141 53 174 71
<< pdiffc >>
rect 37 189 58 207
rect 47 98 64 116
rect 22 53 39 70
<< mvndiffc >>
rect 268 182 302 203
rect 268 17 302 37
<< nsubdiff >>
rect 18 36 68 47
rect 18 19 22 36
rect 39 19 68 36
rect 18 7 68 19
<< mvpsubdiff >>
rect 169 5 185 22
rect 205 5 221 22
<< nsubdiffcont >>
rect 22 19 39 36
<< mvpsubdiffcont >>
rect 185 5 205 22
<< poly >>
rect 87 192 114 200
rect 87 182 92 192
rect 5 167 18 182
rect 68 175 92 182
rect 109 182 114 192
rect 109 175 131 182
rect 68 167 131 175
rect 182 167 195 182
rect 87 138 114 146
rect 87 137 92 138
rect 5 122 18 137
rect 68 122 92 137
rect 87 121 92 122
rect 109 137 114 138
rect 216 162 260 172
rect 109 122 131 137
rect 182 122 195 137
rect 216 132 221 162
rect 241 132 260 162
rect 216 122 260 132
rect 310 162 354 172
rect 310 132 329 162
rect 349 132 354 162
rect 310 122 354 132
rect 109 121 114 122
rect 87 113 114 121
rect 5 77 18 92
rect 68 84 131 92
rect 68 77 92 84
rect 87 67 92 77
rect 109 77 131 84
rect 182 77 195 92
rect 216 87 260 97
rect 109 67 114 77
rect 87 59 114 67
rect 216 57 221 87
rect 241 57 260 87
rect 216 47 260 57
rect 310 87 354 97
rect 310 57 329 87
rect 349 57 354 87
rect 310 47 354 57
<< polycont >>
rect 92 175 109 192
rect 92 121 109 138
rect 221 132 241 162
rect 329 132 349 162
rect 92 67 109 84
rect 221 57 241 87
rect 329 57 349 87
<< locali >>
rect 3 207 66 215
rect 3 189 37 207
rect 58 189 66 207
rect 92 192 109 201
rect 3 78 22 189
rect 131 188 139 206
rect 176 188 194 206
rect 92 166 109 175
rect 92 138 109 147
rect 127 143 135 161
rect 152 143 160 161
rect 39 98 47 116
rect 64 98 73 116
rect 92 112 109 121
rect 177 116 194 188
rect 260 203 310 207
rect 260 182 268 203
rect 302 182 310 203
rect 216 162 246 172
rect 324 162 354 172
rect 216 132 221 162
rect 241 132 329 162
rect 349 132 354 162
rect 216 122 354 132
rect 131 98 139 116
rect 176 98 194 116
rect 3 70 39 78
rect 3 19 22 70
rect 56 41 73 98
rect 92 84 109 93
rect 216 87 354 97
rect 216 71 221 87
rect 92 58 109 67
rect 133 53 141 71
rect 174 57 221 71
rect 241 57 329 87
rect 349 57 354 87
rect 174 53 246 57
rect 133 41 150 53
rect 216 47 246 53
rect 324 47 354 57
rect 56 24 150 41
rect 3 11 39 19
rect 173 5 185 22
rect 205 5 217 22
rect 260 17 268 37
rect 302 17 310 37
<< viali >>
rect 92 175 109 192
rect 135 143 152 161
rect 92 121 109 138
rect 268 182 302 203
rect 329 132 349 162
rect 22 36 39 53
rect 92 67 109 84
rect 185 5 205 22
rect 268 17 302 37
<< metal1 >>
rect 173 203 310 212
rect 77 192 112 201
rect 77 175 92 192
rect 109 175 112 192
rect 77 166 112 175
rect 173 182 268 203
rect 302 182 310 203
rect 173 177 310 182
rect 173 169 208 177
rect 132 161 208 169
rect 42 138 112 147
rect 42 121 92 138
rect 109 121 112 138
rect 132 143 135 161
rect 152 143 208 161
rect 132 134 208 143
rect 42 112 112 121
rect 77 84 112 93
rect 77 67 92 84
rect 109 67 112 84
rect 7 53 42 62
rect 77 58 112 67
rect 7 36 22 53
rect 39 36 42 53
rect 7 27 42 36
rect 173 31 208 134
rect 324 162 364 172
rect 324 132 329 162
rect 349 132 364 162
rect 324 122 364 132
rect 260 37 310 40
rect 173 22 217 31
rect 173 5 185 22
rect 205 5 217 22
rect 173 -4 217 5
rect 260 17 268 37
rect 302 17 310 37
rect 260 -4 310 17
<< labels >>
flabel mvndiff 265 102 305 117 0 FreeSans 80 0 0 0 SM
flabel metal1 329 127 359 167 0 FreeSans 80 0 0 0 Vbias
port 1 nsew
flabel metal1 178 139 203 164 0 FreeSans 64 0 0 0 VGND
port 4 nsew
flabel metal1 265 1 305 35 0 FreeSans 64 0 0 0 Iout
port 5 nsew
flabel metal1 82 63 107 88 0 FreeSans 64 0 0 0 Sn
port 6 nsew
flabel metal1 47 117 72 142 0 FreeSans 64 0 0 0 Cn
port 7 nsew
flabel metal1 82 171 107 196 0 FreeSans 64 0 0 0 Rn
port 8 nsew
flabel metal1 12 32 37 57 0 FreeSans 64 0 0 0 VPWR
port 9 nsew
flabel locali 92 25 122 40 0 FreeSans 80 0 0 0 Ien
flabel locali 133 190 167 204 0 FreeSans 80 0 0 0 PDM
flabel pdiff 26 145 60 159 0 FreeSans 80 0 0 0 PUM
<< properties >>
string FIXED_BBOX 0 0 393 232
<< end >>
