magic
tech sky130A
timestamp 1756902890
<< metal2 >>
rect 173 3651 217 3669
rect -28 3436 0 3450
rect -28 3204 -14 3218
rect -28 2972 -14 2986
rect -28 2740 -14 2754
rect -28 2508 -14 2522
rect -28 2276 -14 2290
rect -28 2044 -14 2058
rect -28 1812 -14 1826
rect -28 1580 -14 1594
rect -28 1348 -14 1362
rect -28 1116 -14 1130
rect -28 884 -14 898
rect -28 652 -14 666
rect -28 420 -14 434
rect -28 188 -14 202
rect 0 -44 39 77
<< metal3 >>
rect 722 4026 760 4029
rect 722 3994 725 4026
rect 757 3994 760 4026
rect 722 3991 760 3994
rect 1115 4026 1153 4029
rect 1115 3994 1118 4026
rect 1150 3994 1153 4026
rect 1115 3991 1153 3994
rect 1508 4026 1546 4029
rect 1508 3994 1511 4026
rect 1543 3994 1546 4026
rect 1508 3991 1546 3994
rect 1901 4026 1939 4029
rect 1901 3994 1904 4026
rect 1936 3994 1939 4026
rect 1901 3991 1939 3994
rect 2294 4026 2332 4029
rect 2294 3994 2297 4026
rect 2329 3994 2332 4026
rect 2294 3991 2332 3994
rect 2687 4026 2725 4029
rect 2687 3994 2690 4026
rect 2722 3994 2725 4026
rect 2687 3991 2725 3994
rect 3080 4026 3118 4029
rect 3080 3994 3083 4026
rect 3115 3994 3118 4026
rect 3080 3991 3118 3994
rect 3473 4026 3511 4029
rect 3473 3994 3476 4026
rect 3508 3994 3511 4026
rect 3473 3991 3511 3994
rect 3866 4026 3904 4029
rect 3866 3994 3869 4026
rect 3901 3994 3904 4026
rect 3866 3991 3904 3994
rect 4259 4026 4297 4029
rect 4259 3994 4262 4026
rect 4294 3994 4297 4026
rect 4259 3991 4297 3994
rect 4652 4026 4690 4029
rect 4652 3994 4655 4026
rect 4687 3994 4690 4026
rect 4652 3991 4690 3994
rect 5045 4026 5083 4029
rect 5045 3994 5048 4026
rect 5080 3994 5083 4026
rect 5045 3991 5083 3994
rect 5438 4026 5476 4029
rect 5438 3994 5441 4026
rect 5473 3994 5476 4026
rect 5438 3991 5476 3994
rect 5831 4026 5869 4029
rect 5831 3994 5834 4026
rect 5866 3994 5869 4026
rect 5831 3991 5869 3994
rect 6224 4026 6262 4029
rect 6224 3994 6227 4026
rect 6259 3994 6262 4026
rect 6224 3991 6262 3994
rect 6617 4026 6655 4029
rect 6617 3994 6620 4026
rect 6652 3994 6655 4026
rect 6617 3991 6655 3994
rect 173 3958 217 3961
rect 173 3864 176 3958
rect 214 3864 217 3958
rect 0 3828 38 3831
rect 0 3734 3 3828
rect 35 3734 38 3828
rect 0 3731 38 3734
rect 0 3700 30 3731
rect 173 3700 217 3864
rect 566 3958 610 3961
rect 566 3864 569 3958
rect 607 3864 610 3958
rect 393 3828 431 3831
rect 393 3734 396 3828
rect 428 3734 431 3828
rect 393 3731 431 3734
rect 393 3700 423 3731
rect 462 3700 492 3753
rect 566 3700 610 3864
rect 726 3700 756 3991
rect 959 3958 1003 3961
rect 959 3864 962 3958
rect 1000 3864 1003 3958
rect 786 3828 824 3831
rect 786 3734 789 3828
rect 821 3734 824 3828
rect 786 3731 824 3734
rect 786 3700 816 3731
rect 855 3700 885 3753
rect 959 3700 1003 3864
rect 1119 3700 1149 3991
rect 1352 3958 1396 3961
rect 1352 3864 1355 3958
rect 1393 3864 1396 3958
rect 1179 3828 1217 3831
rect 1179 3734 1182 3828
rect 1214 3734 1217 3828
rect 1179 3731 1217 3734
rect 1179 3700 1209 3731
rect 1248 3700 1278 3753
rect 1352 3700 1396 3864
rect 1512 3700 1542 3991
rect 1745 3958 1789 3961
rect 1745 3864 1748 3958
rect 1786 3864 1789 3958
rect 1572 3828 1610 3831
rect 1572 3734 1575 3828
rect 1607 3734 1610 3828
rect 1572 3731 1610 3734
rect 1572 3700 1602 3731
rect 1641 3700 1671 3753
rect 1745 3700 1789 3864
rect 1905 3700 1935 3991
rect 2138 3958 2182 3961
rect 2138 3864 2141 3958
rect 2179 3864 2182 3958
rect 1965 3828 2003 3831
rect 1965 3734 1968 3828
rect 2000 3734 2003 3828
rect 1965 3731 2003 3734
rect 1965 3700 1995 3731
rect 2034 3700 2064 3753
rect 2138 3700 2182 3864
rect 2298 3700 2328 3991
rect 2531 3958 2575 3961
rect 2531 3864 2534 3958
rect 2572 3864 2575 3958
rect 2358 3828 2396 3831
rect 2358 3734 2361 3828
rect 2393 3734 2396 3828
rect 2358 3731 2396 3734
rect 2358 3700 2388 3731
rect 2427 3700 2457 3753
rect 2531 3700 2575 3864
rect 2691 3700 2721 3991
rect 2924 3958 2968 3961
rect 2924 3864 2927 3958
rect 2965 3864 2968 3958
rect 2751 3828 2789 3831
rect 2751 3734 2754 3828
rect 2786 3734 2789 3828
rect 2751 3731 2789 3734
rect 2751 3700 2781 3731
rect 2820 3700 2850 3753
rect 2924 3700 2968 3864
rect 3084 3700 3114 3991
rect 3317 3958 3361 3961
rect 3317 3864 3320 3958
rect 3358 3864 3361 3958
rect 3144 3828 3182 3831
rect 3144 3734 3147 3828
rect 3179 3734 3182 3828
rect 3144 3731 3182 3734
rect 3144 3700 3174 3731
rect 3213 3700 3243 3753
rect 3317 3700 3361 3864
rect 3477 3700 3507 3991
rect 3710 3958 3754 3961
rect 3710 3864 3713 3958
rect 3751 3864 3754 3958
rect 3537 3828 3575 3831
rect 3537 3734 3540 3828
rect 3572 3734 3575 3828
rect 3537 3731 3575 3734
rect 3537 3700 3567 3731
rect 3606 3700 3636 3753
rect 3710 3700 3754 3864
rect 3870 3700 3900 3991
rect 4103 3958 4147 3961
rect 4103 3864 4106 3958
rect 4144 3864 4147 3958
rect 3930 3828 3968 3831
rect 3930 3734 3933 3828
rect 3965 3734 3968 3828
rect 3930 3731 3968 3734
rect 3930 3700 3960 3731
rect 3999 3700 4029 3753
rect 4103 3700 4147 3864
rect 4263 3700 4293 3991
rect 4496 3958 4540 3961
rect 4496 3864 4499 3958
rect 4537 3864 4540 3958
rect 4323 3828 4361 3831
rect 4323 3734 4326 3828
rect 4358 3734 4361 3828
rect 4323 3731 4361 3734
rect 4323 3700 4353 3731
rect 4392 3700 4422 3753
rect 4496 3700 4540 3864
rect 4656 3700 4686 3991
rect 4889 3958 4933 3961
rect 4889 3864 4892 3958
rect 4930 3864 4933 3958
rect 4716 3828 4754 3831
rect 4716 3734 4719 3828
rect 4751 3734 4754 3828
rect 4716 3731 4754 3734
rect 4716 3700 4746 3731
rect 4785 3700 4815 3753
rect 4889 3700 4933 3864
rect 5049 3700 5079 3991
rect 5282 3958 5326 3961
rect 5282 3864 5285 3958
rect 5323 3864 5326 3958
rect 5109 3828 5147 3831
rect 5109 3734 5112 3828
rect 5144 3734 5147 3828
rect 5109 3731 5147 3734
rect 5109 3700 5139 3731
rect 5178 3700 5208 3753
rect 5282 3700 5326 3864
rect 5442 3700 5472 3991
rect 5675 3958 5719 3961
rect 5675 3864 5678 3958
rect 5716 3864 5719 3958
rect 5502 3828 5540 3831
rect 5502 3734 5505 3828
rect 5537 3734 5540 3828
rect 5502 3731 5540 3734
rect 5502 3700 5532 3731
rect 5571 3700 5601 3753
rect 5675 3700 5719 3864
rect 5835 3700 5865 3991
rect 6068 3958 6112 3961
rect 6068 3864 6071 3958
rect 6109 3864 6112 3958
rect 5895 3828 5933 3831
rect 5895 3734 5898 3828
rect 5930 3734 5933 3828
rect 5895 3731 5933 3734
rect 5895 3700 5925 3731
rect 5964 3700 5994 3753
rect 6068 3700 6112 3864
rect 6228 3700 6258 3991
rect 6461 3958 6505 3961
rect 6461 3864 6464 3958
rect 6502 3864 6505 3958
rect 6288 3828 6326 3831
rect 6288 3734 6291 3828
rect 6323 3734 6326 3828
rect 6288 3731 6326 3734
rect 6288 3700 6318 3731
rect 6461 3700 6505 3864
rect 6621 3700 6651 3991
rect 6854 3958 6898 3961
rect 6854 3864 6857 3958
rect 6895 3864 6898 3958
rect 6681 3828 6719 3831
rect 6681 3734 6684 3828
rect 6716 3734 6719 3828
rect 6681 3731 6719 3734
rect 6681 3700 6711 3731
rect 6854 3700 6898 3864
<< via3 >>
rect 725 3994 757 4026
rect 1118 3994 1150 4026
rect 1511 3994 1543 4026
rect 1904 3994 1936 4026
rect 2297 3994 2329 4026
rect 2690 3994 2722 4026
rect 3083 3994 3115 4026
rect 3476 3994 3508 4026
rect 3869 3994 3901 4026
rect 4262 3994 4294 4026
rect 4655 3994 4687 4026
rect 5048 3994 5080 4026
rect 5441 3994 5473 4026
rect 5834 3994 5866 4026
rect 6227 3994 6259 4026
rect 6620 3994 6652 4026
rect 176 3864 214 3958
rect 3 3734 35 3828
rect 569 3864 607 3958
rect 396 3734 428 3828
rect 962 3864 1000 3958
rect 789 3734 821 3828
rect 1355 3864 1393 3958
rect 1182 3734 1214 3828
rect 1748 3864 1786 3958
rect 1575 3734 1607 3828
rect 2141 3864 2179 3958
rect 1968 3734 2000 3828
rect 2534 3864 2572 3958
rect 2361 3734 2393 3828
rect 2927 3864 2965 3958
rect 2754 3734 2786 3828
rect 3320 3864 3358 3958
rect 3147 3734 3179 3828
rect 3713 3864 3751 3958
rect 3540 3734 3572 3828
rect 4106 3864 4144 3958
rect 3933 3734 3965 3828
rect 4499 3864 4537 3958
rect 4326 3734 4358 3828
rect 4892 3864 4930 3958
rect 4719 3734 4751 3828
rect 5285 3864 5323 3958
rect 5112 3734 5144 3828
rect 5678 3864 5716 3958
rect 5505 3734 5537 3828
rect 6071 3864 6109 3958
rect 5898 3734 5930 3828
rect 6464 3864 6502 3958
rect 6291 3734 6323 3828
rect 6857 3864 6895 3958
rect 6684 3734 6716 3828
<< metal4 >>
rect 722 4026 760 4029
rect 722 4021 725 4026
rect -30 3994 725 4021
rect 757 4021 760 4026
rect 1115 4026 1153 4029
rect 1115 4021 1118 4026
rect 757 3994 1118 4021
rect 1150 4021 1153 4026
rect 1508 4026 1546 4029
rect 1508 4021 1511 4026
rect 1150 3994 1511 4021
rect 1543 4021 1546 4026
rect 1901 4026 1939 4029
rect 1901 4021 1904 4026
rect 1543 3994 1904 4021
rect 1936 4021 1939 4026
rect 2294 4026 2332 4029
rect 2294 4021 2297 4026
rect 1936 3994 2297 4021
rect 2329 4021 2332 4026
rect 2687 4026 2725 4029
rect 2687 4021 2690 4026
rect 2329 3994 2690 4021
rect 2722 4021 2725 4026
rect 3080 4026 3118 4029
rect 3080 4021 3083 4026
rect 2722 3994 3083 4021
rect 3115 4021 3118 4026
rect 3473 4026 3511 4029
rect 3473 4021 3476 4026
rect 3115 3994 3476 4021
rect 3508 4021 3511 4026
rect 3866 4026 3904 4029
rect 3866 4021 3869 4026
rect 3508 3994 3869 4021
rect 3901 4021 3904 4026
rect 4259 4026 4297 4029
rect 4259 4021 4262 4026
rect 3901 3994 4262 4021
rect 4294 4021 4297 4026
rect 4652 4026 4690 4029
rect 4652 4021 4655 4026
rect 4294 3994 4655 4021
rect 4687 4021 4690 4026
rect 5045 4026 5083 4029
rect 5045 4021 5048 4026
rect 4687 3994 5048 4021
rect 5080 4021 5083 4026
rect 5438 4026 5476 4029
rect 5438 4021 5441 4026
rect 5080 3994 5441 4021
rect 5473 4021 5476 4026
rect 5831 4026 5869 4029
rect 5831 4021 5834 4026
rect 5473 3994 5834 4021
rect 5866 4021 5869 4026
rect 6224 4026 6262 4029
rect 6224 4021 6227 4026
rect 5866 3994 6227 4021
rect 6259 4021 6262 4026
rect 6617 4026 6655 4029
rect 6617 4021 6620 4026
rect 6259 3994 6620 4021
rect 6652 4021 6655 4026
rect 6652 3994 7074 4021
rect -30 3991 7074 3994
rect -30 3958 7074 3961
rect -30 3864 176 3958
rect 214 3864 569 3958
rect 607 3864 962 3958
rect 1000 3864 1355 3958
rect 1393 3864 1748 3958
rect 1786 3864 2141 3958
rect 2179 3864 2534 3958
rect 2572 3864 2927 3958
rect 2965 3864 3320 3958
rect 3358 3864 3713 3958
rect 3751 3864 4106 3958
rect 4144 3864 4499 3958
rect 4537 3864 4892 3958
rect 4930 3864 5285 3958
rect 5323 3864 5678 3958
rect 5716 3864 6071 3958
rect 6109 3864 6464 3958
rect 6502 3864 6857 3958
rect 6895 3864 7074 3958
rect -30 3861 7074 3864
rect -30 3828 7074 3831
rect -30 3734 3 3828
rect 35 3734 396 3828
rect 428 3734 789 3828
rect 821 3734 1182 3828
rect 1214 3734 1575 3828
rect 1607 3734 1968 3828
rect 2000 3734 2361 3828
rect 2393 3734 2754 3828
rect 2786 3734 3147 3828
rect 3179 3734 3540 3828
rect 3572 3734 3933 3828
rect 3965 3734 4326 3828
rect 4358 3734 4719 3828
rect 4751 3734 5112 3828
rect 5144 3734 5505 3828
rect 5537 3734 5898 3828
rect 5930 3734 6291 3828
rect 6323 3734 6684 3828
rect 6716 3734 7074 3828
rect -30 3731 7074 3734
rect 393 -152 6681 48
use row15x  XIR
array 1 1 7074 15 0 232
timestamp 1756902890
transform 1 0 0 0 1 0
box -28 -55 7074 243
<< labels >>
flabel metal2 -28 3436 -14 3450 0 FreeSans 40 0 0 0 Rn[0]
port 0 nsew
flabel metal2 -28 3204 -14 3218 0 FreeSans 40 0 0 0 Rn[1]
port 1 nsew
flabel metal2 -28 2972 -14 2986 0 FreeSans 40 0 0 0 Rn[2]
port 2 nsew
flabel metal2 -28 2740 -14 2754 0 FreeSans 40 0 0 0 Rn[3]
port 3 nsew
flabel metal2 -28 2508 -14 2522 0 FreeSans 40 0 0 0 Rn[4]
port 4 nsew
flabel metal2 -28 2276 -14 2290 0 FreeSans 40 0 0 0 Rn[5]
port 5 nsew
flabel metal2 -28 2044 -14 2058 0 FreeSans 40 0 0 0 Rn[6]
port 6 nsew
flabel metal2 -28 1812 -14 1826 0 FreeSans 40 0 0 0 Rn[7]
port 7 nsew
flabel metal2 -28 1580 -14 1594 0 FreeSans 40 0 0 0 Rn[8]
port 8 nsew
flabel metal2 -28 1348 -14 1362 0 FreeSans 40 0 0 0 Rn[9]
port 9 nsew
flabel metal2 -28 1116 -14 1130 0 FreeSans 40 0 0 0 Rn[10]
port 10 nsew
flabel metal2 -28 884 -14 898 0 FreeSans 40 0 0 0 Rn[11]
port 11 nsew
flabel metal2 -28 652 -14 666 0 FreeSans 40 0 0 0 Rn[12]
port 12 nsew
flabel metal2 -28 420 -14 434 0 FreeSans 40 0 0 0 Rn[13]
port 13 nsew
flabel metal2 -28 188 -14 202 0 FreeSans 40 0 0 0 Rn[14]
port 14 nsew
flabel metal3 462 3738 492 3753 0 FreeSans 40 0 0 0 Cn[0]
port 100 nsew
flabel metal3 855 3738 885 3753 0 FreeSans 40 0 0 0 Cn[1]
port 101 nsew
flabel metal3 1248 3738 1278 3753 0 FreeSans 40 0 0 0 Cn[2]
port 102 nsew
flabel metal3 1641 3738 1671 3753 0 FreeSans 40 0 0 0 Cn[3]
port 103 nsew
flabel metal3 2034 3738 2064 3753 0 FreeSans 40 0 0 0 Cn[4]
port 104 nsew
flabel metal3 2427 3738 2457 3753 0 FreeSans 40 0 0 0 Cn[5]
port 105 nsew
flabel metal3 2820 3738 2850 3753 0 FreeSans 40 0 0 0 Cn[6]
port 106 nsew
flabel metal3 3213 3738 3243 3753 0 FreeSans 40 0 0 0 Cn[7]
port 107 nsew
flabel metal3 3606 3738 3636 3753 0 FreeSans 40 0 0 0 Cn[8]
port 108 nsew
flabel metal3 3999 3738 4029 3753 0 FreeSans 40 0 0 0 Cn[9]
port 109 nsew
flabel metal3 4392 3738 4422 3753 0 FreeSans 40 0 0 0 Cn[10]
port 110 nsew
flabel metal3 4785 3738 4815 3753 0 FreeSans 40 0 0 0 Cn[11]
port 111 nsew
flabel metal3 5178 3738 5208 3753 0 FreeSans 40 0 0 0 Cn[12]
port 112 nsew
flabel metal3 5571 3738 5601 3753 0 FreeSans 40 0 0 0 Cn[13]
port 113 nsew
flabel metal3 5964 3738 5994 3753 0 FreeSans 40 0 0 0 Cn[14]
port 114 nsew
flabel metal4 -30 3861 0 3961 0 FreeSans 80 90 0 0 VGND
port 200 nsew
flabel metal4 -30 3731 0 3831 0 FreeSans 80 90 0 0 VPWR
port 201 nsew
flabel metal4 -30 3991 0 4021 0 FreeSans 80 90 0 0 Vbias
port 202 nsew
flabel metal4 6581 -152 6681 -52 0 FreeSans 80 0 0 0 Iout
port 203 nsew
<< end >>
