* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias bias[2] bias[1] bias[0] data[0] data[1]
+ data[2] data[3] data[4] data[5] data[6] data[7]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t1409 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1408 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t194 VGND.t1979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t381 VPWR.t383 VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t91 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t1837 XThR.XTBN.Y a_n997_2667# VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t735 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t1805 VPWR.t1804 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t2327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t11 XThC.XTBN.Y.t4 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t189 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t363 VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t49 XThC.XTBN.Y.t5 XThC.Tn[5].t11 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t785 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t204 VGND.t2054 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t2329 VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t687 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t135 VGND.t1363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t219 VGND.t2188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t3 XThC.XTB5.Y VPWR.t784 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t191 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t203 VGND.t2053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t3 VPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t379 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t192 VGND.t1731 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t1668 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t7 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1976 VGND.t1978 VGND.t1977 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t2634 VGND.t2633 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t7 XThR.XTBN.Y a_n1049_5611# VPWR.t1283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t544 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t51 XThC.XTBN.Y.t8 XThC.Tn[2].t7 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t395 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t502 VGND.t501 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t81 VGND.t743 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t1621 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t1620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t378 VPWR.t376 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t193 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t1852 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1851 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t2540 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t2539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t498 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t1378 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t1377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t195 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t550 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t549 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1260 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t373 VPWR.t375 VPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t11 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t2542 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t2541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t1911 VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t7 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t1558 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.XTB5.Y XThC.XTB7.B VGND.t248 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t3 XThC.XTBN.Y.t9 VPWR.t415 VPWR.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t365 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t1504 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t1503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t1560 VPWR.t1559 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t1347 XThR.XTBN.Y XThR.Tn[9].t11 VPWR.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1854 VPWR.t1853 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t1856 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t2331 VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t2687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t1407 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1406 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t737 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t736 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t372 VPWR.t370 XA.XIR[2].XIC_15.icell.PUM VPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.XTB7.Y VPWR.t773 VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t2025 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t2636 VGND.t2635 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t3 XThR.XTBN.Y VPWR.t1346 VPWR.t1345 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t989 VGND.t988 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.XTBN.Y.t10 VGND.t53 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t2544 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t2543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t1516 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t1515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t109 VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t183 VGND.t1690 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t197 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t1836 XThR.XTBN.Y XThR.Tn[5].t11 VGND.t1819 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t2546 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t2545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t2548 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t2547 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t808 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t807 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t689 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t230 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t1562 VPWR.t1561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t1254 XThR.XTB6.Y a_n1049_5611# VPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t1164 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t2550 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t2549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t1623 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t1622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 a_n1049_7787# XThR.XTB2.Y VPWR.t411 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 VGND.t546 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X96 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t1402 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X97 VGND.t2552 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t2551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X98 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t836 VPWR.t835 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X99 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t1449 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X100 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t368 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 VGND.t2295 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t2294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X102 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t991 VGND.t990 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X103 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1564 VPWR.t1563 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X104 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t1404 VGND.t1403 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X105 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t1137 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t1858 VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X107 VGND.t17 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X108 VPWR.t1710 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X109 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X110 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 VPWR.t1268 data[4].t0 a_n1335_4229# VPWR.t1267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X112 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1405 VPWR.t1404 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X113 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t133 VGND.t1357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X114 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X115 VGND.t1835 XThR.XTBN.Y XThR.Tn[7].t7 VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X116 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X117 a_n1319_5317# XThR.XTB7.A VPWR.t775 VPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X118 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t1138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X119 VPWR.t1175 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t1174 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X120 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X121 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t598 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X122 XThC.Tn[9].t7 XThC.XTB2.Y VPWR.t1868 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 XA.XIR[15].XIC[4].icell.Ien VPWR.t365 VPWR.t367 VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X124 VGND.t2297 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t2296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X125 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t53 VGND.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X126 VGND.t2299 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t2298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X127 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t362 VPWR.t364 VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X128 XThC.Tn[5].t10 XThC.XTBN.Y.t11 VGND.t54 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X130 VGND.t2301 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t2300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X131 VGND.t2303 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t2302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t1518 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t1517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X133 VPWR.t1013 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t1012 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X134 VPWR.t1693 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t1692 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VGND.t1975 VGND.t1973 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X136 XThR.Tn[9].t7 XThR.XTB2.Y a_n997_3755# VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X137 XThC.Tn[0].t2 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t200 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X139 XThC.Tn[5].t6 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X140 VGND.t543 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X141 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X142 VGND.t2305 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t2304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X143 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t7 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X144 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X145 XThC.Tn[7].t7 XThC.XTBN.Y.t14 VGND.t319 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X146 XThC.Tn[2].t6 XThC.XTBN.Y.t15 VGND.t320 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 VGND.t2518 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X148 a_n997_1579# XThR.XTBN.Y VGND.t1833 VGND.t1817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X149 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t287 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X150 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t289 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t360 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t69 VGND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X153 VGND.t2008 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t2007 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X154 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X155 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X156 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t2674 VGND.t2673 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t636 VGND.t635 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X159 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X160 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t1141 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t28 VGND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X162 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t19 VGND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t1536 VGND.t1535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X164 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t1695 VPWR.t1694 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X166 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t167 VGND.t1655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X167 XA.XIR[15].XIC[0].icell.Ien VPWR.t357 VPWR.t359 VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X168 VGND.t2307 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t2306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X169 VGND.t1692 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t1691 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X170 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t354 VPWR.t356 VPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X171 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X172 VGND.t338 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t337 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X173 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t1807 VPWR.t1806 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X174 VGND.t321 XThC.XTBN.Y.t16 XThC.Tn[1].t7 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VGND.t2309 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t2308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X176 VPWR.t1697 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t1696 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X177 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t1095 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X178 XA.XIR[2].XIC_15.icell.PUM VPWR.t352 XA.XIR[2].XIC_15.icell.Ien VPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X180 VPWR.t609 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t608 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X181 VPWR.t1015 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t1014 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VGND.t2311 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t2310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X183 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t202 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X184 VPWR.t351 VPWR.t349 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X185 VPWR.t580 XThC.XTBN.Y.t17 XThC.Tn[10].t0 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VGND.t1832 XThR.XTBN.Y XThR.Tn[3].t6 VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t61 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X188 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t1891 VPWR.t1890 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X189 XThR.Tn[0].t6 XThR.XTBN.Y a_n1049_8581# VPWR.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t1779 VPWR.t1778 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X191 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t106 VGND.t1004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X192 VPWR.t1440 VGND.t2688 XA.XIR[0].XIC[8].icell.PUM VPWR.t1439 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X193 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X194 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XThC.Tn[12].t2 XThC.XTB5.Y VPWR.t783 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X196 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t852 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X197 XThR.Tn[11].t9 XThR.XTBN.Y VPWR.t1343 VPWR.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t980 VPWR.t979 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X199 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X200 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t786 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t1143 VGND.t1142 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t1334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X203 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t291 VGND.t290 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X204 VGND.t691 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t690 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t1768 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XThR.Tn[2].t11 XThR.XTBN.Y VGND.t1831 VGND.t1782 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VGND.t693 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X208 VGND.t1972 VGND.t1970 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1971 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X209 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t1699 VPWR.t1698 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X210 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1225 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X211 VPWR.t1342 XThR.XTBN.Y XThR.Tn[12].t11 VPWR.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X212 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t638 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X213 XThC.XTB7.A data[0].t0 VPWR.t985 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 VPWR.t611 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X215 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t1096 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X216 VGND.t2313 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t2312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X217 XA.XIR[0].XIC[13].icell.PDM VGND.t1967 VGND.t1969 VGND.t1968 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X218 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t2534 VGND.t2533 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 VGND.t204 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t1625 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t1624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t2315 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t2314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X222 XThC.Tn[9].t11 XThC.XTB2.Y a_7875_9569# VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 VGND.t70 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X224 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X225 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X226 VGND.t1627 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t1626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t1380 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t208 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 a_n1319_5611# XThR.XTB6.A VPWR.t393 VPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X230 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t1781 VPWR.t1780 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X231 VGND.t1830 XThR.XTBN.Y a_n997_3979# VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X232 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t21 VGND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X233 VPWR.t582 XThC.XTBN.Y.t18 XThC.Tn[14].t11 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 VGND.t2317 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t2316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X235 VPWR.t1701 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t1700 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X236 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t1450 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X237 VGND.t2319 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t2318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X238 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t1393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X239 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t1123 VPWR.t1122 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X241 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X242 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t1893 VPWR.t1892 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X243 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X244 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t163 VGND.t1582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X245 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t838 VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X246 VGND.t661 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X247 VGND.t2016 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t2015 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X248 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t293 VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 VPWR.t1463 XThR.XTB4.Y.t2 a_n1049_6699# VPWR.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X250 VGND.t210 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X251 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t26 VGND.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X252 VPWR.t1438 VGND.t2689 XA.XIR[0].XIC[3].icell.PUM VPWR.t1437 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X253 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X254 VPWR.t661 XThC.XTB6.Y a_5949_9615# VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VPWR.t418 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X256 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X257 VPWR.t1206 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t1205 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X258 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t1125 VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X259 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X260 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t245 VGND.t2630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X261 VGND.t663 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X262 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X263 VGND.t1520 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t1519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t2373 XThR.XTB7.B a_n1335_8107# VGND.t2367 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VPWR.t1109 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t1108 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X266 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t1458 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X267 VPWR.t348 VPWR.t346 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t347 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X268 VGND.t1522 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t1521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X269 VGND.t665 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X270 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t1111 VPWR.t1110 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X271 XThC.XTB4.Y.t0 XThC.XTB7.B VPWR.t508 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X272 VGND.t1966 VGND.t1964 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1965 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X273 VGND.t613 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X274 VPWR.t345 VPWR.t343 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X275 XThR.Tn[2].t2 XThR.XTB3.Y.t3 VGND.t1151 VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X276 VGND.t1829 XThR.XTBN.Y a_n997_2891# VGND.t1778 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 VPWR.t613 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X278 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t138 VGND.t1367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X279 VPWR.t892 XThR.XTB5.Y XThR.Tn[12].t3 VPWR.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t1194 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X281 VGND.t1556 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t667 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X283 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t2581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X284 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t25 VGND.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X285 VGND.t1828 XThR.XTBN.Y XThR.Tn[6].t11 VGND.t1827 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1578 VGND.t1577 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X287 VPWR.t1341 XThR.XTBN.Y XThR.Tn[9].t10 VPWR.t1327 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t171 VGND.t1664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X289 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t1783 VPWR.t1782 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X290 VGND.t1963 VGND.t1961 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X291 XA.XIR[14].XIC_15.icell.PUM VPWR.t341 XA.XIR[14].XIC_15.icell.Ien VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X292 a_n997_715# XThR.XTBN.Y VGND.t1826 VGND.t1825 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X293 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X294 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t1395 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XThC.Tn[1].t6 XThC.XTBN.Y.t19 VGND.t322 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 VPWR.t1208 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t1207 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X297 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X298 XThR.Tn[14].t3 XThR.XTB7.Y VPWR.t1151 VPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t389 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X300 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t254 VGND.t2685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X301 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t198 VGND.t2035 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t212 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X303 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t255 VGND.t2686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X304 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t1455 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X305 VGND.t669 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X306 VGND.t671 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X308 VPWR.t1113 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t1112 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X309 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X310 VPWR.t890 XThR.XTB5.Y a_n1049_6405# VPWR.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X311 VPWR.t1240 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1239 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X312 XThR.XTB7.B data[6].t0 VPWR.t528 VPWR.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X313 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t600 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X314 VPWR.t1669 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t129 VGND.t1353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X316 VGND.t673 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t672 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X317 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t1913 VPWR.t1912 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X318 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t338 VPWR.t340 VPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 VGND.t44 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t1459 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X321 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t1660 VGND.t1659 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X322 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t128 VGND.t1352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X323 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t1713 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t169 VGND.t1657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X325 VGND.t675 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X326 XA.XIR[15].XIC[13].icell.Ien VPWR.t335 VPWR.t337 VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X327 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t140 VGND.t1369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X328 VPWR.t556 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X329 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X330 VPWR.t1915 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X331 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X332 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t7 VPWR.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X333 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t32 VGND.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X334 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t1769 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X335 VGND.t323 XThC.XTBN.Y.t20 XThC.Tn[4].t11 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X336 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t1653 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X337 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t112 VGND.t1106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X338 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t42 VGND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t333 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X340 VGND.t1960 VGND.t1958 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1959 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X341 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X342 VGND.t2352 data[1].t1 a_8739_10571# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 XA.XIR[0].XIC[1].icell.PDM VGND.t1955 VGND.t1957 VGND.t1956 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X344 VPWR.t409 XThR.XTB2.Y XThR.Tn[9].t3 VPWR.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND.t1824 XThR.XTBN.Y XThR.Tn[7].t6 VGND.t1823 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VGND.t2018 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t2017 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X347 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t174 VGND.t1668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X348 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X349 XThR.Tn[13].t11 XThR.XTBN.Y VPWR.t1340 VPWR.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X350 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X351 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t124 VGND.t1158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X352 VGND.t677 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X353 VGND.t1954 VGND.t1952 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t1917 VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X355 VPWR.t1403 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1402 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X356 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t330 VPWR.t332 VPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X357 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t1703 VPWR.t1702 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 VPWR.t1895 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t1894 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X359 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t1097 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X360 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t327 VPWR.t329 VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X361 VPWR.t558 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t557 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X362 VGND.t232 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X363 VGND.t1673 XThR.XTB6.Y XThR.Tn[5].t3 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X365 XThR.Tn[9].t6 XThR.XTB2.Y a_n997_3755# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 VGND.t679 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X367 XThR.XTB6.Y XThR.XTB6.A VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X368 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t216 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X369 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t39 VGND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X370 a_n997_1579# XThR.XTBN.Y VGND.t1822 VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 VGND.t548 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X372 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t116 VGND.t1123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X373 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t2637 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X374 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t2638 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 VPWR.t1809 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t1808 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X376 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t325 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X377 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t2356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X378 VPWR.t1785 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t1784 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X379 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t428 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X380 XA.XIR[15].XIC[6].icell.Ien VPWR.t322 VPWR.t324 VPWR.t323 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X381 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t218 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X382 VGND.t681 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X383 VPWR.t1705 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t1704 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X384 VPWR.t1919 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t1170 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X386 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t1860 VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X387 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t308 VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X388 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t2583 VGND.t2582 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t1172 VGND.t1171 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t2536 VGND.t2535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 VPWR.t944 XThR.XTBN.A XThR.XTBN.Y VPWR.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X392 VPWR.t560 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X393 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X394 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t1452 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X395 VPWR.t1811 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t1810 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X396 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t241 VGND.t2438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X397 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t500 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X398 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t1453 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t320 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 a_3523_10575# XThC.XTB7.B VGND.t246 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X401 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t626 VGND.t625 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X402 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t628 VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t1456 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t27 VGND.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X405 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t1261 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X406 VPWR.t583 XThC.XTBN.Y.t21 XThC.Tn[13].t11 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X408 VGND.t683 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X409 VGND.t2010 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t2009 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X410 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t1707 VPWR.t1706 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X411 XThC.Tn[5].t3 XThC.XTB6.Y VGND.t402 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t542 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X414 VGND.t1174 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X415 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t2639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X416 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t1813 VPWR.t1812 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X417 VPWR.t1815 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t1814 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X418 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t1985 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X419 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t7 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 VPWR.t1492 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t1491 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X421 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t2332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X422 VPWR.t615 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t614 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X423 XA.XIR[15].XIC[1].icell.Ien VPWR.t317 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X424 VGND.t685 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X425 VGND.t927 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t926 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t314 VPWR.t316 VPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X427 VGND.t1694 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X428 VGND.t340 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t10 VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 XThC.Tn[4].t10 XThC.XTBN.Y.t22 VGND.t324 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VPWR.t1127 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t1126 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X432 a_n1049_5317# XThR.XTB7.Y VPWR.t1149 VPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t1494 VPWR.t1493 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X434 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t48 VGND.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X435 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t2585 VGND.t2584 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X436 VGND.t929 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t928 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VGND.t1951 VGND.t1949 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VPWR.t1921 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X439 VPWR.t828 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t827 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 XThC.XTB6.Y XThC.XTB7.B VGND.t244 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VPWR.t313 VPWR.t311 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X442 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t1175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X443 VPWR.t1017 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t1016 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X444 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t1176 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X445 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t1376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X447 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t2168 VGND.t2167 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X448 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t150 VGND.t1461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X450 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X451 XThC.Tn[13].t3 XThC.XTB6.Y VPWR.t660 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X452 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t86 VGND.t761 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X453 VGND.t325 XThC.XTBN.Y.t24 XThC.Tn[0].t7 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 XThR.Tn[3].t10 XThR.XTBN.Y a_n1049_6699# VPWR.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t2340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X456 VGND.t234 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X457 VGND.t2026 XThR.XTB4.Y.t3 XThR.Tn[3].t11 VGND.t1348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t2640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X459 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t2170 VGND.t2169 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X460 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t787 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t97 VGND.t895 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X462 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X463 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t2342 VGND.t2341 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t2 VGND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X465 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t1178 VGND.t1177 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X466 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t54 VGND.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X467 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t369 VGND.t368 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X468 VGND.t931 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t930 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X469 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t1709 VPWR.t1708 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X470 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X471 VGND.t933 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t932 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X472 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t220 VGND.t2264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X473 XThR.Tn[11].t10 XThR.XTB4.Y.t4 VPWR.t1464 VPWR.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X474 VGND.t342 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X475 VGND.t267 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 XThC.Tn[14].t7 XThC.XTB7.Y a_10915_9569# VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 VPWR.t1129 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t1128 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X478 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t1817 VPWR.t1816 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X479 VGND.t19 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X480 VPWR.t1714 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t1713 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X481 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t2333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X482 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t1166 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X483 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t1179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X484 VPWR.t310 VPWR.t308 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X485 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t824 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X486 VGND.t2249 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VPWR.t1867 XThC.XTB2.Y XThC.Tn[9].t6 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X488 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t562 VPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X489 VGND.t1382 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t1381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X490 VGND.t935 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t934 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X491 VGND.t1181 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t1180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X492 VPWR.t888 XThR.XTB5.Y XThR.Tn[12].t2 VPWR.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VGND.t550 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X494 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t3 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X495 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X496 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t1923 VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X498 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t2675 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X499 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t2676 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 VPWR.t1147 XThR.XTB7.Y XThR.Tn[14].t2 VPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t2172 VGND.t2171 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X502 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t2071 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X503 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t788 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X504 XThR.Tn[8].t3 XThR.XTB1.Y.t4 a_n997_3979# VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t1770 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X506 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t2344 VGND.t2343 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 VGND.t695 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t1183 VGND.t1182 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 VPWR.t1019 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t1018 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X510 VPWR.t1622 data[2].t0 XThC.XTB7.B VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X511 VGND.t1948 VGND.t1946 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1947 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X512 VPWR.t554 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t553 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X513 VGND.t2520 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t2519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X514 XThC.Tn[13].t6 XThC.XTB6.Y a_10051_9569# VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X515 XThR.Tn[4].t11 XThR.XTBN.Y a_n1049_6405# VPWR.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t1738 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X517 VGND.t937 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t936 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X518 XThC.Tn[8].t3 XThC.XTBN.Y.t25 VPWR.t585 VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X519 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t2073 VGND.t2072 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X520 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t371 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X523 VGND.t1629 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1628 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X524 VGND.t939 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X525 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t1897 VPWR.t1896 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X526 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t2335 VGND.t2334 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X528 VGND.t615 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t941 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t940 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X530 VGND.t943 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 XThC.Tn[8].t10 XThC.XTB1.Y.t4 a_7651_9569# VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 XThC.Tn[13].t10 XThC.XTBN.Y.t26 VPWR.t586 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X533 VGND.t1384 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t1383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X534 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t619 VPWR.t618 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X535 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t95 VGND.t893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X536 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t96 VGND.t894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 VPWR.t1436 VGND.t2690 XA.XIR[0].XIC[9].icell.PUM VPWR.t1435 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X538 VGND.t401 XThC.XTB6.Y XThC.Tn[5].t2 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t501 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X540 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t305 VPWR.t307 VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X541 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t1300 VGND.t1299 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X542 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t1302 VGND.t1301 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t2074 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X544 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t1226 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X545 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t523 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 VGND.t945 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X548 VGND.t2012 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t2011 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X549 a_n1049_5611# XThR.XTB6.Y VPWR.t1253 VPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 XA.XIR[13].XIC_15.icell.PUM VPWR.t303 XA.XIR[13].XIC_15.icell.Ien VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X551 XThR.Tn[10].t6 XThR.XTB3.Y.t4 a_n997_2891# VGND.t1492 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X552 VGND.t947 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t946 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X553 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1460 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X554 VGND.t72 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X555 VGND.t552 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VPWR.t588 XThC.XTBN.Y.t27 XThC.Tn[7].t2 VPWR.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t2677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X558 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t2173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 VPWR.t1472 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X560 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t301 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X561 VPWR.t407 XThR.XTB2.Y XThR.Tn[9].t2 VPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X563 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X564 VGND.t949 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X565 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t1925 VPWR.t1924 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X566 VGND.t1524 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X567 VPWR.t1058 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t1057 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X568 VPWR.t1021 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t1020 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X569 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t2375 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X570 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1242 VPWR.t1241 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X571 VGND.t951 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X572 VGND.t617 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t616 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X573 XA.XIR[15].XIC_15.icell.Ien VPWR.t298 VPWR.t300 VPWR.t299 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X574 VPWR.t1474 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1473 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X575 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X576 VPWR.t566 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X577 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t7 VPWR.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X578 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t2046 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X579 XThC.Tn[0].t6 XThC.XTBN.Y.t29 VGND.t326 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 VGND.t2466 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t2465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X581 VPWR.t297 VPWR.t295 XA.XIR[9].XIC_15.icell.PUM VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X582 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t2377 VGND.t2376 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X583 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t2379 VGND.t2378 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X584 VGND.t2468 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t2467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X585 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t3 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X586 XThR.Tn[0].t0 XThR.XTB1.Y.t5 VGND.t186 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X587 VGND.t1821 XThR.XTBN.Y XThR.Tn[5].t10 VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X588 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t50 VGND.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X589 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t568 VPWR.t567 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X590 VGND.t2470 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t2469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X591 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t1502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X593 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t1147 VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X594 VGND.t2472 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t2471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X595 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X596 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t2038 VGND.t2037 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X597 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t16 VGND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X598 VGND.t1185 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t1184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X599 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t2678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X600 VGND.t1820 XThR.XTBN.Y XThR.Tn[4].t7 VGND.t1819 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X601 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t1304 VGND.t1303 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X602 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X603 VGND.t1187 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t1186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t7 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X605 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t432 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 VGND.t2474 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t2473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X607 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t82 VGND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X608 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t293 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X609 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X610 VGND.t2476 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t2475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X611 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t2380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X612 VGND.t2014 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t2013 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X613 VGND.t2224 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t2223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X614 VGND.t2478 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t2477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X615 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1244 VPWR.t1243 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X616 VGND.t21 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X617 VPWR.t1060 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t1059 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X618 VGND.t2480 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t2479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X619 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X620 VGND.t93 XThC.XTBN.Y.t31 a_8739_9569# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X621 VGND.t76 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X622 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X623 VGND.t2482 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t2481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X624 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t1716 VPWR.t1715 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X625 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t1482 VPWR.t1481 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X626 VGND.t2484 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t2483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X627 VGND.t344 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X628 VGND.t269 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X629 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1246 VPWR.t1245 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X630 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t1149 VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t111 VGND.t1105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X632 a_9827_9569# XThC.XTBN.Y.t32 VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X633 VGND.t2486 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t2485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X634 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t33 VGND.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X635 VPWR.t1594 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t1593 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X636 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t2047 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X637 VPWR.t1740 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t1739 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X638 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t1189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X639 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t187 VGND.t1711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X640 VPWR.t1718 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t1717 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X641 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t1661 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X642 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t1306 VGND.t1305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X643 VPWR.t292 VPWR.t290 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X644 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t1190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X645 VGND.t2076 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X646 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t2382 VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X647 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t186 VGND.t1710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X648 XThR.XTB7.A data[5].t1 VPWR.t850 VPWR.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X649 VGND.t2522 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t2521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X650 VPWR.t452 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X651 VGND.t2436 XThC.XTBN.A XThC.XTBN.Y.t3 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X652 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t789 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X653 VPWR.t1737 XThR.XTB7.B XThR.XTB1.Y.t2 VPWR.t1736 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X654 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t6 VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t1984 VGND.t1983 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X656 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t1720 VPWR.t1719 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X657 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t60 VGND.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X658 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t1192 VGND.t1191 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t287 VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t107 VGND.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X661 VPWR.t1596 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t1595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X662 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t1168 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X663 XThC.Tn[7].t1 XThC.XTBN.Y.t33 VPWR.t439 VPWR.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X664 VGND.t2372 XThR.XTB7.B a_n1335_7243# VGND.t2371 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X665 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t1169 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X666 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X667 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t2384 VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X668 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t1194 VGND.t1193 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[12].XIC_15.icell.PUM VPWR.t285 XA.XIR[12].XIC_15.icell.Ien VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t2049 VGND.t2048 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X672 VGND.t2204 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t2203 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t602 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X674 VGND.t554 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X675 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t100 VGND.t900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X676 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1401 VPWR.t1400 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X677 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t249 VGND.t2642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X678 XThC.Tn[11].t8 XThC.XTB4.Y.t6 VPWR.t1670 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X679 VGND.t556 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X680 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t210 VGND.t2133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t282 VPWR.t284 VPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X682 a_n997_1803# XThR.XTBN.Y VGND.t1818 VGND.t1817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X683 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X684 XThR.Tn[3].t9 XThR.XTBN.Y a_n1049_6699# VPWR.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X685 VPWR.t663 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X686 VGND.t1816 XThR.XTBN.Y XThR.Tn[3].t5 VGND.t1780 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X687 VGND.t2488 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t2487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X688 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t1476 VPWR.t1475 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X689 VGND.t1196 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X690 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t1198 VGND.t1197 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X691 XThC.Tn[2].t2 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X692 VPWR.t1153 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t1152 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X693 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t1496 VPWR.t1495 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X694 VPWR.t1545 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X695 VPWR.t454 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X696 XThR.Tn[11].t11 XThR.XTB4.Y.t5 VPWR.t1465 VPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X697 VPWR.t281 VPWR.t279 XA.XIR[8].XIC_15.icell.PUM VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 VPWR.t1866 XThC.XTB2.Y a_3773_9615# VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t492 VPWR.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t277 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X701 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t1982 VGND.t1981 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X702 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t1843 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X703 VGND.t2490 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t2489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X704 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t2040 VGND.t2039 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 VGND.t619 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t618 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X706 VGND.t1945 VGND.t1943 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X707 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t406 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t149 VGND.t1405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X710 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1399 VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X711 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X712 VGND.t1200 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t1199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X713 VPWR.t1263 XThC.XTB6.A a_5949_10571# VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X714 VPWR.t1598 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t1597 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X715 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t1554 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X717 VGND.t898 XThR.XTB3.Y.t5 XThR.Tn[2].t1 VGND.t897 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X718 VPWR.t1616 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t1615 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X719 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1662 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X720 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t1227 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X721 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X722 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t2051 VGND.t2050 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t125 VGND.t1160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X724 XThC.XTBN.Y.t1 XThC.XTBN.A VPWR.t1747 VPWR.t1746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X725 VGND.t1309 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t1308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X726 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t1642 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X727 VGND.t2137 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t2136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X728 VGND.t1311 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t1310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X729 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t1478 VPWR.t1477 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X730 XThR.Tn[8].t0 XThR.XTB1.Y.t7 a_n997_3979# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 XA.XIR[6].XIC_15.icell.PUM VPWR.t275 XA.XIR[6].XIC_15.icell.Ien VPWR.t276 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X732 VGND.t2234 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t2233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X733 VGND.t1313 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t1312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X734 VGND.t2139 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t2138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t1315 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t1314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X736 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t1023 VPWR.t1022 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X737 VGND.t1202 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t1201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 VGND.t74 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X739 VGND.t78 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X740 VGND.t96 XThC.XTBN.Y.t35 a_9827_9569# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X741 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t391 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VPWR.t665 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t664 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X743 VPWR.t772 XThC.XTB7.Y XThC.Tn[14].t3 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X744 XThR.Tn[4].t10 XThR.XTBN.Y a_n1049_6405# VPWR.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X745 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X746 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t2587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X747 VGND.t1317 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t1316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X748 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t1480 VPWR.t1479 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X749 VGND.t1319 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t1318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X750 VPWR.t1209 XThR.XTB4.Y.t6 a_n1049_6699# VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X751 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t570 VPWR.t569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X752 VGND.t1321 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t1320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X753 VPWR.t1155 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t1154 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X754 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t1618 VPWR.t1617 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X755 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t667 VPWR.t666 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X756 VGND.t1323 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t1322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X757 VPWR.t1547 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t1546 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X758 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t208 VGND.t2075 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X759 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t1484 VPWR.t1483 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X760 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t1203 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X761 VPWR.t1062 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t1061 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X762 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X763 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t1204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X764 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t1157 VPWR.t1156 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X765 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X766 VGND.t1325 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t1324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X767 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t71 VGND.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X768 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t153 VGND.t1490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X769 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t312 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X770 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1397 VPWR.t1396 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X771 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t2374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 VGND.t1327 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t1326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X773 VPWR.t1337 XThR.XTBN.Y XThR.Tn[8].t7 VPWR.t1336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X774 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t385 VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X775 XThR.Tn[10].t11 XThR.XTB3.Y.t6 a_n997_2891# VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X776 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t1819 VPWR.t1818 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X777 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t1771 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X778 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t506 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X779 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t244 VGND.t2606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X780 VGND.t1329 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t1328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X781 VGND.t1942 VGND.t1940 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X782 VGND.t1331 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t1330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X783 VPWR.t1262 XThC.XTB6.A XThC.XTB2.Y VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X784 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t1560 VGND.t1559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X785 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t1562 VGND.t1561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X786 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t75 VGND.t658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X787 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t387 VPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X788 VGND.t1333 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t1332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X789 VGND.t2226 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t2225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X790 VGND.t2109 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t2108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X791 XThR.XTB3.Y.t0 XThR.XTB7.A VPWR.t774 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X792 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t132 VGND.t1356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X793 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X794 VGND.t80 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X795 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X796 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t1206 VGND.t1205 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X797 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t1501 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X798 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X799 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X800 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t1081 VPWR.t1080 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X801 VGND.t442 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X802 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t14 VGND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X803 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t1159 VPWR.t1158 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 XThR.Tn[0].t10 XThR.XTBN.Y VGND.t1815 VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X805 VPWR.t886 XThR.XTB5.Y a_n1049_6405# VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X806 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t1549 VPWR.t1548 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 VGND.t444 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X808 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t247 VGND.t2632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X809 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t2042 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X810 XThC.Tn[10].t10 XThC.XTB3.Y.t4 VPWR.t1711 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X812 VPWR.t1335 XThR.XTBN.Y XThR.Tn[10].t10 VPWR.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X814 VPWR.t1196 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t1195 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X815 VPWR.t441 XThC.XTBN.Y.t36 XThC.Tn[13].t9 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X816 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X817 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t2052 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X818 a_3773_9615# XThC.XTB2.Y VPWR.t1865 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XThC.Tn[5].t1 XThC.XTB6.Y VGND.t400 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X820 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t202 VGND.t2045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X821 XThC.Tn[2].t10 XThC.XTB3.Y.t5 VGND.t2336 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 VPWR.t1064 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t1063 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X823 VPWR.t1395 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1394 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X824 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t105 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X825 VGND.t2524 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t2523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X826 VPWR.t1899 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t1898 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t137 VGND.t1366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X828 VPWR.t962 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t961 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X829 VGND.t1814 XThR.XTBN.Y a_n997_3755# VGND.t1803 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X830 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t430 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X831 VPWR.t1498 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t1497 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t409 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X833 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t1208 VGND.t1207 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X834 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t2589 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X835 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t1083 VPWR.t1082 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X836 VGND.t446 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X837 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X838 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t227 VGND.t2353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X839 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t1564 VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X840 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t34 VGND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X841 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t1732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X842 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t123 VGND.t1156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X843 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t1525 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X844 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t78 VGND.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 VGND.t2619 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t2618 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X846 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t1210 VGND.t1209 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X847 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t80 VGND.t742 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t919 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X849 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X850 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t61 VGND.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X853 a_5155_9615# XThC.XTB5.Y VPWR.t782 VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X854 XA.XIR[5].XIC_15.icell.PUM VPWR.t273 XA.XIR[5].XIC_15.icell.Ien VPWR.t274 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X855 VPWR.t1198 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t1197 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X856 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t2680 VGND.t2679 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X857 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t851 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X858 VGND.t2236 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t2235 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X859 XA.XIR[9].XIC_15.icell.PUM VPWR.t271 XA.XIR[9].XIC_15.icell.Ien VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X860 VGND.t2251 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t2250 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X861 VPWR.t1393 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X862 VPWR.t1901 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t1900 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X863 VGND.t1212 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X864 XThC.Tn[8].t7 XThC.XTB1.Y.t7 VPWR.t1500 VPWR.t1499 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X865 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t1551 VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X866 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t1066 VPWR.t1065 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X867 VGND.t756 XThR.XTB5.Y XThR.Tn[4].t3 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X868 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t7 VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X869 VGND.t1214 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t1213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X870 VPWR.t1068 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1067 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X871 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X872 VPWR.t1391 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1390 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X873 XThR.XTB5.Y XThR.XTB5.A VGND.t1491 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X874 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t1566 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X875 VPWR.t1903 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t1902 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X876 VPWR.t1085 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X877 VPWR.t964 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t963 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X878 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t1772 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X879 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t1666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X880 VPWR.t270 VPWR.t268 XA.XIR[1].XIC_15.icell.PUM VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X881 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t2134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X882 VPWR.t267 VPWR.t265 XA.XIR[5].XIC_15.icell.PUM VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X883 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X884 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t2682 VGND.t2681 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X885 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t1087 VPWR.t1086 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X886 VGND.t448 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X887 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t179 VGND.t1678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X888 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 VGND.t450 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X890 VGND.t1217 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t1216 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X891 VGND.t452 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X892 VGND.t1526 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t1525 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VPWR.t264 VPWR.t262 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X894 XThC.Tn[14].t6 XThC.XTB7.Y a_10915_9569# VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X895 XThC.XTB3.Y.t2 XThC.XTB7.A a_4387_10575# VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X896 a_n997_1803# XThR.XTBN.Y VGND.t1813 VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X897 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t434 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X898 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1070 VPWR.t1069 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X899 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t2591 VGND.t2590 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X900 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t3 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X901 VGND.t2238 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t176 VGND.t1674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X903 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t373 VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 VGND.t454 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X905 VGND.t82 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 VPWR.t1723 XThC.XTB5.A XThC.XTB1.Y.t1 VPWR.t1722 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X907 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t1218 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X908 VGND.t84 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X909 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t1219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X910 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t1360 VGND.t1359 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X911 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 VGND.t456 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X913 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t1553 VPWR.t1552 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X914 VGND.t458 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X915 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1072 VPWR.t1071 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X916 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X917 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t260 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X918 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1389 VPWR.t1388 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X919 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t57 VGND.t537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X920 VGND.t2337 XThC.XTB3.Y.t6 XThC.Tn[2].t11 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X921 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1215 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X922 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t4 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t647 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X924 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X925 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t1540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X926 a_n1319_6405# XThR.XTB5.A VPWR.t1135 VPWR.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X927 VPWR.t623 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t622 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X928 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t1538 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t826 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X930 VPWR.t259 VPWR.t257 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X931 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t94 VGND.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X932 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t1502 VPWR.t1501 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X933 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t1161 VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X934 VGND.t460 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X935 VGND.t462 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X936 XThR.Tn[12].t10 XThR.XTBN.Y VPWR.t1333 VPWR.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X937 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t2145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X938 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t254 VPWR.t256 VPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X939 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t30 VGND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X940 XThC.Tn[11].t3 XThC.XTBN.Y.t39 VPWR.t445 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X941 VGND.t1715 data[4].t2 XThR.XTB5.A VGND.t1714 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X942 XThR.XTBN.Y XThR.XTBN.A VGND.t904 VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X943 VGND.t1351 data[3].t0 XThC.XTBN.A VGND.t1350 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X944 VGND.t464 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X945 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t1221 VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X946 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t649 VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X947 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t7 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X948 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X949 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t211 VGND.t2144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X950 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t1223 VGND.t1222 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t55 VGND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X952 a_n997_2667# XThR.XTBN.Y VGND.t1811 VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X953 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t252 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t253 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X954 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t83 VGND.t758 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X955 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t1441 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X956 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t1362 VGND.t1361 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X957 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t1539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X958 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t1844 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X959 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t1505 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t1611 VGND.t1610 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 VPWR.t625 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X962 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t651 VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 VGND.t558 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t189 VGND.t1716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X966 XThC.Tn[4].t6 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X967 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t1541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X968 VGND.t1225 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t1224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 VPWR.t456 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t455 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X970 VPWR.t1331 XThR.XTBN.Y XThR.Tn[8].t6 VPWR.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X971 VGND.t271 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X972 VGND.t346 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X974 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t525 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X975 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t249 VPWR.t251 VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X976 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t9 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X977 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X978 VGND.t466 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X979 VPWR.t781 XThC.XTB5.Y XThC.Tn[12].t1 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t1226 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X981 VPWR.t1180 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t1179 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X982 VPWR.t248 VPWR.t246 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t247 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X983 VGND.t2440 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t2439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X984 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t1905 VPWR.t1904 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X985 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t966 VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X986 VGND.t1597 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t1596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X987 VGND.t1810 XThR.XTBN.Y XThR.Tn[1].t11 VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X988 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t377 VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X989 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t921 VGND.t920 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X990 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t669 VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X991 VPWR.t1434 VGND.t2691 XA.XIR[0].XIC[7].icell.PUM VPWR.t1433 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X992 VPWR.t245 VPWR.t243 XA.XIR[4].XIC_15.icell.PUM VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X993 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t1163 VPWR.t1162 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X994 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X995 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t2183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X996 VGND.t2442 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t2441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X997 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t1988 VGND.t1987 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X998 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t1500 VGND.t1499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 a_9827_9569# XThC.XTBN.Y.t41 VGND.t97 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1000 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t1845 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1001 XThR.Tn[9].t9 XThR.XTBN.Y VPWR.t1329 VPWR.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1002 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t653 VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1003 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t923 VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1004 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t2070 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1006 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t173 VGND.t1667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1007 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t1514 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1008 XThC.Tn[1].t2 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1009 VGND.t2621 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t2620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1010 XThR.Tn[0].t9 XThR.XTBN.Y VGND.t1809 VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1011 XThC.Tn[13].t5 XThC.XTB6.Y a_10051_9569# VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1012 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1013 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t1986 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1014 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t1672 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1015 VPWR.t1328 XThR.XTBN.Y XThR.Tn[10].t9 VPWR.t1327 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1016 VPWR.t671 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1017 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1018 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t1613 VGND.t1612 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t240 VPWR.t242 VPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1020 XA.XIR[0].XIC[12].icell.PDM VGND.t1937 VGND.t1939 VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1021 VGND.t2141 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t2140 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 VGND.t2240 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2239 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 VGND.t2444 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t2443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1024 VGND.t2446 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t2445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1025 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t1907 VPWR.t1906 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1026 VPWR.t771 XThC.XTB7.Y a_6243_9615# VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t209 VGND.t2120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1028 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t1228 VGND.t1227 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1029 VGND.t2242 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1030 VGND.t1599 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t1598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1031 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t1620 VPWR.t1619 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1032 VGND.t2253 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t2252 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VPWR.t1432 VGND.t2692 XA.XIR[0].XIC[11].icell.PUM VPWR.t1431 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1034 VGND.t2206 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t2205 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t1296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1036 VGND.t1230 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t1229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 VGND.t98 XThC.XTBN.Y.t43 a_8963_9569# VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1038 VGND.t2448 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t2447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1039 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t1555 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1040 VPWR.t494 XThR.XTB1.Y.t8 XThR.Tn[8].t1 VPWR.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1041 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t238 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1042 VGND.t2450 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t2449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1043 VGND.t2452 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t2451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1044 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t1909 VPWR.t1908 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1045 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t237 VGND.t2402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1046 VGND.t2228 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t2227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1047 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t1089 VPWR.t1088 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1048 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t968 VPWR.t967 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 VGND.t2111 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t2110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1050 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t925 VGND.t924 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1051 XThR.XTBN.A data[7].t0 VPWR.t1079 VPWR.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1052 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t673 VPWR.t672 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t1224 VPWR.t1223 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1054 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t38 VGND.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1055 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1056 VPWR.t1430 VGND.t2693 XA.XIR[0].XIC[2].icell.PUM VPWR.t1429 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1057 VPWR.t405 XThR.XTB2.Y a_n1049_7787# VPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1058 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1059 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1060 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t973 VPWR.t972 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1061 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t2184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1062 VPWR.t1182 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t1181 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1063 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t58 VGND.t538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1065 XA.XIR[0].XIC[10].icell.PDM VGND.t1934 VGND.t1936 VGND.t1935 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1066 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t980 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1067 VGND.t2454 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t2453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1068 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t6 VPWR.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1069 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t155 VGND.t1506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1070 VGND.t1991 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1071 XThC.Tn[8].t6 XThC.XTB1.Y.t10 VPWR.t1504 VPWR.t1503 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1072 VPWR.t1046 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1073 VPWR.t237 VPWR.t235 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1074 VGND.t1933 VGND.t1931 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1932 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1075 VGND.t2078 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1076 XThR.Tn[0].t1 XThR.XTB1.Y.t9 VGND.t187 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1077 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1078 VGND.t2456 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t2455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1079 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 VPWR.t597 XThR.XTB3.Y.t8 XThR.Tn[10].t1 VPWR.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1081 VGND.t2526 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t2525 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1082 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1083 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t22 VGND.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1085 VPWR.t1864 XThC.XTB2.Y a_3773_9615# VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1086 VGND.t2230 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t2229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 VGND.t1808 XThR.XTBN.Y XThR.Tn[4].t6 VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1088 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t233 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1089 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t40 VGND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1090 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t1298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1092 VPWR.t447 XThC.XTBN.Y.t44 XThC.Tn[9].t3 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1093 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1094 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t799 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1095 VGND.t99 XThC.XTBN.Y.t45 XThC.Tn[5].t9 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1096 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t1543 VGND.t1542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1097 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1098 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t170 VGND.t1663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1099 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t41 VGND.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1100 VGND.t1806 XThR.XTBN.Y a_n997_1579# VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1101 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t1526 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1102 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t230 VGND.t2358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1103 VGND.t2458 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t2457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1104 VGND.t2460 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t2459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1105 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t1 VPWR.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1106 VGND.t273 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1107 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1108 VGND.t348 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1109 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t641 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1110 VPWR.t1184 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t1183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1111 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1112 XThC.Tn[12].t6 XThC.XTB5.Y a_9827_9569# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1114 VPWR.t1048 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t1047 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1115 XThR.XTB6.A data[5].t2 VPWR.t996 VPWR.t995 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1116 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t235 VGND.t2400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1117 VPWR.t232 VPWR.t230 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1118 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t1498 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1119 VPWR.t627 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1120 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t7 VPWR.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1121 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1186 VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1122 VGND.t2462 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t2461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1123 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t201 VGND.t2044 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1124 XA.XIR[15].XIC[12].icell.Ien VPWR.t227 VPWR.t229 VPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1125 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t157 VGND.t1508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1126 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t5 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1127 VPWR.t840 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1128 VPWR.t846 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1129 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t800 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1130 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t1233 VGND.t1232 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1131 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t982 VGND.t981 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1132 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t791 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1133 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t802 VGND.t801 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1134 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t92 VGND.t810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1135 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t98 VGND.t896 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1136 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t1235 VGND.t1234 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t1773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t159 VGND.t1510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1139 a_6243_9615# XThC.XTB7.Y VPWR.t770 VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1140 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t225 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1141 VGND.t1930 VGND.t1928 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1142 XThC.Tn[10].t11 XThC.XTBN.Y.t47 VPWR.t1869 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1143 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1144 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t1545 VGND.t1544 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1146 VGND.t2113 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1147 XA.XIR[1].XIC_15.icell.PUM VPWR.t223 XA.XIR[1].XIC_15.icell.Ien VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1148 XThC.Tn[10].t5 XThC.XTB3.Y.t8 a_8739_9569# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1149 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t644 VGND.t643 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 VGND.t531 XThC.XTB7.Y XThC.Tn[6].t3 VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1151 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t93 VGND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1152 VGND.t1237 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t1236 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1153 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t1239 VGND.t1238 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 XThR.Tn[11].t8 XThR.XTBN.Y VPWR.t1325 VPWR.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1155 VGND.t2208 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t2207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1156 VPWR.t1870 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 VGND.t1241 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t1240 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XA.XIR[15].XIC[10].icell.Ien VPWR.t220 VPWR.t222 VPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1159 VGND.t2464 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t2463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1160 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t458 VPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1188 VPWR.t1187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1162 VGND.t1243 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t1242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1163 VPWR.t970 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1164 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1165 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t217 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VPWR.t848 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1167 VGND.t2407 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t2406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1168 VGND.t2409 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t2408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1169 VGND.t1601 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1170 VGND.t2411 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t2410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1171 VGND.t1375 XThC.XTB7.A XThC.XTB7.Y VGND.t1374 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1172 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t804 VGND.t803 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1173 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1387 VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1174 VPWR.t842 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1175 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t6 VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t9 VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1177 a_n997_2667# XThR.XTBN.Y VGND.t1805 VGND.t1760 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1178 VPWR.t629 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t628 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1179 VPWR.t998 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1180 a_7875_9569# XThC.XTBN.Y.t49 VGND.t2650 VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1181 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t984 VGND.t983 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1182 VGND.t2528 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t2527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1183 VGND.t1804 XThR.XTBN.Y a_n997_3979# VGND.t1803 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1184 VGND.t2538 Vbias.t1 Vbias.t2 VGND.t2537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X1185 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t975 VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1186 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t250 VGND.t2643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1187 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1188 XThC.Tn[14].t10 XThC.XTBN.Y.t50 VPWR.t1871 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1189 a_n1049_6699# XThR.XTB4.Y.t7 VPWR.t1210 VPWR.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t3 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1191 VGND.t2413 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t2412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1192 VGND.t2080 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1193 VGND.t2415 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t2414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1194 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t460 VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1195 XThC.Tn[2].t9 XThC.XTB3.Y.t9 VGND.t1365 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1196 XThC.Tn[9].t2 XThC.XTBN.Y.t52 VPWR.t1872 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1197 XThC.Tn[5].t8 XThC.XTBN.Y.t53 VGND.t2651 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1199 VGND.t2417 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t2416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1200 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t1110 VGND.t1109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1201 VGND.t86 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1202 XA.XIR[15].XIC[5].icell.Ien VPWR.t214 VPWR.t216 VPWR.t215 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1203 VGND.t1927 VGND.t1925 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1926 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1204 VPWR.t989 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1205 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t1244 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1206 XThC.Tn[0].t0 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t1873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1207 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1208 VPWR.t952 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t951 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1209 VPWR.t1000 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1210 XThR.Tn[12].t1 XThR.XTB5.Y VPWR.t884 VPWR.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1211 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t1556 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1212 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t1527 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1213 VGND.t2419 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t2418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1214 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t212 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1215 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t59 VGND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1216 VGND.t2232 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t2231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1217 XThR.Tn[6].t10 XThR.XTBN.Y VGND.t1802 VGND.t1801 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1218 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t6 VPWR.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1219 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 VGND.t1800 XThR.XTBN.Y a_n997_2891# VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 VGND.t2370 XThR.XTB7.B XThR.XTB7.Y VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1222 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1385 VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1223 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t91 VGND.t809 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1224 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1225 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t1547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1226 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t631 VPWR.t630 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1227 VPWR.t633 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t632 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1228 VGND.t1246 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t1245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1229 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t605 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1230 VPWR.t1002 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 a_n997_2667# XThR.XTB4.Y.t8 XThR.Tn[11].t4 VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1232 VPWR.t211 VPWR.t209 XA.XIR[12].XIC_15.icell.PUM VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1233 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t89 VGND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1234 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t1050 VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1235 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t206 VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1236 VGND.t2421 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t2420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1237 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t1153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1238 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t18 VGND.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1239 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t1112 VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1240 VGND.t2423 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t2422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1241 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t203 VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1242 VGND.t2652 XThC.XTBN.Y.t55 XThC.Tn[1].t5 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1243 a_n1049_6405# XThR.XTB5.Y VPWR.t882 VPWR.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1244 VGND.t2425 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t2424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1245 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t462 VPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1246 VPWR.t916 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t915 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1247 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t985 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1248 VGND.t1924 VGND.t1922 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1249 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t1247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1250 VGND.t1249 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t1248 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1251 VPWR.t1052 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t1051 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1252 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t1617 VGND.t1616 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1253 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t1774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 VPWR.t1883 XThR.XTB1.Y.t10 XThR.Tn[8].t8 VPWR.t1882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1255 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t130 VGND.t1354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1257 VPWR.t1323 XThR.XTBN.Y XThR.Tn[7].t2 VPWR.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t201 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 VGND.t2648 XThC.XTB2.Y XThC.Tn[1].t11 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1260 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t199 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1261 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t45 VGND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1262 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t1548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1263 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t1874 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1264 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t646 VGND.t645 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1265 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t635 VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1266 VGND.t41 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 XThR.Tn[1].t6 XThR.XTBN.Y a_n1049_7787# VPWR.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1268 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t1619 VGND.t1618 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1269 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t178 VGND.t1677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1270 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1271 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 VGND.t2623 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t2622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1273 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t29 VGND.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1274 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t918 VPWR.t917 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1275 VGND.t2427 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t2426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1276 VGND.t2429 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t2428 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1277 VGND.t1921 VGND.t1919 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1920 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1278 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t1054 VPWR.t1053 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1279 VGND.t350 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1280 VGND.t906 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t905 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1281 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t637 VPWR.t636 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1282 XThR.Tn[9].t1 XThR.XTB2.Y VPWR.t403 VPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1283 XThR.Tn[7].t5 XThR.XTBN.Y VGND.t1798 VGND.t1797 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1284 VPWR.t971 data[1].t2 XThC.XTB6.A VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1285 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1645 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1286 VPWR.t920 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t919 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1287 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t1442 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1288 VPWR.t198 VPWR.t196 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1289 VGND.t2653 XThC.XTBN.Y.t57 a_7875_9569# VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1290 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1291 VPWR.t1321 XThR.XTBN.Y XThR.Tn[13].t10 VPWR.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1292 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t844 VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1293 VPWR.t195 VPWR.t193 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1294 VGND.t2255 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t2254 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1295 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1296 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t215 VGND.t2162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1297 VGND.t2431 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t2430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1298 VPWR.t823 XThR.XTB3.Y.t9 XThR.Tn[10].t3 VPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1299 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t954 VPWR.t953 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1300 VGND.t560 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1301 XThC.Tn[3].t2 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1303 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1304 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t1458 VPWR.t1457 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1305 XThR.Tn[5].t2 XThR.XTB6.Y VGND.t1672 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1306 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1307 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1308 VPWR.t1735 XThR.XTB7.B XThR.XTB4.Y.t0 VPWR.t1734 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1309 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t913 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1310 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t792 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1311 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t2084 VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1312 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1217 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1313 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t1251 VGND.t1250 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t1775 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t2617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1316 VGND.t1433 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t1432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1317 VGND.t2625 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t2624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 VPWR.t1056 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t1055 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1319 VGND.t1918 VGND.t1916 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1320 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t904 VPWR.t903 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1321 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1322 VGND.t1734 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t1733 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1323 VGND.t1435 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t1434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1324 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t590 VPWR.t589 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1325 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1326 VGND.t1993 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1327 VGND.t1437 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t1436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1328 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t2020 VGND.t2019 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1329 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t1253 VGND.t1252 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 VGND.t2257 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t2256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1331 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t675 VPWR.t674 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1332 VGND.t2210 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1333 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 VGND.t1439 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t1438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1335 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t956 VPWR.t955 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1336 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t147 VGND.t1397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1337 VPWR.t906 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1338 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1339 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1275 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1340 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1341 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t477 VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1342 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t479 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t1520 VPWR.t1519 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1344 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t10 VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1345 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t945 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1346 VGND.t1441 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t1440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1347 VGND.t1443 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t1442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1348 VGND.t2143 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t2142 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1349 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1350 VGND.t1255 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t1254 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1351 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1352 XThC.Tn[1].t4 XThC.XTBN.Y.t59 VGND.t2654 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1353 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1354 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 VPWR.t192 VPWR.t190 XA.XIR[15].XIC_15.icell.PUM VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1356 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1218 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1357 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t986 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1358 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t1460 VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1359 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t9 VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1360 VPWR.t1383 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1361 VGND.t1445 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t1444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1362 VGND.t1995 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1363 XA.XIR[15].XIC[14].icell.Ien VPWR.t187 VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1364 VGND.t1447 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t1446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1365 VPWR.t1099 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t1098 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1366 VGND.t2082 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1367 VPWR.t717 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t716 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1368 VPWR.t186 VPWR.t184 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 XThR.Tn[13].t5 XThR.XTB6.Y a_n997_1579# VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1370 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t5 VPWR.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1371 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t1162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1372 VPWR.t958 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1373 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t2021 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1374 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t1550 VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1375 VGND.t1449 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t1448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1376 VGND.t1451 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t1450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1377 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t191 VGND.t1730 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1378 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t2023 VGND.t2022 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1379 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t199 VGND.t2036 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1380 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1381 VGND.t1453 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t1452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1382 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t960 VPWR.t959 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1383 VGND.t1455 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t1454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1384 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t1387 VGND.t1386 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1385 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1386 VGND.t2181 data[2].t1 XThC.XTB7.B VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1388 VGND.t1796 XThR.XTBN.Y XThR.Tn[2].t10 VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1389 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t1552 VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1390 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t47 VGND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1391 a_n1049_5317# XThR.XTB7.Y VPWR.t1145 VPWR.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1392 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1393 VGND.t2655 XThC.XTBN.Y.t60 XThC.Tn[4].t9 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1394 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t1529 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1395 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1396 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t1257 VGND.t1256 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1397 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t200 VGND.t2043 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1398 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t214 VGND.t2161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1399 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t1530 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 VGND.t1457 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1401 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t436 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1402 VGND.t155 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1403 VGND.t157 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t216 VGND.t2179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1405 XThR.Tn[3].t1 XThR.XTB4.Y.t9 VGND.t1579 VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1406 VGND.t159 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1407 VPWR.t1381 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1408 VGND.t2115 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t2114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1409 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1410 VPWR.t719 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1411 VPWR.t769 XThC.XTB7.Y a_6243_9615# VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1412 VPWR.t659 XThC.XTB6.Y XThC.Tn[13].t2 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VPWR.t183 VPWR.t181 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1414 VGND.t1373 data[1].t3 XThC.XTB5.A VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1415 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t279 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1416 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1190 VPWR.t1189 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1417 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t915 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1418 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t1462 VPWR.t1461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1419 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t178 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 VGND.t161 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1421 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t85 VGND.t760 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1422 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t67 VGND.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1423 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1101 VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1424 VPWR.t530 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t529 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1425 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t1389 VGND.t1388 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1426 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1427 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t73 VGND.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1428 VGND.t2657 XThC.XTBN.Y.t61 XThC.Tn[7].t6 VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1429 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1554 VGND.t1553 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1430 VPWR.t1510 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1509 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1431 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t2024 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1432 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t121 VGND.t1154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1433 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t1258 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1434 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t281 VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1435 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t1776 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1436 XThR.Tn[12].t0 XThR.XTB5.Y VPWR.t880 VPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1437 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 a_10915_9569# XThC.XTBN.Y.t62 VGND.t2659 VGND.t2658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1439 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t217 VGND.t2180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1440 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1777 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1441 XThR.Tn[6].t9 XThR.XTBN.Y VGND.t1794 VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 VPWR.t806 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t805 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1443 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t2628 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1444 XThC.Tn[9].t5 XThC.XTB2.Y VPWR.t1863 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 VGND.t2530 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t2529 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1446 a_n997_2667# XThR.XTB4.Y.t10 XThR.Tn[11].t5 VGND.t978 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 VGND.t2627 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t2626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1448 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t381 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t333 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1450 VGND.t163 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1451 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t1192 VPWR.t1191 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1452 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t236 VGND.t2401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1453 VGND.t1260 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1454 VPWR.t1522 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t1521 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1455 VPWR.t532 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t531 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1456 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t908 VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1457 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t175 VPWR.t177 VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1458 VPWR.t1512 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1511 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1459 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t1261 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1460 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t946 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1461 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1462 VGND.t2368 XThR.XTB7.B a_n1335_8331# VGND.t2367 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1463 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t283 VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1465 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t917 VGND.t916 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1466 VGND.t2259 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t2258 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t1507 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1468 VPWR.t1875 XThC.XTBN.Y.t63 XThC.Tn[9].t1 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1469 XA.XIR[15].XIC_15.icell.PUM VPWR.t173 XA.XIR[15].XIC_15.icell.Ien VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t76 VGND.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1471 a_10051_9569# XThC.XTBN.Y.t64 VGND.t2385 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1472 VGND.t562 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1473 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t231 VGND.t2359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1474 VPWR.t1319 XThR.XTBN.Y XThR.Tn[7].t1 VPWR.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1475 VPWR.t808 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t807 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1476 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1557 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1477 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t171 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1478 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t101 VGND.t911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1479 VPWR.t1821 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t1820 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1480 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1481 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1482 XThC.Tn[11].t9 XThC.XTB4.Y.t8 VPWR.t1850 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1483 VGND.t1792 XThR.XTBN.Y XThR.Tn[1].t10 VGND.t1748 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1484 XThR.Tn[1].t5 XThR.XTBN.Y a_n1049_7787# VPWR.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1485 a_7651_9569# XThC.XTBN.Y.t65 VGND.t2386 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1486 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1487 VGND.t165 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1488 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1103 VPWR.t1102 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1489 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1220 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1490 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t510 VPWR.t509 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1491 VGND.t167 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1492 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t1263 VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 VPWR.t810 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1494 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1495 VPWR.t910 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1496 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1497 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t1390 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1498 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t1496 VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1499 a_n1049_5611# XThR.XTB6.Y VPWR.t1252 VPWR.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1500 XThR.Tn[9].t0 XThR.XTB2.Y VPWR.t401 VPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1501 VPWR.t170 VPWR.t168 XA.XIR[11].XIC_15.icell.PUM VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1502 VGND.t169 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1503 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1504 XThC.Tn[4].t8 XThC.XTBN.Y.t66 VGND.t2387 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 VGND.t1997 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1506 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t335 VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1507 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t383 VGND.t382 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1508 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t1847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 VPWR.t1317 XThR.XTBN.Y XThR.Tn[13].t9 VPWR.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1510 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t2593 VGND.t2592 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1379 VPWR.t1378 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1512 VGND.t1915 VGND.t1913 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1513 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t605 VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t233 VGND.t2361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1515 VPWR.t534 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1516 VGND.t1265 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t1264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 VPWR.t1514 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1513 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1518 VPWR.t1823 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t1822 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1276 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1521 VGND.t2672 XThR.XTB1.Y.t11 XThR.Tn[0].t11 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1522 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t1 VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1523 XThR.Tn[5].t9 XThR.XTBN.Y VGND.t1791 VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1524 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1525 XA.XIR[0].XIC[8].icell.PDM VGND.t1910 VGND.t1912 VGND.t1911 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1526 XA.XIR[0].XIC[14].icell.PDM VGND.t1907 VGND.t1909 VGND.t1908 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1527 VGND.t2366 XThR.XTB7.B XThR.XTB6.Y VGND.t2364 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1528 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t2388 XThC.XTBN.Y.t67 XThC.Tn[0].t5 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 VGND.t171 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1532 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t912 VPWR.t911 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1533 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t512 VPWR.t511 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1534 VGND.t173 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 VGND.t1641 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t1640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1536 VGND.t1011 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t1010 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1537 VGND.t2117 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t2116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1538 VGND.t2389 XThC.XTBN.Y.t68 XThC.Tn[3].t7 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 VGND.t175 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1540 VGND.t1603 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t1602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t2057 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t2056 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1542 VPWR.t1825 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1543 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1544 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1545 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t798 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1546 XThC.Tn[7].t5 XThC.XTBN.Y.t69 VGND.t2391 VGND.t2390 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 VPWR.t1741 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 VGND.t177 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1549 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t1105 VPWR.t1104 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1550 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t721 VPWR.t720 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1551 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t165 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1552 VGND.t179 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1553 VGND.t698 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1554 VGND.t1267 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t1266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1555 VGND.t908 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t907 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1556 VPWR.t399 XThR.XTB2.Y a_n1049_7787# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1557 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t514 VPWR.t513 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1558 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t2595 VGND.t2594 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VGND.t700 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1560 VGND.t702 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1561 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t115 VGND.t1122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1562 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1563 VGND.t2393 XThC.XTBN.Y.t71 a_10915_9569# VGND.t2392 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1564 VPWR.t1428 VGND.t2694 XA.XIR[0].XIC[4].icell.PUM VPWR.t1427 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1565 VPWR.t1627 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1566 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1567 VPWR.t1377 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t1013 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1569 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t223 VGND.t2267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1570 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t1171 VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1571 XThC.Tn[11].t10 XThC.XTB4.Y.t9 a_8963_9569# VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1572 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1573 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t1014 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1574 VPWR.t723 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t722 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1575 VGND.t2629 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1576 VGND.t704 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1577 XThR.Tn[14].t11 XThR.XTBN.Y VPWR.t1316 VPWR.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1578 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1579 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t163 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1580 a_7875_9569# XThC.XTBN.Y.t72 VGND.t2394 VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1581 VPWR.t1251 XThR.XTB6.Y XThR.Tn[13].t3 VPWR.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1582 VGND.t2532 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t2531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t793 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1584 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1585 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t182 VGND.t1689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1586 XA.XIR[0].XIC[3].icell.PDM VGND.t1904 VGND.t1906 VGND.t1905 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t1015 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t384 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1589 XThC.Tn[11].t11 XThC.XTB4.Y.t11 a_8963_9569# VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1590 VGND.t706 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1591 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t914 VPWR.t913 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1592 VGND.t708 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1593 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t725 VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1594 VGND.t1903 VGND.t1901 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1902 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1595 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t161 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1596 XThC.Tn[0].t8 XThC.XTB1.Y.t12 VGND.t1000 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1597 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t44 VGND.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1598 VGND.t2395 XThC.XTBN.Y.t73 a_10051_9569# VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1599 VGND.t2661 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t2660 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1600 VPWR.t1629 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t1628 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1601 VGND.t2119 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t2118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1602 XThR.XTB1.Y.t0 XThR.XTB5.A VPWR.t1133 VPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1603 VPWR.t1426 VGND.t2695 XA.XIR[0].XIC[0].icell.PUM VPWR.t1425 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1605 XThR.Tn[13].t4 XThR.XTB6.Y a_n997_1579# VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1606 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1607 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1608 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t1017 VGND.t1016 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1609 VGND.t576 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1610 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 VGND.t2396 XThC.XTBN.Y.t74 a_7651_9569# VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1612 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1516 VPWR.t1515 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1613 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t212 VGND.t2146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1614 XThC.XTBN.Y.t2 XThC.XTBN.A VGND.t2434 VGND.t2433 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1615 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t1631 VPWR.t1630 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t158 VPWR.t160 VPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1617 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t2086 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1618 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t166 VGND.t1654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1619 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1620 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1621 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1622 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1624 XA.XIR[0].XIC[7].icell.PDM VGND.t1898 VGND.t1900 VGND.t1899 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1625 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t6 VPWR.t1313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1626 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t1019 VGND.t1018 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t1090 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1629 VPWR.t1743 XThC.XTBN.Y.t75 XThC.Tn[7].t0 VPWR.t1742 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1630 VPWR.t1375 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1374 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1631 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t1529 VGND.t1528 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1632 XA.XIR[15].XIC[8].icell.Ien VPWR.t155 VPWR.t157 VPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1633 VPWR.t727 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t726 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 VGND.t1790 XThR.XTBN.Y a_n997_1803# VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1635 VPWR.t592 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t591 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1636 XThR.Tn[3].t4 XThR.XTBN.Y VGND.t1788 VGND.t1742 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1637 VGND.t2496 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t2495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1638 VPWR.t478 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 VPWR.t1176 XThC.XTB4.Y.t12 XThC.Tn[11].t4 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1640 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1641 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1642 VGND.t710 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t709 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1643 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t607 VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1644 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t1524 VPWR.t1523 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1645 VGND.t222 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t221 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1646 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t1531 VGND.t1530 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t726 VGND.t725 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1648 VPWR.t1424 VGND.t2696 Vbias.t5 VPWR.t1264 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X1649 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1518 VPWR.t1517 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1650 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t224 VGND.t2320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1651 VGND.t1021 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t1020 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1652 XThC.Tn[0].t4 XThC.XTBN.Y.t76 VGND.t2397 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1653 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t253 VGND.t2684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1654 VPWR.t1633 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t1632 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1655 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t63 VGND.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 XThC.Tn[3].t6 XThC.XTBN.Y.t77 VGND.t2398 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1657 VGND.t1269 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t1268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1658 VGND.t910 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t909 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1659 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t1228 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1661 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t948 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t797 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1663 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t949 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[8].XIC_15.icell.PUM VPWR.t153 XA.XIR[8].XIC_15.icell.Ien VPWR.t154 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t1885 VPWR.t1884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1666 VGND.t1736 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t1735 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1668 VPWR.t152 VPWR.t150 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1669 VGND.t712 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1670 VGND.t1605 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t1604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1671 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t2088 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1672 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t812 VPWR.t811 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1673 VPWR.t594 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1674 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t1233 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1675 VGND.t714 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1676 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t1485 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 XThC.XTB1.Y.t2 XThC.XTB5.A a_3299_10575# VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1678 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t1635 VPWR.t1634 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1679 VPWR.t1373 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1372 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1680 VGND.t1349 XThR.XTB3.Y.t10 XThR.Tn[2].t3 VGND.t1348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1681 XA.XIR[15].XIC[3].icell.Ien VPWR.t147 VPWR.t149 VPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1682 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t1533 VGND.t1532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1683 VGND.t716 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1684 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t1107 VPWR.t1106 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1685 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t794 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1686 VPWR.t729 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t728 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1687 VPWR.t596 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1688 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1689 VPWR.t894 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t893 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t2197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1691 VPWR.t516 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t515 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 VPWR.t480 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1693 VGND.t876 XThC.XTBN.Y.t78 XThC.Tn[6].t10 VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1694 VGND.t718 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1695 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t164 VGND.t1584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1696 XThC.Tn[10].t6 XThC.XTB3.Y.t11 VPWR.t1091 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1697 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t728 VGND.t727 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1698 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t358 VGND.t357 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1699 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t518 VPWR.t517 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1700 VGND.t1897 VGND.t1895 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1896 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1701 VGND.t720 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1702 VGND.t722 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 XThC.Tn[14].t2 XThC.XTB7.Y VPWR.t768 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1704 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t433 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1705 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1706 VGND.t1023 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 VGND.t1001 XThC.XTB1.Y.t13 XThC.Tn[0].t9 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1708 VGND.t578 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1710 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 VGND.t1271 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t1270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1713 XThR.Tn[8].t5 XThR.XTBN.Y VPWR.t1315 VPWR.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1714 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t84 VGND.t759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1715 VGND.t1273 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t1272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1716 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t193 VGND.t1741 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t259 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1718 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t2028 VGND.t2027 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1719 VGND.t2663 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t2662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 VGND.t2212 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t2211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t814 VPWR.t813 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1722 VGND.t2214 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t2213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 VGND.t1275 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t1274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1724 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t855 VPWR.t854 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1725 VGND.t2059 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t2058 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1726 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1727 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t5 VPWR.t1313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1728 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1637 VPWR.t1636 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1729 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t261 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1730 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1731 VGND.t1277 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t1276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1732 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t36 VGND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1733 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t356 VGND.t355 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1734 XThR.XTBN.A data[7].t1 VGND.t422 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1735 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t731 VPWR.t730 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1736 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1737 XThC.Tn[14].t1 XThC.XTB7.Y VPWR.t767 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1738 VPWR.t1467 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t1466 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1739 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t1534 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1740 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t1444 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1741 VPWR.t1423 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1742 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t1025 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1743 VGND.t224 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1744 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t1585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 XThC.XTB2.Y XThC.XTB7.B VPWR.t504 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1746 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1748 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1747 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t154 VGND.t1505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1748 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t896 VPWR.t895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1749 XThR.Tn[5].t8 XThR.XTBN.Y VGND.t1787 VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1750 VGND.t564 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1751 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t512 VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1752 VGND.t1279 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t1278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1753 VGND.t2498 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 XThR.Tn[10].t8 XThR.XTBN.Y VPWR.t1312 VPWR.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 VPWR.t857 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t856 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1756 Vbias.t3 bias[1].t0 VPWR.t1131 VPWR.t1130 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X1757 VGND.t2500 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t2499 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1758 a_5949_9615# XThC.XTB6.Y VPWR.t658 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1759 VGND.t1281 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t1280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1760 VGND.t1283 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t1282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t118 VGND.t1135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1762 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t514 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1763 VPWR.t1092 XThC.XTB3.Y.t12 XThC.Tn[10].t7 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1764 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t2030 VGND.t2029 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1765 VGND.t1894 VGND.t1892 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1766 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t99 VGND.t899 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1767 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t151 VGND.t1462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XThC.Tn[13].t8 XThC.XTBN.Y.t79 VPWR.t932 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1769 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t1027 VGND.t1026 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1770 a_n997_3755# XThR.XTBN.Y VGND.t1786 VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1771 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t181 VGND.t1680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1772 VPWR.t1310 XThR.XTBN.Y XThR.Tn[14].t10 VPWR.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1773 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t87 VGND.t769 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1774 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t1445 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1775 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t126 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t263 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t1029 VGND.t1028 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 VPWR.t1469 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t1468 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1781 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1782 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t898 VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1783 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t141 VGND.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1784 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t1042 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1785 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t65 VGND.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1786 XThR.Tn[7].t4 XThR.XTBN.Y VGND.t1785 VGND.t1784 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1787 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t134 VGND.t1358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1788 VPWR.t146 VPWR.t144 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1789 VGND.t1337 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t1336 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1790 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t747 VPWR.t746 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1791 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1792 VGND.t1031 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t1030 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 XThC.XTB4.Y.t1 XThC.XTB7.B VGND.t243 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1794 VPWR.t1250 XThR.XTB6.Y XThR.Tn[13].t2 VPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1795 VPWR.t1621 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1221 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1797 VPWR.t1173 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1798 VGND.t1285 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t1284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1799 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t1791 VPWR.t1790 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1800 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t703 VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 VPWR.t1270 data[4].t3 XThR.XTB7.A VPWR.t1269 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1802 VGND.t1643 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1803 VGND.t1287 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t1286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1804 VGND.t1033 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t1032 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1805 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t1035 VGND.t1034 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t516 VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XThC.Tn[6].t9 XThC.XTBN.Y.t80 VGND.t878 VGND.t877 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1808 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t2032 VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1809 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t1827 VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1810 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t1115 VPWR.t1114 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 VPWR.t1421 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t1420 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1812 VPWR.t1639 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t1638 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 XThR.Tn[5].t1 XThR.XTB6.Y VGND.t1671 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1814 VPWR.t859 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t858 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1815 VPWR.t780 XThC.XTB5.Y a_5155_9615# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1816 VPWR.t143 VPWR.t141 XA.XIR[3].XIC_15.icell.PUM VPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1817 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t2565 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1818 VPWR.t140 VPWR.t138 XA.XIR[7].XIC_15.icell.PUM VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1819 VGND.t1289 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t1288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1820 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t1849 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1821 XThR.Tn[4].t2 XThR.XTB5.Y VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1822 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1177 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1823 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t5 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1824 VGND.t1291 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t1290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1825 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t435 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1826 VGND.t1037 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t1036 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t72 VGND.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1828 VGND.t879 XThC.XTBN.Y.t82 XThC.Tn[2].t5 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1829 VGND.t1039 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t1038 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1830 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t136 VGND.t1364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1831 VPWR.t991 XThC.XTB1.Y.t14 XThC.Tn[8].t5 VPWR.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1832 VGND.t2608 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t2607 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1833 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1834 a_10915_9569# XThC.XTBN.Y.t83 VGND.t881 VGND.t880 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1835 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t749 VPWR.t748 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1836 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1278 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1837 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t1229 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 VPWR.t1761 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1760 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1839 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t900 VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1840 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t799 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1841 VGND.t1293 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t1292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1842 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t705 VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1843 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t1537 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1844 VGND.t1295 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t1294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1845 VGND.t1645 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1846 VGND.t1738 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t1737 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t1607 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t1829 VPWR.t1828 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1849 VGND.t1631 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1850 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t2200 VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t2033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1852 XThR.Tn[3].t3 XThR.XTBN.Y VGND.t1783 VGND.t1782 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1853 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t1487 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1854 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t1793 VPWR.t1792 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1855 VGND.t1464 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t1463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1856 VGND.t1466 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t1465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t707 VPWR.t706 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1858 VGND.t1468 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t1467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1859 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t136 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1860 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t5 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1861 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t1831 VPWR.t1830 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1862 a_4387_10575# XThC.XTB7.B VGND.t241 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1863 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t520 VPWR.t519 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1864 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t143 VGND.t1372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1865 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t1117 VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1866 VPWR.t1419 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t1418 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1867 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t1641 VPWR.t1640 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1868 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1869 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t162 VGND.t1581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1870 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1871 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t416 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t2596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 a_10051_9569# XThC.XTBN.Y.t84 VGND.t882 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1876 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t2512 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1877 XThC.XTB1.Y.t0 XThC.XTB7.B VPWR.t503 VPWR.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1878 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t8 VPWR.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1879 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t160 VGND.t1512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1880 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t175 VGND.t1669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 VGND.t1470 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t1469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1882 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t133 VPWR.t135 VPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1883 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1884 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t4 VPWR.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1885 a_7651_9569# XThC.XTBN.Y.t85 VGND.t884 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1886 VGND.t1891 VGND.t1889 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1890 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1887 VGND.t1999 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1888 VPWR.t1094 XThC.XTB7.A a_6243_10571# VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1889 VPWR.t132 VPWR.t130 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1890 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t766 VGND.t765 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1891 VPWR.t1763 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1892 XThC.Tn[10].t1 XThC.XTB3.Y.t13 a_8739_9569# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1893 VGND.t1472 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t1471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1894 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t226 VGND.t2351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1895 VGND.t2665 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t2664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1896 VGND.t1781 XThR.XTBN.Y XThR.Tn[2].t9 VGND.t1780 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1897 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t1588 VGND.t1587 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1898 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t1590 VGND.t1589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t239 VGND.t2432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1900 XThR.XTB5.A data[5].t3 VGND.t2187 VGND.t2186 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1901 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t105 VGND.t1003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1902 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t128 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1903 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t2202 VGND.t2201 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t992 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1905 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XThR.Tn[12].t9 XThR.XTBN.Y VPWR.t1307 VPWR.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1907 VGND.t1042 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t1041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1908 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t2568 VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XThR.Tn[12].t5 XThR.XTB5.Y a_n997_1803# VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1911 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t127 VGND.t1335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1912 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1913 XThR.Tn[3].t2 XThR.XTB4.Y.t11 VGND.t1580 VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1914 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t188 VGND.t1712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1915 VGND.t1779 XThR.XTBN.Y a_n997_2667# VGND.t1778 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1916 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t1044 VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1917 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1918 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t108 VGND.t1006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1919 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t1159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1920 VGND.t1474 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t1473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1921 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t125 VPWR.t127 VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1922 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t1446 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1923 VGND.t131 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1924 VGND.t488 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1925 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t2597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1926 a_5155_9615# XThC.XTB5.Y VPWR.t779 VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1927 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1928 VPWR.t778 XThC.XTB5.Y XThC.Tn[12].t0 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1929 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t1163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1930 VPWR.t751 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t750 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1931 XA.XIR[7].XIC_15.icell.PUM VPWR.t123 XA.XIR[7].XIC_15.icell.Ien VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1932 VPWR.t679 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t678 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1933 VPWR.t122 VPWR.t120 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VGND.t1339 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t1338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1935 XThC.Tn[5].t4 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1936 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t62 VGND.t566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1937 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t994 VGND.t993 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1938 VGND.t541 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1939 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t9 VPWR.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1940 VPWR.t1584 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t1583 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1941 VPWR.t902 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1942 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t251 VGND.t2644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1943 XThC.Tn[2].t4 XThC.XTBN.Y.t87 VGND.t885 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1944 VPWR.t522 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t521 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1945 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t1045 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t1046 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1947 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t5 VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1948 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t768 VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1949 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t996 VGND.t995 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t1073 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1951 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t168 VGND.t1656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1952 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t1009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1953 VPWR.t1733 XThR.XTB7.B XThR.XTB2.Y VPWR.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1954 Vbias.t0 bias[2].t0 VPWR.t978 VPWR.t977 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1955 XThC.Tn[8].t8 XThC.XTB1.Y.t15 a_7651_9569# VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t1592 VGND.t1591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1957 VGND.t2610 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t2609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t24 VGND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t1048 VGND.t1047 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t2357 XThC.XTB5.A XThC.XTB5.Y VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t1888 VGND.t1886 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 VGND.t1494 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t800 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1966 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t2570 VGND.t2569 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t2164 VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 VPWR.t753 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t752 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1969 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t801 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[4].XIC_15.icell.PUM VPWR.t118 XA.XIR[4].XIC_15.icell.Ien VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t2151 VGND.t2150 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t77 VGND.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1973 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t1050 VGND.t1049 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[15].XIC[9].icell.Ien VPWR.t115 VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1975 VGND.t1633 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1632 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1976 XThR.Tn[9].t8 XThR.XTBN.Y VPWR.t1301 VPWR.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 VGND.t886 XThC.XTBN.Y.t89 a_9827_9569# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1978 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t1586 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t1585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 VGND.t580 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t579 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1981 VGND.t1052 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t1051 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t1119 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t1476 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t1475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1984 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t755 VPWR.t754 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1985 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t112 VPWR.t114 VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1986 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1987 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t110 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t111 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1988 XThC.Tn[0].t10 XThC.XTB1.Y.t16 VGND.t1002 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t1478 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t1477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 VGND.t1480 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t1479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1991 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1992 VGND.t1647 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1993 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t4 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t998 VGND.t997 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1995 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1371 VPWR.t1370 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VGND.t1482 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t1481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1997 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t1795 VPWR.t1794 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1998 VPWR.t1588 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t1587 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1999 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t1594 VGND.t1593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2000 VGND.t2061 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t2060 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2001 VPWR.t711 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t2148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2003 XThR.Tn[14].t9 XThR.XTBN.Y VPWR.t1304 VPWR.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1568 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1567 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 VPWR.t109 VPWR.t107 XA.XIR[0].XIC_15.icell.PUM VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2006 VPWR.t681 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t680 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2007 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2008 a_n997_3755# XThR.XTBN.Y VGND.t1777 VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 XThR.Tn[8].t9 XThR.XTB1.Y.t13 VPWR.t1887 VPWR.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2010 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t1595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t713 VPWR.t712 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2012 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t2166 VGND.t2165 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2013 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t165 VGND.t1639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 VGND.t1484 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t1483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2015 a_n1049_7787# XThR.XTB2.Y VPWR.t397 VPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t68 VGND.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t2001 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t2000 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2018 VPWR.t816 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2019 a_n1331_2891# data[5].t4 VGND.t149 VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND.t1486 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t1485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2021 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t818 VPWR.t817 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2022 VPWR.t106 VPWR.t104 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t226 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2024 VPWR.t757 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t756 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2025 XThR.XTB7.B data[6].t1 VGND.t1709 VGND.t1708 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 XThR.Tn[2].t5 XThR.XTBN.Y a_n1049_7493# VPWR.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2027 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t2599 VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t2601 VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2029 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1369 VPWR.t1368 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2030 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t158 VGND.t1509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2031 VGND.t2216 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 VGND.t2063 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t2062 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2033 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t1054 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VGND.t1488 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t1487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2036 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 VPWR.t934 XThC.XTBN.Y.t90 XThC.Tn[8].t2 VPWR.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2038 XThR.Tn[10].t5 XThR.XTB3.Y.t12 VPWR.t976 VPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2039 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t999 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t1234 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XThR.Tn[4].t5 XThR.XTBN.Y VGND.t1776 VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2043 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t102 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1367 VPWR.t1366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t146 VGND.t1396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t2365 XThR.XTB7.B XThR.XTB5.Y VGND.t2364 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t1407 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t1406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t133 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2049 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2050 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t759 VPWR.t758 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2051 VGND.t490 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 VPWR.t683 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t682 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t496 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2054 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t359 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2055 VPWR.t820 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t819 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 VPWR.t1833 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t1832 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t2571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t46 VGND.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2060 VPWR.t1765 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1764 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2061 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t5 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 XThC.Tn[4].t4 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2063 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t685 VPWR.t684 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2064 VGND.t1409 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t1408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2065 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t206 VGND.t2068 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2066 VGND.t1411 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t1410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t66 VGND.t574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2068 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t99 VPWR.t101 VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 VGND.t2502 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t2501 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 VGND.t1413 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t1412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2071 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t467 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2072 VPWR.t1026 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2073 VGND.t1774 XThR.XTBN.Y a_n997_1579# VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2074 VPWR.t1212 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t1211 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2075 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t1057 VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2076 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1074 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2077 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2078 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1749 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t2603 VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t177 VGND.t1675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t117 VGND.t1124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2082 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t5 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2083 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t4 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t97 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t161 VGND.t1513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2087 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t1836 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t2153 VGND.t2152 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[0].XIC[5].icell.PDM VGND.t1883 VGND.t1885 VGND.t1884 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 VPWR.t1835 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t1834 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2091 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t1166 VGND.t1165 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t102 VGND.t912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2093 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t2514 VGND.t2513 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2094 VGND.t582 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t761 VPWR.t760 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2096 XThR.XTBN.Y XThR.XTBN.A VPWR.t942 VPWR.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2097 VGND.t1415 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t1414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2098 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t485 VPWR.t484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 VPWR.t982 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t981 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2100 VGND.t135 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2101 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2102 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t1230 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2103 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2104 VGND.t492 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2105 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t94 VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VPWR.t1214 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t1213 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2107 XA.XIR[0].XIC_15.icell.PUM VPWR.t92 XA.XIR[0].XIC_15.icell.Ien VPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2109 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t1590 VPWR.t1589 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2110 VGND.t1417 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t1416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 VGND.t1740 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t1739 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2112 VGND.t1609 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t1608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t1300 XThR.XTBN.Y XThR.Tn[11].t7 VPWR.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1570 VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2115 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t387 VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t1470 data[1].t4 XThC.XTB7.A VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 VPWR.t1028 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2118 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1767 VPWR.t1766 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2119 a_8739_9569# XThC.XTBN.Y.t92 VGND.t2131 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 VGND.t902 XThR.XTBN.A XThR.XTBN.Y VGND.t901 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XThC.Tn[6].t2 XThC.XTB7.Y VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t470 VGND.t469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1075 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t4 XThR.XTB5.Y a_n997_1803# VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t1059 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t1058 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t1419 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t1418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2130 VGND.t2612 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t2611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 VGND.t228 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t1421 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t1420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 a_n997_3979# XThR.XTBN.Y VGND.t1773 VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 XThC.XTB7.Y XThC.XTB7.B VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 XA.XIR[0].XIC[0].icell.PDM VGND.t1880 VGND.t1882 VGND.t1881 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2136 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t89 VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2137 VGND.t1423 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t1422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2138 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t1592 VPWR.t1591 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2139 VGND.t1425 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t1424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2140 XThC.Tn[8].t1 XThC.XTBN.Y.t93 VPWR.t1539 VPWR.t1538 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2141 VGND.t2122 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2121 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2142 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t2516 VGND.t2515 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2143 VGND.t1635 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t1634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 VGND.t1427 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t1426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2145 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t1121 VPWR.t1120 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2147 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t1061 VGND.t1060 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2148 VGND.t2190 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t2189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2150 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t466 VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2151 a_n1049_6699# XThR.XTB4.Y.t12 VPWR.t1199 VPWR.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2152 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t11 VGND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2153 VPWR.t1681 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t1680 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2154 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t388 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2155 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t1235 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2156 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t1007 VPWR.t1006 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2157 VGND.t1429 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t1428 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2158 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t87 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2159 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t229 VGND.t2355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2160 VGND.t2667 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t2666 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t85 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1572 VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2163 VGND.t1431 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t1430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t2269 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t2268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VGND.t2065 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t2064 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t2572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2167 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t1125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 VGND.t1064 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t1063 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2171 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t1401 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t1167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t764 data[1].t5 XThC.XTB6.A VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 VPWR.t763 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2176 VPWR.t84 VPWR.t82 XA.XIR[14].XIC_15.icell.PUM VPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2177 a_n997_2891# XThR.XTBN.Y VGND.t1771 VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 VGND.t2271 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t2270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2179 VGND.t2273 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t2272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2180 VGND.t2003 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t2002 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2181 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t1837 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 VPWR.t709 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t708 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2183 VPWR.t81 VPWR.t79 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2184 VGND.t2275 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t2274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2185 VGND.t1879 VGND.t1877 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2186 VGND.t1115 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t78 VPWR.t76 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VPWR.t822 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t821 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2189 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2190 XThR.Tn[11].t0 XThR.XTB4.Y.t13 a_n997_2667# VGND.t1492 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2191 VGND.t2277 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t2276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2192 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t2574 VGND.t2573 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2193 VPWR.t776 XThC.XTB5.Y a_5155_9615# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2195 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t35 VGND.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t1705 VGND.t1704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t1703 VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 VGND.t2279 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t2278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2199 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t1231 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2201 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t468 VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t1169 VGND.t1168 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2203 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t390 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2204 VGND.t1718 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t1717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t2174 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t1769 XThR.XTBN.Y XThR.Tn[0].t8 VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2207 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t2576 VGND.t2575 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2208 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t732 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 a_n1049_6405# XThR.XTB5.Y VPWR.t878 VPWR.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2210 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t52 VGND.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2211 XThR.Tn[8].t10 XThR.XTB1.Y.t14 VPWR.t1889 VPWR.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t6 VGND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2213 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2214 VGND.t2281 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t2280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t520 VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t7 VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t1067 VGND.t1066 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t2283 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t2282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t1488 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t494 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 VGND.t137 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t1126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2223 VGND.t2285 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t2284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2224 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2225 VGND.t139 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 VGND.t496 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2227 VPWR.t536 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2228 VGND.t2132 XThC.XTBN.Y.t94 a_8739_9569# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t765 VPWR.t764 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2230 VGND.t2287 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t2286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2231 VPWR.t75 VPWR.t73 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 XThC.Tn[1].t10 XThC.XTB2.Y VGND.t2647 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 VGND.t526 XThC.XTB7.Y XThC.Tn[6].t1 VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2235 VPWR.t639 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t638 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 VPWR.t72 VPWR.t70 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2237 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2238 VGND.t2289 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t2288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2239 VGND.t2291 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t2290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2240 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t1683 VPWR.t1682 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[2].t4 XThR.XTBN.Y a_n1049_7493# VPWR.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t1070 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t1069 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2243 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t70 VGND.t597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2244 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t487 VPWR.t486 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t148 VGND.t1398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2246 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t472 VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XThR.Tn[13].t8 XThR.XTBN.Y VPWR.t1298 VPWR.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2248 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1076 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2249 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t2578 VGND.t2577 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2250 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t715 VPWR.t714 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t142 VGND.t1371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2252 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1077 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t1701 VGND.t1700 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XThR.Tn[10].t0 XThR.XTB3.Y.t13 VPWR.t490 VPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t1750 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2256 XThR.Tn[4].t4 XThR.XTBN.Y VGND.t1767 VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 VPWR.t923 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t922 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2258 VGND.t1876 VGND.t1874 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2259 VGND.t1670 XThR.XTB6.Y XThR.Tn[5].t0 VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 VGND.t2669 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t2668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2261 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 VGND.t2293 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t2292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t1 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t424 VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t74 VGND.t621 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2266 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t143 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t1072 VGND.t1071 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t4 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 VGND.t2192 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t2191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2270 VGND.t771 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t1685 VPWR.t1684 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t131 VGND.t1355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t2194 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t2193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t773 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t984 VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 VPWR.t830 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t829 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2277 VGND.t1074 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t1073 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t67 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2279 VGND.t775 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VPWR.t1574 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1573 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t2124 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t1447 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2283 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t482 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t1699 VGND.t1698 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2286 VGND.t1076 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t1075 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t195 VGND.t1980 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 VGND.t1341 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VPWR.t601 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2290 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t184 VGND.t1696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2291 VPWR.t641 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t640 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2292 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t2579 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2293 VPWR.t470 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2294 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t832 VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2295 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2296 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t489 VPWR.t488 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2297 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t240 VGND.t2437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2298 VGND.t777 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t776 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2299 VGND.t1117 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t1116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 VPWR.t925 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t924 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2301 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VPWR.t66 VPWR.t64 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2303 VGND.t1119 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t1118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VGND.t779 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2305 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t572 VPWR.t571 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2306 XThR.Tn[4].t1 XThR.XTB5.Y VGND.t748 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2307 VPWR.t1296 XThR.XTBN.Y XThR.Tn[14].t8 VPWR.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2308 VPWR.t1687 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t1686 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2309 XThC.Tn[13].t1 XThC.XTB6.Y VPWR.t657 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2310 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2311 VGND.t398 XThC.XTB6.Y XThC.Tn[5].t0 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2312 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t146 VGND.t145 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2313 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t43 VGND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2314 VPWR.t1294 XThR.XTBN.Y XThR.Tn[11].t6 VPWR.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 VGND.t781 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2316 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t1689 VPWR.t1688 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2317 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t838 VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2318 VGND.t1873 VGND.t1871 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2319 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2320 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t234 VGND.t2399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2321 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2322 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XThC.Tn[9].t8 XThC.XTB2.Y a_7875_9569# VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t1078 VGND.t1077 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2325 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 VGND.t1695 XThC.XTB6.A XThC.XTB6.Y VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 VGND.t2646 XThC.XTB2.Y XThC.Tn[1].t9 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t1489 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t103 VGND.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2330 VGND.t783 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2331 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t62 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2332 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2333 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t238 VGND.t2405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t785 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 VGND.t787 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t2218 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2337 VGND.t1649 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2339 VPWR.t1143 XThR.XTB7.Y a_n1049_5317# VPWR.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 VPWR.t643 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t642 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2341 VGND.t1080 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t1079 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 VPWR.t656 XThC.XTB6.Y XThC.Tn[13].t0 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2343 VPWR.t472 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2344 a_n997_3979# XThR.XTBN.Y VGND.t1765 VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t538 VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2346 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t861 VPWR.t860 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t645 VPWR.t644 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2348 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t205 VGND.t2055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2349 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t59 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 VGND.t789 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t791 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t218 VGND.t2185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t1568 XThR.XTB4.Y.t14 XThR.Tn[3].t0 VGND.t897 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t222 VGND.t2266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t987 VPWR.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t1 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 VPWR.t1365 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1364 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2358 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t840 VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t12 VGND.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t474 VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2361 VGND.t793 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VGND.t1870 VGND.t1868 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2363 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t574 VPWR.t573 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2364 VPWR.t1797 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t1796 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2365 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2366 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t196 VGND.t2006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t1081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2368 VPWR.t540 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t7 VPWR.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 XA.XIR[0].XIC[11].icell.PDM VGND.t1865 VGND.t1867 VGND.t1866 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2372 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t1083 VGND.t1082 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2373 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t197 VGND.t2034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2374 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t23 VGND.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XThC.Tn[3].t0 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t213 VGND.t2147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t57 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 VPWR.t1265 bias[0].t0 Vbias.t4 VPWR.t1264 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X2379 XThC.XTB5.A data[0].t3 VGND.t1658 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VGND.t2504 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t2503 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2381 VPWR.t1200 XThR.XTB4.Y.t15 XThR.Tn[11].t1 VPWR.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2382 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t1707 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2383 XA.XIR[0].XIC[2].icell.PDM VGND.t1862 VGND.t1864 VGND.t1863 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2384 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t232 VGND.t2360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2385 VGND.t2614 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t2613 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2386 VGND.t1763 XThR.XTBN.Y a_n997_715# VGND.t1762 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 a_n997_2891# XThR.XTBN.Y VGND.t1761 VGND.t1760 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2388 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t314 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2389 VGND.t1861 VGND.t1859 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2390 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t542 VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2391 VPWR.t1030 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t1029 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2392 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t647 VPWR.t646 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2393 VPWR.t1363 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1362 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2394 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t54 VPWR.t56 VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2395 VPWR.t1799 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t1798 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2396 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2397 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2398 XThR.Tn[11].t2 XThR.XTB4.Y.t16 a_n997_2667# VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2399 VPWR.t53 VPWR.t51 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2400 VGND.t1637 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t1636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2401 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2402 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t49 VGND.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2403 VPWR.t1862 XThC.XTB2.Y XThC.Tn[9].t4 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2404 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t1032 VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2405 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t11 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2406 VGND.t1085 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t1084 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2407 VGND.t1343 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1342 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2408 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t152 VGND.t1489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2409 VPWR.t1541 XThC.XTBN.Y.t100 XThC.Tn[8].t0 VPWR.t1540 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2410 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t252 VGND.t2649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2411 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t2243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2412 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t2244 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2413 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t1511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2414 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2415 VPWR.t693 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t692 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2416 XA.XIR[0].XIC[6].icell.PDM VGND.t1856 VGND.t1858 VGND.t1857 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2417 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2418 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t8 VPWR.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2419 XA.XIR[15].XIC[7].icell.Ien VPWR.t48 VPWR.t50 VPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2420 XThR.Tn[7].t0 XThR.XTBN.Y VPWR.t1291 VPWR.t1290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2421 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t1087 VGND.t1086 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2422 VPWR.t544 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2423 VGND.t1855 VGND.t1853 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1854 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2424 VPWR.t1600 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t1599 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2425 XThC.Tn[9].t0 XThC.XTBN.Y.t101 VPWR.t1542 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2426 XThR.Tn[1].t9 XThR.XTBN.Y VGND.t1759 VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2427 VPWR.t47 VPWR.t45 XA.XIR[13].XIC_15.icell.PUM VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2428 VGND.t795 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t794 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2429 VGND.t2005 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t2004 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t2510 VGND.t2509 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t316 VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t1089 VGND.t1088 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2434 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1665 VPWR.t1664 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t1034 VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2436 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t2323 VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2437 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t145 VGND.t1392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2438 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t428 VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2439 VPWR.t1543 XThC.XTBN.Y.t102 XThC.Tn[11].t2 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2440 VPWR.t1361 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2441 VPWR.t1249 XThR.XTB6.Y a_n1049_5611# VPWR.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2442 VGND.t1091 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2443 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t2 VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2444 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t1127 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2445 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t172 VGND.t1665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2446 VPWR.t1801 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t1800 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2447 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2448 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t43 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2449 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t51 VGND.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2450 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t1129 VGND.t1128 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t1131 VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t1232 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2453 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t2511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2454 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t2176 VGND.t2175 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2456 VGND.t953 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2457 XA.XIR[15].XIC[11].icell.Ien VPWR.t40 VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2458 VGND.t1651 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 VGND.t1093 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[11].XIC_15.icell.PUM VPWR.t38 XA.XIR[11].XIC_15.icell.Ien VPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2461 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t1132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2462 VGND.t955 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2463 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t927 VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2464 VGND.t1720 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t1719 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 VGND.t1095 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2466 XThC.Tn[2].t0 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2467 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2468 VPWR.t1602 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t1601 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 VPWR.t695 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t694 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2470 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t1650 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2471 VGND.t2363 XThR.XTB7.B XThR.XTB4.Y.t1 VGND.t2362 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2472 VPWR.t37 VPWR.t35 XA.XIR[10].XIC_15.icell.PUM VPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2473 VGND.t957 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2474 XA.XIR[15].XIC[2].icell.Ien VPWR.t32 VPWR.t34 VPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2475 VGND.t959 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2476 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t1691 VPWR.t1690 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2477 VGND.t415 XThR.XTB1.Y.t16 XThR.Tn[0].t2 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2478 VPWR.t420 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2479 VPWR.t546 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2480 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t863 VPWR.t862 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2481 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t190 VGND.t1729 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2482 VPWR.t1604 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2483 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2484 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t595 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2485 VGND.t2616 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t2615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2486 VGND.t961 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2487 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t29 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2488 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t120 VGND.t1152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2489 a_8739_9569# XThC.XTBN.Y.t104 VGND.t1681 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2490 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t2178 VGND.t2177 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2491 XThC.Tn[6].t0 XThC.XTB7.Y VGND.t524 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2492 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t1036 VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2493 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t2325 VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t298 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2495 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2496 VGND.t963 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2497 VGND.t1683 XThC.XTBN.Y.t105 XThC.Tn[7].t4 VGND.t1682 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2498 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t1255 VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2499 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t929 VPWR.t928 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2500 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t2246 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2501 VGND.t2261 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t2260 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2502 XThC.Tn[12].t4 XThC.XTB5.Y a_9827_9569# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2503 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t110 VGND.t1008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2504 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t66 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1751 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2507 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t5 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2508 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t225 VGND.t2321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2509 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t1490 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2510 VGND.t965 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2511 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t27 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2512 VGND.t967 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2513 VGND.t498 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 VGND.t568 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2515 XThR.Tn[13].t1 XThR.XTB6.Y VPWR.t1248 VPWR.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2516 VGND.t969 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2517 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t931 VPWR.t930 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2518 VGND.t2671 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t2670 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2519 VGND.t971 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2520 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t576 VPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2521 VGND.t2220 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2522 VPWR.t422 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2523 VGND.t2067 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t2066 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t1004 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2525 VGND.t1684 XThC.XTBN.Y.t107 a_7875_9569# VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2526 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1097 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2528 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t733 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2529 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1359 VPWR.t1358 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2530 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2531 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t126 VGND.t1307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2532 VGND.t973 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2533 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t1803 VPWR.t1802 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t548 VPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2535 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t104 VGND.t987 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2536 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t649 VPWR.t648 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2537 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t300 VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2538 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2539 VPWR.t1417 VGND.t2700 XA.XIR[0].XIC[12].icell.PUM VPWR.t1416 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2540 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2541 a_8963_9569# XThC.XTBN.Y.t108 VGND.t1685 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2542 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t2326 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2543 VGND.t352 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t351 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2545 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t68 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2546 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2547 VPWR.t26 VPWR.t24 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2548 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t1752 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2552 VPWR.t578 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2553 VGND.t2506 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t2505 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2554 XThC.Tn[11].t1 XThC.XTBN.Y.t109 VPWR.t1256 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2555 VPWR.t1576 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2556 VGND.t975 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2557 XThR.Tn[6].t5 XThR.XTBN.Y a_n1049_5317# VPWR.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2558 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1272 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2559 VPWR.t1178 XThC.XTB4.Y.t16 XThC.Tn[11].t6 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2560 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t1732 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2561 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2562 VGND.t977 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2563 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t431 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t735 VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t1100 VGND.t1099 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 VGND.t2196 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t2195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2568 VGND.t850 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2569 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t739 VPWR.t738 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1357 VPWR.t1356 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2571 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t1102 VGND.t1101 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2572 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t113 VGND.t1107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2573 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t242 VGND.t2604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2574 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t139 VGND.t1368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2575 VPWR.t1415 VGND.t2701 XA.XIR[0].XIC[10].icell.PUM VPWR.t1414 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2576 VPWR.t874 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2577 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2578 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t842 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2579 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2580 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2581 VGND.t1757 XThR.XTBN.Y a_n997_1803# VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2582 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2583 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t834 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2584 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1624 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2586 XA.XIR[10].XIC_15.icell.PUM VPWR.t22 XA.XIR[10].XIC_15.icell.Ien VPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2587 a_3773_9615# XThC.XTB2.Y VPWR.t1861 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2588 VPWR.t21 VPWR.t19 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2589 VGND.t852 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2590 VGND.t1345 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1344 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 VGND.t1722 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t1721 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2592 VPWR.t865 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t864 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2593 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t1237 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2594 VPWR.t1201 XThR.XTB4.Y.t17 XThR.Tn[11].t3 VPWR.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2595 a_n997_715# XThR.XTBN.Y VGND.t1755 VGND.t1754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2596 VGND.t854 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2597 VPWR.t677 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2598 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1273 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2599 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t687 VPWR.t686 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2600 XThR.Tn[14].t1 XThR.XTB7.Y VPWR.t1141 VPWR.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2601 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t890 VGND.t889 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2602 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t651 VPWR.t650 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2603 VGND.t856 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2604 VGND.t1686 XThC.XTBN.Y.t110 XThC.Tn[3].t5 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2605 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t1606 VPWR.t1605 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2606 VGND.t1121 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t1120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2607 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t1104 VGND.t1103 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2608 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2609 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t1583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2610 VPWR.t867 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t866 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2611 XThC.Tn[1].t8 XThC.XTB2.Y VGND.t2645 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2612 VPWR.t1355 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1354 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2613 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2614 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1755 VPWR.t1754 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2615 VPWR.t1745 XThC.XTBN.A XThC.XTBN.Y.t0 VPWR.t1744 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2616 VPWR.t1578 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2617 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2618 VPWR.t741 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t740 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2619 VGND.t858 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2620 VPWR.t18 VPWR.t16 XA.XIR[6].XIC_15.icell.PUM VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2621 VGND.t860 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2622 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2623 XThR.Tn[2].t0 XThR.XTB3.Y.t16 VGND.t504 VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2624 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2625 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t1840 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2626 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t180 VGND.t1679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2627 VGND.t862 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2628 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t743 VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2629 VGND.t1852 VGND.t1850 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 VGND.t864 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t863 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2631 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t738 VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2632 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t2 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2633 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t221 VGND.t2265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2634 a_3299_10575# XThC.XTB7.B VGND.t238 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2635 VGND.t2091 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t2090 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2636 VGND.t1753 XThR.XTBN.Y XThR.Tn[6].t8 VGND.t1752 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 VPWR.t1413 VGND.t2702 XA.XIR[0].XIC[5].icell.PUM VPWR.t1412 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2638 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t1533 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2639 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2640 VPWR.t1757 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1756 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2641 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2642 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t13 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2643 VGND.t866 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VGND.t868 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2645 VGND.t586 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 VGND.t1653 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2647 VGND.t870 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2648 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t1009 VPWR.t1008 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2649 VGND.t2126 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2650 VGND.t872 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2651 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2652 VGND.t1724 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t1723 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2653 VPWR.t1257 XThC.XTBN.Y.t111 XThC.Tn[10].t8 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2654 VGND.t1571 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2655 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t2092 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2656 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2657 VGND.t1687 XThC.XTBN.Y.t112 a_8963_9569# VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2658 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t689 VPWR.t688 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2659 VGND.t874 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2660 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t506 VGND.t505 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2661 VPWR.t1721 XThC.XTB5.A a_5155_10571# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2662 VPWR.t766 XThC.XTB7.Y XThC.Tn[14].t0 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2663 XThR.Tn[1].t8 XThR.XTBN.Y VGND.t1751 VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2664 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t424 VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t653 VPWR.t652 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2666 VGND.t812 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t811 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2667 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t1011 VPWR.t1010 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2668 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t1038 VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2669 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t119 VGND.t1144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2670 VPWR.t1093 XThC.XTB7.A XThC.XTB3.Y.t1 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2671 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1759 VPWR.t1758 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2672 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2673 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t185 VGND.t1697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2674 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t20 VGND.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2675 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2676 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2677 XThR.Tn[8].t4 XThR.XTBN.Y VPWR.t1289 VPWR.t1288 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2678 VPWR.t426 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2679 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2680 XThR.Tn[5].t4 XThR.XTBN.Y a_n1049_5611# VPWR.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2681 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t4 VGND.t978 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2682 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2683 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t1732 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2684 VPWR.t12 VPWR.t10 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t11 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2685 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t13 VGND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2686 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t144 VGND.t1385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2687 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t4 VPWR.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2688 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t1 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2689 VPWR.t1731 XThR.XTB7.B XThR.XTB3.Y.t2 VPWR.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2690 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t2094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2691 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1753 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2692 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t875 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2693 VGND.t814 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2694 VPWR.t876 XThC.XTB3.Y.t16 XThC.Tn[10].t2 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2695 VPWR.t1258 XThC.XTBN.Y.t114 XThC.Tn[14].t9 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2696 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t1608 VPWR.t1607 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2697 VGND.t1849 VGND.t1847 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1848 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2698 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t1238 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2699 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t2096 VGND.t2095 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2700 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t156 VGND.t1507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2701 VGND.t588 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2702 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t56 VGND.t521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2703 VGND.t1749 XThR.XTBN.Y XThR.Tn[0].t7 VGND.t1748 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2704 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t88 VGND.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2705 VGND.t744 XThC.XTB3.Y.t17 XThC.Tn[2].t8 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2706 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t1565 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2707 XThR.Tn[10].t7 XThR.XTBN.Y VPWR.t1285 VPWR.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2708 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t508 VGND.t507 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t2098 VGND.t2097 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2710 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2711 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t114 VGND.t1113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2712 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t1712 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2713 VGND.t816 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2714 VPWR.t655 XThC.XTB6.Y a_5949_9615# VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2715 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t35 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2716 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t37 VGND.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2717 VGND.t1747 XThR.XTBN.Y a_n997_3755# VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2718 VPWR.t1024 data[3].t1 XThC.XTBN.A VPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2719 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t243 VGND.t2605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2720 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t993 VPWR.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2721 XThC.Tn[3].t4 XThC.XTBN.Y.t115 VGND.t1688 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2722 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1353 VPWR.t1352 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2723 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t17 VGND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2724 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t1134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2725 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2726 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t795 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2727 VPWR.t936 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t935 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2728 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t15 VGND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2729 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1580 VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2730 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2731 VPWR.t1610 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t1609 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2732 VPWR.t1725 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t1724 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2733 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2156 VGND.t2155 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2734 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2735 XThR.Tn[13].t0 XThR.XTB6.Y VPWR.t1247 VPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2736 VPWR.t1667 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2737 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t207 VGND.t2069 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2738 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t994 VPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2739 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2741 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t1842 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t740 VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2743 VGND.t1846 VGND.t1844 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2744 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t2346 VGND.t2345 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2745 VGND.t818 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2746 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t2158 VGND.t2157 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2747 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t8 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2748 VPWR.t873 XThC.XTB1.Y.t18 XThC.Tn[8].t4 VPWR.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2749 VGND.t2404 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2750 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t246 VGND.t2631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2751 VGND.t746 XThR.XTB5.Y XThR.Tn[4].t0 VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2752 XThC.Tn[10].t9 XThC.XTBN.Y.t116 VPWR.t1259 VPWR.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2753 VGND.t2556 XThC.XTBN.Y.t117 XThC.Tn[6].t8 VGND.t2555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2754 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2755 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2756 VPWR.t697 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t696 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2757 VPWR.t938 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t937 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2758 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t1678 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2759 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t1625 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[3].XIC_15.icell.PUM VPWR.t8 XA.XIR[3].XIC_15.icell.Ien VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t2248 VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2763 VGND.t820 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2764 VGND.t2128 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t2127 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t2100 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t2099 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t1726 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t1725 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 VGND.t2263 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t2262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VGND.t1728 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t1727 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2769 VPWR.t1727 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t1726 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2770 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t869 VPWR.t868 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2771 VPWR.t1679 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2772 VPWR.t1535 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2773 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t699 VPWR.t698 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2774 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t2101 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2775 VGND.t2103 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t2102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1202 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2777 VGND.t822 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2778 XThR.Tn[6].t4 XThR.XTBN.Y a_n1049_5317# VPWR.t1283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2779 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t6 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t7 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2780 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t4 VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2781 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1351 VPWR.t1350 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2782 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1582 VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2783 VGND.t824 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2784 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t745 VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2785 VGND.t2558 XThC.XTBN.Y.t118 a_10915_9569# VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2786 VPWR.t1612 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t1611 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2787 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t691 VPWR.t690 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2788 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t2160 VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2789 VGND.t2222 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t2221 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2790 VGND.t826 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2791 VPWR.t1729 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t1728 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2792 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t1789 VPWR.t1788 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2793 VPWR.t1537 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1536 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 VPWR.t1411 VGND.t2703 XA.XIR[0].XIC[14].icell.PUM VPWR.t1410 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2795 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t2104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2797 XThC.Tn[1].t0 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2798 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t122 VGND.t1155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2799 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t892 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2800 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t2349 VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2801 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t2130 VGND.t2129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2802 VGND.t828 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2803 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t248 VGND.t2641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2804 XThC.Tn[14].t8 XThC.XTBN.Y.t120 VPWR.t1786 VPWR.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2805 VGND.t830 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2806 VGND.t832 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2807 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t2105 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2808 VGND.t354 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2809 VGND.t1745 XThR.XTBN.Y a_n997_715# VGND.t1744 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2810 VPWR.t5 VPWR.t3 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2811 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t701 VPWR.t700 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2812 VPWR.t940 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t939 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2813 VPWR.t1139 XThR.XTB7.Y XThR.Tn[14].t0 VPWR.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2814 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2815 VGND.t1843 VGND.t1841 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2816 VGND.t834 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2817 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t64 VGND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2818 XThR.XTB6.A data[5].t5 VGND.t656 VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2819 XThR.Tn[0].t3 XThR.XTBN.Y a_n1049_8581# VPWR.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2820 VGND.t590 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t845 VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2822 a_5949_9615# XThC.XTB6.Y VPWR.t654 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2823 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t847 VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2824 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t90 VGND.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2825 VGND.t592 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 VGND.t2508 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t2507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2827 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t871 VPWR.t870 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2828 VGND.t2559 XThC.XTBN.Y.t121 a_10051_9569# VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2829 VGND.t836 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2830 VGND.t2554 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t2553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 VGND.t1573 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2832 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t2106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2833 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t2107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2834 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2835 XA.XIR[0].XIC[9].icell.PDM VGND.t1838 VGND.t1840 VGND.t1839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2836 VPWR.t1787 XThC.XTBN.Y.t122 XThC.Tn[11].t0 VPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2837 VGND.t2560 XThC.XTBN.Y.t123 a_7651_9569# VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2838 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1349 VPWR.t1348 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2839 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t79 VGND.t741 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2840 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t1614 VPWR.t1613 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2841 XThR.Tn[2].t8 XThR.XTBN.Y VGND.t1743 VGND.t1742 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2842 VPWR.t1137 XThR.XTB7.Y a_n1049_5317# VPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2843 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t2683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2844 VGND.t2492 Vbias.t260 XA.XIR[15].XIC_15.icell.SM VGND.t2491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2845 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t3 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2847 VGND.t570 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t569 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2848 VGND.t2339 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t2338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2849 VPWR.t1281 XThR.XTBN.Y XThR.Tn[12].t8 VPWR.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2850 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t2347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2851 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2852 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t420 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2853 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t228 VGND.t2354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2854 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t2562 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2855 VPWR.t2 VPWR.t0 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2856 VGND.t1347 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2857 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t31 VGND.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2858 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t2564 VGND.t2563 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2859 VGND.t2494 Vbias.t261 XA.XIR[13].XIC[2].icell.SM VGND.t2493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2860 VPWR.t803 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t802 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n2839 VGND.n7 32072.7
R1 VGND.n3017 VGND.n3016 21075.4
R2 VGND.n2875 VGND.n2843 13477
R3 VGND.n2843 VGND.n2842 11635.6
R4 VGND.n3010 VGND.n3009 9309.26
R5 VGND.n2908 VGND.n2875 9223.7
R6 VGND.n2909 VGND.n2908 9223.7
R7 VGND.n2962 VGND.n34 9223.7
R8 VGND.n2995 VGND.n2962 9223.7
R9 VGND.n2996 VGND.n2995 7447.41
R10 VGND.n1508 VGND.n1507 7387.65
R11 VGND.n1507 VGND.n1506 7387.65
R12 VGND.n2833 VGND.n147 7387.65
R13 VGND.n3015 VGND.n3014 7387.65
R14 VGND.n3014 VGND.n3013 7387.65
R15 VGND.n3013 VGND.n3012 7387.65
R16 VGND.n3012 VGND.n3011 7387.65
R17 VGND.n3011 VGND.n3010 7387.65
R18 VGND.n2838 VGND.n2833 7048.53
R19 VGND.n1510 VGND.t1350 6324.96
R20 VGND.n3016 VGND.n3015 5925.05
R21 VGND.n2909 VGND.n34 5231.11
R22 VGND.n1290 VGND.t1028 5131.29
R23 VGND.n3009 VGND.n3008 5074.71
R24 VGND.n2842 VGND.n7 4937.78
R25 VGND.n3016 VGND.n7 4804.6
R26 VGND.n1110 VGND.n578 4542.17
R27 VGND.n2839 VGND.n2838 4343.1
R28 VGND.n3009 VGND 4240.58
R29 VGND.n2414 VGND.n273 4110.84
R30 VGND.n1294 VGND.n1292 3417.39
R31 VGND.n1294 VGND.n1293 3417.39
R32 VGND.n1512 VGND.n1511 3417.39
R33 VGND.n960 VGND.n580 3417.39
R34 VGND.n635 VGND.n177 3417.39
R35 VGND.n2832 VGND.n114 3417.39
R36 VGND.n2841 VGND.n2840 3417.39
R37 VGND.n2415 VGND.n2414 3331.79
R38 VGND.n2416 VGND.n2415 3331.79
R39 VGND.n2417 VGND.n2416 3331.79
R40 VGND.n2418 VGND.n2417 3331.79
R41 VGND.n2419 VGND.n2418 3331.79
R42 VGND.n2420 VGND.n2419 3331.79
R43 VGND.n2421 VGND.n2420 3331.79
R44 VGND.n2422 VGND.n2421 3331.79
R45 VGND.n2423 VGND.n2422 3331.79
R46 VGND.n2424 VGND.n2423 3331.79
R47 VGND.n2425 VGND.n2424 3331.79
R48 VGND.n2426 VGND.n2425 3331.79
R49 VGND.n2427 VGND.n2426 3331.79
R50 VGND.n2427 VGND.n32 3331.79
R51 VGND.n2998 VGND.n32 3331.79
R52 VGND.n2998 VGND.n2997 3331.79
R53 VGND.n1293 VGND.n578 3273.91
R54 VGND.n961 VGND.n579 3265.22
R55 VGND.n2839 VGND.n114 2756.52
R56 VGND.n2875 VGND.t1795 2655.17
R57 VGND.n2908 VGND.t1819 2655.17
R58 VGND.n2997 VGND.n2996 2602.7
R59 VGND.n2833 VGND.n2832 2517.39
R60 VGND.n2836 VGND.n5 2229.43
R61 VGND.n3018 VGND.n5 2229.43
R62 VGND.n3018 VGND.n6 2229.43
R63 VGND.n2836 VGND.n6 2229.43
R64 VGND.n1292 VGND.n1291 2130.43
R65 VGND.n2842 VGND.n2841 2082.61
R66 VGND VGND.n34 1997.7
R67 VGND.n2962 VGND 1997.7
R68 VGND.n2995 VGND 1997.7
R69 VGND.n1505 VGND.n147 1831.57
R70 VGND.t1752 VGND.n2909 1807.04
R71 VGND.n2993 VGND.t421 1785.51
R72 VGND.n1506 VGND.n580 1691.3
R73 VGND.n2921 VGND.t45 1618.39
R74 VGND.t1492 VGND.n2961 1618.39
R75 VGND.t750 VGND.n2994 1618.39
R76 VGND.n2843 VGND.t1768 1517.24
R77 VGND.n1509 VGND.n1508 1513.49
R78 VGND.n1510 VGND.n1509 1370.36
R79 VGND.n1291 VGND.n1290 1286.96
R80 VGND.n1509 VGND.t1839 1270.28
R81 VGND.n1083 VGND.t399 1268.93
R82 VGND.n1083 VGND.t94 1268.93
R83 VGND.n146 VGND.t242 1253.59
R84 VGND.t50 VGND.n146 1253.59
R85 VGND.n614 VGND.t48 1253.59
R86 VGND.t247 VGND.n614 1253.59
R87 VGND.n1021 VGND.t763 1253.59
R88 VGND.n1021 VGND.t883 1253.59
R89 VGND.n1052 VGND.t52 1253.59
R90 VGND.n1052 VGND.t92 1253.59
R91 VGND.n176 VGND.t245 1253.59
R92 VGND.t237 VGND.n176 1253.59
R93 VGND.n1505 VGND.t1884 1237.71
R94 VGND.n2838 VGND.n2837 1217.3
R95 VGND.n2921 VGND.t1714 1213.79
R96 VGND.n1111 VGND.n1110 1198.25
R97 VGND.n3008 VGND.n3007 1198.25
R98 VGND.n2651 VGND.n33 1180.79
R99 VGND.n3000 VGND.n2999 1180.79
R100 VGND.n2490 VGND.n2489 1180.79
R101 VGND.n2429 VGND.n2428 1180.79
R102 VGND.n2312 VGND.n261 1180.79
R103 VGND.n2126 VGND.n262 1180.79
R104 VGND.n2121 VGND.n263 1180.79
R105 VGND.n2337 VGND.n264 1180.79
R106 VGND.n1952 VGND.n265 1180.79
R107 VGND.n1947 VGND.n266 1180.79
R108 VGND.n2362 VGND.n267 1180.79
R109 VGND.n1778 VGND.n268 1180.79
R110 VGND.n1773 VGND.n269 1180.79
R111 VGND.n2387 VGND.n270 1180.79
R112 VGND.n1604 VGND.n271 1180.79
R113 VGND.n2407 VGND.n272 1180.79
R114 VGND.n1232 VGND.n273 1180.79
R115 VGND.n2413 VGND.n2412 1180.79
R116 VGND.n1289 VGND.n1288 1180.46
R117 VGND.n720 VGND.n679 1180.46
R118 VGND.n725 VGND.n724 1180.46
R119 VGND.n730 VGND.n729 1180.46
R120 VGND.n735 VGND.n734 1180.46
R121 VGND.n740 VGND.n739 1180.46
R122 VGND.n745 VGND.n744 1180.46
R123 VGND.n750 VGND.n749 1180.46
R124 VGND.n755 VGND.n754 1180.46
R125 VGND.n760 VGND.n759 1180.46
R126 VGND.n765 VGND.n764 1180.46
R127 VGND.n770 VGND.n769 1180.46
R128 VGND.n775 VGND.n774 1180.46
R129 VGND.n780 VGND.n779 1180.46
R130 VGND.n782 VGND.n781 1180.46
R131 VGND.n1229 VGND.n1228 1180.46
R132 VGND.n1227 VGND.n1226 1180.46
R133 VGND.n1210 VGND.n1209 1180.46
R134 VGND.n1208 VGND.n1207 1180.46
R135 VGND.n1197 VGND.n1196 1180.46
R136 VGND.n1195 VGND.n1194 1180.46
R137 VGND.n1178 VGND.n1177 1180.46
R138 VGND.n1176 VGND.n1175 1180.46
R139 VGND.n1165 VGND.n1164 1180.46
R140 VGND.n1163 VGND.n1162 1180.46
R141 VGND.n1146 VGND.n1145 1180.46
R142 VGND.n1144 VGND.n1143 1180.46
R143 VGND.n1133 VGND.n1132 1180.46
R144 VGND.n1131 VGND.n1130 1180.46
R145 VGND.n1123 VGND.n1122 1180.46
R146 VGND.n2578 VGND.n2577 1180.46
R147 VGND.n2706 VGND.n2705 1180.46
R148 VGND.n2704 VGND.n2703 1180.46
R149 VGND.n2698 VGND.n2697 1180.46
R150 VGND.n2696 VGND.n2695 1180.46
R151 VGND.n2690 VGND.n2689 1180.46
R152 VGND.n2688 VGND.n2687 1180.46
R153 VGND.n2682 VGND.n2681 1180.46
R154 VGND.n2680 VGND.n2679 1180.46
R155 VGND.n2674 VGND.n2673 1180.46
R156 VGND.n2672 VGND.n2671 1180.46
R157 VGND.n2666 VGND.n2665 1180.46
R158 VGND.n2664 VGND.n2663 1180.46
R159 VGND.n2658 VGND.n2657 1180.46
R160 VGND.n2656 VGND.n2655 1180.46
R161 VGND.n234 VGND.n233 1180.46
R162 VGND.n2719 VGND.n2718 1180.46
R163 VGND.n2724 VGND.n2723 1180.46
R164 VGND.n2729 VGND.n2728 1180.46
R165 VGND.n2734 VGND.n2733 1180.46
R166 VGND.n2739 VGND.n2738 1180.46
R167 VGND.n2744 VGND.n2743 1180.46
R168 VGND.n2749 VGND.n2748 1180.46
R169 VGND.n2754 VGND.n2753 1180.46
R170 VGND.n2759 VGND.n2758 1180.46
R171 VGND.n2764 VGND.n2763 1180.46
R172 VGND.n2769 VGND.n2768 1180.46
R173 VGND.n2774 VGND.n2773 1180.46
R174 VGND.n2779 VGND.n2778 1180.46
R175 VGND.n2781 VGND.n2780 1180.46
R176 VGND.n2515 VGND.n2514 1180.46
R177 VGND.n2513 VGND.n2512 1180.46
R178 VGND.n2508 VGND.n2507 1180.46
R179 VGND.n2433 VGND.n244 1180.46
R180 VGND.n2438 VGND.n2437 1180.46
R181 VGND.n2443 VGND.n2442 1180.46
R182 VGND.n2448 VGND.n2447 1180.46
R183 VGND.n2453 VGND.n2452 1180.46
R184 VGND.n2458 VGND.n2457 1180.46
R185 VGND.n2463 VGND.n2462 1180.46
R186 VGND.n2468 VGND.n2467 1180.46
R187 VGND.n2473 VGND.n2472 1180.46
R188 VGND.n2478 VGND.n2477 1180.46
R189 VGND.n2483 VGND.n2482 1180.46
R190 VGND.n2488 VGND.n2487 1180.46
R191 VGND.n2831 VGND.n2830 1180.46
R192 VGND.n371 VGND.n182 1180.46
R193 VGND.n373 VGND.n372 1180.46
R194 VGND.n2171 VGND.n2170 1180.46
R195 VGND.n2173 VGND.n2172 1180.46
R196 VGND.n2197 VGND.n2196 1180.46
R197 VGND.n2199 VGND.n2198 1180.46
R198 VGND.n2223 VGND.n2222 1180.46
R199 VGND.n2225 VGND.n2224 1180.46
R200 VGND.n2249 VGND.n2248 1180.46
R201 VGND.n2251 VGND.n2250 1180.46
R202 VGND.n2280 VGND.n2279 1180.46
R203 VGND.n2285 VGND.n2284 1180.46
R204 VGND.n2290 VGND.n2289 1180.46
R205 VGND.n2292 VGND.n2291 1180.46
R206 VGND.n1428 VGND.n1427 1180.46
R207 VGND.n1430 VGND.n1429 1180.46
R208 VGND.n2158 VGND.n2157 1180.46
R209 VGND.n2160 VGND.n2159 1180.46
R210 VGND.n2184 VGND.n2183 1180.46
R211 VGND.n2186 VGND.n2185 1180.46
R212 VGND.n2210 VGND.n2209 1180.46
R213 VGND.n2212 VGND.n2211 1180.46
R214 VGND.n2236 VGND.n2235 1180.46
R215 VGND.n2238 VGND.n2237 1180.46
R216 VGND.n2262 VGND.n2261 1180.46
R217 VGND.n2269 VGND.n2268 1180.46
R218 VGND.n2267 VGND.n2266 1180.46
R219 VGND.n2307 VGND.n2306 1180.46
R220 VGND.n2309 VGND.n2308 1180.46
R221 VGND.n1442 VGND.n1441 1180.46
R222 VGND.n1494 VGND.n1493 1180.46
R223 VGND.n1492 VGND.n1491 1180.46
R224 VGND.n1487 VGND.n1486 1180.46
R225 VGND.n1482 VGND.n1481 1180.46
R226 VGND.n1477 VGND.n1476 1180.46
R227 VGND.n1472 VGND.n1471 1180.46
R228 VGND.n1467 VGND.n1466 1180.46
R229 VGND.n1462 VGND.n1461 1180.46
R230 VGND.n1457 VGND.n1456 1180.46
R231 VGND.n1452 VGND.n1451 1180.46
R232 VGND.n1447 VGND.n1446 1180.46
R233 VGND.n2137 VGND.n2136 1180.46
R234 VGND.n2135 VGND.n2134 1180.46
R235 VGND.n2130 VGND.n2129 1180.46
R236 VGND.n1504 VGND.n1503 1180.46
R237 VGND.n626 VGND.n619 1180.46
R238 VGND.n628 VGND.n627 1180.46
R239 VGND.n1997 VGND.n1996 1180.46
R240 VGND.n1999 VGND.n1998 1180.46
R241 VGND.n2023 VGND.n2022 1180.46
R242 VGND.n2025 VGND.n2024 1180.46
R243 VGND.n2049 VGND.n2048 1180.46
R244 VGND.n2051 VGND.n2050 1180.46
R245 VGND.n2075 VGND.n2074 1180.46
R246 VGND.n2077 VGND.n2076 1180.46
R247 VGND.n2106 VGND.n2105 1180.46
R248 VGND.n2111 VGND.n2110 1180.46
R249 VGND.n2116 VGND.n2115 1180.46
R250 VGND.n2118 VGND.n2117 1180.46
R251 VGND.n652 VGND.n651 1180.46
R252 VGND.n654 VGND.n653 1180.46
R253 VGND.n1984 VGND.n1983 1180.46
R254 VGND.n1986 VGND.n1985 1180.46
R255 VGND.n2010 VGND.n2009 1180.46
R256 VGND.n2012 VGND.n2011 1180.46
R257 VGND.n2036 VGND.n2035 1180.46
R258 VGND.n2038 VGND.n2037 1180.46
R259 VGND.n2062 VGND.n2061 1180.46
R260 VGND.n2064 VGND.n2063 1180.46
R261 VGND.n2088 VGND.n2087 1180.46
R262 VGND.n2095 VGND.n2094 1180.46
R263 VGND.n2093 VGND.n2092 1180.46
R264 VGND.n2332 VGND.n2331 1180.46
R265 VGND.n2334 VGND.n2333 1180.46
R266 VGND.n959 VGND.n958 1180.46
R267 VGND.n954 VGND.n953 1180.46
R268 VGND.n949 VGND.n948 1180.46
R269 VGND.n944 VGND.n943 1180.46
R270 VGND.n939 VGND.n938 1180.46
R271 VGND.n934 VGND.n933 1180.46
R272 VGND.n929 VGND.n928 1180.46
R273 VGND.n924 VGND.n923 1180.46
R274 VGND.n919 VGND.n918 1180.46
R275 VGND.n914 VGND.n913 1180.46
R276 VGND.n909 VGND.n908 1180.46
R277 VGND.n904 VGND.n903 1180.46
R278 VGND.n1963 VGND.n1962 1180.46
R279 VGND.n1961 VGND.n1960 1180.46
R280 VGND.n1956 VGND.n1955 1180.46
R281 VGND.n1395 VGND.n1394 1180.46
R282 VGND.n1400 VGND.n1399 1180.46
R283 VGND.n1402 VGND.n1401 1180.46
R284 VGND.n1823 VGND.n1822 1180.46
R285 VGND.n1825 VGND.n1824 1180.46
R286 VGND.n1849 VGND.n1848 1180.46
R287 VGND.n1851 VGND.n1850 1180.46
R288 VGND.n1875 VGND.n1874 1180.46
R289 VGND.n1877 VGND.n1876 1180.46
R290 VGND.n1901 VGND.n1900 1180.46
R291 VGND.n1903 VGND.n1902 1180.46
R292 VGND.n1932 VGND.n1931 1180.46
R293 VGND.n1937 VGND.n1936 1180.46
R294 VGND.n1942 VGND.n1941 1180.46
R295 VGND.n1944 VGND.n1943 1180.46
R296 VGND.n1380 VGND.n1379 1180.46
R297 VGND.n1382 VGND.n1381 1180.46
R298 VGND.n1810 VGND.n1809 1180.46
R299 VGND.n1812 VGND.n1811 1180.46
R300 VGND.n1836 VGND.n1835 1180.46
R301 VGND.n1838 VGND.n1837 1180.46
R302 VGND.n1862 VGND.n1861 1180.46
R303 VGND.n1864 VGND.n1863 1180.46
R304 VGND.n1888 VGND.n1887 1180.46
R305 VGND.n1890 VGND.n1889 1180.46
R306 VGND.n1914 VGND.n1913 1180.46
R307 VGND.n1921 VGND.n1920 1180.46
R308 VGND.n1919 VGND.n1918 1180.46
R309 VGND.n2357 VGND.n2356 1180.46
R310 VGND.n2359 VGND.n2358 1180.46
R311 VGND.n1312 VGND.n1311 1180.46
R312 VGND.n1364 VGND.n1363 1180.46
R313 VGND.n1362 VGND.n1361 1180.46
R314 VGND.n1357 VGND.n1356 1180.46
R315 VGND.n1352 VGND.n1351 1180.46
R316 VGND.n1347 VGND.n1346 1180.46
R317 VGND.n1342 VGND.n1341 1180.46
R318 VGND.n1337 VGND.n1336 1180.46
R319 VGND.n1332 VGND.n1331 1180.46
R320 VGND.n1327 VGND.n1326 1180.46
R321 VGND.n1322 VGND.n1321 1180.46
R322 VGND.n1317 VGND.n1316 1180.46
R323 VGND.n1789 VGND.n1788 1180.46
R324 VGND.n1787 VGND.n1786 1180.46
R325 VGND.n1782 VGND.n1781 1180.46
R326 VGND.n1517 VGND.n1516 1180.46
R327 VGND.n1522 VGND.n1521 1180.46
R328 VGND.n1524 VGND.n1523 1180.46
R329 VGND.n1649 VGND.n1648 1180.46
R330 VGND.n1651 VGND.n1650 1180.46
R331 VGND.n1675 VGND.n1674 1180.46
R332 VGND.n1677 VGND.n1676 1180.46
R333 VGND.n1701 VGND.n1700 1180.46
R334 VGND.n1703 VGND.n1702 1180.46
R335 VGND.n1727 VGND.n1726 1180.46
R336 VGND.n1729 VGND.n1728 1180.46
R337 VGND.n1758 VGND.n1757 1180.46
R338 VGND.n1763 VGND.n1762 1180.46
R339 VGND.n1768 VGND.n1767 1180.46
R340 VGND.n1770 VGND.n1769 1180.46
R341 VGND.n1537 VGND.n1536 1180.46
R342 VGND.n1539 VGND.n1538 1180.46
R343 VGND.n1636 VGND.n1635 1180.46
R344 VGND.n1638 VGND.n1637 1180.46
R345 VGND.n1662 VGND.n1661 1180.46
R346 VGND.n1664 VGND.n1663 1180.46
R347 VGND.n1688 VGND.n1687 1180.46
R348 VGND.n1690 VGND.n1689 1180.46
R349 VGND.n1714 VGND.n1713 1180.46
R350 VGND.n1716 VGND.n1715 1180.46
R351 VGND.n1740 VGND.n1739 1180.46
R352 VGND.n1747 VGND.n1746 1180.46
R353 VGND.n1745 VGND.n1744 1180.46
R354 VGND.n2382 VGND.n2381 1180.46
R355 VGND.n2384 VGND.n2383 1180.46
R356 VGND.n1296 VGND.n1295 1180.46
R357 VGND.n1550 VGND.n1549 1180.46
R358 VGND.n1555 VGND.n1554 1180.46
R359 VGND.n1560 VGND.n1559 1180.46
R360 VGND.n1565 VGND.n1564 1180.46
R361 VGND.n1570 VGND.n1569 1180.46
R362 VGND.n1575 VGND.n1574 1180.46
R363 VGND.n1580 VGND.n1579 1180.46
R364 VGND.n1585 VGND.n1584 1180.46
R365 VGND.n1590 VGND.n1589 1180.46
R366 VGND.n1595 VGND.n1594 1180.46
R367 VGND.n1600 VGND.n1599 1180.46
R368 VGND.n1615 VGND.n1614 1180.46
R369 VGND.n1613 VGND.n1612 1180.46
R370 VGND.n1608 VGND.n1607 1180.46
R371 VGND.n835 VGND.n834 1180.46
R372 VGND.n840 VGND.n839 1180.46
R373 VGND.n892 VGND.n891 1180.46
R374 VGND.n890 VGND.n889 1180.46
R375 VGND.n885 VGND.n884 1180.46
R376 VGND.n880 VGND.n879 1180.46
R377 VGND.n875 VGND.n874 1180.46
R378 VGND.n870 VGND.n869 1180.46
R379 VGND.n865 VGND.n864 1180.46
R380 VGND.n860 VGND.n859 1180.46
R381 VGND.n855 VGND.n854 1180.46
R382 VGND.n850 VGND.n849 1180.46
R383 VGND.n845 VGND.n844 1180.46
R384 VGND.n2402 VGND.n2401 1180.46
R385 VGND.n2404 VGND.n2403 1180.46
R386 VGND.n2961 VGND.t1713 1180.08
R387 VGND.n1511 VGND.n1510 1169.57
R388 VGND.n3013 VGND.t32 1146.36
R389 VGND.n3015 VGND.t31 1112.64
R390 VGND.n3014 VGND.t534 1112.64
R391 VGND.n2996 VGND 1055.35
R392 VGND.n1506 VGND.n1505 1052.29
R393 VGND.t46 VGND.n961 1032.59
R394 VGND.t201 VGND.n2578 988.926
R395 VGND.n2705 VGND.t1056 988.926
R396 VGND.n2704 VGND.t1034 988.926
R397 VGND.n2697 VGND.t199 988.926
R398 VGND.n2696 VGND.t188 988.926
R399 VGND.n2689 VGND.t1103 988.926
R400 VGND.n2688 VGND.t1220 988.926
R401 VGND.n2681 VGND.t1197 988.926
R402 VGND.n2680 VGND.t1099 988.926
R403 VGND.n2673 VGND.t1018 988.926
R404 VGND.n2672 VGND.t1262 988.926
R405 VGND.n2665 VGND.t217 988.926
R406 VGND.n2664 VGND.t1086 988.926
R407 VGND.n2657 VGND.t1250 988.926
R408 VGND.n2656 VGND.t1182 988.926
R409 VGND.n233 VGND.t983 988.926
R410 VGND.t637 VGND.n2719 988.926
R411 VGND.t2348 VGND.n2724 988.926
R412 VGND.t1544 VGND.n2729 988.926
R413 VGND.t1612 VGND.n2734 988.926
R414 VGND.t311 VGND.n2739 988.926
R415 VGND.t2569 VGND.n2744 988.926
R416 VGND.t727 VGND.n2749 988.926
R417 VGND.t2050 VGND.n2754 988.926
R418 VGND.t394 VGND.n2759 988.926
R419 VGND.t2324 VGND.n2764 988.926
R420 VGND.t2022 VGND.n2769 988.926
R421 VGND.t100 VGND.n2774 988.926
R422 VGND.t145 VGND.n2779 988.926
R423 VGND.n2780 VGND.t382 988.926
R424 VGND.n2514 VGND.t471 988.926
R425 VGND.n2513 VGND.t645 988.926
R426 VGND.n2508 VGND.t1987 988.926
R427 VGND.t1168 VGND.n2433 988.926
R428 VGND.t2152 VGND.n2438 988.926
R429 VGND.t434 VGND.n2443 988.926
R430 VGND.t2673 VGND.n2448 988.926
R431 VGND.t739 VGND.n2453 988.926
R432 VGND.t125 VGND.n2458 988.926
R433 VGND.t408 VGND.n2463 988.926
R434 VGND.t2039 VGND.n2468 988.926
R435 VGND.t2509 VGND.n2473 988.926
R436 VGND.t606 VGND.n2478 988.926
R437 VGND.t2072 VGND.n2483 988.926
R438 VGND.t430 VGND.n2488 988.926
R439 VGND.n2831 VGND.t280 988.926
R440 VGND.t2169 VGND.n371 988.926
R441 VGND.n372 VGND.t58 988.926
R442 VGND.t1551 VGND.n2171 988.926
R443 VGND.n2172 VGND.t1618 988.926
R444 VGND.t922 VGND.n2197 988.926
R445 VGND.n2198 VGND.t2575 988.926
R446 VGND.t995 VGND.n2223 988.926
R447 VGND.n2224 VGND.t650 988.926
R448 VGND.t362 VGND.n2249 988.926
R449 VGND.n2250 VGND.t2157 988.926
R450 VGND.t1530 VGND.n2280 988.926
R451 VGND.t106 VGND.n2285 988.926
R452 VGND.t734 VGND.n2290 988.926
R453 VGND.n2291 VGND.t513 988.926
R454 VGND.t2381 VGND.n1428 988.926
R455 VGND.n1429 VGND.t65 988.926
R456 VGND.t1700 VGND.n2158 988.926
R457 VGND.n2159 VGND.t1303 988.926
R458 VGND.t2341 VGND.n2184 988.926
R459 VGND.n2185 VGND.t290 988.926
R460 VGND.t482 VGND.n2210 988.926
R461 VGND.n2211 VGND.t801 988.926
R462 VGND.t1140 VGND.n2236 988.926
R463 VGND.n2237 VGND.t2602 988.926
R464 VGND.t1591 VGND.n2262 988.926
R465 VGND.n2268 VGND.t1563 988.926
R466 VGND.n2267 VGND.t2328 988.926
R467 VGND.t2029 VGND.n2307 988.926
R468 VGND.n2308 VGND.t374 988.926
R469 VGND.t767 VGND.n1442 988.926
R470 VGND.n1493 VGND.t1361 988.926
R471 VGND.n1492 VGND.t1981 988.926
R472 VGND.n1487 VGND.t2201 988.926
R473 VGND.n1482 VGND.t262 988.926
R474 VGND.n1477 VGND.t334 988.926
R475 VGND.n1472 VGND.t507 988.926
R476 VGND.n1467 VGND.t315 988.926
R477 VGND.n1462 VGND.t916 988.926
R478 VGND.n1457 VGND.t370 988.926
R479 VGND.n1452 VGND.t307 988.926
R480 VGND.n1447 VGND.t2515 988.926
R481 VGND.n2136 VGND.t113 988.926
R482 VGND.n2135 VGND.t2533 988.926
R483 VGND.n2130 VGND.t423 988.926
R484 VGND.n1504 VGND.t981 988.926
R485 VGND.t635 VGND.n626 988.926
R486 VGND.n627 VGND.t2345 988.926
R487 VGND.t1542 VGND.n1997 988.926
R488 VGND.n1998 VGND.t1610 988.926
R489 VGND.t309 VGND.n2023 988.926
R490 VGND.n2024 VGND.t2567 988.926
R491 VGND.t725 VGND.n2049 988.926
R492 VGND.n2050 VGND.t2048 988.926
R493 VGND.t391 VGND.n2075 988.926
R494 VGND.n2076 VGND.t2322 988.926
R495 VGND.t2019 VGND.n2106 988.926
R496 VGND.t2334 VGND.n2111 988.926
R497 VGND.t142 VGND.n2116 988.926
R498 VGND.n2117 VGND.t380 988.926
R499 VGND.t282 VGND.n652 988.926
R500 VGND.n653 VGND.t2171 988.926
R501 VGND.t56 VGND.n1984 988.926
R502 VGND.n1985 VGND.t1553 988.926
R503 VGND.t2083 VGND.n2010 988.926
R504 VGND.n2011 VGND.t924 988.926
R505 VGND.t2577 VGND.n2036 988.926
R506 VGND.n2037 VGND.t997 988.926
R507 VGND.t652 VGND.n2062 988.926
R508 VGND.n2063 VGND.t364 988.926
R509 VGND.t2159 VGND.n2088 988.926
R510 VGND.n2094 VGND.t1532 988.926
R511 VGND.n2093 VGND.t108 988.926
R512 VGND.t889 VGND.n2332 988.926
R513 VGND.n2333 VGND.t515 988.926
R514 VGND.n959 VGND.t2383 988.926
R515 VGND.n954 VGND.t67 988.926
R516 VGND.n949 VGND.t1698 988.926
R517 VGND.n944 VGND.t1305 988.926
R518 VGND.n939 VGND.t2343 988.926
R519 VGND.n934 VGND.t292 988.926
R520 VGND.n929 VGND.t484 988.926
R521 VGND.n924 VGND.t803 988.926
R522 VGND.n919 VGND.t1142 988.926
R523 VGND.n914 VGND.t386 988.926
R524 VGND.n909 VGND.t1593 988.926
R525 VGND.n904 VGND.t1565 988.926
R526 VGND.n1962 VGND.t2330 988.926
R527 VGND.n1961 VGND.t2031 988.926
R528 VGND.n1956 VGND.t376 988.926
R529 VGND.t2376 VGND.n1395 988.926
R530 VGND.t1128 VGND.n1400 988.926
R531 VGND.n1401 VGND.t1704 988.926
R532 VGND.t1299 VGND.n1823 988.926
R533 VGND.n1824 VGND.t625 988.926
R534 VGND.t288 VGND.n1849 988.926
R535 VGND.n1850 VGND.t478 988.926
R536 VGND.t6 VGND.n1875 988.926
R537 VGND.n1876 VGND.t1136 988.926
R538 VGND.t2600 VGND.n1901 988.926
R539 VGND.n1902 VGND.t1589 988.926
R540 VGND.t1561 VGND.n1932 988.926
R541 VGND.t846 VGND.n1937 988.926
R542 VGND.t258 VGND.n1942 988.926
R543 VGND.n1943 VGND.t372 988.926
R544 VGND.t765 VGND.n1380 988.926
R545 VGND.n1381 VGND.t1359 988.926
R546 VGND.t1983 VGND.n1810 988.926
R547 VGND.n1811 VGND.t2199 988.926
R548 VGND.t260 VGND.n1836 988.926
R549 VGND.n1837 VGND.t332 988.926
R550 VGND.t505 VGND.n1862 988.926
R551 VGND.n1863 VGND.t313 988.926
R552 VGND.t914 VGND.n1888 988.926
R553 VGND.n1889 VGND.t368 988.926
R554 VGND.t305 VGND.n1914 988.926
R555 VGND.n1920 VGND.t2513 988.926
R556 VGND.n1919 VGND.t111 988.926
R557 VGND.t1535 VGND.n2357 988.926
R558 VGND.n2358 VGND.t519 988.926
R559 VGND.t990 VGND.n1312 988.926
R560 VGND.n1363 VGND.t2165 988.926
R561 VGND.n1362 VGND.t355 988.926
R562 VGND.n1357 VGND.t2635 988.926
R563 VGND.n1352 VGND.t2129 988.926
R564 VGND.n1347 VGND.t299 988.926
R565 VGND.n1342 VGND.t2681 988.926
R566 VGND.n1337 VGND.t1148 988.926
R567 VGND.n1332 VGND.t2177 988.926
R568 VGND.n1327 VGND.t2594 988.926
R569 VGND.n1322 VGND.t1388 988.926
R570 VGND.n1317 VGND.t1659 988.926
R571 VGND.n1788 VGND.t839 988.926
R572 VGND.n1787 VGND.t1111 988.926
R573 VGND.n1782 VGND.t2584 988.926
R574 VGND.t278 VGND.n1517 988.926
R575 VGND.t2167 VGND.n1522 988.926
R576 VGND.n1523 VGND.t60 988.926
R577 VGND.t1549 VGND.n1649 988.926
R578 VGND.n1650 VGND.t1616 988.926
R579 VGND.t920 VGND.n1675 988.926
R580 VGND.n1676 VGND.t2573 988.926
R581 VGND.t993 VGND.n1701 988.926
R582 VGND.n1702 VGND.t648 988.926
R583 VGND.t2563 VGND.n1727 988.926
R584 VGND.n1728 VGND.t2155 988.926
R585 VGND.t1528 VGND.n1758 988.926
R586 VGND.t104 VGND.n1763 988.926
R587 VGND.t732 VGND.n1768 988.926
R588 VGND.n1769 VGND.t511 988.926
R589 VGND.t988 VGND.n1537 988.926
R590 VGND.n1538 VGND.t2163 988.926
R591 VGND.t357 VGND.n1636 988.926
R592 VGND.n1637 VGND.t2633 988.926
R593 VGND.t2247 VGND.n1662 988.926
R594 VGND.n1663 VGND.t297 988.926
R595 VGND.t2679 VGND.n1688 988.926
R596 VGND.n1689 VGND.t1146 988.926
R597 VGND.t2175 VGND.n1714 988.926
R598 VGND.n1715 VGND.t2592 988.926
R599 VGND.t1386 VGND.n1740 988.926
R600 VGND.n1746 VGND.t1577 988.926
R601 VGND.n1745 VGND.t837 988.926
R602 VGND.t1109 VGND.n2382 988.926
R603 VGND.n2383 VGND.t2582 988.926
R604 VGND.n1295 VGND.t469 988.926
R605 VGND.t643 VGND.n1550 988.926
R606 VGND.t9 VGND.n1555 988.926
R607 VGND.t1165 VGND.n1560 988.926
R608 VGND.t2150 VGND.n1565 988.926
R609 VGND.t432 VGND.n1570 988.926
R610 VGND.t501 VGND.n1575 988.926
R611 VGND.t737 VGND.n1580 988.926
R612 VGND.t123 VGND.n1585 988.926
R613 VGND.t405 VGND.n1590 988.926
R614 VGND.t2037 VGND.n1595 988.926
R615 VGND.t116 VGND.n1600 988.926
R616 VGND.n1614 VGND.t604 988.926
R617 VGND.n1613 VGND.t2535 988.926
R618 VGND.n1608 VGND.t427 988.926
R619 VGND.t2378 VGND.n835 988.926
R620 VGND.t1130 VGND.n840 988.926
R621 VGND.n891 VGND.t1702 988.926
R622 VGND.n890 VGND.t1301 988.926
R623 VGND.n885 VGND.t627 988.926
R624 VGND.n880 VGND.t286 988.926
R625 VGND.n875 VGND.t476 988.926
R626 VGND.n870 VGND.t4 988.926
R627 VGND.n865 VGND.t1403 988.926
R628 VGND.n860 VGND.t2598 988.926
R629 VGND.n855 VGND.t1587 988.926
R630 VGND.n850 VGND.t1559 988.926
R631 VGND.n845 VGND.t844 988.926
R632 VGND.t2027 VGND.n2402 988.926
R633 VGND.n2403 VGND.t2590 988.926
R634 VGND.n1289 VGND.t1082 988.926
R635 VGND.t1256 VGND.n720 988.926
R636 VGND.t1234 VGND.n725 988.926
R637 VGND.t1077 VGND.n730 988.926
R638 VGND.t1066 VGND.n735 988.926
R639 VGND.t1047 VGND.n740 988.926
R640 VGND.t211 VGND.n745 988.926
R641 VGND.t190 VGND.n750 988.926
R642 VGND.t1043 VGND.n755 988.926
R643 VGND.t1222 VGND.n760 988.926
R644 VGND.t1209 VGND.n765 988.926
R645 VGND.t1101 VGND.n770 988.926
R646 VGND.t1026 VGND.n775 988.926
R647 VGND.t1191 VGND.n780 988.926
R648 VGND.n781 VGND.t2095 988.926
R649 VGND.n1508 VGND.n579 934.784
R650 VGND.n2907 VGND 927.203
R651 VGND.n2910 VGND 927.203
R652 VGND.n962 VGND 918.774
R653 VGND.n113 VGND 910.346
R654 VGND.n2874 VGND 910.346
R655 VGND.n3008 VGND.t1502 909.365
R656 VGND.n2833 VGND.n177 900
R657 VGND.n2578 VGND.t2617 852.769
R658 VGND.n2705 VGND.t1334 852.769
R659 VGND.t1161 VGND.n2704 852.769
R660 VGND.n2697 VGND.t2148 852.769
R661 VGND.t2070 VGND.n2696 852.769
R662 VGND.n2689 VGND.t236 852.769
R663 VGND.t1009 VGND.n2688 852.769
R664 VGND.n2681 VGND.t657 852.769
R665 VGND.t1666 VGND.n2680 852.769
R666 VGND.n2673 VGND.t1583 852.769
R667 VGND.t595 VGND.n2672 852.769
R668 VGND.n2665 VGND.t1732 852.769
R669 VGND.t1157 VGND.n2664 852.769
R670 VGND.n2657 VGND.t1376 852.769
R671 VGND.t599 VGND.n2656 852.769
R672 VGND.t1162 VGND.n33 852.769
R673 VGND.n233 VGND.t1689 852.769
R674 VGND.n2719 VGND.t895 852.769
R675 VGND.n2724 VGND.t1668 852.769
R676 VGND.n2729 VGND.t1371 852.769
R677 VGND.n2734 VGND.t1677 852.769
R678 VGND.n2739 VGND.t184 852.769
R679 VGND.n2744 VGND.t403 852.769
R680 VGND.n2749 VGND.t1656 852.769
R681 VGND.n2754 VGND.t810 852.769
R682 VGND.n2759 VGND.t2054 852.769
R683 VGND.n2764 VGND.t28 852.769
R684 VGND.n2769 VGND.t1663 852.769
R685 VGND.n2774 VGND.t2353 852.769
R686 VGND.n2779 VGND.t0 852.769
R687 VGND.n2780 VGND.t1135 852.769
R688 VGND.n2999 VGND.t2320 852.769
R689 VGND.n2514 VGND.t2606 852.769
R690 VGND.t1008 VGND.n2513 852.769
R691 VGND.t2360 VGND.n2508 852.769
R692 VGND.n2433 VGND.t2180 852.769
R693 VGND.n2438 VGND.t440 852.769
R694 VGND.n2443 VGND.t2034 852.769
R695 VGND.n2448 VGND.t2043 852.769
R696 VGND.n2453 VGND.t1510 852.769
R697 VGND.n2458 VGND.t1106 852.769
R698 VGND.n2463 VGND.t1124 852.769
R699 VGND.n2468 VGND.t150 852.769
R700 VGND.n2473 VGND.t2035 852.769
R701 VGND.n2478 VGND.t1363 852.769
R702 VGND.n2483 VGND.t2631 852.769
R703 VGND.n2488 VGND.t2144 852.769
R704 VGND.n2489 VGND.t723 852.769
R705 VGND.t2400 VGND.n2831 852.769
R706 VGND.n371 VGND.t2354 852.769
R707 VGND.n372 VGND.t115 852.769
R708 VGND.n2171 VGND.t1370 852.769
R709 VGND.n2172 VGND.t2045 852.769
R710 VGND.n2197 VGND.t1113 852.769
R711 VGND.n2198 VGND.t1505 852.769
R712 VGND.n2223 VGND.t659 852.769
R713 VGND.n2224 VGND.t900 852.769
R714 VGND.n2249 VGND.t336 852.769
R715 VGND.n2250 VGND.t1980 852.769
R716 VGND.n2280 VGND.t1710 852.769
R717 VGND.n2285 VGND.t251 852.769
R718 VGND.n2290 VGND.t152 852.769
R719 VGND.n2291 VGND.t2162 852.769
R720 VGND.n2428 VGND.t29 852.769
R721 VGND.n1428 VGND.t1353 852.769
R722 VGND.n1429 VGND.t276 852.769
R723 VGND.n2158 VGND.t566 852.769
R724 VGND.n2159 VGND.t1716 852.769
R725 VGND.n2184 VGND.t183 852.769
R726 VGND.n2185 VGND.t1712 852.769
R727 VGND.n2210 VGND.t888 852.769
R728 VGND.n2211 VGND.t2642 852.769
R729 VGND.n2236 VGND.t2605 852.769
R730 VGND.n2237 VGND.t2146 852.769
R731 VGND.n2262 VGND.t2359 852.769
R732 VGND.n2268 VGND.t1385 852.769
R733 VGND.t1489 VGND.n2267 852.769
R734 VGND.n2307 VGND.t1696 852.769
R735 VGND.n2308 VGND.t22 852.769
R736 VGND.t1123 VGND.n261 852.769
R737 VGND.n1442 VGND.t2055 852.769
R738 VGND.n1493 VGND.t797 852.769
R739 VGND.t2044 VGND.n1492 852.769
R740 VGND.t1655 VGND.n1487 852.769
R741 VGND.t2068 VGND.n1482 852.769
R742 VGND.t2358 VGND.n1477 852.769
R743 VGND.t404 VGND.n1472 852.769
R744 VGND.t120 VGND.n1467 852.769
R745 VGND.t1006 VGND.n1462 852.769
R746 VGND.t2632 VGND.n1457 852.769
R747 VGND.t2133 VGND.n1452 852.769
R748 VGND.t1669 VGND.n1447 852.769
R749 VGND.n2136 VGND.t1654 852.769
R750 VGND.t911 VGND.n2135 852.769
R751 VGND.t987 VGND.n2130 852.769
R752 VGND.t2649 VGND.n262 852.769
R753 VGND.t8 VGND.n1504 852.769
R754 VGND.n626 VGND.t2438 852.769
R755 VGND.n627 VGND.t2685 852.769
R756 VGND.n1997 VGND.t220 852.769
R757 VGND.n1998 VGND.t539 852.769
R758 VGND.n2023 VGND.t1367 852.769
R759 VGND.n2024 VGND.t2355 852.769
R760 VGND.n2049 VGND.t2351 852.769
R761 VGND.n2050 VGND.t141 852.769
R762 VGND.n2075 VGND.t572 852.769
R763 VGND.n2076 VGND.t1507 852.769
R764 VGND.n2106 VGND.t2402 852.769
R765 VGND.n2111 VGND.t658 852.769
R766 VGND.n2116 VGND.t1005 852.769
R767 VGND.n2117 VGND.t1741 852.769
R768 VGND.t265 VGND.n263 852.769
R769 VGND.n652 VGND.t1160 852.769
R770 VGND.n653 VGND.t397 852.769
R771 VGND.n1984 VGND.t979 852.769
R772 VGND.n1985 VGND.t2036 852.769
R773 VGND.n2010 VGND.t153 852.769
R774 VGND.n2011 VGND.t255 852.769
R775 VGND.n2036 VGND.t30 852.769
R776 VGND.n2037 VGND.t252 852.769
R777 VGND.n2062 VGND.t1664 852.769
R778 VGND.n2063 VGND.t1509 852.769
R779 VGND.n2088 VGND.t2432 852.769
R780 VGND.n2094 VGND.t1582 852.769
R781 VGND.t806 VGND.n2093 852.769
R782 VGND.n2332 VGND.t796 852.769
R783 VGND.n2333 VGND.t1674 852.769
R784 VGND.t1356 VGND.n264 852.769
R785 VGND.t538 VGND.n959 852.769
R786 VGND.t1155 VGND.n954 852.769
R787 VGND.t88 VGND.n949 852.769
R788 VGND.t235 VGND.n944 852.769
R789 VGND.t598 VGND.n939 852.769
R790 VGND.t1144 VGND.n934 852.769
R791 VGND.t1584 VGND.n929 852.769
R792 VGND.t760 VGND.n924 852.769
R793 VGND.t1105 VGND.n919 852.769
R794 VGND.t2185 VGND.n914 852.769
R795 VGND.t597 VGND.n909 852.769
R796 VGND.t396 VGND.n904 852.769
R797 VGND.n1962 VGND.t1352 852.769
R798 VGND.t1004 VGND.n1961 852.769
R799 VGND.t127 VGND.n1956 852.769
R800 VGND.t25 VGND.n265 852.769
R801 VGND.n1395 VGND.t2630 852.769
R802 VGND.n1400 VGND.t1639 852.769
R803 VGND.n1401 VGND.t1512 852.769
R804 VGND.n1823 VGND.t537 852.769
R805 VGND.n1824 VGND.t2641 852.769
R806 VGND.n1849 VGND.t1372 852.769
R807 VGND.n1850 VGND.t1678 852.769
R808 VGND.n1875 VGND.t185 852.769
R809 VGND.n1876 VGND.t1697 852.769
R810 VGND.n1901 VGND.t1122 852.769
R811 VGND.n1902 VGND.t620 852.769
R812 VGND.n1932 VGND.t1679 852.769
R813 VGND.n1937 VGND.t87 852.769
R814 VGND.n1942 VGND.t1398 852.769
R815 VGND.n1943 VGND.t327 852.769
R816 VGND.t1369 VGND.n266 852.769
R817 VGND.n1380 VGND.t2437 852.769
R818 VGND.n1381 VGND.t2643 852.769
R819 VGND.n1810 VGND.t1506 852.769
R820 VGND.n1811 VGND.t1357 852.769
R821 VGND.n1836 VGND.t594 852.769
R822 VGND.n1837 VGND.t250 852.769
R823 VGND.n1862 VGND.t1007 852.769
R824 VGND.n1863 VGND.t129 852.769
R825 VGND.n1888 VGND.t1581 852.769
R826 VGND.n1889 VGND.t2075 852.769
R827 VGND.n1914 VGND.t1711 852.769
R828 VGND.n1920 VGND.t601 852.769
R829 VGND.t2267 VGND.n1919 852.769
R830 VGND.n2357 VGND.t1154 852.769
R831 VGND.n2358 VGND.t1729 852.769
R832 VGND.t2006 VGND.n267 852.769
R833 VGND.n1312 VGND.t1490 852.769
R834 VGND.n1363 VGND.t1152 852.769
R835 VGND.t147 VGND.n1362 852.769
R836 VGND.t593 VGND.n1357 852.769
R837 VGND.t1461 VGND.n1352 852.769
R838 VGND.t2266 VGND.n1347 852.769
R839 VGND.t1730 VGND.n1342 852.769
R840 VGND.t1508 VGND.n1337 852.769
R841 VGND.t1657 VGND.n1332 852.769
R842 VGND.t574 VGND.n1327 852.769
R843 VGND.t2644 VGND.n1322 852.769
R844 VGND.t151 VGND.n1317 852.769
R845 VGND.n1788 VGND.t1979 852.769
R846 VGND.t2069 VGND.n1787 852.769
R847 VGND.t182 VGND.n1782 852.769
R848 VGND.t1366 VGND.n268 852.769
R849 VGND.n1517 VGND.t621 852.769
R850 VGND.n1522 VGND.t887 852.769
R851 VGND.n1523 VGND.t2120 852.769
R852 VGND.n1649 VGND.t1690 852.769
R853 VGND.n1650 VGND.t696 852.769
R854 VGND.n1675 VGND.t1667 852.769
R855 VGND.n1676 VGND.t743 852.769
R856 VGND.n1701 VGND.t2265 852.769
R857 VGND.n1702 VGND.t1364 852.769
R858 VGND.n1727 VGND.t1405 852.769
R859 VGND.n1728 VGND.t119 852.769
R860 VGND.n1758 VGND.t573 852.769
R861 VGND.n1763 VGND.t2361 852.769
R862 VGND.n1768 VGND.t277 852.769
R863 VGND.n1769 VGND.t1392 852.769
R864 VGND.t2399 VGND.n269 852.769
R865 VGND.n1537 VGND.t15 852.769
R866 VGND.n1538 VGND.t26 852.769
R867 VGND.n1636 VGND.t912 852.769
R868 VGND.n1637 VGND.t896 852.769
R869 VGND.n1662 VGND.t128 852.769
R870 VGND.n1663 VGND.t1675 852.769
R871 VGND.n1688 VGND.t253 852.769
R872 VGND.n1689 VGND.t1156 852.769
R873 VGND.n1714 VGND.t2188 852.769
R874 VGND.n1715 VGND.t1462 852.769
R875 VGND.n1740 VGND.t2684 852.769
R876 VGND.n1746 VGND.t741 852.769
R877 VGND.t1107 VGND.n1745 852.769
R878 VGND.n2382 VGND.t1665 852.769
R879 VGND.n2383 VGND.t540 852.769
R880 VGND.t894 VGND.n270 852.769
R881 VGND.n1295 VGND.t2321 852.769
R882 VGND.n1550 VGND.t2161 852.769
R883 VGND.n1555 VGND.t181 852.769
R884 VGND.n1560 VGND.t254 852.769
R885 VGND.n1565 VGND.t27 852.769
R886 VGND.n1570 VGND.t1354 852.769
R887 VGND.n1575 VGND.t2686 852.769
R888 VGND.n1580 VGND.t2053 852.769
R889 VGND.n1585 VGND.t23 852.769
R890 VGND.n1590 VGND.t499 852.769
R891 VGND.n1595 VGND.t742 852.769
R892 VGND.n1600 VGND.t1396 852.769
R893 VGND.n1614 VGND.t1680 852.769
R894 VGND.t571 VGND.n1613 852.769
R895 VGND.t521 VGND.n1608 852.769
R896 VGND.t1368 VGND.n271 852.769
R897 VGND.n835 VGND.t759 852.769
R898 VGND.n840 VGND.t757 852.769
R899 VGND.n891 VGND.t2264 852.769
R900 VGND.t2147 VGND.n890 852.769
R901 VGND.t2179 VGND.n885 852.769
R902 VGND.t761 VGND.n880 852.769
R903 VGND.t2405 VGND.n875 852.769
R904 VGND.t1513 VGND.n870 852.769
R905 VGND.t275 VGND.n865 852.769
R906 VGND.t596 VGND.n860 852.769
R907 VGND.t1731 VGND.n855 852.769
R908 VGND.t809 VGND.n850 852.769
R909 VGND.t758 VGND.n845 852.769
R910 VGND.n2402 VGND.t565 852.769
R911 VGND.n2403 VGND.t1003 852.769
R912 VGND.t769 VGND.n272 852.769
R913 VGND.t180 VGND.n1289 852.769
R914 VGND.n720 VGND.t1335 852.769
R915 VGND.n725 VGND.t1358 852.769
R916 VGND.n730 VGND.t219 852.769
R917 VGND.n735 VGND.t249 852.769
R918 VGND.n740 VGND.t899 852.769
R919 VGND.n745 VGND.t89 852.769
R920 VGND.n750 VGND.t893 852.769
R921 VGND.n755 VGND.t2604 852.769
R922 VGND.n760 VGND.t2401 852.769
R923 VGND.n765 VGND.t1397 852.769
R924 VGND.n770 VGND.t1307 852.769
R925 VGND.n775 VGND.t1355 852.769
R926 VGND.n780 VGND.t63 852.769
R927 VGND.n781 VGND.t1158 852.769
R928 VGND.n2413 VGND.t140 852.769
R929 VGND.n1507 VGND 851.341
R930 VGND.n2841 VGND.t1232 809.773
R931 VGND.n2840 VGND.t1881 809.773
R932 VGND.t1956 VGND.n114 809.773
R933 VGND.n2832 VGND.t1863 809.773
R934 VGND.t1905 VGND.n177 809.773
R935 VGND.t1977 VGND.n635 809.773
R936 VGND.t1857 VGND.n580 809.773
R937 VGND.n960 VGND.t1899 809.773
R938 VGND.t1911 VGND.n579 809.773
R939 VGND.n1511 VGND.t1935 809.773
R940 VGND.t1866 VGND.n1512 809.773
R941 VGND.n1293 VGND.t1938 809.773
R942 VGND.t1968 VGND.n1294 809.773
R943 VGND.n1292 VGND.t1908 809.773
R944 VGND.n1290 VGND.t1177 809.773
R945 VGND.t1768 VGND.t1750 708.047
R946 VGND.t1750 VGND.t1748 708.047
R947 VGND.t1748 VGND.t1758 708.047
R948 VGND.t1758 VGND.t40 708.047
R949 VGND.t40 VGND.t37 708.047
R950 VGND.t37 VGND.t43 708.047
R951 VGND.t43 VGND.t34 708.047
R952 VGND.t2367 VGND.t31 708.047
R953 VGND.t1795 VGND.t1782 708.047
R954 VGND.t1782 VGND.t1780 708.047
R955 VGND.t1780 VGND.t1742 708.047
R956 VGND.t1742 VGND.t1348 708.047
R957 VGND.t1348 VGND.t503 708.047
R958 VGND.t503 VGND.t897 708.047
R959 VGND.t897 VGND.t1150 708.047
R960 VGND.t1819 VGND.t1766 708.047
R961 VGND.t1766 VGND.t1807 708.047
R962 VGND.t1807 VGND.t1775 708.047
R963 VGND.t1775 VGND.t755 708.047
R964 VGND.t755 VGND.t751 708.047
R965 VGND.t751 VGND.t745 708.047
R966 VGND.t745 VGND.t747 708.047
R967 VGND.t2364 VGND.t32 708.047
R968 VGND.t1803 VGND.t1764 708.047
R969 VGND.t1772 VGND.t1803 708.047
R970 VGND.t1746 VGND.t1772 708.047
R971 VGND.t36 VGND.t1746 708.047
R972 VGND.t42 VGND.t36 708.047
R973 VGND.t39 VGND.t42 708.047
R974 VGND.t45 VGND.t39 708.047
R975 VGND.t1760 VGND.t1799 708.047
R976 VGND.t1799 VGND.t1770 708.047
R977 VGND.t1770 VGND.t1778 708.047
R978 VGND.t1778 VGND.t978 708.047
R979 VGND.t978 VGND.t1569 708.047
R980 VGND.t1569 VGND.t486 708.047
R981 VGND.t486 VGND.t1492 708.047
R982 VGND.t1812 VGND.t1756 708.047
R983 VGND.t1756 VGND.t1817 708.047
R984 VGND.t1817 VGND.t1789 708.047
R985 VGND.t1789 VGND.t753 708.047
R986 VGND.t753 VGND.t749 708.047
R987 VGND.t749 VGND.t754 708.047
R988 VGND.t754 VGND.t750 708.047
R989 VGND.n2994 VGND.n2993 708.047
R990 VGND.t2433 VGND.t1374 691.188
R991 VGND.t901 VGND.t535 691.188
R992 VGND.n2837 VGND.t2537 685.545
R993 VGND.n3017 VGND.t2537 685.545
R994 VGND.n2840 VGND.n2839 660.87
R995 VGND.t2656 VGND.t527 657.471
R996 VGND.t2390 VGND.t525 657.471
R997 VGND.t1682 VGND.t523 657.471
R998 VGND.t318 VGND.t875 657.471
R999 VGND.t1823 VGND.t1801 657.471
R1000 VGND.t1797 VGND.t1503 657.471
R1001 VGND.t1834 VGND.t1499 657.471
R1002 VGND.t1784 VGND.t1493 657.471
R1003 VGND.t875 VGND.t877 654.197
R1004 VGND.t1801 VGND.t1827 654.197
R1005 VGND.n962 VGND 640.614
R1006 VGND VGND.n113 640.614
R1007 VGND VGND.n2874 640.614
R1008 VGND VGND.n2907 640.614
R1009 VGND.n2910 VGND 632.184
R1010 VGND.t1062 VGND.t203 630.62
R1011 VGND.t1244 VGND.t1058 630.62
R1012 VGND.t1236 VGND.t1231 630.62
R1013 VGND.t2106 VGND.t1216 630.62
R1014 VGND.t196 VGND.t1054 630.62
R1015 VGND.t1218 VGND.t1036 630.62
R1016 VGND.t1022 VGND.t198 630.62
R1017 VGND.t2094 VGND.t192 630.62
R1018 VGND.t2090 VGND.t1024 630.62
R1019 VGND.t1219 VGND.t1038 630.62
R1020 VGND.t1199 VGND.t2092 630.62
R1021 VGND.t1097 VGND.t1184 630.62
R1022 VGND.t1020 VGND.t1015 630.62
R1023 VGND.t1188 VGND.t1264 630.62
R1024 VGND.t1248 VGND.t214 630.62
R1025 VGND.t1090 VGND.t1012 630.62
R1026 VGND.t1459 VGND.t2231 630.62
R1027 VGND.t1555 VGND.t1126 630.62
R1028 VGND.t1706 VGND.t2666 630.62
R1029 VGND.t1541 VGND.t2664 630.62
R1030 VGND.t623 VGND.t2229 630.62
R1031 VGND.t437 VGND.t589 630.62
R1032 VGND.t474 VGND.t587 630.62
R1033 VGND.t2 VGND.t2227 630.62
R1034 VGND.t1134 VGND.t2225 630.62
R1035 VGND.t2597 VGND.t591 630.62
R1036 VGND.t2042 VGND.t2662 630.62
R1037 VGND.t1662 VGND.t2660 630.62
R1038 VGND.t842 VGND.t585 630.62
R1039 VGND.t257 VGND.t2670 630.62
R1040 VGND.t379 VGND.t2668 630.62
R1041 VGND.t2223 VGND.t1098 630.62
R1042 VGND.t986 VGND.t2123 630.62
R1043 VGND.t1733 VGND.t640 630.62
R1044 VGND.t231 VGND.t55 630.62
R1045 VGND.t1164 VGND.t229 630.62
R1046 VGND.t1615 VGND.t2121 630.62
R1047 VGND.t285 VGND.t2239 630.62
R1048 VGND.t2572 VGND.t2237 630.62
R1049 VGND.t992 VGND.t1739 630.62
R1050 VGND.t647 VGND.t1737 630.62
R1051 VGND.t366 VGND.t2241 630.62
R1052 VGND.t1586 VGND.t2127 630.62
R1053 VGND.t1534 VGND.t2125 630.62
R1054 VGND.t103 VGND.t2235 630.62
R1055 VGND.t891 VGND.t2233 630.62
R1056 VGND.t426 VGND.t233 630.62
R1057 VGND.t1203 VGND.t1735 630.62
R1058 VGND.t2258 VGND.t2375 630.62
R1059 VGND.t1132 VGND.t1628 630.62
R1060 VGND.t360 VGND.t1636 630.62
R1061 VGND.t1634 VGND.t1547 630.62
R1062 VGND.t629 VGND.t2256 630.62
R1063 VGND.t1624 VGND.t439 630.62
R1064 VGND.t480 VGND.t1622 630.62
R1065 VGND.t2254 VGND.t799 630.62
R1066 VGND.t1138 VGND.t2252 630.62
R1067 VGND.t1626 VGND.t389 630.62
R1068 VGND.t1297 VGND.t1632 630.62
R1069 VGND.t1630 VGND.t1538 630.62
R1070 VGND.t848 VGND.t1620 630.62
R1071 VGND.t416 VGND.t2262 630.62
R1072 VGND.t385 VGND.t2260 630.62
R1073 VGND.t2250 VGND.t2104 630.62
R1074 VGND.t632 VGND.t2203 630.62
R1075 VGND.t2088 VGND.t2195 630.62
R1076 VGND.t575 VGND.t11 630.62
R1077 VGND.t2639 VGND.t2209 630.62
R1078 VGND.t1383 VGND.t2245 630.62
R1079 VGND.t330 VGND.t2191 630.62
R1080 VGND.t2189 VGND.t2677 630.62
R1081 VGND.t1395 VGND.t1381 630.62
R1082 VGND.t1379 VGND.t1401 630.62
R1083 VGND.t413 VGND.t2193 630.62
R1084 VGND.t2207 VGND.t303 630.62
R1085 VGND.t1575 VGND.t2205 630.62
R1086 VGND.t581 VGND.t610 630.62
R1087 VGND.t579 VGND.t2184 630.62
R1088 VGND.t2588 VGND.t577 630.62
R1089 VGND.t1377 VGND.t1053 630.62
R1090 VGND.t980 VGND.t1646 630.62
R1091 VGND.t634 VGND.t2140 630.62
R1092 VGND.t1557 VGND.t2347 630.62
R1093 VGND.t1652 VGND.t2198 630.62
R1094 VGND.t1644 VGND.t2135 630.62
R1095 VGND.t2136 VGND.t419 630.62
R1096 VGND.t2013 VGND.t2566 630.62
R1097 VGND.t1642 VGND.t724 630.62
R1098 VGND.t1640 VGND.t2047 630.62
R1099 VGND.t2138 VGND.t2561 630.62
R1100 VGND.t1650 VGND.t1391 630.62
R1101 VGND.t1648 VGND.t2024 630.62
R1102 VGND.t2011 VGND.t2333 630.62
R1103 VGND.t2009 VGND.t730 630.62
R1104 VGND.t2007 VGND.t518 630.62
R1105 VGND.t2142 VGND.t1175 630.62
R1106 VGND.t1600 VGND.t1458 630.62
R1107 VGND.t1125 VGND.t69 630.62
R1108 VGND.t359 VGND.t1608 630.62
R1109 VGND.t1606 VGND.t1540 630.62
R1110 VGND.t622 VGND.t1598 630.62
R1111 VGND.t1725 VGND.t436 630.62
R1112 VGND.t473 VGND.t1723 630.62
R1113 VGND.t1596 VGND.t1 630.62
R1114 VGND.t1133 VGND.t73 630.62
R1115 VGND.t1727 VGND.t2596 630.62
R1116 VGND.t2041 VGND.t1604 630.62
R1117 VGND.t1602 VGND.t1661 630.62
R1118 VGND.t841 VGND.t1721 630.62
R1119 VGND.t256 VGND.t1719 630.62
R1120 VGND.t378 VGND.t1717 630.62
R1121 VGND.t71 VGND.t1096 630.62
R1122 VGND.t2380 VGND.t1996 630.62
R1123 VGND.t64 VGND.t1523 630.62
R1124 VGND.t2004 VGND.t1707 630.62
R1125 VGND.t1548 VGND.t2002 630.62
R1126 VGND.t1994 VGND.t2340 630.62
R1127 VGND.t296 VGND.t1519 630.62
R1128 VGND.t1517 VGND.t481 630.62
R1129 VGND.t800 VGND.t1992 630.62
R1130 VGND.t1990 VGND.t1139 630.62
R1131 VGND.t390 VGND.t1521 630.62
R1132 VGND.t2000 VGND.t1298 630.62
R1133 VGND.t1539 VGND.t1998 630.62
R1134 VGND.t1515 VGND.t2327 630.62
R1135 VGND.t353 VGND.t417 630.62
R1136 VGND.t510 VGND.t351 630.62
R1137 VGND.t1525 VGND.t2107 630.62
R1138 VGND.t618 VGND.t633 630.62
R1139 VGND.t1120 VGND.t2089 630.62
R1140 VGND.t221 VGND.t14 630.62
R1141 VGND.t2081 VGND.t2640 630.62
R1142 VGND.t616 VGND.t2246 630.62
R1143 VGND.t1116 VGND.t331 630.62
R1144 VGND.t1114 VGND.t2678 630.62
R1145 VGND.t614 VGND.t1145 630.62
R1146 VGND.t612 VGND.t2174 630.62
R1147 VGND.t1118 VGND.t414 630.62
R1148 VGND.t2079 VGND.t304 630.62
R1149 VGND.t2077 VGND.t1576 630.62
R1150 VGND.t227 VGND.t611 630.62
R1151 VGND.t225 VGND.t1108 630.62
R1152 VGND.t223 VGND.t2589 630.62
R1153 VGND.t807 VGND.t1055 630.62
R1154 VGND.t630 VGND.t343 630.62
R1155 VGND.t2087 VGND.t497 630.62
R1156 VGND.t13 VGND.t1266 630.62
R1157 VGND.t349 VGND.t2638 630.62
R1158 VGND.t2243 VGND.t341 630.62
R1159 VGND.t493 VGND.t328 630.62
R1160 VGND.t2676 VGND.t491 630.62
R1161 VGND.t339 VGND.t1394 630.62
R1162 VGND.t1400 VGND.t337 630.62
R1163 VGND.t495 VGND.t412 630.62
R1164 VGND.t302 VGND.t347 630.62
R1165 VGND.t345 VGND.t1574 630.62
R1166 VGND.t609 VGND.t489 630.62
R1167 VGND.t2183 VGND.t487 630.62
R1168 VGND.t2586 VGND.t1268 630.62
R1169 VGND.t2338 VGND.t1046 630.62
R1170 VGND.t1514 VGND.t1338 630.62
R1171 VGND.t2687 VGND.t557 630.62
R1172 VGND.t1346 VGND.t2350 630.62
R1173 VGND.t2197 VGND.t1344 630.62
R1174 VGND.t1336 VGND.t2134 630.62
R1175 VGND.t418 VGND.t553 630.62
R1176 VGND.t551 VGND.t2565 630.62
R1177 VGND.t798 VGND.t563 630.62
R1178 VGND.t561 VGND.t2046 630.62
R1179 VGND.t393 VGND.t555 630.62
R1180 VGND.t1342 VGND.t1390 630.62
R1181 VGND.t2021 VGND.t1340 630.62
R1182 VGND.t549 VGND.t2332 630.62
R1183 VGND.t547 VGND.t144 630.62
R1184 VGND.t517 VGND.t545 630.62
R1185 VGND.t559 VGND.t1170 630.62
R1186 VGND.t468 VGND.t2517 630.62
R1187 VGND.t642 VGND.t2501 630.62
R1188 VGND.t2525 VGND.t1986 630.62
R1189 VGND.t2523 VGND.t584 630.62
R1190 VGND.t90 VGND.t2149 630.62
R1191 VGND.t2497 VGND.t919 630.62
R1192 VGND.t2495 VGND.t500 630.62
R1193 VGND.t2507 VGND.t736 630.62
R1194 VGND.t2505 VGND.t122 630.62
R1195 VGND.t2499 VGND.t410 630.62
R1196 VGND.t2521 VGND.t2154 630.62
R1197 VGND.t2519 VGND.t2511 630.62
R1198 VGND.t2531 VGND.t603 630.62
R1199 VGND.t2529 VGND.t2074 630.62
R1200 VGND.t2527 VGND.t2581 630.62
R1201 VGND.t2503 VGND.t1261 630.62
R1202 VGND.t1460 VGND.t2626 630.62
R1203 VGND.t1127 VGND.t694 630.62
R1204 VGND.t361 VGND.t2613 630.62
R1205 VGND.t2611 VGND.t1546 630.62
R1206 VGND.t624 VGND.t2624 630.62
R1207 VGND.t690 VGND.t438 630.62
R1208 VGND.t475 VGND.t688 630.62
R1209 VGND.t2622 VGND.t3 630.62
R1210 VGND.t1402 VGND.t2620 630.62
R1211 VGND.t692 VGND.t388 630.62
R1212 VGND.t1296 VGND.t2609 630.62
R1213 VGND.t2607 VGND.t1567 630.62
R1214 VGND.t843 VGND.t686 630.62
R1215 VGND.t2033 VGND.t2403 630.62
R1216 VGND.t384 VGND.t2615 630.62
R1217 VGND.t2618 VGND.t2101 630.62
R1218 VGND.t16 VGND.t467 630.62
R1219 VGND.t641 VGND.t2215 630.62
R1220 VGND.t2110 VGND.t1989 630.62
R1221 VGND.t583 VGND.t2108 630.62
R1222 VGND.t2553 VGND.t264 630.62
R1223 VGND.t918 VGND.t2211 630.62
R1224 VGND.t2118 VGND.t509 630.62
R1225 VGND.t317 VGND.t2221 630.62
R1226 VGND.t2219 VGND.t121 630.62
R1227 VGND.t407 VGND.t2213 630.62
R1228 VGND.t20 VGND.t2326 630.62
R1229 VGND.t118 VGND.t18 630.62
R1230 VGND.t2116 VGND.t602 630.62
R1231 VGND.t2114 VGND.t2071 630.62
R1232 VGND.t2580 VGND.t2112 630.62
R1233 VGND.t2217 VGND.t1258 630.62
R1234 VGND.t985 VGND.t2064 630.62
R1235 VGND.t85 VGND.t639 630.62
R1236 VGND.t62 VGND.t2015 630.62
R1237 VGND.t1163 VGND.t1572 630.62
R1238 VGND.t1614 VGND.t2062 630.62
R1239 VGND.t420 VGND.t81 630.62
R1240 VGND.t2571 VGND.t79 630.62
R1241 VGND.t729 VGND.t2060 630.62
R1242 VGND.t2052 VGND.t2058 630.62
R1243 VGND.t2562 VGND.t83 630.62
R1244 VGND.t1585 VGND.t1570 630.62
R1245 VGND.t1527 VGND.t2066 630.62
R1246 VGND.t102 VGND.t77 630.62
R1247 VGND.t75 VGND.t731 630.62
R1248 VGND.t2017 VGND.t425 630.62
R1249 VGND.t2056 VGND.t1190 630.62
R1250 VGND.t631 VGND.t268 630.62
R1251 VGND.t2086 VGND.t567 630.62
R1252 VGND.t12 VGND.t907 630.62
R1253 VGND.t905 VGND.t2637 630.62
R1254 VGND.t266 VGND.t2244 630.62
R1255 VGND.t136 VGND.t329 630.62
R1256 VGND.t134 VGND.t2675 630.62
R1257 VGND.t1693 VGND.t1393 630.62
R1258 VGND.t1691 VGND.t1399 630.62
R1259 VGND.t138 VGND.t411 630.62
R1260 VGND.t272 VGND.t301 630.62
R1261 VGND.t270 VGND.t2025 630.62
R1262 VGND.t132 VGND.t608 630.62
R1263 VGND.t130 VGND.t2182 630.62
R1264 VGND.t2587 VGND.t909 630.62
R1265 VGND.t569 VGND.t1045 630.62
R1266 VGND.t1084 VGND.t284 630.62
R1267 VGND.t2173 VGND.t1259 630.62
R1268 VGND.t1985 VGND.t1180 630.62
R1269 VGND.t1167 VGND.t207 630.62
R1270 VGND.t2085 VGND.t1073 630.62
R1271 VGND.t294 VGND.t1240 630.62
R1272 VGND.t2579 VGND.t1229 630.62
R1273 VGND.t999 VGND.t1069 630.62
R1274 VGND.t654 VGND.t1051 630.62
R1275 VGND.t367 VGND.t1242 630.62
R1276 VGND.t1595 VGND.t194 630.62
R1277 VGND.t2512 VGND.t2102 630.62
R1278 VGND.t110 VGND.t1224 630.62
R1279 VGND.t892 VGND.t1211 630.62
R1280 VGND.t429 VGND.t1186 630.62
R1281 VGND.t1030 VGND.t1215 630.62
R1282 VGND.n990 VGND.n962 599.125
R1283 VGND.n113 VGND.n112 599.125
R1284 VGND.n2874 VGND.n2873 599.125
R1285 VGND.n2907 VGND.n2906 599.125
R1286 VGND.n2911 VGND.n2910 599.125
R1287 VGND.n2922 VGND.n2921 599.125
R1288 VGND.n2994 VGND.n2992 599.125
R1289 VGND.n2961 VGND.n2960 599.125
R1290 VGND.t148 VGND 581.61
R1291 VGND.t34 VGND 573.181
R1292 VGND.t1150 VGND 573.181
R1293 VGND.t747 VGND 573.181
R1294 VGND VGND.t1495 573.181
R1295 VGND.t903 VGND 564.751
R1296 VGND.n3012 VGND 564.751
R1297 VGND.n3011 VGND 564.751
R1298 VGND.n3010 VGND 556.322
R1299 VGND VGND.t239 539.465
R1300 VGND.t2186 VGND 539.465
R1301 VGND.n1122 VGND.t1207 500.166
R1302 VGND.t2097 VGND.n1131 500.166
R1303 VGND.n1132 VGND.t1088 500.166
R1304 VGND.t1205 VGND.n1144 500.166
R1305 VGND.n1145 VGND.t1193 500.166
R1306 VGND.t1171 VGND.n1163 500.166
R1307 VGND.n1164 VGND.t1016 500.166
R1308 VGND.t1252 VGND.n1176 500.166
R1309 VGND.n1177 VGND.t215 500.166
R1310 VGND.t1071 VGND.n1195 500.166
R1311 VGND.n1196 VGND.t1060 500.166
R1312 VGND.t1227 VGND.n1208 500.166
R1313 VGND.n1209 VGND.t205 500.166
R1314 VGND.t1049 VGND.n1227 500.166
R1315 VGND.n1228 VGND.t1238 500.166
R1316 VGND.t399 VGND.n578 494.779
R1317 VGND.t877 VGND.t2555 481.877
R1318 VGND.t2555 VGND.t46 481.877
R1319 VGND.t1793 VGND.t1752 481.877
R1320 VGND.t1827 VGND.t1793 481.877
R1321 VGND.t1350 VGND 452.382
R1322 VGND.n1122 VGND.t1153 431.301
R1323 VGND.n1131 VGND.t600 431.301
R1324 VGND.n1132 VGND.t805 431.301
R1325 VGND.n1144 VGND.t1159 431.301
R1326 VGND.n1145 VGND.t2145 431.301
R1327 VGND.n1163 VGND.t2683 431.301
R1328 VGND.n1164 VGND.t295 431.301
R1329 VGND.n1176 VGND.t1676 431.301
R1330 VGND.n1177 VGND.t762 431.301
R1331 VGND.n1195 VGND.t274 431.301
R1332 VGND.n1196 VGND.t1511 431.301
R1333 VGND.n1208 VGND.t2374 431.301
R1334 VGND.n1209 VGND.t24 431.301
R1335 VGND.n1227 VGND.t2356 431.301
R1336 VGND.n1228 VGND.t1638 431.301
R1337 VGND.t913 VGND.n273 431.301
R1338 VGND.t94 VGND 419.68
R1339 VGND.n635 VGND.n147 413.043
R1340 VGND.t1893 VGND.t1232 408.469
R1341 VGND.t1842 VGND.t201 408.469
R1342 VGND.t1056 VGND.t1848 408.469
R1343 VGND.t1854 VGND.t1034 408.469
R1344 VGND.t199 VGND.t1941 408.469
R1345 VGND.t1947 VGND.t188 408.469
R1346 VGND.t1103 VGND.t1860 408.469
R1347 VGND.t1902 VGND.t1220 408.469
R1348 VGND.t1197 VGND.t1917 408.469
R1349 VGND.t1953 VGND.t1099 408.469
R1350 VGND.t1018 VGND.t1875 408.469
R1351 VGND.t1920 VGND.t1262 408.469
R1352 VGND.t217 VGND.t1959 408.469
R1353 VGND.t1971 VGND.t1086 408.469
R1354 VGND.t1250 VGND.t1887 408.469
R1355 VGND.t1182 VGND.t1929 408.469
R1356 VGND.t1487 VGND.t1881 408.469
R1357 VGND.t983 VGND.t2316 408.469
R1358 VGND.t2551 VGND.t637 408.469
R1359 VGND.t813 VGND.t2348 408.469
R1360 VGND.t2447 VGND.t1544 408.469
R1361 VGND.t1328 VGND.t1612 408.469
R1362 VGND.t873 VGND.t311 408.469
R1363 VGND.t1463 VGND.t2569 408.469
R1364 VGND.t705 VGND.t727 408.469
R1365 VGND.t2481 VGND.t2050 408.469
R1366 VGND.t964 VGND.t394 408.469
R1367 VGND.t176 VGND.t2324 408.469
R1368 VGND.t2473 VGND.t2022 408.469
R1369 VGND.t930 VGND.t100 408.469
R1370 VGND.t2280 VGND.t145 408.469
R1371 VGND.t382 VGND.t1456 408.469
R1372 VGND.t2418 VGND.t1956 408.469
R1373 VGND.t471 VGND.t774 408.469
R1374 VGND.t645 VGND.t1428 408.469
R1375 VGND.t1471 VGND.t1987 408.469
R1376 VGND.t2318 VGND.t1168 408.469
R1377 VGND.t833 VGND.t2152 408.469
R1378 VGND.t1467 VGND.t434 408.469
R1379 VGND.t2449 VGND.t2673 408.469
R1380 VGND.t1330 VGND.t739 408.469
R1381 VGND.t811 VGND.t125 408.469
R1382 VGND.t1270 VGND.t408 408.469
R1383 VGND.t1316 VGND.t2039 408.469
R1384 VGND.t865 VGND.t2509 408.469
R1385 VGND.t968 VGND.t606 408.469
R1386 VGND.t154 VGND.t2072 408.469
R1387 VGND.t2475 VGND.t430 408.469
R1388 VGND.t1863 VGND.t703 408.469
R1389 VGND.t857 VGND.t280 408.469
R1390 VGND.t960 VGND.t2169 408.469
R1391 VGND.t58 VGND.t2288 408.469
R1392 VGND.t2465 VGND.t1551 408.469
R1393 VGND.t1618 VGND.t672 408.469
R1394 VGND.t2276 VGND.t922 408.469
R1395 VGND.t2575 VGND.t1448 408.469
R1396 VGND.t2461 VGND.t995 408.469
R1397 VGND.t650 VGND.t2304 408.469
R1398 VGND.t1408 VGND.t362 408.469
R1399 VGND.t2157 VGND.t2455 408.469
R1400 VGND.t2296 VGND.t1530 408.469
R1401 VGND.t2493 VGND.t106 408.469
R1402 VGND.t1278 VGND.t734 408.469
R1403 VGND.t513 VGND.t459 408.469
R1404 VGND.t1324 VGND.t1905 408.469
R1405 VGND.t1288 VGND.t2381 408.469
R1406 VGND.t65 VGND.t717 408.469
R1407 VGND.t160 VGND.t1700 408.469
R1408 VGND.t1303 VGND.t859 408.469
R1409 VGND.t788 VGND.t2341 408.469
R1410 VGND.t290 VGND.t1450 408.469
R1411 VGND.t2467 VGND.t482 408.469
R1412 VGND.t801 VGND.t674 408.469
R1413 VGND.t2278 VGND.t1140 408.469
R1414 VGND.t2602 VGND.t2422 408.469
R1415 VGND.t666 VGND.t1591 408.469
R1416 VGND.t1563 VGND.t2270 408.469
R1417 VGND.t2328 VGND.t1412 408.469
R1418 VGND.t461 VGND.t2029 408.469
R1419 VGND.t374 VGND.t2300 408.469
R1420 VGND.t827 VGND.t1977 408.469
R1421 VGND.t2441 VGND.t767 408.469
R1422 VGND.t1361 VGND.t447 408.469
R1423 VGND.t1981 VGND.t2485 408.469
R1424 VGND.t2201 VGND.t1290 408.469
R1425 VGND.t262 VGND.t699 408.469
R1426 VGND.t334 VGND.t2469 408.469
R1427 VGND.t507 VGND.t861 408.469
R1428 VGND.t315 VGND.t792 408.469
R1429 VGND.t916 VGND.t1452 408.469
R1430 VGND.t370 VGND.t928 408.469
R1431 VGND.t307 VGND.t780 408.469
R1432 VGND.t2515 VGND.t1446 408.469
R1433 VGND.t113 VGND.t2424 408.469
R1434 VGND.t2533 VGND.t2302 408.469
R1435 VGND.t423 VGND.t2274 408.469
R1436 VGND.t1884 VGND.t1477 408.469
R1437 VGND.t2308 VGND.t981 408.469
R1438 VGND.t2541 VGND.t635 408.469
R1439 VGND.t2345 VGND.t867 408.469
R1440 VGND.t465 VGND.t1542 408.469
R1441 VGND.t1610 VGND.t1308 408.469
R1442 VGND.t853 VGND.t309 408.469
R1443 VGND.t2567 VGND.t1284 408.469
R1444 VGND.t170 VGND.t725 408.469
R1445 VGND.t2048 VGND.t948 408.469
R1446 VGND.t952 VGND.t391 408.469
R1447 VGND.t2322 VGND.t164 408.469
R1448 VGND.t944 VGND.t2019 408.469
R1449 VGND.t682 VGND.t2334 408.469
R1450 VGND.t2268 VGND.t142 408.469
R1451 VGND.t380 VGND.t1440 408.469
R1452 VGND.t2408 VGND.t1857 408.469
R1453 VGND.t2286 VGND.t282 408.469
R1454 VGND.t2171 VGND.t1416 408.469
R1455 VGND.t1294 VGND.t56 408.469
R1456 VGND.t1553 VGND.t2310 408.469
R1457 VGND.t819 VGND.t2083 408.469
R1458 VGND.t924 VGND.t1286 408.469
R1459 VGND.t2439 VGND.t2577 408.469
R1460 VGND.t997 VGND.t1314 408.469
R1461 VGND.t855 VGND.t652 408.469
R1462 VGND.t364 VGND.t711 408.469
R1463 VGND.t2487 VGND.t2159 408.469
R1464 VGND.t1532 VGND.t851 408.469
R1465 VGND.t108 VGND.t954 408.469
R1466 VGND.t1442 VGND.t889 408.469
R1467 VGND.t515 VGND.t946 408.469
R1468 VGND.t1899 VGND.t168 408.469
R1469 VGND.t2383 VGND.t974 408.469
R1470 VGND.t67 VGND.t794 408.469
R1471 VGND.t1698 VGND.t2272 408.469
R1472 VGND.t1305 VGND.t936 408.469
R1473 VGND.t2343 VGND.t662 408.469
R1474 VGND.t292 VGND.t1422 408.469
R1475 VGND.t484 VGND.t1434 408.469
R1476 VGND.t803 VGND.t2453 408.469
R1477 VGND.t1142 VGND.t2549 408.469
R1478 VGND.t386 VGND.t1483 408.469
R1479 VGND.t1593 VGND.t2443 408.469
R1480 VGND.t1565 VGND.t2543 408.469
R1481 VGND.t2330 VGND.t831 408.469
R1482 VGND.t2031 VGND.t719 408.469
R1483 VGND.t376 VGND.t449 408.469
R1484 VGND.t2489 VGND.t1911 408.469
R1485 VGND.t1280 VGND.t2376 408.469
R1486 VGND.t709 VGND.t1128 408.469
R1487 VGND.t1704 VGND.t1444 408.469
R1488 VGND.t976 VGND.t1299 408.469
R1489 VGND.t625 VGND.t776 408.469
R1490 VGND.t1436 VGND.t288 408.469
R1491 VGND.t478 VGND.t938 408.469
R1492 VGND.t664 VGND.t6 408.469
R1493 VGND.t1136 VGND.t1426 408.469
R1494 VGND.t2412 VGND.t2600 408.469
R1495 VGND.t1589 VGND.t2314 408.469
R1496 VGND.t1418 VGND.t1561 408.469
R1497 VGND.t1485 VGND.t846 408.469
R1498 VGND.t451 VGND.t258 408.469
R1499 VGND.t372 VGND.t2545 408.469
R1500 VGND.t817 VGND.t1839 408.469
R1501 VGND.t463 VGND.t765 408.469
R1502 VGND.t1359 VGND.t445 408.469
R1503 VGND.t950 VGND.t1983 408.469
R1504 VGND.t2199 VGND.t1282 408.469
R1505 VGND.t166 VGND.t260 408.469
R1506 VGND.t332 VGND.t940 408.469
R1507 VGND.t849 VGND.t505 408.469
R1508 VGND.t313 VGND.t778 408.469
R1509 VGND.t1438 VGND.t914 408.469
R1510 VGND.t368 VGND.t680 408.469
R1511 VGND.t770 VGND.t305 408.469
R1512 VGND.t2513 VGND.t1432 408.469
R1513 VGND.t111 VGND.t2414 408.469
R1514 VGND.t2547 VGND.t1535 408.469
R1515 VGND.t519 VGND.t1420 408.469
R1516 VGND.t2416 VGND.t1935 408.469
R1517 VGND.t2292 VGND.t990 408.469
R1518 VGND.t2165 VGND.t1424 408.469
R1519 VGND.t355 VGND.t1469 408.469
R1520 VGND.t2635 VGND.t2312 408.469
R1521 VGND.t2129 VGND.t829 408.469
R1522 VGND.t299 VGND.t1292 408.469
R1523 VGND.t2681 VGND.t2445 408.469
R1524 VGND.t1148 VGND.t1326 408.469
R1525 VGND.t2177 VGND.t869 408.469
R1526 VGND.t2594 VGND.t721 408.469
R1527 VGND.t1388 VGND.t1310 408.469
R1528 VGND.t1659 VGND.t863 408.469
R1529 VGND.t839 VGND.t962 408.469
R1530 VGND.t1111 VGND.t1454 408.469
R1531 VGND.t2584 VGND.t2471 408.469
R1532 VGND.t815 VGND.t1866 408.469
R1533 VGND.t455 VGND.t278 408.469
R1534 VGND.t441 VGND.t2167 408.469
R1535 VGND.t60 VGND.t942 408.469
R1536 VGND.t1276 VGND.t1549 408.469
R1537 VGND.t1616 VGND.t162 408.469
R1538 VGND.t934 VGND.t920 408.469
R1539 VGND.t2573 VGND.t972 408.469
R1540 VGND.t772 VGND.t993 408.469
R1541 VGND.t648 VGND.t2430 408.469
R1542 VGND.t676 VGND.t2563 408.469
R1543 VGND.t2155 VGND.t2290 408.469
R1544 VGND.t2428 VGND.t1528 408.469
R1545 VGND.t2463 VGND.t104 408.469
R1546 VGND.t2539 VGND.t732 408.469
R1547 VGND.t511 VGND.t1414 408.469
R1548 VGND.t1938 VGND.t457 408.469
R1549 VGND.t1475 VGND.t988 408.469
R1550 VGND.t2163 VGND.t1465 408.469
R1551 VGND.t707 VGND.t357 408.469
R1552 VGND.t2633 VGND.t821 408.469
R1553 VGND.t966 VGND.t2247 408.469
R1554 VGND.t297 VGND.t697 408.469
R1555 VGND.t1318 VGND.t2679 408.469
R1556 VGND.t1146 VGND.t932 408.469
R1557 VGND.t790 VGND.t2175 408.469
R1558 VGND.t2592 VGND.t156 408.469
R1559 VGND.t684 VGND.t1386 408.469
R1560 VGND.t1577 VGND.t782 408.469
R1561 VGND.t837 VGND.t2284 408.469
R1562 VGND.t2457 VGND.t1109 408.469
R1563 VGND.t2582 VGND.t668 408.469
R1564 VGND.t2294 VGND.t1968 408.469
R1565 VGND.t469 VGND.t2406 408.469
R1566 VGND.t2451 VGND.t643 408.469
R1567 VGND.t1332 VGND.t9 408.469
R1568 VGND.t1479 VGND.t1165 408.469
R1569 VGND.t1272 VGND.t2150 408.469
R1570 VGND.t1320 VGND.t432 408.469
R1571 VGND.t823 VGND.t501 408.469
R1572 VGND.t970 VGND.t737 408.469
R1573 VGND.t701 VGND.t123 408.469
R1574 VGND.t2477 VGND.t405 408.469
R1575 VGND.t958 VGND.t2037 408.469
R1576 VGND.t172 VGND.t116 408.469
R1577 VGND.t604 VGND.t158 408.469
R1578 VGND.t2535 VGND.t670 408.469
R1579 VGND.t427 VGND.t784 408.469
R1580 VGND.t1430 VGND.t1908 408.469
R1581 VGND.t678 VGND.t2378 408.469
R1582 VGND.t660 VGND.t1130 408.469
R1583 VGND.t1702 VGND.t835 408.469
R1584 VGND.t1301 VGND.t2410 408.469
R1585 VGND.t627 VGND.t453 408.469
R1586 VGND.t286 VGND.t825 408.469
R1587 VGND.t476 VGND.t1481 408.469
R1588 VGND.t4 VGND.t1274 408.469
R1589 VGND.t1403 VGND.t1322 408.469
R1590 VGND.t2598 VGND.t871 408.469
R1591 VGND.t1587 VGND.t715 408.469
R1592 VGND.t1559 VGND.t1312 408.469
R1593 VGND.t844 VGND.t2479 408.469
R1594 VGND.t786 VGND.t2027 408.469
R1595 VGND.t2590 VGND.t174 408.469
R1596 VGND.t1177 VGND.t2483 408.469
R1597 VGND.t713 VGND.t1082 408.469
R1598 VGND.t178 VGND.t1256 408.469
R1599 VGND.t2426 VGND.t1234 408.469
R1600 VGND.t956 VGND.t1077 408.469
R1601 VGND.t2282 VGND.t1066 408.469
R1602 VGND.t2420 VGND.t1047 408.469
R1603 VGND.t926 VGND.t211 408.469
R1604 VGND.t2306 VGND.t190 408.469
R1605 VGND.t1410 VGND.t1043 408.469
R1606 VGND.t2459 VGND.t1222 408.469
R1607 VGND.t2298 VGND.t1209 408.469
R1608 VGND.t1406 VGND.t1101 408.469
R1609 VGND.t1473 VGND.t1026 408.469
R1610 VGND.t443 VGND.t1191 408.469
R1611 VGND.t2095 VGND.t2491 408.469
R1612 VGND.t1825 VGND.t1744 397.848
R1613 VGND.t1744 VGND.t1754 397.848
R1614 VGND.t1754 VGND.t1762 397.848
R1615 VGND.t1762 VGND.t1497 397.848
R1616 VGND.t1497 VGND.t1498 397.848
R1617 VGND.t1498 VGND.t1501 397.848
R1618 VGND.t1501 VGND.t1502 397.848
R1619 VGND.t2362 VGND.t534 396.17
R1620 VGND.t1713 VGND.t1708 396.17
R1621 VGND.n2997 VGND.n33 394.137
R1622 VGND.n2999 VGND.n2998 394.137
R1623 VGND.n2489 VGND.n32 394.137
R1624 VGND.n2428 VGND.n2427 394.137
R1625 VGND.n2426 VGND.n261 394.137
R1626 VGND.n2425 VGND.n262 394.137
R1627 VGND.n2424 VGND.n263 394.137
R1628 VGND.n2423 VGND.n264 394.137
R1629 VGND.n2422 VGND.n265 394.137
R1630 VGND.n2421 VGND.n266 394.137
R1631 VGND.n2420 VGND.n267 394.137
R1632 VGND.n2419 VGND.n268 394.137
R1633 VGND.n2418 VGND.n269 394.137
R1634 VGND.n2417 VGND.n270 394.137
R1635 VGND.n2416 VGND.n271 394.137
R1636 VGND.n2415 VGND.n272 394.137
R1637 VGND.n2414 VGND.n2413 394.137
R1638 VGND.n147 VGND.t242 387.421
R1639 VGND.n1506 VGND.t48 387.421
R1640 VGND.n1508 VGND.t763 387.421
R1641 VGND.n1510 VGND.t52 387.421
R1642 VGND.n2833 VGND.t245 387.421
R1643 VGND.t1714 VGND.t655 362.452
R1644 VGND.t655 VGND.t2186 345.594
R1645 VGND VGND.t50 328.616
R1646 VGND VGND.t247 328.616
R1647 VGND.t883 VGND 328.616
R1648 VGND.t92 VGND 328.616
R1649 VGND VGND.t237 328.616
R1650 VGND.t2105 VGND.t1213 318.947
R1651 VGND.t2099 VGND.t1040 318.947
R1652 VGND.t1025 VGND.t1032 318.947
R1653 VGND.t1010 VGND.t1189 318.947
R1654 VGND.t2093 VGND.t1201 318.947
R1655 VGND.t1092 VGND.t1013 318.947
R1656 VGND.t1204 VGND.t1079 318.947
R1657 VGND.t1195 VGND.t1179 318.947
R1658 VGND.t1081 VGND.t1173 318.947
R1659 VGND.t1094 VGND.t1014 318.947
R1660 VGND.t1176 VGND.t1254 318.947
R1661 VGND.t1245 VGND.t213 318.947
R1662 VGND.t1068 VGND.t1075 318.947
R1663 VGND.t1063 VGND.t1247 318.947
R1664 VGND.t1226 VGND.t1041 318.947
R1665 VGND.t209 VGND.t1065 318.947
R1666 VGND.t2371 VGND.t2362 311.877
R1667 VGND.t1708 VGND.t148 311.877
R1668 VGND VGND.t2367 303.449
R1669 VGND VGND.t2371 295.019
R1670 VGND.n70 VGND.t1753 287.832
R1671 VGND VGND.t530 286.591
R1672 VGND.n964 VGND.t2657 282.327
R1673 VGND.n62 VGND.t1785 282.327
R1674 VGND.n969 VGND.t319 281.13
R1675 VGND.n73 VGND.t1824 281.13
R1676 VGND.n126 VGND.t320 280.978
R1677 VGND.n126 VGND.t1688 280.978
R1678 VGND.n594 VGND.t2387 280.978
R1679 VGND.n594 VGND.t2651 280.978
R1680 VGND.n974 VGND.t47 280.978
R1681 VGND.n156 VGND.t2397 280.978
R1682 VGND.n156 VGND.t2654 280.978
R1683 VGND.n96 VGND.t1769 280.978
R1684 VGND.n96 VGND.t1810 280.978
R1685 VGND.n2855 VGND.t1796 280.978
R1686 VGND.n2855 VGND.t1832 280.978
R1687 VGND.n2887 VGND.t1820 280.978
R1688 VGND.n2887 VGND.t1836 280.978
R1689 VGND.t2435 VGND 278.161
R1690 VGND.n2993 VGND 271.014
R1691 VGND.n3019 VGND.n4 259.389
R1692 VGND.n2835 VGND.n4 259.389
R1693 VGND.n3020 VGND.n3 252.988
R1694 VGND VGND.t2364 252.875
R1695 VGND VGND.t2369 252.875
R1696 VGND.t1764 VGND 252.875
R1697 VGND VGND.t1760 252.875
R1698 VGND VGND.t1812 252.875
R1699 VGND.n676 VGND.t2484 241.393
R1700 VGND.n2574 VGND.t1894 241.393
R1701 VGND.n229 VGND.t1488 241.393
R1702 VGND.n239 VGND.t2419 241.393
R1703 VGND.n179 VGND.t704 241.393
R1704 VGND.n1419 VGND.t1325 241.393
R1705 VGND.n637 VGND.t828 241.393
R1706 VGND.n616 VGND.t1478 241.393
R1707 VGND.n643 VGND.t2409 241.393
R1708 VGND.n659 VGND.t169 241.393
R1709 VGND.n668 VGND.t2490 241.393
R1710 VGND.n1371 VGND.t818 241.393
R1711 VGND.n1303 VGND.t2417 241.393
R1712 VGND.n572 VGND.t816 241.393
R1713 VGND.n568 VGND.t458 241.393
R1714 VGND.n671 VGND.t2295 241.393
R1715 VGND.n825 VGND.t1431 241.393
R1716 VGND.n815 VGND.t1897 241.393
R1717 VGND.n1287 VGND.t714 241.284
R1718 VGND.n683 VGND.t179 241.284
R1719 VGND.n723 VGND.t2427 241.284
R1720 VGND.n728 VGND.t957 241.284
R1721 VGND.n733 VGND.t2283 241.284
R1722 VGND.n738 VGND.t2421 241.284
R1723 VGND.n743 VGND.t927 241.284
R1724 VGND.n748 VGND.t2307 241.284
R1725 VGND.n753 VGND.t1411 241.284
R1726 VGND.n758 VGND.t2460 241.284
R1727 VGND.n763 VGND.t2299 241.284
R1728 VGND.n768 VGND.t1407 241.284
R1729 VGND.n773 VGND.t1474 241.284
R1730 VGND.n778 VGND.t444 241.284
R1731 VGND.n1230 VGND.t1933 241.284
R1732 VGND.n1225 VGND.t1891 241.284
R1733 VGND.n794 VGND.t1975 241.284
R1734 VGND.n1206 VGND.t1966 241.284
R1735 VGND.n1198 VGND.t1927 241.284
R1736 VGND.n1193 VGND.t1879 241.284
R1737 VGND.n802 VGND.t1963 241.284
R1738 VGND.n1174 VGND.t1924 241.284
R1739 VGND.n1166 VGND.t1915 241.284
R1740 VGND.n1161 VGND.t1873 241.284
R1741 VGND.n810 VGND.t1951 241.284
R1742 VGND.n1142 VGND.t1945 241.284
R1743 VGND.n1134 VGND.t1870 241.284
R1744 VGND.n1129 VGND.t1852 241.284
R1745 VGND.n1124 VGND.t1846 241.284
R1746 VGND.n2576 VGND.t1843 241.284
R1747 VGND.n2572 VGND.t1849 241.284
R1748 VGND.n2702 VGND.t1855 241.284
R1749 VGND.n2627 VGND.t1942 241.284
R1750 VGND.n2694 VGND.t1948 241.284
R1751 VGND.n2631 VGND.t1861 241.284
R1752 VGND.n2686 VGND.t1903 241.284
R1753 VGND.n2635 VGND.t1918 241.284
R1754 VGND.n2678 VGND.t1954 241.284
R1755 VGND.n2639 VGND.t1876 241.284
R1756 VGND.n2670 VGND.t1921 241.284
R1757 VGND.n2643 VGND.t1960 241.284
R1758 VGND.n2662 VGND.t1972 241.284
R1759 VGND.n2647 VGND.t1888 241.284
R1760 VGND.n2654 VGND.t1930 241.284
R1761 VGND.n232 VGND.t2317 241.284
R1762 VGND.n2717 VGND.t2552 241.284
R1763 VGND.n2722 VGND.t814 241.284
R1764 VGND.n2727 VGND.t2448 241.284
R1765 VGND.n2732 VGND.t1329 241.284
R1766 VGND.n2737 VGND.t874 241.284
R1767 VGND.n2742 VGND.t1464 241.284
R1768 VGND.n2747 VGND.t706 241.284
R1769 VGND.n2752 VGND.t2482 241.284
R1770 VGND.n2757 VGND.t965 241.284
R1771 VGND.n2762 VGND.t177 241.284
R1772 VGND.n2767 VGND.t2474 241.284
R1773 VGND.n2772 VGND.t931 241.284
R1774 VGND.n2777 VGND.t2281 241.284
R1775 VGND.n227 VGND.t1457 241.284
R1776 VGND.n242 VGND.t775 241.284
R1777 VGND.n2511 VGND.t1429 241.284
R1778 VGND.n2506 VGND.t1472 241.284
R1779 VGND.n246 VGND.t2319 241.284
R1780 VGND.n2436 VGND.t834 241.284
R1781 VGND.n2441 VGND.t1468 241.284
R1782 VGND.n2446 VGND.t2450 241.284
R1783 VGND.n2451 VGND.t1331 241.284
R1784 VGND.n2456 VGND.t812 241.284
R1785 VGND.n2461 VGND.t1271 241.284
R1786 VGND.n2466 VGND.t1317 241.284
R1787 VGND.n2471 VGND.t866 241.284
R1788 VGND.n2476 VGND.t969 241.284
R1789 VGND.n2481 VGND.t155 241.284
R1790 VGND.n2486 VGND.t2476 241.284
R1791 VGND.n2829 VGND.t858 241.284
R1792 VGND.n366 VGND.t961 241.284
R1793 VGND.n370 VGND.t2289 241.284
R1794 VGND.n2169 VGND.t2466 241.284
R1795 VGND.n364 VGND.t673 241.284
R1796 VGND.n2195 VGND.t2277 241.284
R1797 VGND.n356 VGND.t1449 241.284
R1798 VGND.n2221 VGND.t2462 241.284
R1799 VGND.n348 VGND.t2305 241.284
R1800 VGND.n2247 VGND.t1409 241.284
R1801 VGND.n340 VGND.t2456 241.284
R1802 VGND.n2278 VGND.t2297 241.284
R1803 VGND.n2283 VGND.t2494 241.284
R1804 VGND.n2288 VGND.t1279 241.284
R1805 VGND.n332 VGND.t460 241.284
R1806 VGND.n1426 VGND.t1289 241.284
R1807 VGND.n1423 VGND.t718 241.284
R1808 VGND.n2156 VGND.t161 241.284
R1809 VGND.n379 VGND.t860 241.284
R1810 VGND.n2182 VGND.t789 241.284
R1811 VGND.n360 VGND.t1451 241.284
R1812 VGND.n2208 VGND.t2468 241.284
R1813 VGND.n352 VGND.t675 241.284
R1814 VGND.n2234 VGND.t2279 241.284
R1815 VGND.n344 VGND.t2423 241.284
R1816 VGND.n2260 VGND.t667 241.284
R1817 VGND.n336 VGND.t2271 241.284
R1818 VGND.n2265 VGND.t1413 241.284
R1819 VGND.n2305 VGND.t462 241.284
R1820 VGND.n2310 VGND.t2301 241.284
R1821 VGND.n1440 VGND.t2442 241.284
R1822 VGND.n634 VGND.t448 241.284
R1823 VGND.n1490 VGND.t2486 241.284
R1824 VGND.n1485 VGND.t1291 241.284
R1825 VGND.n1480 VGND.t700 241.284
R1826 VGND.n1475 VGND.t2470 241.284
R1827 VGND.n1470 VGND.t862 241.284
R1828 VGND.n1465 VGND.t793 241.284
R1829 VGND.n1460 VGND.t1453 241.284
R1830 VGND.n1455 VGND.t929 241.284
R1831 VGND.n1450 VGND.t781 241.284
R1832 VGND.n1445 VGND.t1447 241.284
R1833 VGND.n393 VGND.t2425 241.284
R1834 VGND.n2133 VGND.t2303 241.284
R1835 VGND.n2128 VGND.t2275 241.284
R1836 VGND.n1502 VGND.t2309 241.284
R1837 VGND.n621 VGND.t2542 241.284
R1838 VGND.n625 VGND.t868 241.284
R1839 VGND.n1995 VGND.t466 241.284
R1840 VGND.n431 VGND.t1309 241.284
R1841 VGND.n2021 VGND.t854 241.284
R1842 VGND.n423 VGND.t1285 241.284
R1843 VGND.n2047 VGND.t171 241.284
R1844 VGND.n415 VGND.t949 241.284
R1845 VGND.n2073 VGND.t953 241.284
R1846 VGND.n407 VGND.t165 241.284
R1847 VGND.n2104 VGND.t945 241.284
R1848 VGND.n2109 VGND.t683 241.284
R1849 VGND.n2114 VGND.t2269 241.284
R1850 VGND.n2119 VGND.t1441 241.284
R1851 VGND.n650 VGND.t2287 241.284
R1852 VGND.n647 VGND.t1417 241.284
R1853 VGND.n1982 VGND.t1295 241.284
R1854 VGND.n435 VGND.t2311 241.284
R1855 VGND.n2008 VGND.t820 241.284
R1856 VGND.n427 VGND.t1287 241.284
R1857 VGND.n2034 VGND.t2440 241.284
R1858 VGND.n419 VGND.t1315 241.284
R1859 VGND.n2060 VGND.t856 241.284
R1860 VGND.n411 VGND.t712 241.284
R1861 VGND.n2086 VGND.t2488 241.284
R1862 VGND.n403 VGND.t852 241.284
R1863 VGND.n2091 VGND.t955 241.284
R1864 VGND.n2330 VGND.t1443 241.284
R1865 VGND.n2335 VGND.t947 241.284
R1866 VGND.n957 VGND.t975 241.284
R1867 VGND.n952 VGND.t795 241.284
R1868 VGND.n947 VGND.t2273 241.284
R1869 VGND.n942 VGND.t937 241.284
R1870 VGND.n937 VGND.t663 241.284
R1871 VGND.n932 VGND.t1423 241.284
R1872 VGND.n927 VGND.t1435 241.284
R1873 VGND.n922 VGND.t2454 241.284
R1874 VGND.n917 VGND.t2550 241.284
R1875 VGND.n912 VGND.t1484 241.284
R1876 VGND.n907 VGND.t2444 241.284
R1877 VGND.n902 VGND.t2544 241.284
R1878 VGND.n449 VGND.t832 241.284
R1879 VGND.n1959 VGND.t720 241.284
R1880 VGND.n1954 VGND.t450 241.284
R1881 VGND.n1393 VGND.t1281 241.284
R1882 VGND.n1398 VGND.t710 241.284
R1883 VGND.n666 VGND.t1445 241.284
R1884 VGND.n1821 VGND.t977 241.284
R1885 VGND.n487 VGND.t777 241.284
R1886 VGND.n1847 VGND.t1437 241.284
R1887 VGND.n479 VGND.t939 241.284
R1888 VGND.n1873 VGND.t665 241.284
R1889 VGND.n471 VGND.t1427 241.284
R1890 VGND.n1899 VGND.t2413 241.284
R1891 VGND.n463 VGND.t2315 241.284
R1892 VGND.n1930 VGND.t1419 241.284
R1893 VGND.n1935 VGND.t1486 241.284
R1894 VGND.n1940 VGND.t452 241.284
R1895 VGND.n1945 VGND.t2546 241.284
R1896 VGND.n1378 VGND.t464 241.284
R1897 VGND.n1375 VGND.t446 241.284
R1898 VGND.n1808 VGND.t951 241.284
R1899 VGND.n491 VGND.t1283 241.284
R1900 VGND.n1834 VGND.t167 241.284
R1901 VGND.n483 VGND.t941 241.284
R1902 VGND.n1860 VGND.t850 241.284
R1903 VGND.n475 VGND.t779 241.284
R1904 VGND.n1886 VGND.t1439 241.284
R1905 VGND.n467 VGND.t681 241.284
R1906 VGND.n1912 VGND.t771 241.284
R1907 VGND.n459 VGND.t1433 241.284
R1908 VGND.n1917 VGND.t2415 241.284
R1909 VGND.n2355 VGND.t2548 241.284
R1910 VGND.n2360 VGND.t1421 241.284
R1911 VGND.n1310 VGND.t2293 241.284
R1912 VGND.n1307 VGND.t1425 241.284
R1913 VGND.n1360 VGND.t1470 241.284
R1914 VGND.n1355 VGND.t2313 241.284
R1915 VGND.n1350 VGND.t830 241.284
R1916 VGND.n1345 VGND.t1293 241.284
R1917 VGND.n1340 VGND.t2446 241.284
R1918 VGND.n1335 VGND.t1327 241.284
R1919 VGND.n1330 VGND.t870 241.284
R1920 VGND.n1325 VGND.t722 241.284
R1921 VGND.n1320 VGND.t1311 241.284
R1922 VGND.n1315 VGND.t864 241.284
R1923 VGND.n505 VGND.t963 241.284
R1924 VGND.n1785 VGND.t1455 241.284
R1925 VGND.n1780 VGND.t2472 241.284
R1926 VGND.n1515 VGND.t456 241.284
R1927 VGND.n1520 VGND.t442 241.284
R1928 VGND.n577 VGND.t943 241.284
R1929 VGND.n1647 VGND.t1277 241.284
R1930 VGND.n543 VGND.t163 241.284
R1931 VGND.n1673 VGND.t935 241.284
R1932 VGND.n535 VGND.t973 241.284
R1933 VGND.n1699 VGND.t773 241.284
R1934 VGND.n527 VGND.t2431 241.284
R1935 VGND.n1725 VGND.t677 241.284
R1936 VGND.n519 VGND.t2291 241.284
R1937 VGND.n1756 VGND.t2429 241.284
R1938 VGND.n1761 VGND.t2464 241.284
R1939 VGND.n1766 VGND.t2540 241.284
R1940 VGND.n1771 VGND.t1415 241.284
R1941 VGND.n1535 VGND.t1476 241.284
R1942 VGND.n566 VGND.t1466 241.284
R1943 VGND.n1634 VGND.t708 241.284
R1944 VGND.n547 VGND.t822 241.284
R1945 VGND.n1660 VGND.t967 241.284
R1946 VGND.n539 VGND.t698 241.284
R1947 VGND.n1686 VGND.t1319 241.284
R1948 VGND.n531 VGND.t933 241.284
R1949 VGND.n1712 VGND.t791 241.284
R1950 VGND.n523 VGND.t157 241.284
R1951 VGND.n1738 VGND.t685 241.284
R1952 VGND.n515 VGND.t783 241.284
R1953 VGND.n1743 VGND.t2285 241.284
R1954 VGND.n2380 VGND.t2458 241.284
R1955 VGND.n2385 VGND.t669 241.284
R1956 VGND.n674 VGND.t2407 241.284
R1957 VGND.n1548 VGND.t2452 241.284
R1958 VGND.n1553 VGND.t1333 241.284
R1959 VGND.n1558 VGND.t1480 241.284
R1960 VGND.n1563 VGND.t1273 241.284
R1961 VGND.n1568 VGND.t1321 241.284
R1962 VGND.n1573 VGND.t824 241.284
R1963 VGND.n1578 VGND.t971 241.284
R1964 VGND.n1583 VGND.t702 241.284
R1965 VGND.n1588 VGND.t2478 241.284
R1966 VGND.n1593 VGND.t959 241.284
R1967 VGND.n1598 VGND.t173 241.284
R1968 VGND.n561 VGND.t159 241.284
R1969 VGND.n1611 VGND.t671 241.284
R1970 VGND.n1606 VGND.t785 241.284
R1971 VGND.n833 VGND.t679 241.284
R1972 VGND.n838 VGND.t661 241.284
R1973 VGND.n830 VGND.t836 241.284
R1974 VGND.n888 VGND.t2411 241.284
R1975 VGND.n883 VGND.t454 241.284
R1976 VGND.n878 VGND.t826 241.284
R1977 VGND.n873 VGND.t1482 241.284
R1978 VGND.n868 VGND.t1275 241.284
R1979 VGND.n863 VGND.t1323 241.284
R1980 VGND.n858 VGND.t872 241.284
R1981 VGND.n853 VGND.t716 241.284
R1982 VGND.n848 VGND.t1313 241.284
R1983 VGND.n843 VGND.t2480 241.284
R1984 VGND.n2400 VGND.t787 241.284
R1985 VGND.n2405 VGND.t175 241.284
R1986 VGND.n719 VGND.t2492 241.284
R1987 VGND.t203 VGND.t1893 222.15
R1988 VGND.t2617 VGND.t1062 222.15
R1989 VGND.t1058 VGND.t1842 222.15
R1990 VGND.t1334 VGND.t1244 222.15
R1991 VGND.t1848 VGND.t1236 222.15
R1992 VGND.t1231 VGND.t1161 222.15
R1993 VGND.t1216 VGND.t1854 222.15
R1994 VGND.t2148 VGND.t2106 222.15
R1995 VGND.t1941 VGND.t196 222.15
R1996 VGND.t1054 VGND.t2070 222.15
R1997 VGND.t1036 VGND.t1947 222.15
R1998 VGND.t236 VGND.t1218 222.15
R1999 VGND.t1860 VGND.t1022 222.15
R2000 VGND.t198 VGND.t1009 222.15
R2001 VGND.t192 VGND.t1902 222.15
R2002 VGND.t657 VGND.t2094 222.15
R2003 VGND.t1917 VGND.t2090 222.15
R2004 VGND.t1024 VGND.t1666 222.15
R2005 VGND.t1038 VGND.t1953 222.15
R2006 VGND.t1583 VGND.t1219 222.15
R2007 VGND.t1875 VGND.t1199 222.15
R2008 VGND.t2092 VGND.t595 222.15
R2009 VGND.t1184 VGND.t1920 222.15
R2010 VGND.t1732 VGND.t1097 222.15
R2011 VGND.t1959 VGND.t1020 222.15
R2012 VGND.t1015 VGND.t1157 222.15
R2013 VGND.t1264 VGND.t1971 222.15
R2014 VGND.t1376 VGND.t1188 222.15
R2015 VGND.t1887 VGND.t1248 222.15
R2016 VGND.t214 VGND.t599 222.15
R2017 VGND.t1929 VGND.t1090 222.15
R2018 VGND.t1012 VGND.t1162 222.15
R2019 VGND.t2231 VGND.t1487 222.15
R2020 VGND.t1689 VGND.t1459 222.15
R2021 VGND.t2316 VGND.t1555 222.15
R2022 VGND.t1126 VGND.t895 222.15
R2023 VGND.t2666 VGND.t2551 222.15
R2024 VGND.t1668 VGND.t1706 222.15
R2025 VGND.t2664 VGND.t813 222.15
R2026 VGND.t1371 VGND.t1541 222.15
R2027 VGND.t2229 VGND.t2447 222.15
R2028 VGND.t1677 VGND.t623 222.15
R2029 VGND.t589 VGND.t1328 222.15
R2030 VGND.t184 VGND.t437 222.15
R2031 VGND.t587 VGND.t873 222.15
R2032 VGND.t403 VGND.t474 222.15
R2033 VGND.t2227 VGND.t1463 222.15
R2034 VGND.t1656 VGND.t2 222.15
R2035 VGND.t2225 VGND.t705 222.15
R2036 VGND.t810 VGND.t1134 222.15
R2037 VGND.t591 VGND.t2481 222.15
R2038 VGND.t2054 VGND.t2597 222.15
R2039 VGND.t2662 VGND.t964 222.15
R2040 VGND.t28 VGND.t2042 222.15
R2041 VGND.t2660 VGND.t176 222.15
R2042 VGND.t1663 VGND.t1662 222.15
R2043 VGND.t585 VGND.t2473 222.15
R2044 VGND.t2353 VGND.t842 222.15
R2045 VGND.t2670 VGND.t930 222.15
R2046 VGND.t0 VGND.t257 222.15
R2047 VGND.t2668 VGND.t2280 222.15
R2048 VGND.t1135 VGND.t379 222.15
R2049 VGND.t1456 VGND.t2223 222.15
R2050 VGND.t1098 VGND.t2320 222.15
R2051 VGND.t2123 VGND.t2418 222.15
R2052 VGND.t2606 VGND.t986 222.15
R2053 VGND.t774 VGND.t1733 222.15
R2054 VGND.t640 VGND.t1008 222.15
R2055 VGND.t1428 VGND.t231 222.15
R2056 VGND.t55 VGND.t2360 222.15
R2057 VGND.t229 VGND.t1471 222.15
R2058 VGND.t2180 VGND.t1164 222.15
R2059 VGND.t2121 VGND.t2318 222.15
R2060 VGND.t440 VGND.t1615 222.15
R2061 VGND.t2239 VGND.t833 222.15
R2062 VGND.t2034 VGND.t285 222.15
R2063 VGND.t2237 VGND.t1467 222.15
R2064 VGND.t2043 VGND.t2572 222.15
R2065 VGND.t1739 VGND.t2449 222.15
R2066 VGND.t1510 VGND.t992 222.15
R2067 VGND.t1737 VGND.t1330 222.15
R2068 VGND.t1106 VGND.t647 222.15
R2069 VGND.t2241 VGND.t811 222.15
R2070 VGND.t1124 VGND.t366 222.15
R2071 VGND.t2127 VGND.t1270 222.15
R2072 VGND.t150 VGND.t1586 222.15
R2073 VGND.t2125 VGND.t1316 222.15
R2074 VGND.t2035 VGND.t1534 222.15
R2075 VGND.t2235 VGND.t865 222.15
R2076 VGND.t1363 VGND.t103 222.15
R2077 VGND.t2233 VGND.t968 222.15
R2078 VGND.t2631 VGND.t891 222.15
R2079 VGND.t233 VGND.t154 222.15
R2080 VGND.t2144 VGND.t426 222.15
R2081 VGND.t1735 VGND.t2475 222.15
R2082 VGND.t723 VGND.t1203 222.15
R2083 VGND.t703 VGND.t2258 222.15
R2084 VGND.t2375 VGND.t2400 222.15
R2085 VGND.t1628 VGND.t857 222.15
R2086 VGND.t2354 VGND.t1132 222.15
R2087 VGND.t1636 VGND.t960 222.15
R2088 VGND.t115 VGND.t360 222.15
R2089 VGND.t2288 VGND.t1634 222.15
R2090 VGND.t1547 VGND.t1370 222.15
R2091 VGND.t2256 VGND.t2465 222.15
R2092 VGND.t2045 VGND.t629 222.15
R2093 VGND.t672 VGND.t1624 222.15
R2094 VGND.t439 VGND.t1113 222.15
R2095 VGND.t1622 VGND.t2276 222.15
R2096 VGND.t1505 VGND.t480 222.15
R2097 VGND.t1448 VGND.t2254 222.15
R2098 VGND.t799 VGND.t659 222.15
R2099 VGND.t2252 VGND.t2461 222.15
R2100 VGND.t900 VGND.t1138 222.15
R2101 VGND.t2304 VGND.t1626 222.15
R2102 VGND.t389 VGND.t336 222.15
R2103 VGND.t1632 VGND.t1408 222.15
R2104 VGND.t1980 VGND.t1297 222.15
R2105 VGND.t2455 VGND.t1630 222.15
R2106 VGND.t1538 VGND.t1710 222.15
R2107 VGND.t1620 VGND.t2296 222.15
R2108 VGND.t251 VGND.t848 222.15
R2109 VGND.t2262 VGND.t2493 222.15
R2110 VGND.t152 VGND.t416 222.15
R2111 VGND.t2260 VGND.t1278 222.15
R2112 VGND.t2162 VGND.t385 222.15
R2113 VGND.t459 VGND.t2250 222.15
R2114 VGND.t2104 VGND.t29 222.15
R2115 VGND.t2203 VGND.t1324 222.15
R2116 VGND.t1353 VGND.t632 222.15
R2117 VGND.t2195 VGND.t1288 222.15
R2118 VGND.t276 VGND.t2088 222.15
R2119 VGND.t717 VGND.t575 222.15
R2120 VGND.t11 VGND.t566 222.15
R2121 VGND.t2209 VGND.t160 222.15
R2122 VGND.t1716 VGND.t2639 222.15
R2123 VGND.t859 VGND.t1383 222.15
R2124 VGND.t2245 VGND.t183 222.15
R2125 VGND.t2191 VGND.t788 222.15
R2126 VGND.t1712 VGND.t330 222.15
R2127 VGND.t1450 VGND.t2189 222.15
R2128 VGND.t2677 VGND.t888 222.15
R2129 VGND.t1381 VGND.t2467 222.15
R2130 VGND.t2642 VGND.t1395 222.15
R2131 VGND.t674 VGND.t1379 222.15
R2132 VGND.t1401 VGND.t2605 222.15
R2133 VGND.t2193 VGND.t2278 222.15
R2134 VGND.t2146 VGND.t413 222.15
R2135 VGND.t2422 VGND.t2207 222.15
R2136 VGND.t303 VGND.t2359 222.15
R2137 VGND.t2205 VGND.t666 222.15
R2138 VGND.t1385 VGND.t1575 222.15
R2139 VGND.t2270 VGND.t581 222.15
R2140 VGND.t610 VGND.t1489 222.15
R2141 VGND.t1412 VGND.t579 222.15
R2142 VGND.t2184 VGND.t1696 222.15
R2143 VGND.t577 VGND.t461 222.15
R2144 VGND.t22 VGND.t2588 222.15
R2145 VGND.t2300 VGND.t1377 222.15
R2146 VGND.t1053 VGND.t1123 222.15
R2147 VGND.t1646 VGND.t827 222.15
R2148 VGND.t2055 VGND.t980 222.15
R2149 VGND.t2140 VGND.t2441 222.15
R2150 VGND.t797 VGND.t634 222.15
R2151 VGND.t447 VGND.t1557 222.15
R2152 VGND.t2347 VGND.t2044 222.15
R2153 VGND.t2485 VGND.t1652 222.15
R2154 VGND.t2198 VGND.t1655 222.15
R2155 VGND.t1290 VGND.t1644 222.15
R2156 VGND.t2135 VGND.t2068 222.15
R2157 VGND.t699 VGND.t2136 222.15
R2158 VGND.t419 VGND.t2358 222.15
R2159 VGND.t2469 VGND.t2013 222.15
R2160 VGND.t2566 VGND.t404 222.15
R2161 VGND.t861 VGND.t1642 222.15
R2162 VGND.t724 VGND.t120 222.15
R2163 VGND.t792 VGND.t1640 222.15
R2164 VGND.t2047 VGND.t1006 222.15
R2165 VGND.t1452 VGND.t2138 222.15
R2166 VGND.t2561 VGND.t2632 222.15
R2167 VGND.t928 VGND.t1650 222.15
R2168 VGND.t1391 VGND.t2133 222.15
R2169 VGND.t780 VGND.t1648 222.15
R2170 VGND.t2024 VGND.t1669 222.15
R2171 VGND.t1446 VGND.t2011 222.15
R2172 VGND.t2333 VGND.t1654 222.15
R2173 VGND.t2424 VGND.t2009 222.15
R2174 VGND.t730 VGND.t911 222.15
R2175 VGND.t2302 VGND.t2007 222.15
R2176 VGND.t518 VGND.t987 222.15
R2177 VGND.t2274 VGND.t2142 222.15
R2178 VGND.t1175 VGND.t2649 222.15
R2179 VGND.t1477 VGND.t1600 222.15
R2180 VGND.t1458 VGND.t8 222.15
R2181 VGND.t69 VGND.t2308 222.15
R2182 VGND.t2438 VGND.t1125 222.15
R2183 VGND.t1608 VGND.t2541 222.15
R2184 VGND.t2685 VGND.t359 222.15
R2185 VGND.t867 VGND.t1606 222.15
R2186 VGND.t1540 VGND.t220 222.15
R2187 VGND.t1598 VGND.t465 222.15
R2188 VGND.t539 VGND.t622 222.15
R2189 VGND.t1308 VGND.t1725 222.15
R2190 VGND.t436 VGND.t1367 222.15
R2191 VGND.t1723 VGND.t853 222.15
R2192 VGND.t2355 VGND.t473 222.15
R2193 VGND.t1284 VGND.t1596 222.15
R2194 VGND.t1 VGND.t2351 222.15
R2195 VGND.t73 VGND.t170 222.15
R2196 VGND.t141 VGND.t1133 222.15
R2197 VGND.t948 VGND.t1727 222.15
R2198 VGND.t2596 VGND.t572 222.15
R2199 VGND.t1604 VGND.t952 222.15
R2200 VGND.t1507 VGND.t2041 222.15
R2201 VGND.t164 VGND.t1602 222.15
R2202 VGND.t1661 VGND.t2402 222.15
R2203 VGND.t1721 VGND.t944 222.15
R2204 VGND.t658 VGND.t841 222.15
R2205 VGND.t1719 VGND.t682 222.15
R2206 VGND.t1005 VGND.t256 222.15
R2207 VGND.t1717 VGND.t2268 222.15
R2208 VGND.t1741 VGND.t378 222.15
R2209 VGND.t1440 VGND.t71 222.15
R2210 VGND.t1096 VGND.t265 222.15
R2211 VGND.t1996 VGND.t2408 222.15
R2212 VGND.t1160 VGND.t2380 222.15
R2213 VGND.t1523 VGND.t2286 222.15
R2214 VGND.t397 VGND.t64 222.15
R2215 VGND.t1416 VGND.t2004 222.15
R2216 VGND.t1707 VGND.t979 222.15
R2217 VGND.t2002 VGND.t1294 222.15
R2218 VGND.t2036 VGND.t1548 222.15
R2219 VGND.t2310 VGND.t1994 222.15
R2220 VGND.t2340 VGND.t153 222.15
R2221 VGND.t1519 VGND.t819 222.15
R2222 VGND.t255 VGND.t296 222.15
R2223 VGND.t1286 VGND.t1517 222.15
R2224 VGND.t481 VGND.t30 222.15
R2225 VGND.t1992 VGND.t2439 222.15
R2226 VGND.t252 VGND.t800 222.15
R2227 VGND.t1314 VGND.t1990 222.15
R2228 VGND.t1139 VGND.t1664 222.15
R2229 VGND.t1521 VGND.t855 222.15
R2230 VGND.t1509 VGND.t390 222.15
R2231 VGND.t711 VGND.t2000 222.15
R2232 VGND.t1298 VGND.t2432 222.15
R2233 VGND.t1998 VGND.t2487 222.15
R2234 VGND.t1582 VGND.t1539 222.15
R2235 VGND.t851 VGND.t1515 222.15
R2236 VGND.t2327 VGND.t806 222.15
R2237 VGND.t954 VGND.t353 222.15
R2238 VGND.t417 VGND.t796 222.15
R2239 VGND.t351 VGND.t1442 222.15
R2240 VGND.t1674 VGND.t510 222.15
R2241 VGND.t946 VGND.t1525 222.15
R2242 VGND.t2107 VGND.t1356 222.15
R2243 VGND.t168 VGND.t618 222.15
R2244 VGND.t633 VGND.t538 222.15
R2245 VGND.t974 VGND.t1120 222.15
R2246 VGND.t2089 VGND.t1155 222.15
R2247 VGND.t794 VGND.t221 222.15
R2248 VGND.t14 VGND.t88 222.15
R2249 VGND.t2272 VGND.t2081 222.15
R2250 VGND.t2640 VGND.t235 222.15
R2251 VGND.t936 VGND.t616 222.15
R2252 VGND.t2246 VGND.t598 222.15
R2253 VGND.t662 VGND.t1116 222.15
R2254 VGND.t331 VGND.t1144 222.15
R2255 VGND.t1422 VGND.t1114 222.15
R2256 VGND.t2678 VGND.t1584 222.15
R2257 VGND.t1434 VGND.t614 222.15
R2258 VGND.t1145 VGND.t760 222.15
R2259 VGND.t2453 VGND.t612 222.15
R2260 VGND.t2174 VGND.t1105 222.15
R2261 VGND.t2549 VGND.t1118 222.15
R2262 VGND.t414 VGND.t2185 222.15
R2263 VGND.t1483 VGND.t2079 222.15
R2264 VGND.t304 VGND.t597 222.15
R2265 VGND.t2443 VGND.t2077 222.15
R2266 VGND.t1576 VGND.t396 222.15
R2267 VGND.t2543 VGND.t227 222.15
R2268 VGND.t611 VGND.t1352 222.15
R2269 VGND.t831 VGND.t225 222.15
R2270 VGND.t1108 VGND.t1004 222.15
R2271 VGND.t719 VGND.t223 222.15
R2272 VGND.t2589 VGND.t127 222.15
R2273 VGND.t449 VGND.t807 222.15
R2274 VGND.t1055 VGND.t25 222.15
R2275 VGND.t343 VGND.t2489 222.15
R2276 VGND.t2630 VGND.t630 222.15
R2277 VGND.t497 VGND.t1280 222.15
R2278 VGND.t1639 VGND.t2087 222.15
R2279 VGND.t1266 VGND.t709 222.15
R2280 VGND.t1512 VGND.t13 222.15
R2281 VGND.t1444 VGND.t349 222.15
R2282 VGND.t2638 VGND.t537 222.15
R2283 VGND.t341 VGND.t976 222.15
R2284 VGND.t2641 VGND.t2243 222.15
R2285 VGND.t776 VGND.t493 222.15
R2286 VGND.t328 VGND.t1372 222.15
R2287 VGND.t491 VGND.t1436 222.15
R2288 VGND.t1678 VGND.t2676 222.15
R2289 VGND.t938 VGND.t339 222.15
R2290 VGND.t1394 VGND.t185 222.15
R2291 VGND.t337 VGND.t664 222.15
R2292 VGND.t1697 VGND.t1400 222.15
R2293 VGND.t1426 VGND.t495 222.15
R2294 VGND.t412 VGND.t1122 222.15
R2295 VGND.t347 VGND.t2412 222.15
R2296 VGND.t620 VGND.t302 222.15
R2297 VGND.t2314 VGND.t345 222.15
R2298 VGND.t1574 VGND.t1679 222.15
R2299 VGND.t489 VGND.t1418 222.15
R2300 VGND.t87 VGND.t609 222.15
R2301 VGND.t487 VGND.t1485 222.15
R2302 VGND.t1398 VGND.t2183 222.15
R2303 VGND.t1268 VGND.t451 222.15
R2304 VGND.t327 VGND.t2586 222.15
R2305 VGND.t2545 VGND.t2338 222.15
R2306 VGND.t1046 VGND.t1369 222.15
R2307 VGND.t1338 VGND.t817 222.15
R2308 VGND.t2437 VGND.t1514 222.15
R2309 VGND.t557 VGND.t463 222.15
R2310 VGND.t2643 VGND.t2687 222.15
R2311 VGND.t445 VGND.t1346 222.15
R2312 VGND.t2350 VGND.t1506 222.15
R2313 VGND.t1344 VGND.t950 222.15
R2314 VGND.t1357 VGND.t2197 222.15
R2315 VGND.t1282 VGND.t1336 222.15
R2316 VGND.t2134 VGND.t594 222.15
R2317 VGND.t553 VGND.t166 222.15
R2318 VGND.t250 VGND.t418 222.15
R2319 VGND.t940 VGND.t551 222.15
R2320 VGND.t2565 VGND.t1007 222.15
R2321 VGND.t563 VGND.t849 222.15
R2322 VGND.t129 VGND.t798 222.15
R2323 VGND.t778 VGND.t561 222.15
R2324 VGND.t2046 VGND.t1581 222.15
R2325 VGND.t555 VGND.t1438 222.15
R2326 VGND.t2075 VGND.t393 222.15
R2327 VGND.t680 VGND.t1342 222.15
R2328 VGND.t1390 VGND.t1711 222.15
R2329 VGND.t1340 VGND.t770 222.15
R2330 VGND.t601 VGND.t2021 222.15
R2331 VGND.t1432 VGND.t549 222.15
R2332 VGND.t2332 VGND.t2267 222.15
R2333 VGND.t2414 VGND.t547 222.15
R2334 VGND.t144 VGND.t1154 222.15
R2335 VGND.t545 VGND.t2547 222.15
R2336 VGND.t1729 VGND.t517 222.15
R2337 VGND.t1420 VGND.t559 222.15
R2338 VGND.t1170 VGND.t2006 222.15
R2339 VGND.t2517 VGND.t2416 222.15
R2340 VGND.t1490 VGND.t468 222.15
R2341 VGND.t2501 VGND.t2292 222.15
R2342 VGND.t1152 VGND.t642 222.15
R2343 VGND.t1424 VGND.t2525 222.15
R2344 VGND.t1986 VGND.t147 222.15
R2345 VGND.t1469 VGND.t2523 222.15
R2346 VGND.t584 VGND.t593 222.15
R2347 VGND.t2312 VGND.t90 222.15
R2348 VGND.t2149 VGND.t1461 222.15
R2349 VGND.t829 VGND.t2497 222.15
R2350 VGND.t919 VGND.t2266 222.15
R2351 VGND.t1292 VGND.t2495 222.15
R2352 VGND.t500 VGND.t1730 222.15
R2353 VGND.t2445 VGND.t2507 222.15
R2354 VGND.t736 VGND.t1508 222.15
R2355 VGND.t1326 VGND.t2505 222.15
R2356 VGND.t122 VGND.t1657 222.15
R2357 VGND.t869 VGND.t2499 222.15
R2358 VGND.t410 VGND.t574 222.15
R2359 VGND.t721 VGND.t2521 222.15
R2360 VGND.t2154 VGND.t2644 222.15
R2361 VGND.t1310 VGND.t2519 222.15
R2362 VGND.t2511 VGND.t151 222.15
R2363 VGND.t863 VGND.t2531 222.15
R2364 VGND.t603 VGND.t1979 222.15
R2365 VGND.t962 VGND.t2529 222.15
R2366 VGND.t2074 VGND.t2069 222.15
R2367 VGND.t1454 VGND.t2527 222.15
R2368 VGND.t2581 VGND.t182 222.15
R2369 VGND.t2471 VGND.t2503 222.15
R2370 VGND.t1261 VGND.t1366 222.15
R2371 VGND.t2626 VGND.t815 222.15
R2372 VGND.t621 VGND.t1460 222.15
R2373 VGND.t694 VGND.t455 222.15
R2374 VGND.t887 VGND.t1127 222.15
R2375 VGND.t2613 VGND.t441 222.15
R2376 VGND.t2120 VGND.t361 222.15
R2377 VGND.t942 VGND.t2611 222.15
R2378 VGND.t1546 VGND.t1690 222.15
R2379 VGND.t2624 VGND.t1276 222.15
R2380 VGND.t696 VGND.t624 222.15
R2381 VGND.t162 VGND.t690 222.15
R2382 VGND.t438 VGND.t1667 222.15
R2383 VGND.t688 VGND.t934 222.15
R2384 VGND.t743 VGND.t475 222.15
R2385 VGND.t972 VGND.t2622 222.15
R2386 VGND.t3 VGND.t2265 222.15
R2387 VGND.t2620 VGND.t772 222.15
R2388 VGND.t1364 VGND.t1402 222.15
R2389 VGND.t2430 VGND.t692 222.15
R2390 VGND.t388 VGND.t1405 222.15
R2391 VGND.t2609 VGND.t676 222.15
R2392 VGND.t119 VGND.t1296 222.15
R2393 VGND.t2290 VGND.t2607 222.15
R2394 VGND.t1567 VGND.t573 222.15
R2395 VGND.t686 VGND.t2428 222.15
R2396 VGND.t2361 VGND.t843 222.15
R2397 VGND.t2403 VGND.t2463 222.15
R2398 VGND.t277 VGND.t2033 222.15
R2399 VGND.t2615 VGND.t2539 222.15
R2400 VGND.t1392 VGND.t384 222.15
R2401 VGND.t1414 VGND.t2618 222.15
R2402 VGND.t2101 VGND.t2399 222.15
R2403 VGND.t457 VGND.t16 222.15
R2404 VGND.t467 VGND.t15 222.15
R2405 VGND.t2215 VGND.t1475 222.15
R2406 VGND.t26 VGND.t641 222.15
R2407 VGND.t1465 VGND.t2110 222.15
R2408 VGND.t1989 VGND.t912 222.15
R2409 VGND.t2108 VGND.t707 222.15
R2410 VGND.t896 VGND.t583 222.15
R2411 VGND.t821 VGND.t2553 222.15
R2412 VGND.t264 VGND.t128 222.15
R2413 VGND.t2211 VGND.t966 222.15
R2414 VGND.t1675 VGND.t918 222.15
R2415 VGND.t697 VGND.t2118 222.15
R2416 VGND.t509 VGND.t253 222.15
R2417 VGND.t2221 VGND.t1318 222.15
R2418 VGND.t1156 VGND.t317 222.15
R2419 VGND.t932 VGND.t2219 222.15
R2420 VGND.t121 VGND.t2188 222.15
R2421 VGND.t2213 VGND.t790 222.15
R2422 VGND.t1462 VGND.t407 222.15
R2423 VGND.t156 VGND.t20 222.15
R2424 VGND.t2326 VGND.t2684 222.15
R2425 VGND.t18 VGND.t684 222.15
R2426 VGND.t741 VGND.t118 222.15
R2427 VGND.t782 VGND.t2116 222.15
R2428 VGND.t602 VGND.t1107 222.15
R2429 VGND.t2284 VGND.t2114 222.15
R2430 VGND.t2071 VGND.t1665 222.15
R2431 VGND.t2112 VGND.t2457 222.15
R2432 VGND.t540 VGND.t2580 222.15
R2433 VGND.t668 VGND.t2217 222.15
R2434 VGND.t1258 VGND.t894 222.15
R2435 VGND.t2064 VGND.t2294 222.15
R2436 VGND.t2321 VGND.t985 222.15
R2437 VGND.t2406 VGND.t85 222.15
R2438 VGND.t639 VGND.t2161 222.15
R2439 VGND.t2015 VGND.t2451 222.15
R2440 VGND.t181 VGND.t62 222.15
R2441 VGND.t1572 VGND.t1332 222.15
R2442 VGND.t254 VGND.t1163 222.15
R2443 VGND.t2062 VGND.t1479 222.15
R2444 VGND.t27 VGND.t1614 222.15
R2445 VGND.t81 VGND.t1272 222.15
R2446 VGND.t1354 VGND.t420 222.15
R2447 VGND.t79 VGND.t1320 222.15
R2448 VGND.t2686 VGND.t2571 222.15
R2449 VGND.t2060 VGND.t823 222.15
R2450 VGND.t2053 VGND.t729 222.15
R2451 VGND.t2058 VGND.t970 222.15
R2452 VGND.t23 VGND.t2052 222.15
R2453 VGND.t83 VGND.t701 222.15
R2454 VGND.t499 VGND.t2562 222.15
R2455 VGND.t1570 VGND.t2477 222.15
R2456 VGND.t742 VGND.t1585 222.15
R2457 VGND.t2066 VGND.t958 222.15
R2458 VGND.t1396 VGND.t1527 222.15
R2459 VGND.t77 VGND.t172 222.15
R2460 VGND.t1680 VGND.t102 222.15
R2461 VGND.t158 VGND.t75 222.15
R2462 VGND.t731 VGND.t571 222.15
R2463 VGND.t670 VGND.t2017 222.15
R2464 VGND.t425 VGND.t521 222.15
R2465 VGND.t784 VGND.t2056 222.15
R2466 VGND.t1190 VGND.t1368 222.15
R2467 VGND.t268 VGND.t1430 222.15
R2468 VGND.t759 VGND.t631 222.15
R2469 VGND.t567 VGND.t678 222.15
R2470 VGND.t757 VGND.t2086 222.15
R2471 VGND.t907 VGND.t660 222.15
R2472 VGND.t2264 VGND.t12 222.15
R2473 VGND.t835 VGND.t905 222.15
R2474 VGND.t2637 VGND.t2147 222.15
R2475 VGND.t2410 VGND.t266 222.15
R2476 VGND.t2244 VGND.t2179 222.15
R2477 VGND.t453 VGND.t136 222.15
R2478 VGND.t329 VGND.t761 222.15
R2479 VGND.t825 VGND.t134 222.15
R2480 VGND.t2675 VGND.t2405 222.15
R2481 VGND.t1481 VGND.t1693 222.15
R2482 VGND.t1393 VGND.t1513 222.15
R2483 VGND.t1274 VGND.t1691 222.15
R2484 VGND.t1399 VGND.t275 222.15
R2485 VGND.t1322 VGND.t138 222.15
R2486 VGND.t411 VGND.t596 222.15
R2487 VGND.t871 VGND.t272 222.15
R2488 VGND.t301 VGND.t1731 222.15
R2489 VGND.t715 VGND.t270 222.15
R2490 VGND.t2025 VGND.t809 222.15
R2491 VGND.t1312 VGND.t132 222.15
R2492 VGND.t608 VGND.t758 222.15
R2493 VGND.t2479 VGND.t130 222.15
R2494 VGND.t2182 VGND.t565 222.15
R2495 VGND.t909 VGND.t786 222.15
R2496 VGND.t1003 VGND.t2587 222.15
R2497 VGND.t174 VGND.t569 222.15
R2498 VGND.t1045 VGND.t769 222.15
R2499 VGND.t2483 VGND.t1084 222.15
R2500 VGND.t284 VGND.t180 222.15
R2501 VGND.t1259 VGND.t713 222.15
R2502 VGND.t1335 VGND.t2173 222.15
R2503 VGND.t1180 VGND.t178 222.15
R2504 VGND.t1358 VGND.t1985 222.15
R2505 VGND.t207 VGND.t2426 222.15
R2506 VGND.t219 VGND.t1167 222.15
R2507 VGND.t1073 VGND.t956 222.15
R2508 VGND.t249 VGND.t2085 222.15
R2509 VGND.t1240 VGND.t2282 222.15
R2510 VGND.t899 VGND.t294 222.15
R2511 VGND.t1229 VGND.t2420 222.15
R2512 VGND.t89 VGND.t2579 222.15
R2513 VGND.t1069 VGND.t926 222.15
R2514 VGND.t893 VGND.t999 222.15
R2515 VGND.t1051 VGND.t2306 222.15
R2516 VGND.t2604 VGND.t654 222.15
R2517 VGND.t1242 VGND.t1410 222.15
R2518 VGND.t2401 VGND.t367 222.15
R2519 VGND.t194 VGND.t2459 222.15
R2520 VGND.t1397 VGND.t1595 222.15
R2521 VGND.t2102 VGND.t2298 222.15
R2522 VGND.t1307 VGND.t2512 222.15
R2523 VGND.t1224 VGND.t1406 222.15
R2524 VGND.t1355 VGND.t110 222.15
R2525 VGND.t1211 VGND.t1473 222.15
R2526 VGND.t63 VGND.t892 222.15
R2527 VGND.t1186 VGND.t443 222.15
R2528 VGND.t1158 VGND.t429 222.15
R2529 VGND.t2491 VGND.t1030 222.15
R2530 VGND.t1215 VGND.t140 222.15
R2531 VGND.n2834 VGND.n3 218.73
R2532 VGND.n133 VGND.n131 214.365
R2533 VGND.n133 VGND.n132 214.365
R2534 VGND.n123 VGND.n121 214.365
R2535 VGND.n123 VGND.n122 214.365
R2536 VGND.n141 VGND.n139 214.365
R2537 VGND.n141 VGND.n140 214.365
R2538 VGND.n601 VGND.n599 214.365
R2539 VGND.n601 VGND.n600 214.365
R2540 VGND.n591 VGND.n589 214.365
R2541 VGND.n591 VGND.n590 214.365
R2542 VGND.n609 VGND.n607 214.365
R2543 VGND.n609 VGND.n608 214.365
R2544 VGND.n971 VGND.n970 214.365
R2545 VGND.n163 VGND.n161 214.365
R2546 VGND.n163 VGND.n162 214.365
R2547 VGND.n153 VGND.n151 214.365
R2548 VGND.n153 VGND.n152 214.365
R2549 VGND.n171 VGND.n169 214.365
R2550 VGND.n171 VGND.n170 214.365
R2551 VGND.n1096 VGND.n1095 213.613
R2552 VGND.n1098 VGND.n1097 213.613
R2553 VGND.n1068 VGND.n1066 213.613
R2554 VGND.n1068 VGND.n1067 213.613
R2555 VGND.n1071 VGND.n1069 213.613
R2556 VGND.n1071 VGND.n1070 213.613
R2557 VGND.n1006 VGND.n1004 213.613
R2558 VGND.n1006 VGND.n1005 213.613
R2559 VGND.n1009 VGND.n1007 213.613
R2560 VGND.n1009 VGND.n1008 213.613
R2561 VGND.n1037 VGND.n1035 213.613
R2562 VGND.n1037 VGND.n1036 213.613
R2563 VGND.n1040 VGND.n1038 213.613
R2564 VGND.n1040 VGND.n1039 213.613
R2565 VGND.n1110 VGND.t522 212.422
R2566 VGND.n968 VGND.n967 207.965
R2567 VGND.n985 VGND.n965 207.965
R2568 VGND.n98 VGND.n94 207.965
R2569 VGND.n98 VGND.n95 207.965
R2570 VGND.n92 VGND.n90 207.965
R2571 VGND.n92 VGND.n91 207.965
R2572 VGND.n105 VGND.n88 207.965
R2573 VGND.n105 VGND.n89 207.965
R2574 VGND.n2857 VGND.n2853 207.965
R2575 VGND.n2857 VGND.n2854 207.965
R2576 VGND.n2851 VGND.n2849 207.965
R2577 VGND.n2851 VGND.n2850 207.965
R2578 VGND.n2864 VGND.n2847 207.965
R2579 VGND.n2864 VGND.n2848 207.965
R2580 VGND.n2889 VGND.n2885 207.965
R2581 VGND.n2889 VGND.n2886 207.965
R2582 VGND.n2883 VGND.n2881 207.965
R2583 VGND.n2883 VGND.n2882 207.965
R2584 VGND.n2896 VGND.n2879 207.965
R2585 VGND.n2896 VGND.n2880 207.965
R2586 VGND.n67 VGND.n66 207.965
R2587 VGND.n79 VGND.n64 207.965
R2588 VGND.n71 VGND.n69 207.965
R2589 VGND.n984 VGND.n966 207.213
R2590 VGND.n14 VGND.n13 207.213
R2591 VGND.n18 VGND.n12 207.213
R2592 VGND.n43 VGND.n41 207.213
R2593 VGND.n43 VGND.n42 207.213
R2594 VGND.n47 VGND.n39 207.213
R2595 VGND.n47 VGND.n40 207.213
R2596 VGND.n78 VGND.n65 207.213
R2597 VGND.n2931 VGND.n2929 207.213
R2598 VGND.n2931 VGND.n2930 207.213
R2599 VGND.n2935 VGND.n2926 207.213
R2600 VGND.n2935 VGND.n2927 207.213
R2601 VGND.n2971 VGND.n2969 207.213
R2602 VGND.n2971 VGND.n2970 207.213
R2603 VGND.n2975 VGND.n2967 207.213
R2604 VGND.n2975 VGND.n2968 207.213
R2605 VGND.t1896 VGND.t1028 206.59
R2606 VGND.t1207 VGND.t1845 206.59
R2607 VGND.t1851 VGND.t2097 206.59
R2608 VGND.t1088 VGND.t1869 206.59
R2609 VGND.t1944 VGND.t1205 206.59
R2610 VGND.t1193 VGND.t1950 206.59
R2611 VGND.t1872 VGND.t1171 206.59
R2612 VGND.t1016 VGND.t1914 206.59
R2613 VGND.t1923 VGND.t1252 206.59
R2614 VGND.t215 VGND.t1962 206.59
R2615 VGND.t1878 VGND.t1071 206.59
R2616 VGND.t1060 VGND.t1926 206.59
R2617 VGND.t1965 VGND.t1227 206.59
R2618 VGND.t205 VGND.t1974 206.59
R2619 VGND.t1890 VGND.t1049 206.59
R2620 VGND.t1238 VGND.t1932 206.59
R2621 VGND VGND.n2652 194.419
R2622 VGND VGND.n2648 194.419
R2623 VGND VGND.n2660 194.419
R2624 VGND VGND.n2644 194.419
R2625 VGND VGND.n2668 194.419
R2626 VGND VGND.n2640 194.419
R2627 VGND VGND.n2676 194.419
R2628 VGND VGND.n2636 194.419
R2629 VGND VGND.n2684 194.419
R2630 VGND VGND.n2632 194.419
R2631 VGND VGND.n2692 194.419
R2632 VGND VGND.n2628 194.419
R2633 VGND VGND.n2700 194.419
R2634 VGND VGND.n2579 194.419
R2635 VGND VGND.n2570 194.419
R2636 VGND.n676 VGND.n675 194.391
R2637 VGND.n1286 VGND.n678 194.391
R2638 VGND.n684 VGND.n682 194.391
R2639 VGND.n722 VGND.n721 194.391
R2640 VGND.n727 VGND.n726 194.391
R2641 VGND.n732 VGND.n731 194.391
R2642 VGND.n737 VGND.n736 194.391
R2643 VGND.n742 VGND.n741 194.391
R2644 VGND.n747 VGND.n746 194.391
R2645 VGND.n752 VGND.n751 194.391
R2646 VGND.n757 VGND.n756 194.391
R2647 VGND.n762 VGND.n761 194.391
R2648 VGND.n767 VGND.n766 194.391
R2649 VGND.n772 VGND.n771 194.391
R2650 VGND.n777 VGND.n776 194.391
R2651 VGND.n1231 VGND.n787 194.391
R2652 VGND.n1224 VGND.n1223 194.391
R2653 VGND.n793 VGND.n792 194.391
R2654 VGND.n1205 VGND.n1204 194.391
R2655 VGND.n1199 VGND.n795 194.391
R2656 VGND.n1192 VGND.n1191 194.391
R2657 VGND.n801 VGND.n800 194.391
R2658 VGND.n1173 VGND.n1172 194.391
R2659 VGND.n1167 VGND.n803 194.391
R2660 VGND.n1160 VGND.n1159 194.391
R2661 VGND.n809 VGND.n808 194.391
R2662 VGND.n1141 VGND.n1140 194.391
R2663 VGND.n1135 VGND.n811 194.391
R2664 VGND.n1128 VGND.n1127 194.391
R2665 VGND.n1125 VGND.n813 194.391
R2666 VGND.n2574 VGND.n2573 194.391
R2667 VGND.n229 VGND.n228 194.391
R2668 VGND.n231 VGND.n230 194.391
R2669 VGND.n2716 VGND.n2715 194.391
R2670 VGND.n2721 VGND.n2720 194.391
R2671 VGND.n2726 VGND.n2725 194.391
R2672 VGND.n2731 VGND.n2730 194.391
R2673 VGND.n2736 VGND.n2735 194.391
R2674 VGND.n2741 VGND.n2740 194.391
R2675 VGND.n2746 VGND.n2745 194.391
R2676 VGND.n2751 VGND.n2750 194.391
R2677 VGND.n2756 VGND.n2755 194.391
R2678 VGND.n2761 VGND.n2760 194.391
R2679 VGND.n2766 VGND.n2765 194.391
R2680 VGND.n2771 VGND.n2770 194.391
R2681 VGND.n2776 VGND.n2775 194.391
R2682 VGND.n226 VGND.n225 194.391
R2683 VGND.n239 VGND.n238 194.391
R2684 VGND.n241 VGND.n240 194.391
R2685 VGND.n2510 VGND.n2509 194.391
R2686 VGND.n2505 VGND.n243 194.391
R2687 VGND.n247 VGND.n245 194.391
R2688 VGND.n2435 VGND.n2434 194.391
R2689 VGND.n2440 VGND.n2439 194.391
R2690 VGND.n2445 VGND.n2444 194.391
R2691 VGND.n2450 VGND.n2449 194.391
R2692 VGND.n2455 VGND.n2454 194.391
R2693 VGND.n2460 VGND.n2459 194.391
R2694 VGND.n2465 VGND.n2464 194.391
R2695 VGND.n2470 VGND.n2469 194.391
R2696 VGND.n2475 VGND.n2474 194.391
R2697 VGND.n2480 VGND.n2479 194.391
R2698 VGND.n2485 VGND.n2484 194.391
R2699 VGND.n179 VGND.n178 194.391
R2700 VGND.n2828 VGND.n181 194.391
R2701 VGND.n367 VGND.n365 194.391
R2702 VGND.n369 VGND.n368 194.391
R2703 VGND.n2168 VGND.n2167 194.391
R2704 VGND.n363 VGND.n362 194.391
R2705 VGND.n2194 VGND.n2193 194.391
R2706 VGND.n355 VGND.n354 194.391
R2707 VGND.n2220 VGND.n2219 194.391
R2708 VGND.n347 VGND.n346 194.391
R2709 VGND.n2246 VGND.n2245 194.391
R2710 VGND.n339 VGND.n338 194.391
R2711 VGND.n2277 VGND.n2276 194.391
R2712 VGND.n2282 VGND.n2281 194.391
R2713 VGND.n2287 VGND.n2286 194.391
R2714 VGND.n331 VGND.n330 194.391
R2715 VGND.n1419 VGND.n1418 194.391
R2716 VGND.n1425 VGND.n1424 194.391
R2717 VGND.n1422 VGND.n1421 194.391
R2718 VGND.n2155 VGND.n2154 194.391
R2719 VGND.n378 VGND.n377 194.391
R2720 VGND.n2181 VGND.n2180 194.391
R2721 VGND.n359 VGND.n358 194.391
R2722 VGND.n2207 VGND.n2206 194.391
R2723 VGND.n351 VGND.n350 194.391
R2724 VGND.n2233 VGND.n2232 194.391
R2725 VGND.n343 VGND.n342 194.391
R2726 VGND.n2259 VGND.n2258 194.391
R2727 VGND.n335 VGND.n334 194.391
R2728 VGND.n2264 VGND.n2263 194.391
R2729 VGND.n2304 VGND.n2303 194.391
R2730 VGND.n2311 VGND.n326 194.391
R2731 VGND.n637 VGND.n636 194.391
R2732 VGND.n1439 VGND.n1438 194.391
R2733 VGND.n633 VGND.n632 194.391
R2734 VGND.n1489 VGND.n1488 194.391
R2735 VGND.n1484 VGND.n1483 194.391
R2736 VGND.n1479 VGND.n1478 194.391
R2737 VGND.n1474 VGND.n1473 194.391
R2738 VGND.n1469 VGND.n1468 194.391
R2739 VGND.n1464 VGND.n1463 194.391
R2740 VGND.n1459 VGND.n1458 194.391
R2741 VGND.n1454 VGND.n1453 194.391
R2742 VGND.n1449 VGND.n1448 194.391
R2743 VGND.n1444 VGND.n1443 194.391
R2744 VGND.n392 VGND.n391 194.391
R2745 VGND.n2132 VGND.n2131 194.391
R2746 VGND.n2127 VGND.n394 194.391
R2747 VGND.n616 VGND.n615 194.391
R2748 VGND.n1501 VGND.n618 194.391
R2749 VGND.n622 VGND.n620 194.391
R2750 VGND.n624 VGND.n623 194.391
R2751 VGND.n1994 VGND.n1993 194.391
R2752 VGND.n430 VGND.n429 194.391
R2753 VGND.n2020 VGND.n2019 194.391
R2754 VGND.n422 VGND.n421 194.391
R2755 VGND.n2046 VGND.n2045 194.391
R2756 VGND.n414 VGND.n413 194.391
R2757 VGND.n2072 VGND.n2071 194.391
R2758 VGND.n406 VGND.n405 194.391
R2759 VGND.n2103 VGND.n2102 194.391
R2760 VGND.n2108 VGND.n2107 194.391
R2761 VGND.n2113 VGND.n2112 194.391
R2762 VGND.n2120 VGND.n397 194.391
R2763 VGND.n643 VGND.n642 194.391
R2764 VGND.n649 VGND.n648 194.391
R2765 VGND.n646 VGND.n645 194.391
R2766 VGND.n1981 VGND.n1980 194.391
R2767 VGND.n434 VGND.n433 194.391
R2768 VGND.n2007 VGND.n2006 194.391
R2769 VGND.n426 VGND.n425 194.391
R2770 VGND.n2033 VGND.n2032 194.391
R2771 VGND.n418 VGND.n417 194.391
R2772 VGND.n2059 VGND.n2058 194.391
R2773 VGND.n410 VGND.n409 194.391
R2774 VGND.n2085 VGND.n2084 194.391
R2775 VGND.n402 VGND.n401 194.391
R2776 VGND.n2090 VGND.n2089 194.391
R2777 VGND.n2329 VGND.n2328 194.391
R2778 VGND.n2336 VGND.n315 194.391
R2779 VGND.n659 VGND.n658 194.391
R2780 VGND.n956 VGND.n955 194.391
R2781 VGND.n951 VGND.n950 194.391
R2782 VGND.n946 VGND.n945 194.391
R2783 VGND.n941 VGND.n940 194.391
R2784 VGND.n936 VGND.n935 194.391
R2785 VGND.n931 VGND.n930 194.391
R2786 VGND.n926 VGND.n925 194.391
R2787 VGND.n921 VGND.n920 194.391
R2788 VGND.n916 VGND.n915 194.391
R2789 VGND.n911 VGND.n910 194.391
R2790 VGND.n906 VGND.n905 194.391
R2791 VGND.n901 VGND.n900 194.391
R2792 VGND.n448 VGND.n447 194.391
R2793 VGND.n1958 VGND.n1957 194.391
R2794 VGND.n1953 VGND.n450 194.391
R2795 VGND.n668 VGND.n667 194.391
R2796 VGND.n1392 VGND.n1391 194.391
R2797 VGND.n1397 VGND.n1396 194.391
R2798 VGND.n665 VGND.n664 194.391
R2799 VGND.n1820 VGND.n1819 194.391
R2800 VGND.n486 VGND.n485 194.391
R2801 VGND.n1846 VGND.n1845 194.391
R2802 VGND.n478 VGND.n477 194.391
R2803 VGND.n1872 VGND.n1871 194.391
R2804 VGND.n470 VGND.n469 194.391
R2805 VGND.n1898 VGND.n1897 194.391
R2806 VGND.n462 VGND.n461 194.391
R2807 VGND.n1929 VGND.n1928 194.391
R2808 VGND.n1934 VGND.n1933 194.391
R2809 VGND.n1939 VGND.n1938 194.391
R2810 VGND.n1946 VGND.n453 194.391
R2811 VGND.n1371 VGND.n1370 194.391
R2812 VGND.n1377 VGND.n1376 194.391
R2813 VGND.n1374 VGND.n1373 194.391
R2814 VGND.n1807 VGND.n1806 194.391
R2815 VGND.n490 VGND.n489 194.391
R2816 VGND.n1833 VGND.n1832 194.391
R2817 VGND.n482 VGND.n481 194.391
R2818 VGND.n1859 VGND.n1858 194.391
R2819 VGND.n474 VGND.n473 194.391
R2820 VGND.n1885 VGND.n1884 194.391
R2821 VGND.n466 VGND.n465 194.391
R2822 VGND.n1911 VGND.n1910 194.391
R2823 VGND.n458 VGND.n457 194.391
R2824 VGND.n1916 VGND.n1915 194.391
R2825 VGND.n2354 VGND.n2353 194.391
R2826 VGND.n2361 VGND.n303 194.391
R2827 VGND.n1303 VGND.n1302 194.391
R2828 VGND.n1309 VGND.n1308 194.391
R2829 VGND.n1306 VGND.n1305 194.391
R2830 VGND.n1359 VGND.n1358 194.391
R2831 VGND.n1354 VGND.n1353 194.391
R2832 VGND.n1349 VGND.n1348 194.391
R2833 VGND.n1344 VGND.n1343 194.391
R2834 VGND.n1339 VGND.n1338 194.391
R2835 VGND.n1334 VGND.n1333 194.391
R2836 VGND.n1329 VGND.n1328 194.391
R2837 VGND.n1324 VGND.n1323 194.391
R2838 VGND.n1319 VGND.n1318 194.391
R2839 VGND.n1314 VGND.n1313 194.391
R2840 VGND.n504 VGND.n503 194.391
R2841 VGND.n1784 VGND.n1783 194.391
R2842 VGND.n1779 VGND.n506 194.391
R2843 VGND.n572 VGND.n571 194.391
R2844 VGND.n1514 VGND.n1513 194.391
R2845 VGND.n1519 VGND.n1518 194.391
R2846 VGND.n576 VGND.n575 194.391
R2847 VGND.n1646 VGND.n1645 194.391
R2848 VGND.n542 VGND.n541 194.391
R2849 VGND.n1672 VGND.n1671 194.391
R2850 VGND.n534 VGND.n533 194.391
R2851 VGND.n1698 VGND.n1697 194.391
R2852 VGND.n526 VGND.n525 194.391
R2853 VGND.n1724 VGND.n1723 194.391
R2854 VGND.n518 VGND.n517 194.391
R2855 VGND.n1755 VGND.n1754 194.391
R2856 VGND.n1760 VGND.n1759 194.391
R2857 VGND.n1765 VGND.n1764 194.391
R2858 VGND.n1772 VGND.n509 194.391
R2859 VGND.n568 VGND.n567 194.391
R2860 VGND.n1534 VGND.n1533 194.391
R2861 VGND.n565 VGND.n564 194.391
R2862 VGND.n1633 VGND.n1632 194.391
R2863 VGND.n546 VGND.n545 194.391
R2864 VGND.n1659 VGND.n1658 194.391
R2865 VGND.n538 VGND.n537 194.391
R2866 VGND.n1685 VGND.n1684 194.391
R2867 VGND.n530 VGND.n529 194.391
R2868 VGND.n1711 VGND.n1710 194.391
R2869 VGND.n522 VGND.n521 194.391
R2870 VGND.n1737 VGND.n1736 194.391
R2871 VGND.n514 VGND.n513 194.391
R2872 VGND.n1742 VGND.n1741 194.391
R2873 VGND.n2379 VGND.n2378 194.391
R2874 VGND.n2386 VGND.n290 194.391
R2875 VGND.n671 VGND.n670 194.391
R2876 VGND.n673 VGND.n672 194.391
R2877 VGND.n1547 VGND.n1546 194.391
R2878 VGND.n1552 VGND.n1551 194.391
R2879 VGND.n1557 VGND.n1556 194.391
R2880 VGND.n1562 VGND.n1561 194.391
R2881 VGND.n1567 VGND.n1566 194.391
R2882 VGND.n1572 VGND.n1571 194.391
R2883 VGND.n1577 VGND.n1576 194.391
R2884 VGND.n1582 VGND.n1581 194.391
R2885 VGND.n1587 VGND.n1586 194.391
R2886 VGND.n1592 VGND.n1591 194.391
R2887 VGND.n1597 VGND.n1596 194.391
R2888 VGND.n560 VGND.n559 194.391
R2889 VGND.n1610 VGND.n1609 194.391
R2890 VGND.n1605 VGND.n1601 194.391
R2891 VGND.n825 VGND.n824 194.391
R2892 VGND.n832 VGND.n831 194.391
R2893 VGND.n837 VGND.n836 194.391
R2894 VGND.n829 VGND.n828 194.391
R2895 VGND.n887 VGND.n886 194.391
R2896 VGND.n882 VGND.n881 194.391
R2897 VGND.n877 VGND.n876 194.391
R2898 VGND.n872 VGND.n871 194.391
R2899 VGND.n867 VGND.n866 194.391
R2900 VGND.n862 VGND.n861 194.391
R2901 VGND.n857 VGND.n856 194.391
R2902 VGND.n852 VGND.n851 194.391
R2903 VGND.n847 VGND.n846 194.391
R2904 VGND.n842 VGND.n841 194.391
R2905 VGND.n2399 VGND.n2398 194.391
R2906 VGND.n2406 VGND.n278 194.391
R2907 VGND.n815 VGND.n814 194.391
R2908 VGND.n718 VGND.n717 194.391
R2909 VGND.n2564 VGND.n2563 161.308
R2910 VGND.n2561 VGND.n2560 161.308
R2911 VGND.n2558 VGND.n2557 161.308
R2912 VGND.n2555 VGND.n2554 161.308
R2913 VGND.n2552 VGND.n2551 161.308
R2914 VGND.n2549 VGND.n2548 161.308
R2915 VGND.n2546 VGND.n2545 161.308
R2916 VGND.n2543 VGND.n2542 161.308
R2917 VGND.n2540 VGND.n2539 161.308
R2918 VGND.n2537 VGND.n2536 161.308
R2919 VGND.n2534 VGND.n2533 161.308
R2920 VGND.n2531 VGND.n2530 161.308
R2921 VGND.n2528 VGND.n2527 161.308
R2922 VGND.n2525 VGND.n2524 161.308
R2923 VGND.n2522 VGND.n2521 161.308
R2924 VGND.n2563 VGND.t2695 159.978
R2925 VGND.n2560 VGND.t2699 159.978
R2926 VGND.n2557 VGND.t2693 159.978
R2927 VGND.n2554 VGND.t2689 159.978
R2928 VGND.n2551 VGND.t2694 159.978
R2929 VGND.n2548 VGND.t2702 159.978
R2930 VGND.n2545 VGND.t2698 159.978
R2931 VGND.n2542 VGND.t2691 159.978
R2932 VGND.n2539 VGND.t2688 159.978
R2933 VGND.n2536 VGND.t2690 159.978
R2934 VGND.n2533 VGND.t2701 159.978
R2935 VGND.n2530 VGND.t2692 159.978
R2936 VGND.n2527 VGND.t2700 159.978
R2937 VGND.n2524 VGND.t2697 159.978
R2938 VGND.n2521 VGND.t2703 159.978
R2939 VGND.n996 VGND.t2436 159.315
R2940 VGND.n2917 VGND.t904 159.315
R2941 VGND.n1088 VGND.t1351 158.361
R2942 VGND.n2987 VGND.t422 158.361
R2943 VGND.n898 VGND.t2434 157.291
R2944 VGND.n2915 VGND.t902 157.291
R2945 VGND.n582 VGND.t248 156.915
R2946 VGND.n2877 VGND.t2365 156.915
R2947 VGND.n582 VGND.t244 156.915
R2948 VGND.n2877 VGND.t2366 156.915
R2949 VGND.n584 VGND.t2357 154.131
R2950 VGND.n584 VGND.t1695 154.131
R2951 VGND.n996 VGND.t1375 154.131
R2952 VGND.n999 VGND.t1658 154.131
R2953 VGND.n2901 VGND.t33 154.131
R2954 VGND.n2901 VGND.t1491 154.131
R2955 VGND.n2917 VGND.t536 154.131
R2956 VGND.n2947 VGND.t1715 154.131
R2957 VGND.n118 VGND.t243 153.631
R2958 VGND.n1026 VGND.t764 153.631
R2959 VGND.n1057 VGND.t2181 153.631
R2960 VGND.n2869 VGND.t2363 153.631
R2961 VGND.n2949 VGND.t656 153.631
R2962 VGND.n2954 VGND.t1709 153.631
R2963 VGND.n1027 VGND.t1373 152.757
R2964 VGND.n2950 VGND.t2187 152.757
R2965 VGND.n991 VGND.t240 152.381
R2966 VGND.n61 VGND.t2370 152.381
R2967 VGND.n961 VGND.n960 152.174
R2968 VGND.n149 VGND.t246 150.922
R2969 VGND.n149 VGND.t238 150.922
R2970 VGND.n86 VGND.t2373 150.922
R2971 VGND.n86 VGND.t2368 150.922
R2972 VGND.n116 VGND.t2249 150.922
R2973 VGND.n581 VGND.t398 150.922
R2974 VGND.n148 VGND.t2648 150.922
R2975 VGND.n85 VGND.t35 150.922
R2976 VGND.n2844 VGND.t1580 150.922
R2977 VGND.n2876 VGND.t1671 150.922
R2978 VGND.n116 VGND.t744 150.922
R2979 VGND.n581 VGND.t541 150.922
R2980 VGND.n148 VGND.t2076 150.922
R2981 VGND.n85 VGND.t187 150.922
R2982 VGND.n2844 VGND.t1151 150.922
R2983 VGND.n2876 VGND.t748 150.922
R2984 VGND.n117 VGND.t241 147.411
R2985 VGND.n1058 VGND.t2352 147.411
R2986 VGND.n2868 VGND.t2372 147.411
R2987 VGND.n2955 VGND.t149 147.411
R2988 VGND.n899 VGND.t531 146.964
R2989 VGND.n84 VGND.t1496 146.964
R2990 VGND.n2563 VGND.t1880 143.911
R2991 VGND.n2560 VGND.t1955 143.911
R2992 VGND.n2557 VGND.t1862 143.911
R2993 VGND.n2554 VGND.t1904 143.911
R2994 VGND.n2551 VGND.t1976 143.911
R2995 VGND.n2548 VGND.t1883 143.911
R2996 VGND.n2545 VGND.t1856 143.911
R2997 VGND.n2542 VGND.t1898 143.911
R2998 VGND.n2539 VGND.t1910 143.911
R2999 VGND.n2536 VGND.t1838 143.911
R3000 VGND.n2533 VGND.t1934 143.911
R3001 VGND.n2530 VGND.t1865 143.911
R3002 VGND.n2527 VGND.t1937 143.911
R3003 VGND.n2524 VGND.t1967 143.911
R3004 VGND.n2521 VGND.t1907 143.911
R3005 VGND.n1512 VGND.n578 143.478
R3006 VGND VGND.t1825 142.089
R3007 VGND.n822 VGND.t1895 119.309
R3008 VGND.n785 VGND.t1931 119.309
R3009 VGND.n2585 VGND.t1928 119.309
R3010 VGND.n2582 VGND.t1892 119.309
R3011 VGND.n2568 VGND.t1841 119.309
R3012 VGND.n2581 VGND.t1847 119.309
R3013 VGND.n2620 VGND.t1853 119.309
R3014 VGND.n2617 VGND.t1940 119.309
R3015 VGND.n2614 VGND.t1946 119.309
R3016 VGND.n2611 VGND.t1859 119.309
R3017 VGND.n2608 VGND.t1901 119.309
R3018 VGND.n2605 VGND.t1916 119.309
R3019 VGND.n2602 VGND.t1952 119.309
R3020 VGND.n2599 VGND.t1874 119.309
R3021 VGND.n2596 VGND.t1919 119.309
R3022 VGND.n2593 VGND.t1958 119.309
R3023 VGND.n2590 VGND.t1970 119.309
R3024 VGND.n2587 VGND.t1886 119.309
R3025 VGND.n819 VGND.t1844 119.309
R3026 VGND.n816 VGND.t1850 119.309
R3027 VGND.n1136 VGND.t1868 119.309
R3028 VGND.n807 VGND.t1943 119.309
R3029 VGND.n805 VGND.t1949 119.309
R3030 VGND.n1151 VGND.t1871 119.309
R3031 VGND.n1168 VGND.t1913 119.309
R3032 VGND.n799 VGND.t1922 119.309
R3033 VGND.n797 VGND.t1961 119.309
R3034 VGND.n1183 VGND.t1877 119.309
R3035 VGND.n1200 VGND.t1925 119.309
R3036 VGND.n791 VGND.t1964 119.309
R3037 VGND.n789 VGND.t1973 119.309
R3038 VGND.n1215 VGND.t1889 119.309
R3039 VGND.n6 VGND.n4 117.001
R3040 VGND.t2537 VGND.n6 117.001
R3041 VGND.n5 VGND.n3 117.001
R3042 VGND.t2537 VGND.n5 117.001
R3043 VGND.t1213 VGND.t1896 112.356
R3044 VGND.t1153 VGND.t2105 112.356
R3045 VGND.t1845 VGND.t2099 112.356
R3046 VGND.t1040 VGND.t600 112.356
R3047 VGND.t1032 VGND.t1851 112.356
R3048 VGND.t805 VGND.t1025 112.356
R3049 VGND.t1869 VGND.t1010 112.356
R3050 VGND.t1189 VGND.t1159 112.356
R3051 VGND.t1201 VGND.t1944 112.356
R3052 VGND.t2145 VGND.t2093 112.356
R3053 VGND.t1950 VGND.t1092 112.356
R3054 VGND.t1013 VGND.t2683 112.356
R3055 VGND.t1079 VGND.t1872 112.356
R3056 VGND.t295 VGND.t1204 112.356
R3057 VGND.t1914 VGND.t1195 112.356
R3058 VGND.t1179 VGND.t1676 112.356
R3059 VGND.t1173 VGND.t1923 112.356
R3060 VGND.t762 VGND.t1081 112.356
R3061 VGND.t1962 VGND.t1094 112.356
R3062 VGND.t1014 VGND.t274 112.356
R3063 VGND.t1254 VGND.t1878 112.356
R3064 VGND.t1511 VGND.t1176 112.356
R3065 VGND.t1926 VGND.t1245 112.356
R3066 VGND.t213 VGND.t2374 112.356
R3067 VGND.t1075 VGND.t1965 112.356
R3068 VGND.t24 VGND.t1068 112.356
R3069 VGND.t1974 VGND.t1063 112.356
R3070 VGND.t1247 VGND.t2356 112.356
R3071 VGND.t1041 VGND.t1890 112.356
R3072 VGND.t1638 VGND.t1226 112.356
R3073 VGND.t1932 VGND.t209 112.356
R3074 VGND.t1065 VGND.t913 112.356
R3075 VGND.t522 VGND.t532 92.9349
R3076 VGND.t532 VGND.t529 92.9349
R3077 VGND.t529 VGND.t533 92.9349
R3078 VGND.t533 VGND.t2658 92.9349
R3079 VGND.t2658 VGND.t2392 92.9349
R3080 VGND.t2392 VGND.t880 92.9349
R3081 VGND.t880 VGND.t2557 92.9349
R3082 VGND VGND.n578 80.9529
R3083 VGND.n1291 VGND 75.2331
R3084 VGND VGND.n578 75.1009
R3085 VGND.t2557 VGND 70.8076
R3086 VGND.n147 VGND 58.8055
R3087 VGND.n1506 VGND 58.8055
R3088 VGND.n1508 VGND 58.8055
R3089 VGND.n1510 VGND 58.8055
R3090 VGND.n2833 VGND 58.8055
R3091 VGND.n2836 VGND.n2835 53.1823
R3092 VGND.n2837 VGND.n2836 53.1823
R3093 VGND.n3019 VGND.n3018 53.1823
R3094 VGND.n3018 VGND.n3017 53.1823
R3095 VGND.t530 VGND.t2656 50.5752
R3096 VGND.t527 VGND.t2390 50.5752
R3097 VGND.t525 VGND.t1682 50.5752
R3098 VGND.t523 VGND.t318 50.5752
R3099 VGND.t1503 VGND.t1823 50.5752
R3100 VGND.t1499 VGND.t1797 50.5752
R3101 VGND.t1493 VGND.t1834 50.5752
R3102 VGND.t1495 VGND.t1784 50.5752
R3103 VGND VGND.n14 43.2063
R3104 VGND VGND.n43 43.2063
R3105 VGND VGND.n2931 43.2063
R3106 VGND VGND.n2971 43.2063
R3107 VGND.n2835 VGND.n2834 40.6593
R3108 VGND.n675 VGND.t1178 34.8005
R3109 VGND.n675 VGND.t1085 34.8005
R3110 VGND.n678 VGND.t1083 34.8005
R3111 VGND.n678 VGND.t1260 34.8005
R3112 VGND.n682 VGND.t1257 34.8005
R3113 VGND.n682 VGND.t1181 34.8005
R3114 VGND.n721 VGND.t1235 34.8005
R3115 VGND.n721 VGND.t208 34.8005
R3116 VGND.n726 VGND.t1078 34.8005
R3117 VGND.n726 VGND.t1074 34.8005
R3118 VGND.n731 VGND.t1067 34.8005
R3119 VGND.n731 VGND.t1241 34.8005
R3120 VGND.n736 VGND.t1048 34.8005
R3121 VGND.n736 VGND.t1230 34.8005
R3122 VGND.n741 VGND.t212 34.8005
R3123 VGND.n741 VGND.t1070 34.8005
R3124 VGND.n746 VGND.t191 34.8005
R3125 VGND.n746 VGND.t1052 34.8005
R3126 VGND.n751 VGND.t1044 34.8005
R3127 VGND.n751 VGND.t1243 34.8005
R3128 VGND.n756 VGND.t1223 34.8005
R3129 VGND.n756 VGND.t195 34.8005
R3130 VGND.n761 VGND.t1210 34.8005
R3131 VGND.n761 VGND.t2103 34.8005
R3132 VGND.n766 VGND.t1102 34.8005
R3133 VGND.n766 VGND.t1225 34.8005
R3134 VGND.n771 VGND.t1027 34.8005
R3135 VGND.n771 VGND.t1212 34.8005
R3136 VGND.n776 VGND.t1192 34.8005
R3137 VGND.n776 VGND.t1187 34.8005
R3138 VGND.n787 VGND.t1239 34.8005
R3139 VGND.n787 VGND.t210 34.8005
R3140 VGND.n1223 VGND.t1050 34.8005
R3141 VGND.n1223 VGND.t1042 34.8005
R3142 VGND.n792 VGND.t206 34.8005
R3143 VGND.n792 VGND.t1064 34.8005
R3144 VGND.n1204 VGND.t1228 34.8005
R3145 VGND.n1204 VGND.t1076 34.8005
R3146 VGND.n795 VGND.t1061 34.8005
R3147 VGND.n795 VGND.t1246 34.8005
R3148 VGND.n1191 VGND.t1072 34.8005
R3149 VGND.n1191 VGND.t1255 34.8005
R3150 VGND.n800 VGND.t216 34.8005
R3151 VGND.n800 VGND.t1095 34.8005
R3152 VGND.n1172 VGND.t1253 34.8005
R3153 VGND.n1172 VGND.t1174 34.8005
R3154 VGND.n803 VGND.t1017 34.8005
R3155 VGND.n803 VGND.t1196 34.8005
R3156 VGND.n1159 VGND.t1172 34.8005
R3157 VGND.n1159 VGND.t1080 34.8005
R3158 VGND.n808 VGND.t1194 34.8005
R3159 VGND.n808 VGND.t1093 34.8005
R3160 VGND.n1140 VGND.t1206 34.8005
R3161 VGND.n1140 VGND.t1202 34.8005
R3162 VGND.n811 VGND.t1089 34.8005
R3163 VGND.n811 VGND.t1011 34.8005
R3164 VGND.n1127 VGND.t2098 34.8005
R3165 VGND.n1127 VGND.t1033 34.8005
R3166 VGND.n813 VGND.t1208 34.8005
R3167 VGND.n813 VGND.t2100 34.8005
R3168 VGND.n2573 VGND.t1233 34.8005
R3169 VGND.n2573 VGND.t204 34.8005
R3170 VGND.n2652 VGND.t1183 34.8005
R3171 VGND.n2652 VGND.t1091 34.8005
R3172 VGND.n2648 VGND.t1251 34.8005
R3173 VGND.n2648 VGND.t1249 34.8005
R3174 VGND.n2660 VGND.t1087 34.8005
R3175 VGND.n2660 VGND.t1265 34.8005
R3176 VGND.n2644 VGND.t218 34.8005
R3177 VGND.n2644 VGND.t1021 34.8005
R3178 VGND.n2668 VGND.t1263 34.8005
R3179 VGND.n2668 VGND.t1185 34.8005
R3180 VGND.n2640 VGND.t1019 34.8005
R3181 VGND.n2640 VGND.t1200 34.8005
R3182 VGND.n2676 VGND.t1100 34.8005
R3183 VGND.n2676 VGND.t1039 34.8005
R3184 VGND.n2636 VGND.t1198 34.8005
R3185 VGND.n2636 VGND.t2091 34.8005
R3186 VGND.n2684 VGND.t1221 34.8005
R3187 VGND.n2684 VGND.t193 34.8005
R3188 VGND.n2632 VGND.t1104 34.8005
R3189 VGND.n2632 VGND.t1023 34.8005
R3190 VGND.n2692 VGND.t189 34.8005
R3191 VGND.n2692 VGND.t1037 34.8005
R3192 VGND.n2628 VGND.t200 34.8005
R3193 VGND.n2628 VGND.t197 34.8005
R3194 VGND.n2700 VGND.t1035 34.8005
R3195 VGND.n2700 VGND.t1217 34.8005
R3196 VGND.n2579 VGND.t1057 34.8005
R3197 VGND.n2579 VGND.t1237 34.8005
R3198 VGND.n2570 VGND.t202 34.8005
R3199 VGND.n2570 VGND.t1059 34.8005
R3200 VGND.n228 VGND.t1882 34.8005
R3201 VGND.n228 VGND.t2232 34.8005
R3202 VGND.n230 VGND.t984 34.8005
R3203 VGND.n230 VGND.t1556 34.8005
R3204 VGND.n2715 VGND.t638 34.8005
R3205 VGND.n2715 VGND.t2667 34.8005
R3206 VGND.n2720 VGND.t2349 34.8005
R3207 VGND.n2720 VGND.t2665 34.8005
R3208 VGND.n2725 VGND.t1545 34.8005
R3209 VGND.n2725 VGND.t2230 34.8005
R3210 VGND.n2730 VGND.t1613 34.8005
R3211 VGND.n2730 VGND.t590 34.8005
R3212 VGND.n2735 VGND.t312 34.8005
R3213 VGND.n2735 VGND.t588 34.8005
R3214 VGND.n2740 VGND.t2570 34.8005
R3215 VGND.n2740 VGND.t2228 34.8005
R3216 VGND.n2745 VGND.t728 34.8005
R3217 VGND.n2745 VGND.t2226 34.8005
R3218 VGND.n2750 VGND.t2051 34.8005
R3219 VGND.n2750 VGND.t592 34.8005
R3220 VGND.n2755 VGND.t395 34.8005
R3221 VGND.n2755 VGND.t2663 34.8005
R3222 VGND.n2760 VGND.t2325 34.8005
R3223 VGND.n2760 VGND.t2661 34.8005
R3224 VGND.n2765 VGND.t2023 34.8005
R3225 VGND.n2765 VGND.t586 34.8005
R3226 VGND.n2770 VGND.t101 34.8005
R3227 VGND.n2770 VGND.t2671 34.8005
R3228 VGND.n2775 VGND.t146 34.8005
R3229 VGND.n2775 VGND.t2669 34.8005
R3230 VGND.n225 VGND.t383 34.8005
R3231 VGND.n225 VGND.t2224 34.8005
R3232 VGND.n238 VGND.t1957 34.8005
R3233 VGND.n238 VGND.t2124 34.8005
R3234 VGND.n240 VGND.t472 34.8005
R3235 VGND.n240 VGND.t1734 34.8005
R3236 VGND.n2509 VGND.t646 34.8005
R3237 VGND.n2509 VGND.t232 34.8005
R3238 VGND.n243 VGND.t1988 34.8005
R3239 VGND.n243 VGND.t230 34.8005
R3240 VGND.n245 VGND.t1169 34.8005
R3241 VGND.n245 VGND.t2122 34.8005
R3242 VGND.n2434 VGND.t2153 34.8005
R3243 VGND.n2434 VGND.t2240 34.8005
R3244 VGND.n2439 VGND.t435 34.8005
R3245 VGND.n2439 VGND.t2238 34.8005
R3246 VGND.n2444 VGND.t2674 34.8005
R3247 VGND.n2444 VGND.t1740 34.8005
R3248 VGND.n2449 VGND.t740 34.8005
R3249 VGND.n2449 VGND.t1738 34.8005
R3250 VGND.n2454 VGND.t126 34.8005
R3251 VGND.n2454 VGND.t2242 34.8005
R3252 VGND.n2459 VGND.t409 34.8005
R3253 VGND.n2459 VGND.t2128 34.8005
R3254 VGND.n2464 VGND.t2040 34.8005
R3255 VGND.n2464 VGND.t2126 34.8005
R3256 VGND.n2469 VGND.t2510 34.8005
R3257 VGND.n2469 VGND.t2236 34.8005
R3258 VGND.n2474 VGND.t607 34.8005
R3259 VGND.n2474 VGND.t2234 34.8005
R3260 VGND.n2479 VGND.t2073 34.8005
R3261 VGND.n2479 VGND.t234 34.8005
R3262 VGND.n2484 VGND.t431 34.8005
R3263 VGND.n2484 VGND.t1736 34.8005
R3264 VGND.n178 VGND.t1864 34.8005
R3265 VGND.n178 VGND.t2259 34.8005
R3266 VGND.n181 VGND.t281 34.8005
R3267 VGND.n181 VGND.t1629 34.8005
R3268 VGND.n365 VGND.t2170 34.8005
R3269 VGND.n365 VGND.t1637 34.8005
R3270 VGND.n368 VGND.t59 34.8005
R3271 VGND.n368 VGND.t1635 34.8005
R3272 VGND.n2167 VGND.t1552 34.8005
R3273 VGND.n2167 VGND.t2257 34.8005
R3274 VGND.n362 VGND.t1619 34.8005
R3275 VGND.n362 VGND.t1625 34.8005
R3276 VGND.n2193 VGND.t923 34.8005
R3277 VGND.n2193 VGND.t1623 34.8005
R3278 VGND.n354 VGND.t2576 34.8005
R3279 VGND.n354 VGND.t2255 34.8005
R3280 VGND.n2219 VGND.t996 34.8005
R3281 VGND.n2219 VGND.t2253 34.8005
R3282 VGND.n346 VGND.t651 34.8005
R3283 VGND.n346 VGND.t1627 34.8005
R3284 VGND.n2245 VGND.t363 34.8005
R3285 VGND.n2245 VGND.t1633 34.8005
R3286 VGND.n338 VGND.t2158 34.8005
R3287 VGND.n338 VGND.t1631 34.8005
R3288 VGND.n2276 VGND.t1531 34.8005
R3289 VGND.n2276 VGND.t1621 34.8005
R3290 VGND.n2281 VGND.t107 34.8005
R3291 VGND.n2281 VGND.t2263 34.8005
R3292 VGND.n2286 VGND.t735 34.8005
R3293 VGND.n2286 VGND.t2261 34.8005
R3294 VGND.n330 VGND.t514 34.8005
R3295 VGND.n330 VGND.t2251 34.8005
R3296 VGND.n1418 VGND.t1906 34.8005
R3297 VGND.n1418 VGND.t2204 34.8005
R3298 VGND.n1424 VGND.t2382 34.8005
R3299 VGND.n1424 VGND.t2196 34.8005
R3300 VGND.n1421 VGND.t66 34.8005
R3301 VGND.n1421 VGND.t576 34.8005
R3302 VGND.n2154 VGND.t1701 34.8005
R3303 VGND.n2154 VGND.t2210 34.8005
R3304 VGND.n377 VGND.t1304 34.8005
R3305 VGND.n377 VGND.t1384 34.8005
R3306 VGND.n2180 VGND.t2342 34.8005
R3307 VGND.n2180 VGND.t2192 34.8005
R3308 VGND.n358 VGND.t291 34.8005
R3309 VGND.n358 VGND.t2190 34.8005
R3310 VGND.n2206 VGND.t483 34.8005
R3311 VGND.n2206 VGND.t1382 34.8005
R3312 VGND.n350 VGND.t802 34.8005
R3313 VGND.n350 VGND.t1380 34.8005
R3314 VGND.n2232 VGND.t1141 34.8005
R3315 VGND.n2232 VGND.t2194 34.8005
R3316 VGND.n342 VGND.t2603 34.8005
R3317 VGND.n342 VGND.t2208 34.8005
R3318 VGND.n2258 VGND.t1592 34.8005
R3319 VGND.n2258 VGND.t2206 34.8005
R3320 VGND.n334 VGND.t1564 34.8005
R3321 VGND.n334 VGND.t582 34.8005
R3322 VGND.n2263 VGND.t2329 34.8005
R3323 VGND.n2263 VGND.t580 34.8005
R3324 VGND.n2303 VGND.t2030 34.8005
R3325 VGND.n2303 VGND.t578 34.8005
R3326 VGND.n326 VGND.t375 34.8005
R3327 VGND.n326 VGND.t1378 34.8005
R3328 VGND.n636 VGND.t1978 34.8005
R3329 VGND.n636 VGND.t1647 34.8005
R3330 VGND.n1438 VGND.t768 34.8005
R3331 VGND.n1438 VGND.t2141 34.8005
R3332 VGND.n632 VGND.t1362 34.8005
R3333 VGND.n632 VGND.t1558 34.8005
R3334 VGND.n1488 VGND.t1982 34.8005
R3335 VGND.n1488 VGND.t1653 34.8005
R3336 VGND.n1483 VGND.t2202 34.8005
R3337 VGND.n1483 VGND.t1645 34.8005
R3338 VGND.n1478 VGND.t263 34.8005
R3339 VGND.n1478 VGND.t2137 34.8005
R3340 VGND.n1473 VGND.t335 34.8005
R3341 VGND.n1473 VGND.t2014 34.8005
R3342 VGND.n1468 VGND.t508 34.8005
R3343 VGND.n1468 VGND.t1643 34.8005
R3344 VGND.n1463 VGND.t316 34.8005
R3345 VGND.n1463 VGND.t1641 34.8005
R3346 VGND.n1458 VGND.t917 34.8005
R3347 VGND.n1458 VGND.t2139 34.8005
R3348 VGND.n1453 VGND.t371 34.8005
R3349 VGND.n1453 VGND.t1651 34.8005
R3350 VGND.n1448 VGND.t308 34.8005
R3351 VGND.n1448 VGND.t1649 34.8005
R3352 VGND.n1443 VGND.t2516 34.8005
R3353 VGND.n1443 VGND.t2012 34.8005
R3354 VGND.n391 VGND.t114 34.8005
R3355 VGND.n391 VGND.t2010 34.8005
R3356 VGND.n2131 VGND.t2534 34.8005
R3357 VGND.n2131 VGND.t2008 34.8005
R3358 VGND.n394 VGND.t424 34.8005
R3359 VGND.n394 VGND.t2143 34.8005
R3360 VGND.n615 VGND.t1885 34.8005
R3361 VGND.n615 VGND.t1601 34.8005
R3362 VGND.n618 VGND.t982 34.8005
R3363 VGND.n618 VGND.t70 34.8005
R3364 VGND.n620 VGND.t636 34.8005
R3365 VGND.n620 VGND.t1609 34.8005
R3366 VGND.n623 VGND.t2346 34.8005
R3367 VGND.n623 VGND.t1607 34.8005
R3368 VGND.n1993 VGND.t1543 34.8005
R3369 VGND.n1993 VGND.t1599 34.8005
R3370 VGND.n429 VGND.t1611 34.8005
R3371 VGND.n429 VGND.t1726 34.8005
R3372 VGND.n2019 VGND.t310 34.8005
R3373 VGND.n2019 VGND.t1724 34.8005
R3374 VGND.n421 VGND.t2568 34.8005
R3375 VGND.n421 VGND.t1597 34.8005
R3376 VGND.n2045 VGND.t726 34.8005
R3377 VGND.n2045 VGND.t74 34.8005
R3378 VGND.n413 VGND.t2049 34.8005
R3379 VGND.n413 VGND.t1728 34.8005
R3380 VGND.n2071 VGND.t392 34.8005
R3381 VGND.n2071 VGND.t1605 34.8005
R3382 VGND.n405 VGND.t2323 34.8005
R3383 VGND.n405 VGND.t1603 34.8005
R3384 VGND.n2102 VGND.t2020 34.8005
R3385 VGND.n2102 VGND.t1722 34.8005
R3386 VGND.n2107 VGND.t2335 34.8005
R3387 VGND.n2107 VGND.t1720 34.8005
R3388 VGND.n2112 VGND.t143 34.8005
R3389 VGND.n2112 VGND.t1718 34.8005
R3390 VGND.n397 VGND.t381 34.8005
R3391 VGND.n397 VGND.t72 34.8005
R3392 VGND.n642 VGND.t1858 34.8005
R3393 VGND.n642 VGND.t1997 34.8005
R3394 VGND.n648 VGND.t283 34.8005
R3395 VGND.n648 VGND.t1524 34.8005
R3396 VGND.n645 VGND.t2172 34.8005
R3397 VGND.n645 VGND.t2005 34.8005
R3398 VGND.n1980 VGND.t57 34.8005
R3399 VGND.n1980 VGND.t2003 34.8005
R3400 VGND.n433 VGND.t1554 34.8005
R3401 VGND.n433 VGND.t1995 34.8005
R3402 VGND.n2006 VGND.t2084 34.8005
R3403 VGND.n2006 VGND.t1520 34.8005
R3404 VGND.n425 VGND.t925 34.8005
R3405 VGND.n425 VGND.t1518 34.8005
R3406 VGND.n2032 VGND.t2578 34.8005
R3407 VGND.n2032 VGND.t1993 34.8005
R3408 VGND.n417 VGND.t998 34.8005
R3409 VGND.n417 VGND.t1991 34.8005
R3410 VGND.n2058 VGND.t653 34.8005
R3411 VGND.n2058 VGND.t1522 34.8005
R3412 VGND.n409 VGND.t365 34.8005
R3413 VGND.n409 VGND.t2001 34.8005
R3414 VGND.n2084 VGND.t2160 34.8005
R3415 VGND.n2084 VGND.t1999 34.8005
R3416 VGND.n401 VGND.t1533 34.8005
R3417 VGND.n401 VGND.t1516 34.8005
R3418 VGND.n2089 VGND.t109 34.8005
R3419 VGND.n2089 VGND.t354 34.8005
R3420 VGND.n2328 VGND.t890 34.8005
R3421 VGND.n2328 VGND.t352 34.8005
R3422 VGND.n315 VGND.t516 34.8005
R3423 VGND.n315 VGND.t1526 34.8005
R3424 VGND.n658 VGND.t1900 34.8005
R3425 VGND.n658 VGND.t619 34.8005
R3426 VGND.n955 VGND.t2384 34.8005
R3427 VGND.n955 VGND.t1121 34.8005
R3428 VGND.n950 VGND.t68 34.8005
R3429 VGND.n950 VGND.t222 34.8005
R3430 VGND.n945 VGND.t1699 34.8005
R3431 VGND.n945 VGND.t2082 34.8005
R3432 VGND.n940 VGND.t1306 34.8005
R3433 VGND.n940 VGND.t617 34.8005
R3434 VGND.n935 VGND.t2344 34.8005
R3435 VGND.n935 VGND.t1117 34.8005
R3436 VGND.n930 VGND.t293 34.8005
R3437 VGND.n930 VGND.t1115 34.8005
R3438 VGND.n925 VGND.t485 34.8005
R3439 VGND.n925 VGND.t615 34.8005
R3440 VGND.n920 VGND.t804 34.8005
R3441 VGND.n920 VGND.t613 34.8005
R3442 VGND.n915 VGND.t1143 34.8005
R3443 VGND.n915 VGND.t1119 34.8005
R3444 VGND.n910 VGND.t387 34.8005
R3445 VGND.n910 VGND.t2080 34.8005
R3446 VGND.n905 VGND.t1594 34.8005
R3447 VGND.n905 VGND.t2078 34.8005
R3448 VGND.n900 VGND.t1566 34.8005
R3449 VGND.n900 VGND.t228 34.8005
R3450 VGND.n447 VGND.t2331 34.8005
R3451 VGND.n447 VGND.t226 34.8005
R3452 VGND.n1957 VGND.t2032 34.8005
R3453 VGND.n1957 VGND.t224 34.8005
R3454 VGND.n450 VGND.t377 34.8005
R3455 VGND.n450 VGND.t808 34.8005
R3456 VGND.n667 VGND.t1912 34.8005
R3457 VGND.n667 VGND.t344 34.8005
R3458 VGND.n1391 VGND.t2377 34.8005
R3459 VGND.n1391 VGND.t498 34.8005
R3460 VGND.n1396 VGND.t1129 34.8005
R3461 VGND.n1396 VGND.t1267 34.8005
R3462 VGND.n664 VGND.t1705 34.8005
R3463 VGND.n664 VGND.t350 34.8005
R3464 VGND.n1819 VGND.t1300 34.8005
R3465 VGND.n1819 VGND.t342 34.8005
R3466 VGND.n485 VGND.t626 34.8005
R3467 VGND.n485 VGND.t494 34.8005
R3468 VGND.n1845 VGND.t289 34.8005
R3469 VGND.n1845 VGND.t492 34.8005
R3470 VGND.n477 VGND.t479 34.8005
R3471 VGND.n477 VGND.t340 34.8005
R3472 VGND.n1871 VGND.t7 34.8005
R3473 VGND.n1871 VGND.t338 34.8005
R3474 VGND.n469 VGND.t1137 34.8005
R3475 VGND.n469 VGND.t496 34.8005
R3476 VGND.n1897 VGND.t2601 34.8005
R3477 VGND.n1897 VGND.t348 34.8005
R3478 VGND.n461 VGND.t1590 34.8005
R3479 VGND.n461 VGND.t346 34.8005
R3480 VGND.n1928 VGND.t1562 34.8005
R3481 VGND.n1928 VGND.t490 34.8005
R3482 VGND.n1933 VGND.t847 34.8005
R3483 VGND.n1933 VGND.t488 34.8005
R3484 VGND.n1938 VGND.t259 34.8005
R3485 VGND.n1938 VGND.t1269 34.8005
R3486 VGND.n453 VGND.t373 34.8005
R3487 VGND.n453 VGND.t2339 34.8005
R3488 VGND.n1370 VGND.t1840 34.8005
R3489 VGND.n1370 VGND.t1339 34.8005
R3490 VGND.n1376 VGND.t766 34.8005
R3491 VGND.n1376 VGND.t558 34.8005
R3492 VGND.n1373 VGND.t1360 34.8005
R3493 VGND.n1373 VGND.t1347 34.8005
R3494 VGND.n1806 VGND.t1984 34.8005
R3495 VGND.n1806 VGND.t1345 34.8005
R3496 VGND.n489 VGND.t2200 34.8005
R3497 VGND.n489 VGND.t1337 34.8005
R3498 VGND.n1832 VGND.t261 34.8005
R3499 VGND.n1832 VGND.t554 34.8005
R3500 VGND.n481 VGND.t333 34.8005
R3501 VGND.n481 VGND.t552 34.8005
R3502 VGND.n1858 VGND.t506 34.8005
R3503 VGND.n1858 VGND.t564 34.8005
R3504 VGND.n473 VGND.t314 34.8005
R3505 VGND.n473 VGND.t562 34.8005
R3506 VGND.n1884 VGND.t915 34.8005
R3507 VGND.n1884 VGND.t556 34.8005
R3508 VGND.n465 VGND.t369 34.8005
R3509 VGND.n465 VGND.t1343 34.8005
R3510 VGND.n1910 VGND.t306 34.8005
R3511 VGND.n1910 VGND.t1341 34.8005
R3512 VGND.n457 VGND.t2514 34.8005
R3513 VGND.n457 VGND.t550 34.8005
R3514 VGND.n1915 VGND.t112 34.8005
R3515 VGND.n1915 VGND.t548 34.8005
R3516 VGND.n2353 VGND.t1536 34.8005
R3517 VGND.n2353 VGND.t546 34.8005
R3518 VGND.n303 VGND.t520 34.8005
R3519 VGND.n303 VGND.t560 34.8005
R3520 VGND.n1302 VGND.t1936 34.8005
R3521 VGND.n1302 VGND.t2518 34.8005
R3522 VGND.n1308 VGND.t991 34.8005
R3523 VGND.n1308 VGND.t2502 34.8005
R3524 VGND.n1305 VGND.t2166 34.8005
R3525 VGND.n1305 VGND.t2526 34.8005
R3526 VGND.n1358 VGND.t356 34.8005
R3527 VGND.n1358 VGND.t2524 34.8005
R3528 VGND.n1353 VGND.t2636 34.8005
R3529 VGND.n1353 VGND.t91 34.8005
R3530 VGND.n1348 VGND.t2130 34.8005
R3531 VGND.n1348 VGND.t2498 34.8005
R3532 VGND.n1343 VGND.t300 34.8005
R3533 VGND.n1343 VGND.t2496 34.8005
R3534 VGND.n1338 VGND.t2682 34.8005
R3535 VGND.n1338 VGND.t2508 34.8005
R3536 VGND.n1333 VGND.t1149 34.8005
R3537 VGND.n1333 VGND.t2506 34.8005
R3538 VGND.n1328 VGND.t2178 34.8005
R3539 VGND.n1328 VGND.t2500 34.8005
R3540 VGND.n1323 VGND.t2595 34.8005
R3541 VGND.n1323 VGND.t2522 34.8005
R3542 VGND.n1318 VGND.t1389 34.8005
R3543 VGND.n1318 VGND.t2520 34.8005
R3544 VGND.n1313 VGND.t1660 34.8005
R3545 VGND.n1313 VGND.t2532 34.8005
R3546 VGND.n503 VGND.t840 34.8005
R3547 VGND.n503 VGND.t2530 34.8005
R3548 VGND.n1783 VGND.t1112 34.8005
R3549 VGND.n1783 VGND.t2528 34.8005
R3550 VGND.n506 VGND.t2585 34.8005
R3551 VGND.n506 VGND.t2504 34.8005
R3552 VGND.n571 VGND.t1867 34.8005
R3553 VGND.n571 VGND.t2627 34.8005
R3554 VGND.n1513 VGND.t279 34.8005
R3555 VGND.n1513 VGND.t695 34.8005
R3556 VGND.n1518 VGND.t2168 34.8005
R3557 VGND.n1518 VGND.t2614 34.8005
R3558 VGND.n575 VGND.t61 34.8005
R3559 VGND.n575 VGND.t2612 34.8005
R3560 VGND.n1645 VGND.t1550 34.8005
R3561 VGND.n1645 VGND.t2625 34.8005
R3562 VGND.n541 VGND.t1617 34.8005
R3563 VGND.n541 VGND.t691 34.8005
R3564 VGND.n1671 VGND.t921 34.8005
R3565 VGND.n1671 VGND.t689 34.8005
R3566 VGND.n533 VGND.t2574 34.8005
R3567 VGND.n533 VGND.t2623 34.8005
R3568 VGND.n1697 VGND.t994 34.8005
R3569 VGND.n1697 VGND.t2621 34.8005
R3570 VGND.n525 VGND.t649 34.8005
R3571 VGND.n525 VGND.t693 34.8005
R3572 VGND.n1723 VGND.t2564 34.8005
R3573 VGND.n1723 VGND.t2610 34.8005
R3574 VGND.n517 VGND.t2156 34.8005
R3575 VGND.n517 VGND.t2608 34.8005
R3576 VGND.n1754 VGND.t1529 34.8005
R3577 VGND.n1754 VGND.t687 34.8005
R3578 VGND.n1759 VGND.t105 34.8005
R3579 VGND.n1759 VGND.t2404 34.8005
R3580 VGND.n1764 VGND.t733 34.8005
R3581 VGND.n1764 VGND.t2616 34.8005
R3582 VGND.n509 VGND.t512 34.8005
R3583 VGND.n509 VGND.t2619 34.8005
R3584 VGND.n567 VGND.t1939 34.8005
R3585 VGND.n567 VGND.t17 34.8005
R3586 VGND.n1533 VGND.t989 34.8005
R3587 VGND.n1533 VGND.t2216 34.8005
R3588 VGND.n564 VGND.t2164 34.8005
R3589 VGND.n564 VGND.t2111 34.8005
R3590 VGND.n1632 VGND.t358 34.8005
R3591 VGND.n1632 VGND.t2109 34.8005
R3592 VGND.n545 VGND.t2634 34.8005
R3593 VGND.n545 VGND.t2554 34.8005
R3594 VGND.n1658 VGND.t2248 34.8005
R3595 VGND.n1658 VGND.t2212 34.8005
R3596 VGND.n537 VGND.t298 34.8005
R3597 VGND.n537 VGND.t2119 34.8005
R3598 VGND.n1684 VGND.t2680 34.8005
R3599 VGND.n1684 VGND.t2222 34.8005
R3600 VGND.n529 VGND.t1147 34.8005
R3601 VGND.n529 VGND.t2220 34.8005
R3602 VGND.n1710 VGND.t2176 34.8005
R3603 VGND.n1710 VGND.t2214 34.8005
R3604 VGND.n521 VGND.t2593 34.8005
R3605 VGND.n521 VGND.t21 34.8005
R3606 VGND.n1736 VGND.t1387 34.8005
R3607 VGND.n1736 VGND.t19 34.8005
R3608 VGND.n513 VGND.t1578 34.8005
R3609 VGND.n513 VGND.t2117 34.8005
R3610 VGND.n1741 VGND.t838 34.8005
R3611 VGND.n1741 VGND.t2115 34.8005
R3612 VGND.n2378 VGND.t1110 34.8005
R3613 VGND.n2378 VGND.t2113 34.8005
R3614 VGND.n290 VGND.t2583 34.8005
R3615 VGND.n290 VGND.t2218 34.8005
R3616 VGND.n670 VGND.t1969 34.8005
R3617 VGND.n670 VGND.t2065 34.8005
R3618 VGND.n672 VGND.t470 34.8005
R3619 VGND.n672 VGND.t86 34.8005
R3620 VGND.n1546 VGND.t644 34.8005
R3621 VGND.n1546 VGND.t2016 34.8005
R3622 VGND.n1551 VGND.t10 34.8005
R3623 VGND.n1551 VGND.t1573 34.8005
R3624 VGND.n1556 VGND.t1166 34.8005
R3625 VGND.n1556 VGND.t2063 34.8005
R3626 VGND.n1561 VGND.t2151 34.8005
R3627 VGND.n1561 VGND.t82 34.8005
R3628 VGND.n1566 VGND.t433 34.8005
R3629 VGND.n1566 VGND.t80 34.8005
R3630 VGND.n1571 VGND.t502 34.8005
R3631 VGND.n1571 VGND.t2061 34.8005
R3632 VGND.n1576 VGND.t738 34.8005
R3633 VGND.n1576 VGND.t2059 34.8005
R3634 VGND.n1581 VGND.t124 34.8005
R3635 VGND.n1581 VGND.t84 34.8005
R3636 VGND.n1586 VGND.t406 34.8005
R3637 VGND.n1586 VGND.t1571 34.8005
R3638 VGND.n1591 VGND.t2038 34.8005
R3639 VGND.n1591 VGND.t2067 34.8005
R3640 VGND.n1596 VGND.t117 34.8005
R3641 VGND.n1596 VGND.t78 34.8005
R3642 VGND.n559 VGND.t605 34.8005
R3643 VGND.n559 VGND.t76 34.8005
R3644 VGND.n1609 VGND.t2536 34.8005
R3645 VGND.n1609 VGND.t2018 34.8005
R3646 VGND.n1601 VGND.t428 34.8005
R3647 VGND.n1601 VGND.t2057 34.8005
R3648 VGND.n824 VGND.t1909 34.8005
R3649 VGND.n824 VGND.t269 34.8005
R3650 VGND.n831 VGND.t2379 34.8005
R3651 VGND.n831 VGND.t568 34.8005
R3652 VGND.n836 VGND.t1131 34.8005
R3653 VGND.n836 VGND.t908 34.8005
R3654 VGND.n828 VGND.t1703 34.8005
R3655 VGND.n828 VGND.t906 34.8005
R3656 VGND.n886 VGND.t1302 34.8005
R3657 VGND.n886 VGND.t267 34.8005
R3658 VGND.n881 VGND.t628 34.8005
R3659 VGND.n881 VGND.t137 34.8005
R3660 VGND.n876 VGND.t287 34.8005
R3661 VGND.n876 VGND.t135 34.8005
R3662 VGND.n871 VGND.t477 34.8005
R3663 VGND.n871 VGND.t1694 34.8005
R3664 VGND.n866 VGND.t5 34.8005
R3665 VGND.n866 VGND.t1692 34.8005
R3666 VGND.n861 VGND.t1404 34.8005
R3667 VGND.n861 VGND.t139 34.8005
R3668 VGND.n856 VGND.t2599 34.8005
R3669 VGND.n856 VGND.t273 34.8005
R3670 VGND.n851 VGND.t1588 34.8005
R3671 VGND.n851 VGND.t271 34.8005
R3672 VGND.n846 VGND.t1560 34.8005
R3673 VGND.n846 VGND.t133 34.8005
R3674 VGND.n841 VGND.t845 34.8005
R3675 VGND.n841 VGND.t131 34.8005
R3676 VGND.n2398 VGND.t2028 34.8005
R3677 VGND.n2398 VGND.t910 34.8005
R3678 VGND.n278 VGND.t2591 34.8005
R3679 VGND.n278 VGND.t570 34.8005
R3680 VGND.n814 VGND.t1029 34.8005
R3681 VGND.n814 VGND.t1214 34.8005
R3682 VGND.n717 VGND.t2096 34.8005
R3683 VGND.n717 VGND.t1031 34.8005
R3684 VGND.n74 VGND.n72 34.6358
R3685 VGND.n1109 VGND.n1091 34.6358
R3686 VGND.n1105 VGND.n1091 34.6358
R3687 VGND.n1105 VGND.n1104 34.6358
R3688 VGND.n1104 VGND.n1103 34.6358
R3689 VGND.n1103 VGND.n1093 34.6358
R3690 VGND.n1087 VGND.n1061 34.6358
R3691 VGND.n1082 VGND.n1062 34.6358
R3692 VGND.n1078 VGND.n1062 34.6358
R3693 VGND.n1078 VGND.n1077 34.6358
R3694 VGND.n1077 VGND.n1076 34.6358
R3695 VGND.n1076 VGND.n1064 34.6358
R3696 VGND.n130 VGND.n125 34.6358
R3697 VGND.n135 VGND.n134 34.6358
R3698 VGND.n598 VGND.n593 34.6358
R3699 VGND.n603 VGND.n602 34.6358
R3700 VGND.n976 VGND.n975 34.6358
R3701 VGND.n984 VGND.n983 34.6358
R3702 VGND.n980 VGND.n979 34.6358
R3703 VGND.n1020 VGND.n1000 34.6358
R3704 VGND.n1016 VGND.n1000 34.6358
R3705 VGND.n1016 VGND.n1015 34.6358
R3706 VGND.n1015 VGND.n1014 34.6358
R3707 VGND.n1014 VGND.n1002 34.6358
R3708 VGND.n1056 VGND.n1030 34.6358
R3709 VGND.n1051 VGND.n1031 34.6358
R3710 VGND.n1047 VGND.n1031 34.6358
R3711 VGND.n1047 VGND.n1046 34.6358
R3712 VGND.n1046 VGND.n1045 34.6358
R3713 VGND.n1045 VGND.n1033 34.6358
R3714 VGND.n160 VGND.n155 34.6358
R3715 VGND.n165 VGND.n164 34.6358
R3716 VGND.n17 VGND.n16 34.6358
R3717 VGND.n19 VGND.n10 34.6358
R3718 VGND.n23 VGND.n10 34.6358
R3719 VGND.n24 VGND.n23 34.6358
R3720 VGND.n25 VGND.n24 34.6358
R3721 VGND.n25 VGND.n8 34.6358
R3722 VGND.n46 VGND.n45 34.6358
R3723 VGND.n48 VGND.n37 34.6358
R3724 VGND.n52 VGND.n37 34.6358
R3725 VGND.n53 VGND.n52 34.6358
R3726 VGND.n54 VGND.n53 34.6358
R3727 VGND.n54 VGND.n35 34.6358
R3728 VGND.n100 VGND.n99 34.6358
R3729 VGND.n104 VGND.n103 34.6358
R3730 VGND.n2859 VGND.n2858 34.6358
R3731 VGND.n2863 VGND.n2862 34.6358
R3732 VGND.n2891 VGND.n2890 34.6358
R3733 VGND.n2895 VGND.n2894 34.6358
R3734 VGND.n78 VGND.n77 34.6358
R3735 VGND.n2934 VGND.n2928 34.6358
R3736 VGND.n2937 VGND.n2936 34.6358
R3737 VGND.n2937 VGND.n2924 34.6358
R3738 VGND.n2941 VGND.n2924 34.6358
R3739 VGND.n2942 VGND.n2941 34.6358
R3740 VGND.n2943 VGND.n2942 34.6358
R3741 VGND.n2959 VGND.n58 34.6358
R3742 VGND.n2974 VGND.n2973 34.6358
R3743 VGND.n2976 VGND.n2965 34.6358
R3744 VGND.n2980 VGND.n2965 34.6358
R3745 VGND.n2981 VGND.n2980 34.6358
R3746 VGND.n2982 VGND.n2981 34.6358
R3747 VGND.n2982 VGND.n2963 34.6358
R3748 VGND.n2991 VGND.n2986 34.6358
R3749 VGND.n2 VGND.t2538 34.4422
R3750 VGND.n995 VGND.n898 33.1299
R3751 VGND.n2916 VGND.n2915 33.1299
R3752 VGND.n80 VGND.n62 32.377
R3753 VGND.n986 VGND.n985 32.377
R3754 VGND.n106 VGND.n105 32.377
R3755 VGND.n2865 VGND.n2864 32.377
R3756 VGND.n2897 VGND.n2896 32.377
R3757 VGND.n80 VGND.n79 32.377
R3758 VGND.n986 VGND.n964 32.0005
R3759 VGND.n141 VGND.n138 30.4946
R3760 VGND.n609 VGND.n606 30.4946
R3761 VGND.n171 VGND.n168 30.4946
R3762 VGND.n109 VGND.n86 29.8709
R3763 VGND.n1099 VGND.n1098 28.9887
R3764 VGND.n1072 VGND.n1071 28.9887
R3765 VGND.n1010 VGND.n1009 28.9887
R3766 VGND.n1041 VGND.n1040 28.9887
R3767 VGND.n18 VGND.n17 27.8593
R3768 VGND.n47 VGND.n46 27.8593
R3769 VGND.n2935 VGND.n2934 27.8593
R3770 VGND.n2975 VGND.n2974 27.8593
R3771 VGND.n119 VGND.n118 27.0003
R3772 VGND.n2870 VGND.n2869 26.8591
R3773 VGND.n983 VGND.n968 26.3534
R3774 VGND.n103 VGND.n92 26.3534
R3775 VGND.n2862 VGND.n2851 26.3534
R3776 VGND.n2894 VGND.n2883 26.3534
R3777 VGND.n77 VGND.n67 26.3534
R3778 VGND.n142 VGND.n141 25.977
R3779 VGND.n610 VGND.n609 25.977
R3780 VGND.n585 VGND.n582 25.977
R3781 VGND.n172 VGND.n171 25.977
R3782 VGND.n2902 VGND.n2877 25.977
R3783 VGND.n1095 VGND.t2659 24.9236
R3784 VGND.n1095 VGND.t2393 24.9236
R3785 VGND.n1097 VGND.t881 24.9236
R3786 VGND.n1097 VGND.t2558 24.9236
R3787 VGND.n1067 VGND.t95 24.9236
R3788 VGND.n1067 VGND.t96 24.9236
R3789 VGND.n1066 VGND.t2385 24.9236
R3790 VGND.n1066 VGND.t2395 24.9236
R3791 VGND.n1070 VGND.t97 24.9236
R3792 VGND.n1070 VGND.t886 24.9236
R3793 VGND.n1069 VGND.t882 24.9236
R3794 VGND.n1069 VGND.t2559 24.9236
R3795 VGND.n132 VGND.t885 24.9236
R3796 VGND.n132 VGND.t51 24.9236
R3797 VGND.n131 VGND.t2398 24.9236
R3798 VGND.n131 VGND.t1686 24.9236
R3799 VGND.n122 VGND.t1365 24.9236
R3800 VGND.n122 VGND.t879 24.9236
R3801 VGND.n121 VGND.t1537 24.9236
R3802 VGND.n121 VGND.t2389 24.9236
R3803 VGND.n140 VGND.t2336 24.9236
R3804 VGND.n140 VGND.t2337 24.9236
R3805 VGND.n139 VGND.t2628 24.9236
R3806 VGND.n139 VGND.t2629 24.9236
R3807 VGND.n600 VGND.t324 24.9236
R3808 VGND.n600 VGND.t2655 24.9236
R3809 VGND.n599 VGND.t54 24.9236
R3810 VGND.n599 VGND.t99 24.9236
R3811 VGND.n590 VGND.t542 24.9236
R3812 VGND.n590 VGND.t323 24.9236
R3813 VGND.n589 VGND.t400 24.9236
R3814 VGND.n589 VGND.t49 24.9236
R3815 VGND.n608 VGND.t544 24.9236
R3816 VGND.n608 VGND.t543 24.9236
R3817 VGND.n607 VGND.t402 24.9236
R3818 VGND.n607 VGND.t401 24.9236
R3819 VGND.n966 VGND.t2391 24.9236
R3820 VGND.n966 VGND.t1683 24.9236
R3821 VGND.n967 VGND.t524 24.9236
R3822 VGND.n967 VGND.t876 24.9236
R3823 VGND.n965 VGND.t528 24.9236
R3824 VGND.n965 VGND.t526 24.9236
R3825 VGND.n970 VGND.t878 24.9236
R3826 VGND.n970 VGND.t2556 24.9236
R3827 VGND.n1005 VGND.t2386 24.9236
R3828 VGND.n1005 VGND.t2396 24.9236
R3829 VGND.n1004 VGND.t2650 24.9236
R3830 VGND.n1004 VGND.t2653 24.9236
R3831 VGND.n1008 VGND.t884 24.9236
R3832 VGND.n1008 VGND.t2560 24.9236
R3833 VGND.n1007 VGND.t2394 24.9236
R3834 VGND.n1007 VGND.t1684 24.9236
R3835 VGND.n1036 VGND.t2131 24.9236
R3836 VGND.n1036 VGND.t2132 24.9236
R3837 VGND.n1035 VGND.t1685 24.9236
R3838 VGND.n1035 VGND.t1687 24.9236
R3839 VGND.n1039 VGND.t1681 24.9236
R3840 VGND.n1039 VGND.t93 24.9236
R3841 VGND.n1038 VGND.t53 24.9236
R3842 VGND.n1038 VGND.t98 24.9236
R3843 VGND.n162 VGND.t326 24.9236
R3844 VGND.n162 VGND.t2388 24.9236
R3845 VGND.n161 VGND.t322 24.9236
R3846 VGND.n161 VGND.t2652 24.9236
R3847 VGND.n152 VGND.t1002 24.9236
R3848 VGND.n152 VGND.t325 24.9236
R3849 VGND.n151 VGND.t2645 24.9236
R3850 VGND.n151 VGND.t321 24.9236
R3851 VGND.n170 VGND.t1000 24.9236
R3852 VGND.n170 VGND.t1001 24.9236
R3853 VGND.n169 VGND.t2647 24.9236
R3854 VGND.n169 VGND.t2646 24.9236
R3855 VGND.n13 VGND.t1826 24.9236
R3856 VGND.n13 VGND.t1745 24.9236
R3857 VGND.n12 VGND.t1755 24.9236
R3858 VGND.n12 VGND.t1763 24.9236
R3859 VGND.n42 VGND.t1805 24.9236
R3860 VGND.n42 VGND.t1837 24.9236
R3861 VGND.n41 VGND.t1761 24.9236
R3862 VGND.n41 VGND.t1800 24.9236
R3863 VGND.n40 VGND.t1811 24.9236
R3864 VGND.n40 VGND.t1779 24.9236
R3865 VGND.n39 VGND.t1771 24.9236
R3866 VGND.n39 VGND.t1829 24.9236
R3867 VGND.n95 VGND.t1751 24.9236
R3868 VGND.n95 VGND.t1792 24.9236
R3869 VGND.n94 VGND.t1809 24.9236
R3870 VGND.n94 VGND.t1749 24.9236
R3871 VGND.n91 VGND.t1759 24.9236
R3872 VGND.n91 VGND.t41 24.9236
R3873 VGND.n90 VGND.t1815 24.9236
R3874 VGND.n90 VGND.t415 24.9236
R3875 VGND.n89 VGND.t38 24.9236
R3876 VGND.n89 VGND.t44 24.9236
R3877 VGND.n88 VGND.t186 24.9236
R3878 VGND.n88 VGND.t2672 24.9236
R3879 VGND.n2854 VGND.t1783 24.9236
R3880 VGND.n2854 VGND.t1816 24.9236
R3881 VGND.n2853 VGND.t1831 24.9236
R3882 VGND.n2853 VGND.t1781 24.9236
R3883 VGND.n2850 VGND.t1788 24.9236
R3884 VGND.n2850 VGND.t2026 24.9236
R3885 VGND.n2849 VGND.t1743 24.9236
R3886 VGND.n2849 VGND.t1349 24.9236
R3887 VGND.n2848 VGND.t1579 24.9236
R3888 VGND.n2848 VGND.t1568 24.9236
R3889 VGND.n2847 VGND.t504 24.9236
R3890 VGND.n2847 VGND.t898 24.9236
R3891 VGND.n2886 VGND.t1787 24.9236
R3892 VGND.n2886 VGND.t1821 24.9236
R3893 VGND.n2885 VGND.t1767 24.9236
R3894 VGND.n2885 VGND.t1808 24.9236
R3895 VGND.n2882 VGND.t1791 24.9236
R3896 VGND.n2882 VGND.t1673 24.9236
R3897 VGND.n2881 VGND.t1776 24.9236
R3898 VGND.n2881 VGND.t756 24.9236
R3899 VGND.n2880 VGND.t1672 24.9236
R3900 VGND.n2880 VGND.t1670 24.9236
R3901 VGND.n2879 VGND.t752 24.9236
R3902 VGND.n2879 VGND.t746 24.9236
R3903 VGND.n65 VGND.t1798 24.9236
R3904 VGND.n65 VGND.t1835 24.9236
R3905 VGND.n66 VGND.t1802 24.9236
R3906 VGND.n66 VGND.t1504 24.9236
R3907 VGND.n64 VGND.t1500 24.9236
R3908 VGND.n64 VGND.t1494 24.9236
R3909 VGND.n69 VGND.t1794 24.9236
R3910 VGND.n69 VGND.t1828 24.9236
R3911 VGND.n2930 VGND.t1777 24.9236
R3912 VGND.n2930 VGND.t1814 24.9236
R3913 VGND.n2929 VGND.t1765 24.9236
R3914 VGND.n2929 VGND.t1804 24.9236
R3915 VGND.n2927 VGND.t1786 24.9236
R3916 VGND.n2927 VGND.t1747 24.9236
R3917 VGND.n2926 VGND.t1773 24.9236
R3918 VGND.n2926 VGND.t1830 24.9236
R3919 VGND.n2970 VGND.t1822 24.9236
R3920 VGND.n2970 VGND.t1774 24.9236
R3921 VGND.n2969 VGND.t1813 24.9236
R3922 VGND.n2969 VGND.t1757 24.9236
R3923 VGND.n2968 VGND.t1833 24.9236
R3924 VGND.n2968 VGND.t1806 24.9236
R3925 VGND.n2967 VGND.t1818 24.9236
R3926 VGND.n2967 VGND.t1790 24.9236
R3927 VGND.n142 VGND.n116 24.4711
R3928 VGND.n610 VGND.n581 24.4711
R3929 VGND.n585 VGND.n584 24.4711
R3930 VGND.n996 VGND.n995 24.4711
R3931 VGND.n1025 VGND.n999 24.4711
R3932 VGND.n172 VGND.n148 24.4711
R3933 VGND.n106 VGND.n85 24.4711
R3934 VGND.n2865 VGND.n2844 24.4711
R3935 VGND.n2897 VGND.n2876 24.4711
R3936 VGND.n2902 VGND.n2901 24.4711
R3937 VGND.n2917 VGND.n2916 24.4711
R3938 VGND.n2948 VGND.n2947 24.4711
R3939 VGND.n2873 VGND.n2845 23.7181
R3940 VGND.n1111 VGND.n1109 23.7181
R3941 VGND.n1083 VGND.n1061 23.7181
R3942 VGND.n1083 VGND.n1082 23.7181
R3943 VGND.n146 VGND.n115 23.7181
R3944 VGND.n990 VGND.n899 23.7181
R3945 VGND.n1021 VGND.n1020 23.7181
R3946 VGND.n1052 VGND.n1030 23.7181
R3947 VGND.n1052 VGND.n1051 23.7181
R3948 VGND.n3007 VGND.n8 23.7181
R3949 VGND.n2960 VGND.n35 23.7181
R3950 VGND.n2943 VGND.n2922 23.7181
R3951 VGND.n2960 VGND.n2959 23.7181
R3952 VGND.n2992 VGND.n2963 23.7181
R3953 VGND.n2992 VGND.n2991 23.7181
R3954 VGND.n991 VGND.n990 23.3417
R3955 VGND.n2911 VGND.n84 23.3417
R3956 VGND.n2911 VGND.n61 23.3417
R3957 VGND.n1099 VGND.n1096 21.4593
R3958 VGND.n1072 VGND.n1068 21.4593
R3959 VGND.n1010 VGND.n1006 21.4593
R3960 VGND.n1041 VGND.n1037 21.4593
R3961 VGND.n98 VGND.n97 21.0905
R3962 VGND.n2857 VGND.n2856 21.0905
R3963 VGND.n2889 VGND.n2888 21.0905
R3964 VGND.n71 VGND.n70 21.0905
R3965 VGND.n99 VGND.n98 20.3299
R3966 VGND.n2858 VGND.n2857 20.3299
R3967 VGND.n2890 VGND.n2889 20.3299
R3968 VGND.n72 VGND.n71 20.3299
R3969 VGND.n138 VGND.n123 19.9534
R3970 VGND.n606 VGND.n591 19.9534
R3971 VGND.n168 VGND.n153 19.9534
R3972 VGND.n1026 VGND.n1025 19.2005
R3973 VGND.n1057 VGND.n1056 19.2005
R3974 VGND.n2949 VGND.n2948 19.2005
R3975 VGND.n2954 VGND.n58 19.2005
R3976 VGND.t1374 VGND.t2435 16.8587
R3977 VGND.t239 VGND.t2433 16.8587
R3978 VGND.t2369 VGND.t901 16.8587
R3979 VGND.t535 VGND.t903 16.8587
R3980 VGND.n1089 VGND.n1088 16.077
R3981 VGND.n2988 VGND.n2987 16.077
R3982 VGND.n1027 VGND.n1026 15.4358
R3983 VGND.n2950 VGND.n2949 15.4358
R3984 VGND.n118 VGND.n117 14.6829
R3985 VGND.n1058 VGND.n1057 14.6829
R3986 VGND.n2869 VGND.n2868 14.6829
R3987 VGND.n2955 VGND.n2954 14.6829
R3988 VGND.n127 VGND.n126 14.5711
R3989 VGND.n595 VGND.n594 14.5711
R3990 VGND.n974 VGND.n973 14.5711
R3991 VGND.n157 VGND.n156 14.5711
R3992 VGND.n614 VGND.n582 14.3064
R3993 VGND.n2906 VGND.n2877 14.3064
R3994 VGND.n134 VGND.n133 13.9299
R3995 VGND.n602 VGND.n601 13.9299
R3996 VGND.n979 VGND.n971 13.9299
R3997 VGND.n164 VGND.n163 13.9299
R3998 VGND.n1021 VGND.n999 13.5534
R3999 VGND.n2947 VGND.n2922 13.5534
R4000 VGND.n146 VGND.n116 13.177
R4001 VGND.n614 VGND.n581 13.177
R4002 VGND.n176 VGND.n148 13.177
R4003 VGND.n112 VGND.n85 13.177
R4004 VGND.n2873 VGND.n2844 13.177
R4005 VGND.n2906 VGND.n2876 13.177
R4006 VGND.n176 VGND.n149 12.8005
R4007 VGND.n112 VGND.n86 12.8005
R4008 VGND.n3021 VGND.t2696 12.5645
R4009 VGND.n1088 VGND.n1087 10.5417
R4010 VGND.n2987 VGND.n2986 10.5417
R4011 VGND.n1059 VGND.n1058 10.0534
R4012 VGND.n2956 VGND.n2955 10.0534
R4013 VGND.n1100 VGND.n1099 9.3005
R4014 VGND.n1101 VGND.n1093 9.3005
R4015 VGND.n1103 VGND.n1102 9.3005
R4016 VGND.n1104 VGND.n1092 9.3005
R4017 VGND.n1106 VGND.n1105 9.3005
R4018 VGND.n1107 VGND.n1091 9.3005
R4019 VGND.n1109 VGND.n1108 9.3005
R4020 VGND.n1112 VGND.n1111 9.3005
R4021 VGND.n1073 VGND.n1072 9.3005
R4022 VGND.n1074 VGND.n1064 9.3005
R4023 VGND.n1076 VGND.n1075 9.3005
R4024 VGND.n1077 VGND.n1063 9.3005
R4025 VGND.n1079 VGND.n1078 9.3005
R4026 VGND.n1080 VGND.n1062 9.3005
R4027 VGND.n1082 VGND.n1081 9.3005
R4028 VGND.n1085 VGND.n1061 9.3005
R4029 VGND.n1087 VGND.n1086 9.3005
R4030 VGND.n1084 VGND.n1083 9.3005
R4031 VGND.n144 VGND.n116 9.3005
R4032 VGND.n128 VGND.n125 9.3005
R4033 VGND.n130 VGND.n129 9.3005
R4034 VGND.n134 VGND.n124 9.3005
R4035 VGND.n136 VGND.n135 9.3005
R4036 VGND.n138 VGND.n137 9.3005
R4037 VGND.n141 VGND.n120 9.3005
R4038 VGND.n143 VGND.n142 9.3005
R4039 VGND.n119 VGND.n115 9.3005
R4040 VGND.n146 VGND.n145 9.3005
R4041 VGND.n584 VGND.n583 9.3005
R4042 VGND.n587 VGND.n582 9.3005
R4043 VGND.n612 VGND.n581 9.3005
R4044 VGND.n596 VGND.n593 9.3005
R4045 VGND.n598 VGND.n597 9.3005
R4046 VGND.n602 VGND.n592 9.3005
R4047 VGND.n604 VGND.n603 9.3005
R4048 VGND.n606 VGND.n605 9.3005
R4049 VGND.n609 VGND.n588 9.3005
R4050 VGND.n611 VGND.n610 9.3005
R4051 VGND.n586 VGND.n585 9.3005
R4052 VGND.n614 VGND.n613 9.3005
R4053 VGND.n997 VGND.n996 9.3005
R4054 VGND.n988 VGND.n899 9.3005
R4055 VGND.n975 VGND.n972 9.3005
R4056 VGND.n977 VGND.n976 9.3005
R4057 VGND.n979 VGND.n978 9.3005
R4058 VGND.n981 VGND.n980 9.3005
R4059 VGND.n983 VGND.n982 9.3005
R4060 VGND.n984 VGND.n963 9.3005
R4061 VGND.n987 VGND.n986 9.3005
R4062 VGND.n993 VGND.n992 9.3005
R4063 VGND.n995 VGND.n994 9.3005
R4064 VGND.n990 VGND.n989 9.3005
R4065 VGND.n1011 VGND.n1010 9.3005
R4066 VGND.n1012 VGND.n1002 9.3005
R4067 VGND.n1014 VGND.n1013 9.3005
R4068 VGND.n1015 VGND.n1001 9.3005
R4069 VGND.n1017 VGND.n1016 9.3005
R4070 VGND.n1018 VGND.n1000 9.3005
R4071 VGND.n1020 VGND.n1019 9.3005
R4072 VGND.n1023 VGND.n999 9.3005
R4073 VGND.n1025 VGND.n1024 9.3005
R4074 VGND.n1028 VGND.n1027 9.3005
R4075 VGND.n1022 VGND.n1021 9.3005
R4076 VGND.n1042 VGND.n1041 9.3005
R4077 VGND.n1043 VGND.n1033 9.3005
R4078 VGND.n1045 VGND.n1044 9.3005
R4079 VGND.n1046 VGND.n1032 9.3005
R4080 VGND.n1048 VGND.n1047 9.3005
R4081 VGND.n1049 VGND.n1031 9.3005
R4082 VGND.n1051 VGND.n1050 9.3005
R4083 VGND.n1054 VGND.n1030 9.3005
R4084 VGND.n1056 VGND.n1055 9.3005
R4085 VGND.n1053 VGND.n1052 9.3005
R4086 VGND.n174 VGND.n148 9.3005
R4087 VGND.n158 VGND.n155 9.3005
R4088 VGND.n160 VGND.n159 9.3005
R4089 VGND.n164 VGND.n154 9.3005
R4090 VGND.n166 VGND.n165 9.3005
R4091 VGND.n168 VGND.n167 9.3005
R4092 VGND.n171 VGND.n150 9.3005
R4093 VGND.n173 VGND.n172 9.3005
R4094 VGND.n176 VGND.n175 9.3005
R4095 VGND.n3007 VGND.n3006 9.3005
R4096 VGND.n16 VGND.n15 9.3005
R4097 VGND.n17 VGND.n11 9.3005
R4098 VGND.n20 VGND.n19 9.3005
R4099 VGND.n21 VGND.n10 9.3005
R4100 VGND.n23 VGND.n22 9.3005
R4101 VGND.n24 VGND.n9 9.3005
R4102 VGND.n26 VGND.n25 9.3005
R4103 VGND.n27 VGND.n8 9.3005
R4104 VGND.n110 VGND.n86 9.3005
R4105 VGND.n99 VGND.n93 9.3005
R4106 VGND.n101 VGND.n100 9.3005
R4107 VGND.n103 VGND.n102 9.3005
R4108 VGND.n104 VGND.n87 9.3005
R4109 VGND.n107 VGND.n106 9.3005
R4110 VGND.n108 VGND.n85 9.3005
R4111 VGND.n112 VGND.n111 9.3005
R4112 VGND.n2871 VGND.n2845 9.3005
R4113 VGND.n2858 VGND.n2852 9.3005
R4114 VGND.n2860 VGND.n2859 9.3005
R4115 VGND.n2862 VGND.n2861 9.3005
R4116 VGND.n2863 VGND.n2846 9.3005
R4117 VGND.n2866 VGND.n2865 9.3005
R4118 VGND.n2867 VGND.n2844 9.3005
R4119 VGND.n2873 VGND.n2872 9.3005
R4120 VGND.n2901 VGND.n2900 9.3005
R4121 VGND.n2890 VGND.n2884 9.3005
R4122 VGND.n2892 VGND.n2891 9.3005
R4123 VGND.n2894 VGND.n2893 9.3005
R4124 VGND.n2895 VGND.n2878 9.3005
R4125 VGND.n2898 VGND.n2897 9.3005
R4126 VGND.n2899 VGND.n2876 9.3005
R4127 VGND.n2904 VGND.n2877 9.3005
R4128 VGND.n2903 VGND.n2902 9.3005
R4129 VGND.n2906 VGND.n2905 9.3005
R4130 VGND.n2918 VGND.n2917 9.3005
R4131 VGND.n72 VGND.n68 9.3005
R4132 VGND.n75 VGND.n74 9.3005
R4133 VGND.n77 VGND.n76 9.3005
R4134 VGND.n78 VGND.n63 9.3005
R4135 VGND.n81 VGND.n80 9.3005
R4136 VGND.n83 VGND.n82 9.3005
R4137 VGND.n2914 VGND.n2913 9.3005
R4138 VGND.n2916 VGND.n60 9.3005
R4139 VGND.n2912 VGND.n2911 9.3005
R4140 VGND.n2951 VGND.n2950 9.3005
R4141 VGND.n2932 VGND.n2928 9.3005
R4142 VGND.n2934 VGND.n2933 9.3005
R4143 VGND.n2936 VGND.n2925 9.3005
R4144 VGND.n2938 VGND.n2937 9.3005
R4145 VGND.n2939 VGND.n2924 9.3005
R4146 VGND.n2941 VGND.n2940 9.3005
R4147 VGND.n2942 VGND.n2923 9.3005
R4148 VGND.n2944 VGND.n2943 9.3005
R4149 VGND.n2947 VGND.n2946 9.3005
R4150 VGND.n2948 VGND.n2920 9.3005
R4151 VGND.n2945 VGND.n2922 9.3005
R4152 VGND.n45 VGND.n44 9.3005
R4153 VGND.n46 VGND.n38 9.3005
R4154 VGND.n49 VGND.n48 9.3005
R4155 VGND.n50 VGND.n37 9.3005
R4156 VGND.n52 VGND.n51 9.3005
R4157 VGND.n53 VGND.n36 9.3005
R4158 VGND.n55 VGND.n54 9.3005
R4159 VGND.n56 VGND.n35 9.3005
R4160 VGND.n2960 VGND.n57 9.3005
R4161 VGND.n2959 VGND.n2958 9.3005
R4162 VGND.n2957 VGND.n58 9.3005
R4163 VGND.n2973 VGND.n2972 9.3005
R4164 VGND.n2974 VGND.n2966 9.3005
R4165 VGND.n2977 VGND.n2976 9.3005
R4166 VGND.n2978 VGND.n2965 9.3005
R4167 VGND.n2980 VGND.n2979 9.3005
R4168 VGND.n2981 VGND.n2964 9.3005
R4169 VGND.n2983 VGND.n2982 9.3005
R4170 VGND.n2984 VGND.n2963 9.3005
R4171 VGND.n2992 VGND.n2985 9.3005
R4172 VGND.n2991 VGND.n2990 9.3005
R4173 VGND.n2989 VGND.n2986 9.3005
R4174 VGND.n100 VGND.n92 8.28285
R4175 VGND.n2859 VGND.n2851 8.28285
R4176 VGND.n2891 VGND.n2883 8.28285
R4177 VGND.n2712 VGND.n235 7.9105
R4178 VGND.n2714 VGND.n2713 7.9105
R4179 VGND.n2819 VGND.n189 7.9105
R4180 VGND.n2818 VGND.n190 7.9105
R4181 VGND.n2813 VGND.n195 7.9105
R4182 VGND.n2812 VGND.n196 7.9105
R4183 VGND.n2807 VGND.n201 7.9105
R4184 VGND.n2806 VGND.n202 7.9105
R4185 VGND.n2801 VGND.n207 7.9105
R4186 VGND.n2800 VGND.n208 7.9105
R4187 VGND.n2795 VGND.n213 7.9105
R4188 VGND.n2794 VGND.n214 7.9105
R4189 VGND.n2789 VGND.n219 7.9105
R4190 VGND.n2788 VGND.n220 7.9105
R4191 VGND.n2783 VGND.n2782 7.9105
R4192 VGND.n3001 VGND.n3000 7.9105
R4193 VGND.n2517 VGND.n2516 7.9105
R4194 VGND.n2823 VGND.n185 7.9105
R4195 VGND.n2822 VGND.n186 7.9105
R4196 VGND.n2504 VGND.n2503 7.9105
R4197 VGND.n2502 VGND.n248 7.9105
R4198 VGND.n2501 VGND.n249 7.9105
R4199 VGND.n2500 VGND.n250 7.9105
R4200 VGND.n2499 VGND.n251 7.9105
R4201 VGND.n2498 VGND.n252 7.9105
R4202 VGND.n2497 VGND.n253 7.9105
R4203 VGND.n2496 VGND.n254 7.9105
R4204 VGND.n2495 VGND.n255 7.9105
R4205 VGND.n2494 VGND.n256 7.9105
R4206 VGND.n2493 VGND.n257 7.9105
R4207 VGND.n2492 VGND.n258 7.9105
R4208 VGND.n2491 VGND.n2490 7.9105
R4209 VGND.n639 VGND.n180 7.9105
R4210 VGND.n2827 VGND.n2826 7.9105
R4211 VGND.n375 VGND.n374 7.9105
R4212 VGND.n2166 VGND.n2165 7.9105
R4213 VGND.n2175 VGND.n2174 7.9105
R4214 VGND.n2192 VGND.n2191 7.9105
R4215 VGND.n2201 VGND.n2200 7.9105
R4216 VGND.n2218 VGND.n2217 7.9105
R4217 VGND.n2227 VGND.n2226 7.9105
R4218 VGND.n2244 VGND.n2243 7.9105
R4219 VGND.n2253 VGND.n2252 7.9105
R4220 VGND.n2275 VGND.n2274 7.9105
R4221 VGND.n2297 VGND.n328 7.9105
R4222 VGND.n2296 VGND.n329 7.9105
R4223 VGND.n2294 VGND.n2293 7.9105
R4224 VGND.n2430 VGND.n2429 7.9105
R4225 VGND.n1433 VGND.n1420 7.9105
R4226 VGND.n1432 VGND.n1431 7.9105
R4227 VGND.n2153 VGND.n2152 7.9105
R4228 VGND.n2162 VGND.n2161 7.9105
R4229 VGND.n2179 VGND.n2178 7.9105
R4230 VGND.n2188 VGND.n2187 7.9105
R4231 VGND.n2205 VGND.n2204 7.9105
R4232 VGND.n2214 VGND.n2213 7.9105
R4233 VGND.n2231 VGND.n2230 7.9105
R4234 VGND.n2240 VGND.n2239 7.9105
R4235 VGND.n2257 VGND.n2256 7.9105
R4236 VGND.n2271 VGND.n2270 7.9105
R4237 VGND.n2300 VGND.n327 7.9105
R4238 VGND.n2302 VGND.n2301 7.9105
R4239 VGND.n2314 VGND.n324 7.9105
R4240 VGND.n2313 VGND.n2312 7.9105
R4241 VGND.n1437 VGND.n1436 7.9105
R4242 VGND.n1496 VGND.n1495 7.9105
R4243 VGND.n2149 VGND.n381 7.9105
R4244 VGND.n2148 VGND.n382 7.9105
R4245 VGND.n2147 VGND.n383 7.9105
R4246 VGND.n2146 VGND.n384 7.9105
R4247 VGND.n2145 VGND.n385 7.9105
R4248 VGND.n2144 VGND.n386 7.9105
R4249 VGND.n2143 VGND.n387 7.9105
R4250 VGND.n2142 VGND.n388 7.9105
R4251 VGND.n2141 VGND.n389 7.9105
R4252 VGND.n2140 VGND.n390 7.9105
R4253 VGND.n2139 VGND.n2138 7.9105
R4254 VGND.n2318 VGND.n321 7.9105
R4255 VGND.n2317 VGND.n322 7.9105
R4256 VGND.n2126 VGND.n2125 7.9105
R4257 VGND.n1414 VGND.n617 7.9105
R4258 VGND.n1500 VGND.n1499 7.9105
R4259 VGND.n630 VGND.n629 7.9105
R4260 VGND.n1992 VGND.n1991 7.9105
R4261 VGND.n2001 VGND.n2000 7.9105
R4262 VGND.n2018 VGND.n2017 7.9105
R4263 VGND.n2027 VGND.n2026 7.9105
R4264 VGND.n2044 VGND.n2043 7.9105
R4265 VGND.n2053 VGND.n2052 7.9105
R4266 VGND.n2070 VGND.n2069 7.9105
R4267 VGND.n2079 VGND.n2078 7.9105
R4268 VGND.n2101 VGND.n2100 7.9105
R4269 VGND.n2322 VGND.n318 7.9105
R4270 VGND.n2321 VGND.n319 7.9105
R4271 VGND.n399 VGND.n398 7.9105
R4272 VGND.n2122 VGND.n2121 7.9105
R4273 VGND.n1412 VGND.n644 7.9105
R4274 VGND.n656 VGND.n655 7.9105
R4275 VGND.n1979 VGND.n1978 7.9105
R4276 VGND.n1988 VGND.n1987 7.9105
R4277 VGND.n2005 VGND.n2004 7.9105
R4278 VGND.n2014 VGND.n2013 7.9105
R4279 VGND.n2031 VGND.n2030 7.9105
R4280 VGND.n2040 VGND.n2039 7.9105
R4281 VGND.n2057 VGND.n2056 7.9105
R4282 VGND.n2066 VGND.n2065 7.9105
R4283 VGND.n2083 VGND.n2082 7.9105
R4284 VGND.n2097 VGND.n2096 7.9105
R4285 VGND.n2325 VGND.n316 7.9105
R4286 VGND.n2327 VGND.n2326 7.9105
R4287 VGND.n2339 VGND.n312 7.9105
R4288 VGND.n2338 VGND.n2337 7.9105
R4289 VGND.n1409 VGND.n660 7.9105
R4290 VGND.n1408 VGND.n661 7.9105
R4291 VGND.n1975 VGND.n437 7.9105
R4292 VGND.n1974 VGND.n438 7.9105
R4293 VGND.n1973 VGND.n439 7.9105
R4294 VGND.n1972 VGND.n440 7.9105
R4295 VGND.n1971 VGND.n441 7.9105
R4296 VGND.n1970 VGND.n442 7.9105
R4297 VGND.n1969 VGND.n443 7.9105
R4298 VGND.n1968 VGND.n444 7.9105
R4299 VGND.n1967 VGND.n445 7.9105
R4300 VGND.n1966 VGND.n446 7.9105
R4301 VGND.n1965 VGND.n1964 7.9105
R4302 VGND.n2343 VGND.n309 7.9105
R4303 VGND.n2342 VGND.n310 7.9105
R4304 VGND.n1952 VGND.n1951 7.9105
R4305 VGND.n1390 VGND.n1389 7.9105
R4306 VGND.n1405 VGND.n663 7.9105
R4307 VGND.n1404 VGND.n1403 7.9105
R4308 VGND.n1818 VGND.n1817 7.9105
R4309 VGND.n1827 VGND.n1826 7.9105
R4310 VGND.n1844 VGND.n1843 7.9105
R4311 VGND.n1853 VGND.n1852 7.9105
R4312 VGND.n1870 VGND.n1869 7.9105
R4313 VGND.n1879 VGND.n1878 7.9105
R4314 VGND.n1896 VGND.n1895 7.9105
R4315 VGND.n1905 VGND.n1904 7.9105
R4316 VGND.n1927 VGND.n1926 7.9105
R4317 VGND.n2347 VGND.n306 7.9105
R4318 VGND.n2346 VGND.n307 7.9105
R4319 VGND.n455 VGND.n454 7.9105
R4320 VGND.n1948 VGND.n1947 7.9105
R4321 VGND.n1386 VGND.n1372 7.9105
R4322 VGND.n1384 VGND.n1383 7.9105
R4323 VGND.n1805 VGND.n1804 7.9105
R4324 VGND.n1814 VGND.n1813 7.9105
R4325 VGND.n1831 VGND.n1830 7.9105
R4326 VGND.n1840 VGND.n1839 7.9105
R4327 VGND.n1857 VGND.n1856 7.9105
R4328 VGND.n1866 VGND.n1865 7.9105
R4329 VGND.n1883 VGND.n1882 7.9105
R4330 VGND.n1892 VGND.n1891 7.9105
R4331 VGND.n1909 VGND.n1908 7.9105
R4332 VGND.n1923 VGND.n1922 7.9105
R4333 VGND.n2350 VGND.n304 7.9105
R4334 VGND.n2352 VGND.n2351 7.9105
R4335 VGND.n2364 VGND.n300 7.9105
R4336 VGND.n2363 VGND.n2362 7.9105
R4337 VGND.n1368 VGND.n1304 7.9105
R4338 VGND.n1367 VGND.n1365 7.9105
R4339 VGND.n1801 VGND.n493 7.9105
R4340 VGND.n1800 VGND.n494 7.9105
R4341 VGND.n1799 VGND.n495 7.9105
R4342 VGND.n1798 VGND.n496 7.9105
R4343 VGND.n1797 VGND.n497 7.9105
R4344 VGND.n1796 VGND.n498 7.9105
R4345 VGND.n1795 VGND.n499 7.9105
R4346 VGND.n1794 VGND.n500 7.9105
R4347 VGND.n1793 VGND.n501 7.9105
R4348 VGND.n1792 VGND.n502 7.9105
R4349 VGND.n1791 VGND.n1790 7.9105
R4350 VGND.n2368 VGND.n297 7.9105
R4351 VGND.n2367 VGND.n298 7.9105
R4352 VGND.n1778 VGND.n1777 7.9105
R4353 VGND.n1528 VGND.n573 7.9105
R4354 VGND.n1527 VGND.n574 7.9105
R4355 VGND.n1526 VGND.n1525 7.9105
R4356 VGND.n1644 VGND.n1643 7.9105
R4357 VGND.n1653 VGND.n1652 7.9105
R4358 VGND.n1670 VGND.n1669 7.9105
R4359 VGND.n1679 VGND.n1678 7.9105
R4360 VGND.n1696 VGND.n1695 7.9105
R4361 VGND.n1705 VGND.n1704 7.9105
R4362 VGND.n1722 VGND.n1721 7.9105
R4363 VGND.n1731 VGND.n1730 7.9105
R4364 VGND.n1753 VGND.n1752 7.9105
R4365 VGND.n2372 VGND.n294 7.9105
R4366 VGND.n2371 VGND.n295 7.9105
R4367 VGND.n511 VGND.n510 7.9105
R4368 VGND.n1774 VGND.n1773 7.9105
R4369 VGND.n1532 VGND.n1531 7.9105
R4370 VGND.n1541 VGND.n1540 7.9105
R4371 VGND.n1631 VGND.n1630 7.9105
R4372 VGND.n1640 VGND.n1639 7.9105
R4373 VGND.n1657 VGND.n1656 7.9105
R4374 VGND.n1666 VGND.n1665 7.9105
R4375 VGND.n1683 VGND.n1682 7.9105
R4376 VGND.n1692 VGND.n1691 7.9105
R4377 VGND.n1709 VGND.n1708 7.9105
R4378 VGND.n1718 VGND.n1717 7.9105
R4379 VGND.n1735 VGND.n1734 7.9105
R4380 VGND.n1749 VGND.n1748 7.9105
R4381 VGND.n2375 VGND.n291 7.9105
R4382 VGND.n2377 VGND.n2376 7.9105
R4383 VGND.n2389 VGND.n287 7.9105
R4384 VGND.n2388 VGND.n2387 7.9105
R4385 VGND.n1298 VGND.n1297 7.9105
R4386 VGND.n1545 VGND.n1544 7.9105
R4387 VGND.n1627 VGND.n549 7.9105
R4388 VGND.n1626 VGND.n550 7.9105
R4389 VGND.n1625 VGND.n551 7.9105
R4390 VGND.n1624 VGND.n552 7.9105
R4391 VGND.n1623 VGND.n553 7.9105
R4392 VGND.n1622 VGND.n554 7.9105
R4393 VGND.n1621 VGND.n555 7.9105
R4394 VGND.n1620 VGND.n556 7.9105
R4395 VGND.n1619 VGND.n557 7.9105
R4396 VGND.n1618 VGND.n558 7.9105
R4397 VGND.n1617 VGND.n1616 7.9105
R4398 VGND.n2393 VGND.n282 7.9105
R4399 VGND.n2392 VGND.n283 7.9105
R4400 VGND.n1604 VGND.n1603 7.9105
R4401 VGND.n896 VGND.n826 7.9105
R4402 VGND.n895 VGND.n827 7.9105
R4403 VGND.n894 VGND.n893 7.9105
R4404 VGND.n1275 VGND.n688 7.9105
R4405 VGND.n1274 VGND.n689 7.9105
R4406 VGND.n1267 VGND.n694 7.9105
R4407 VGND.n1266 VGND.n695 7.9105
R4408 VGND.n1259 VGND.n700 7.9105
R4409 VGND.n1258 VGND.n701 7.9105
R4410 VGND.n1251 VGND.n706 7.9105
R4411 VGND.n1250 VGND.n707 7.9105
R4412 VGND.n1243 VGND.n712 7.9105
R4413 VGND.n1242 VGND.n713 7.9105
R4414 VGND.n2397 VGND.n2396 7.9105
R4415 VGND.n284 VGND.n279 7.9105
R4416 VGND.n2408 VGND.n2407 7.9105
R4417 VGND.n1117 VGND.n677 7.9105
R4418 VGND.n1285 VGND.n1284 7.9105
R4419 VGND.n1279 VGND.n685 7.9105
R4420 VGND.n1278 VGND.n686 7.9105
R4421 VGND.n1271 VGND.n691 7.9105
R4422 VGND.n1270 VGND.n692 7.9105
R4423 VGND.n1263 VGND.n697 7.9105
R4424 VGND.n1262 VGND.n698 7.9105
R4425 VGND.n1255 VGND.n703 7.9105
R4426 VGND.n1254 VGND.n704 7.9105
R4427 VGND.n1247 VGND.n709 7.9105
R4428 VGND.n1246 VGND.n710 7.9105
R4429 VGND.n1239 VGND.n715 7.9105
R4430 VGND.n1238 VGND.n716 7.9105
R4431 VGND.n1237 VGND.n783 7.9105
R4432 VGND.n2412 VGND.n2411 7.9105
R4433 VGND.n133 VGND.n130 7.90638
R4434 VGND.n126 VGND.n125 7.90638
R4435 VGND.n601 VGND.n598 7.90638
R4436 VGND.n594 VGND.n593 7.90638
R4437 VGND.n976 VGND.n971 7.90638
R4438 VGND.n975 VGND.n974 7.90638
R4439 VGND.n163 VGND.n160 7.90638
R4440 VGND.n156 VGND.n155 7.90638
R4441 VGND.n1098 VGND.n1094 7.4049
R4442 VGND.n1071 VGND.n1065 7.4049
R4443 VGND.n1009 VGND.n1003 7.4049
R4444 VGND.n1040 VGND.n1034 7.4049
R4445 VGND VGND.n149 7.12482
R4446 VGND.n97 VGND.n96 6.85473
R4447 VGND.n2856 VGND.n2855 6.85473
R4448 VGND.n2888 VGND.n2887 6.85473
R4449 VGND.n19 VGND.n18 6.77697
R4450 VGND.n48 VGND.n47 6.77697
R4451 VGND.n2936 VGND.n2935 6.77697
R4452 VGND.n2976 VGND.n2975 6.77697
R4453 VGND.n3020 VGND.n3019 6.4005
R4454 VGND.n969 VGND.n968 5.27109
R4455 VGND.n73 VGND.n67 5.27109
R4456 VGND.n2569 VGND.n2568 4.5005
R4457 VGND.n2624 VGND.n2581 4.5005
R4458 VGND.n2621 VGND.n2620 4.5005
R4459 VGND.n2618 VGND.n2617 4.5005
R4460 VGND.n2615 VGND.n2614 4.5005
R4461 VGND.n2612 VGND.n2611 4.5005
R4462 VGND.n2609 VGND.n2608 4.5005
R4463 VGND.n2606 VGND.n2605 4.5005
R4464 VGND.n2603 VGND.n2602 4.5005
R4465 VGND.n2600 VGND.n2599 4.5005
R4466 VGND.n2597 VGND.n2596 4.5005
R4467 VGND.n2594 VGND.n2593 4.5005
R4468 VGND.n2591 VGND.n2590 4.5005
R4469 VGND.n2588 VGND.n2587 4.5005
R4470 VGND.n2650 VGND.n223 4.5005
R4471 VGND.n2659 VGND.n222 4.5005
R4472 VGND.n2646 VGND.n217 4.5005
R4473 VGND.n2667 VGND.n216 4.5005
R4474 VGND.n2642 VGND.n211 4.5005
R4475 VGND.n2675 VGND.n210 4.5005
R4476 VGND.n2638 VGND.n205 4.5005
R4477 VGND.n2683 VGND.n204 4.5005
R4478 VGND.n2634 VGND.n199 4.5005
R4479 VGND.n2691 VGND.n198 4.5005
R4480 VGND.n2630 VGND.n193 4.5005
R4481 VGND.n2699 VGND.n192 4.5005
R4482 VGND.n2626 VGND.n2625 4.5005
R4483 VGND.n2708 VGND.n2707 4.5005
R4484 VGND.n2523 VGND.n2522 4.5005
R4485 VGND.n2526 VGND.n2525 4.5005
R4486 VGND.n2529 VGND.n2528 4.5005
R4487 VGND.n2532 VGND.n2531 4.5005
R4488 VGND.n2535 VGND.n2534 4.5005
R4489 VGND.n2538 VGND.n2537 4.5005
R4490 VGND.n2541 VGND.n2540 4.5005
R4491 VGND.n2544 VGND.n2543 4.5005
R4492 VGND.n2547 VGND.n2546 4.5005
R4493 VGND.n2550 VGND.n2549 4.5005
R4494 VGND.n2553 VGND.n2552 4.5005
R4495 VGND.n2556 VGND.n2555 4.5005
R4496 VGND.n2559 VGND.n2558 4.5005
R4497 VGND.n2562 VGND.n2561 4.5005
R4498 VGND.n2565 VGND.n2564 4.5005
R4499 VGND.n2575 VGND.n2567 4.5005
R4500 VGND.n2583 VGND.n2582 4.5005
R4501 VGND.n2586 VGND.n2585 4.5005
R4502 VGND.n2651 VGND.n30 4.5005
R4503 VGND.n820 VGND.n819 4.5005
R4504 VGND.n817 VGND.n816 4.5005
R4505 VGND.n1137 VGND.n1136 4.5005
R4506 VGND.n1149 VGND.n807 4.5005
R4507 VGND.n1156 VGND.n805 4.5005
R4508 VGND.n1153 VGND.n1151 4.5005
R4509 VGND.n1169 VGND.n1168 4.5005
R4510 VGND.n1181 VGND.n799 4.5005
R4511 VGND.n1188 VGND.n797 4.5005
R4512 VGND.n1185 VGND.n1183 4.5005
R4513 VGND.n1201 VGND.n1200 4.5005
R4514 VGND.n1213 VGND.n791 4.5005
R4515 VGND.n1219 VGND.n789 4.5005
R4516 VGND.n1216 VGND.n1215 4.5005
R4517 VGND.n786 VGND.n785 4.5005
R4518 VGND.n823 VGND.n822 4.5005
R4519 VGND.n1121 VGND.n1120 4.5005
R4520 VGND.n1126 VGND.n680 4.5005
R4521 VGND.n812 VGND.n681 4.5005
R4522 VGND.n1139 VGND.n1138 4.5005
R4523 VGND.n1148 VGND.n1147 4.5005
R4524 VGND.n1158 VGND.n1157 4.5005
R4525 VGND.n1152 VGND.n804 4.5005
R4526 VGND.n1171 VGND.n1170 4.5005
R4527 VGND.n1180 VGND.n1179 4.5005
R4528 VGND.n1190 VGND.n1189 4.5005
R4529 VGND.n1184 VGND.n796 4.5005
R4530 VGND.n1203 VGND.n1202 4.5005
R4531 VGND.n1212 VGND.n1211 4.5005
R4532 VGND.n1222 VGND.n1221 4.5005
R4533 VGND.n788 VGND.n784 4.5005
R4534 VGND.n1233 VGND.n1232 4.5005
R4535 VGND.n1113 VGND.n1112 4.41365
R4536 VGND VGND.n3005 4.35375
R4537 VGND.n1090 VGND.n1089 4.05427
R4538 VGND.n583 VGND.n0 4.05427
R4539 VGND.n998 VGND.n997 4.05427
R4540 VGND.n1029 VGND.n1028 4.05427
R4541 VGND.n1060 VGND.n1059 4.05427
R4542 VGND VGND.n59 3.99438
R4543 VGND.n2919 VGND 3.99438
R4544 VGND.n2952 VGND 3.99438
R4545 VGND VGND.n2953 3.99437
R4546 VGND VGND.n28 3.99437
R4547 VGND.n1234 VGND.n274 3.77268
R4548 VGND.n3003 VGND.n3002 3.77268
R4549 VGND.n1119 VGND.n1118 3.77268
R4550 VGND.n2711 VGND.n2710 3.77268
R4551 VGND.n1281 VGND.n1280 3.77268
R4552 VGND.n2820 VGND.n188 3.77268
R4553 VGND.n1277 VGND.n687 3.77268
R4554 VGND.n2817 VGND.n2816 3.77268
R4555 VGND.n1272 VGND.n690 3.77268
R4556 VGND.n2815 VGND.n2814 3.77268
R4557 VGND.n1269 VGND.n693 3.77268
R4558 VGND.n2811 VGND.n2810 3.77268
R4559 VGND.n1264 VGND.n696 3.77268
R4560 VGND.n2809 VGND.n2808 3.77268
R4561 VGND.n1261 VGND.n699 3.77268
R4562 VGND.n2805 VGND.n2804 3.77268
R4563 VGND.n1256 VGND.n702 3.77268
R4564 VGND.n2803 VGND.n2802 3.77268
R4565 VGND.n1253 VGND.n705 3.77268
R4566 VGND.n2799 VGND.n2798 3.77268
R4567 VGND.n1248 VGND.n708 3.77268
R4568 VGND.n2797 VGND.n2796 3.77268
R4569 VGND.n1245 VGND.n711 3.77268
R4570 VGND.n2793 VGND.n2792 3.77268
R4571 VGND.n1240 VGND.n714 3.77268
R4572 VGND.n2791 VGND.n2790 3.77268
R4573 VGND.n1220 VGND.n280 3.77268
R4574 VGND.n2787 VGND.n2786 3.77268
R4575 VGND.n1236 VGND.n1235 3.77268
R4576 VGND.n2785 VGND.n2784 3.77268
R4577 VGND.n1283 VGND.n1282 3.77268
R4578 VGND.n2709 VGND.n184 3.77268
R4579 VGND.n2584 VGND.n2583 3.75914
R4580 VGND.n2589 VGND.n2586 3.75914
R4581 VGND.n1217 VGND.n786 3.75914
R4582 VGND.n823 VGND.n821 3.75914
R4583 VGND.n2584 VGND.n2569 3.4105
R4584 VGND.n2624 VGND.n2623 3.4105
R4585 VGND.n2622 VGND.n2621 3.4105
R4586 VGND.n2619 VGND.n2618 3.4105
R4587 VGND.n2616 VGND.n2615 3.4105
R4588 VGND.n2613 VGND.n2612 3.4105
R4589 VGND.n2610 VGND.n2609 3.4105
R4590 VGND.n2607 VGND.n2606 3.4105
R4591 VGND.n2604 VGND.n2603 3.4105
R4592 VGND.n2601 VGND.n2600 3.4105
R4593 VGND.n2598 VGND.n2597 3.4105
R4594 VGND.n2595 VGND.n2594 3.4105
R4595 VGND.n2592 VGND.n2591 3.4105
R4596 VGND.n2589 VGND.n2588 3.4105
R4597 VGND.n3003 VGND.n30 3.4105
R4598 VGND.n2785 VGND.n223 3.4105
R4599 VGND.n2786 VGND.n222 3.4105
R4600 VGND.n2791 VGND.n217 3.4105
R4601 VGND.n2792 VGND.n216 3.4105
R4602 VGND.n2797 VGND.n211 3.4105
R4603 VGND.n2798 VGND.n210 3.4105
R4604 VGND.n2803 VGND.n205 3.4105
R4605 VGND.n2804 VGND.n204 3.4105
R4606 VGND.n2809 VGND.n199 3.4105
R4607 VGND.n2810 VGND.n198 3.4105
R4608 VGND.n2815 VGND.n193 3.4105
R4609 VGND.n2816 VGND.n192 3.4105
R4610 VGND.n2625 VGND.n188 3.4105
R4611 VGND.n2709 VGND.n2708 3.4105
R4612 VGND.n2710 VGND.n2567 3.4105
R4613 VGND.n3002 VGND.n3001 3.4105
R4614 VGND.n2712 VGND.n2711 3.4105
R4615 VGND.n2517 VGND.n236 3.4105
R4616 VGND.n2491 VGND.n31 3.4105
R4617 VGND.n2822 VGND.n2821 3.4105
R4618 VGND.n2820 VGND.n2819 3.4105
R4619 VGND.n375 VGND.n187 3.4105
R4620 VGND.n640 VGND.n639 3.4105
R4621 VGND.n2430 VGND.n260 3.4105
R4622 VGND.n2165 VGND.n2164 3.4105
R4623 VGND.n2503 VGND.n191 3.4105
R4624 VGND.n2818 VGND.n2817 3.4105
R4625 VGND.n2163 VGND.n2162 3.4105
R4626 VGND.n2152 VGND.n2151 3.4105
R4627 VGND.n1434 VGND.n1433 3.4105
R4628 VGND.n2313 VGND.n325 3.4105
R4629 VGND.n2178 VGND.n2177 3.4105
R4630 VGND.n2176 VGND.n2175 3.4105
R4631 VGND.n2502 VGND.n194 3.4105
R4632 VGND.n2814 VGND.n2813 3.4105
R4633 VGND.n2147 VGND.n361 3.4105
R4634 VGND.n2148 VGND.n376 3.4105
R4635 VGND.n2150 VGND.n2149 3.4105
R4636 VGND.n1436 VGND.n1435 3.4105
R4637 VGND.n2125 VGND.n395 3.4105
R4638 VGND.n2146 VGND.n357 3.4105
R4639 VGND.n2189 VGND.n2188 3.4105
R4640 VGND.n2191 VGND.n2190 3.4105
R4641 VGND.n2501 VGND.n197 3.4105
R4642 VGND.n2812 VGND.n2811 3.4105
R4643 VGND.n2017 VGND.n2016 3.4105
R4644 VGND.n2002 VGND.n2001 3.4105
R4645 VGND.n1991 VGND.n1990 3.4105
R4646 VGND.n630 VGND.n380 3.4105
R4647 VGND.n1414 VGND.n638 3.4105
R4648 VGND.n2122 VGND.n396 3.4105
R4649 VGND.n2028 VGND.n2027 3.4105
R4650 VGND.n2145 VGND.n353 3.4105
R4651 VGND.n2204 VGND.n2203 3.4105
R4652 VGND.n2202 VGND.n2201 3.4105
R4653 VGND.n2500 VGND.n200 3.4105
R4654 VGND.n2808 VGND.n2807 3.4105
R4655 VGND.n2030 VGND.n2029 3.4105
R4656 VGND.n2015 VGND.n2014 3.4105
R4657 VGND.n2004 VGND.n2003 3.4105
R4658 VGND.n1989 VGND.n1988 3.4105
R4659 VGND.n1978 VGND.n1977 3.4105
R4660 VGND.n1412 VGND.n1411 3.4105
R4661 VGND.n2338 VGND.n313 3.4105
R4662 VGND.n2041 VGND.n2040 3.4105
R4663 VGND.n2043 VGND.n2042 3.4105
R4664 VGND.n2144 VGND.n349 3.4105
R4665 VGND.n2215 VGND.n2214 3.4105
R4666 VGND.n2217 VGND.n2216 3.4105
R4667 VGND.n2499 VGND.n203 3.4105
R4668 VGND.n2806 VGND.n2805 3.4105
R4669 VGND.n1970 VGND.n416 3.4105
R4670 VGND.n1971 VGND.n420 3.4105
R4671 VGND.n1972 VGND.n424 3.4105
R4672 VGND.n1973 VGND.n428 3.4105
R4673 VGND.n1974 VGND.n432 3.4105
R4674 VGND.n1976 VGND.n1975 3.4105
R4675 VGND.n1410 VGND.n1409 3.4105
R4676 VGND.n1951 VGND.n451 3.4105
R4677 VGND.n1969 VGND.n412 3.4105
R4678 VGND.n2056 VGND.n2055 3.4105
R4679 VGND.n2054 VGND.n2053 3.4105
R4680 VGND.n2143 VGND.n345 3.4105
R4681 VGND.n2230 VGND.n2229 3.4105
R4682 VGND.n2228 VGND.n2227 3.4105
R4683 VGND.n2498 VGND.n206 3.4105
R4684 VGND.n2802 VGND.n2801 3.4105
R4685 VGND.n1880 VGND.n1879 3.4105
R4686 VGND.n1869 VGND.n1868 3.4105
R4687 VGND.n1854 VGND.n1853 3.4105
R4688 VGND.n1843 VGND.n1842 3.4105
R4689 VGND.n1828 VGND.n1827 3.4105
R4690 VGND.n1817 VGND.n1816 3.4105
R4691 VGND.n1404 VGND.n436 3.4105
R4692 VGND.n1389 VGND.n657 3.4105
R4693 VGND.n1948 VGND.n452 3.4105
R4694 VGND.n1895 VGND.n1894 3.4105
R4695 VGND.n1968 VGND.n408 3.4105
R4696 VGND.n2067 VGND.n2066 3.4105
R4697 VGND.n2069 VGND.n2068 3.4105
R4698 VGND.n2142 VGND.n341 3.4105
R4699 VGND.n2241 VGND.n2240 3.4105
R4700 VGND.n2243 VGND.n2242 3.4105
R4701 VGND.n2497 VGND.n209 3.4105
R4702 VGND.n2800 VGND.n2799 3.4105
R4703 VGND.n1893 VGND.n1892 3.4105
R4704 VGND.n1882 VGND.n1881 3.4105
R4705 VGND.n1867 VGND.n1866 3.4105
R4706 VGND.n1856 VGND.n1855 3.4105
R4707 VGND.n1841 VGND.n1840 3.4105
R4708 VGND.n1830 VGND.n1829 3.4105
R4709 VGND.n1815 VGND.n1814 3.4105
R4710 VGND.n1804 VGND.n1803 3.4105
R4711 VGND.n1386 VGND.n1385 3.4105
R4712 VGND.n2363 VGND.n301 3.4105
R4713 VGND.n1908 VGND.n1907 3.4105
R4714 VGND.n1906 VGND.n1905 3.4105
R4715 VGND.n1967 VGND.n404 3.4105
R4716 VGND.n2082 VGND.n2081 3.4105
R4717 VGND.n2080 VGND.n2079 3.4105
R4718 VGND.n2141 VGND.n337 3.4105
R4719 VGND.n2256 VGND.n2255 3.4105
R4720 VGND.n2254 VGND.n2253 3.4105
R4721 VGND.n2496 VGND.n212 3.4105
R4722 VGND.n2796 VGND.n2795 3.4105
R4723 VGND.n1793 VGND.n460 3.4105
R4724 VGND.n1794 VGND.n464 3.4105
R4725 VGND.n1795 VGND.n468 3.4105
R4726 VGND.n1796 VGND.n472 3.4105
R4727 VGND.n1797 VGND.n476 3.4105
R4728 VGND.n1798 VGND.n480 3.4105
R4729 VGND.n1799 VGND.n484 3.4105
R4730 VGND.n1800 VGND.n488 3.4105
R4731 VGND.n1802 VGND.n1801 3.4105
R4732 VGND.n1368 VGND.n570 3.4105
R4733 VGND.n1777 VGND.n507 3.4105
R4734 VGND.n1792 VGND.n456 3.4105
R4735 VGND.n1924 VGND.n1923 3.4105
R4736 VGND.n1926 VGND.n1925 3.4105
R4737 VGND.n1966 VGND.n400 3.4105
R4738 VGND.n2098 VGND.n2097 3.4105
R4739 VGND.n2100 VGND.n2099 3.4105
R4740 VGND.n2140 VGND.n333 3.4105
R4741 VGND.n2272 VGND.n2271 3.4105
R4742 VGND.n2274 VGND.n2273 3.4105
R4743 VGND.n2495 VGND.n215 3.4105
R4744 VGND.n2794 VGND.n2793 3.4105
R4745 VGND.n1752 VGND.n1751 3.4105
R4746 VGND.n1732 VGND.n1731 3.4105
R4747 VGND.n1721 VGND.n1720 3.4105
R4748 VGND.n1706 VGND.n1705 3.4105
R4749 VGND.n1695 VGND.n1694 3.4105
R4750 VGND.n1680 VGND.n1679 3.4105
R4751 VGND.n1669 VGND.n1668 3.4105
R4752 VGND.n1654 VGND.n1653 3.4105
R4753 VGND.n1643 VGND.n1642 3.4105
R4754 VGND.n1526 VGND.n492 3.4105
R4755 VGND.n1529 VGND.n1528 3.4105
R4756 VGND.n1774 VGND.n508 3.4105
R4757 VGND.n2373 VGND.n2372 3.4105
R4758 VGND.n1791 VGND.n293 3.4105
R4759 VGND.n2350 VGND.n2349 3.4105
R4760 VGND.n2348 VGND.n2347 3.4105
R4761 VGND.n1965 VGND.n305 3.4105
R4762 VGND.n2325 VGND.n2324 3.4105
R4763 VGND.n2323 VGND.n2322 3.4105
R4764 VGND.n2139 VGND.n317 3.4105
R4765 VGND.n2300 VGND.n2299 3.4105
R4766 VGND.n2298 VGND.n2297 3.4105
R4767 VGND.n2494 VGND.n218 3.4105
R4768 VGND.n2790 VGND.n2789 3.4105
R4769 VGND.n2375 VGND.n2374 3.4105
R4770 VGND.n1750 VGND.n1749 3.4105
R4771 VGND.n1734 VGND.n1733 3.4105
R4772 VGND.n1719 VGND.n1718 3.4105
R4773 VGND.n1708 VGND.n1707 3.4105
R4774 VGND.n1693 VGND.n1692 3.4105
R4775 VGND.n1682 VGND.n1681 3.4105
R4776 VGND.n1667 VGND.n1666 3.4105
R4777 VGND.n1656 VGND.n1655 3.4105
R4778 VGND.n1641 VGND.n1640 3.4105
R4779 VGND.n1630 VGND.n1629 3.4105
R4780 VGND.n1531 VGND.n1530 3.4105
R4781 VGND.n2388 VGND.n288 3.4105
R4782 VGND.n2376 VGND.n281 3.4105
R4783 VGND.n2371 VGND.n2370 3.4105
R4784 VGND.n2369 VGND.n2368 3.4105
R4785 VGND.n2351 VGND.n296 3.4105
R4786 VGND.n2346 VGND.n2345 3.4105
R4787 VGND.n2344 VGND.n2343 3.4105
R4788 VGND.n2326 VGND.n308 3.4105
R4789 VGND.n2321 VGND.n2320 3.4105
R4790 VGND.n2319 VGND.n2318 3.4105
R4791 VGND.n2301 VGND.n320 3.4105
R4792 VGND.n2296 VGND.n2295 3.4105
R4793 VGND.n2493 VGND.n221 3.4105
R4794 VGND.n2788 VGND.n2787 3.4105
R4795 VGND.n2394 VGND.n2393 3.4105
R4796 VGND.n1617 VGND.n292 3.4105
R4797 VGND.n1618 VGND.n512 3.4105
R4798 VGND.n1619 VGND.n516 3.4105
R4799 VGND.n1620 VGND.n520 3.4105
R4800 VGND.n1621 VGND.n524 3.4105
R4801 VGND.n1622 VGND.n528 3.4105
R4802 VGND.n1623 VGND.n532 3.4105
R4803 VGND.n1624 VGND.n536 3.4105
R4804 VGND.n1625 VGND.n540 3.4105
R4805 VGND.n1626 VGND.n544 3.4105
R4806 VGND.n1628 VGND.n1627 3.4105
R4807 VGND.n1298 VGND.n569 3.4105
R4808 VGND.n1603 VGND.n1602 3.4105
R4809 VGND.n2392 VGND.n2391 3.4105
R4810 VGND.n2390 VGND.n2389 3.4105
R4811 VGND.n510 VGND.n286 3.4105
R4812 VGND.n2367 VGND.n2366 3.4105
R4813 VGND.n2365 VGND.n2364 3.4105
R4814 VGND.n454 VGND.n299 3.4105
R4815 VGND.n2342 VGND.n2341 3.4105
R4816 VGND.n2340 VGND.n2339 3.4105
R4817 VGND.n398 VGND.n311 3.4105
R4818 VGND.n2317 VGND.n2316 3.4105
R4819 VGND.n2315 VGND.n2314 3.4105
R4820 VGND.n2294 VGND.n323 3.4105
R4821 VGND.n2492 VGND.n224 3.4105
R4822 VGND.n2784 VGND.n2783 3.4105
R4823 VGND.n285 VGND.n284 3.4105
R4824 VGND.n2396 VGND.n2395 3.4105
R4825 VGND.n1242 VGND.n1241 3.4105
R4826 VGND.n1244 VGND.n1243 3.4105
R4827 VGND.n1250 VGND.n1249 3.4105
R4828 VGND.n1252 VGND.n1251 3.4105
R4829 VGND.n1258 VGND.n1257 3.4105
R4830 VGND.n1260 VGND.n1259 3.4105
R4831 VGND.n1266 VGND.n1265 3.4105
R4832 VGND.n1268 VGND.n1267 3.4105
R4833 VGND.n1274 VGND.n1273 3.4105
R4834 VGND.n1276 VGND.n1275 3.4105
R4835 VGND.n894 VGND.n548 3.4105
R4836 VGND.n897 VGND.n896 3.4105
R4837 VGND.n2408 VGND.n277 3.4105
R4838 VGND.n895 VGND.n562 3.4105
R4839 VGND.n1544 VGND.n1543 3.4105
R4840 VGND.n1542 VGND.n1541 3.4105
R4841 VGND.n1527 VGND.n563 3.4105
R4842 VGND.n1367 VGND.n1366 3.4105
R4843 VGND.n1384 VGND.n662 3.4105
R4844 VGND.n1406 VGND.n1405 3.4105
R4845 VGND.n1408 VGND.n1407 3.4105
R4846 VGND.n656 VGND.n631 3.4105
R4847 VGND.n1499 VGND.n1498 3.4105
R4848 VGND.n1497 VGND.n1496 3.4105
R4849 VGND.n1432 VGND.n183 3.4105
R4850 VGND.n2826 VGND.n2825 3.4105
R4851 VGND.n2824 VGND.n2823 3.4105
R4852 VGND.n2713 VGND.n184 3.4105
R4853 VGND.n1235 VGND.n784 3.4105
R4854 VGND.n1221 VGND.n1220 3.4105
R4855 VGND.n1212 VGND.n714 3.4105
R4856 VGND.n1202 VGND.n711 3.4105
R4857 VGND.n1184 VGND.n708 3.4105
R4858 VGND.n1189 VGND.n705 3.4105
R4859 VGND.n1180 VGND.n702 3.4105
R4860 VGND.n1170 VGND.n699 3.4105
R4861 VGND.n1152 VGND.n696 3.4105
R4862 VGND.n1157 VGND.n693 3.4105
R4863 VGND.n1148 VGND.n690 3.4105
R4864 VGND.n1138 VGND.n687 3.4105
R4865 VGND.n1281 VGND.n681 3.4105
R4866 VGND.n1282 VGND.n680 3.4105
R4867 VGND.n1234 VGND.n1233 3.4105
R4868 VGND.n1217 VGND.n1216 3.4105
R4869 VGND.n1219 VGND.n1218 3.4105
R4870 VGND.n1214 VGND.n1213 3.4105
R4871 VGND.n1201 VGND.n790 3.4105
R4872 VGND.n1186 VGND.n1185 3.4105
R4873 VGND.n1188 VGND.n1187 3.4105
R4874 VGND.n1182 VGND.n1181 3.4105
R4875 VGND.n1169 VGND.n798 3.4105
R4876 VGND.n1154 VGND.n1153 3.4105
R4877 VGND.n1156 VGND.n1155 3.4105
R4878 VGND.n1150 VGND.n1149 3.4105
R4879 VGND.n1137 VGND.n806 3.4105
R4880 VGND.n818 VGND.n817 3.4105
R4881 VGND.n821 VGND.n820 3.4105
R4882 VGND.n1120 VGND.n1119 3.4105
R4883 VGND.n1237 VGND.n1236 3.4105
R4884 VGND.n1238 VGND.n280 3.4105
R4885 VGND.n1240 VGND.n1239 3.4105
R4886 VGND.n1246 VGND.n1245 3.4105
R4887 VGND.n1248 VGND.n1247 3.4105
R4888 VGND.n1254 VGND.n1253 3.4105
R4889 VGND.n1256 VGND.n1255 3.4105
R4890 VGND.n1262 VGND.n1261 3.4105
R4891 VGND.n1264 VGND.n1263 3.4105
R4892 VGND.n1270 VGND.n1269 3.4105
R4893 VGND.n1272 VGND.n1271 3.4105
R4894 VGND.n1278 VGND.n1277 3.4105
R4895 VGND.n1280 VGND.n1279 3.4105
R4896 VGND.n1284 VGND.n1283 3.4105
R4897 VGND.n1118 VGND.n1117 3.4105
R4898 VGND.n2411 VGND.n274 3.4105
R4899 VGND.n980 VGND.n969 3.01226
R4900 VGND.n74 VGND.n73 3.01226
R4901 VGND.n964 VGND.n899 2.63579
R4902 VGND.n2523 VGND 2.52282
R4903 VGND.n2526 VGND 2.52282
R4904 VGND.n2529 VGND 2.52282
R4905 VGND.n2532 VGND 2.52282
R4906 VGND.n2535 VGND 2.52282
R4907 VGND.n2538 VGND 2.52282
R4908 VGND.n2541 VGND 2.52282
R4909 VGND.n2544 VGND 2.52282
R4910 VGND.n2547 VGND 2.52282
R4911 VGND.n2550 VGND 2.52282
R4912 VGND.n2553 VGND 2.52282
R4913 VGND.n2556 VGND 2.52282
R4914 VGND.n2559 VGND 2.52282
R4915 VGND.n2562 VGND 2.52282
R4916 VGND.n2565 VGND 2.52282
R4917 VGND.n985 VGND.n984 2.25932
R4918 VGND.n105 VGND.n104 2.25932
R4919 VGND.n2864 VGND.n2863 2.25932
R4920 VGND.n2896 VGND.n2895 2.25932
R4921 VGND.n83 VGND.n62 2.25932
R4922 VGND.n79 VGND.n78 2.25932
R4923 VGND.n135 VGND.n123 1.88285
R4924 VGND.n603 VGND.n591 1.88285
R4925 VGND.n165 VGND.n153 1.88285
R4926 VGND.n2566 VGND 1.79514
R4927 VGND.n1114 VGND.n275 1.75987
R4928 VGND.n2566 VGND 1.57193
R4929 VGND.n3004 VGND.n3003 1.54254
R4930 VGND.n3001 VGND.n29 1.54254
R4931 VGND.n2491 VGND.n2432 1.54254
R4932 VGND.n2431 VGND.n2430 1.54254
R4933 VGND.n2313 VGND.n259 1.54254
R4934 VGND.n2125 VGND.n2124 1.54254
R4935 VGND.n2123 VGND.n2122 1.54254
R4936 VGND.n2338 VGND.n314 1.54254
R4937 VGND.n1951 VGND.n1950 1.54254
R4938 VGND.n1949 VGND.n1948 1.54254
R4939 VGND.n2363 VGND.n302 1.54254
R4940 VGND.n1777 VGND.n1776 1.54254
R4941 VGND.n1775 VGND.n1774 1.54254
R4942 VGND.n2388 VGND.n289 1.54254
R4943 VGND.n1603 VGND.n276 1.54254
R4944 VGND.n2409 VGND.n2408 1.54254
R4945 VGND.n1234 VGND.n275 1.54254
R4946 VGND.n2411 VGND.n2410 1.54254
R4947 VGND.n992 VGND.n898 1.50638
R4948 VGND.n2915 VGND.n2914 1.50638
R4949 VGND VGND.n2520 1.3946
R4950 VGND.n2519 VGND 1.3946
R4951 VGND.n2518 VGND 1.3946
R4952 VGND VGND.n237 1.3946
R4953 VGND VGND.n1417 1.3946
R4954 VGND.n1416 VGND 1.3946
R4955 VGND.n1415 VGND 1.3946
R4956 VGND.n1413 VGND 1.3946
R4957 VGND VGND.n641 1.3946
R4958 VGND VGND.n1388 1.3946
R4959 VGND.n1387 VGND 1.3946
R4960 VGND.n1369 VGND 1.3946
R4961 VGND.n1301 VGND 1.3946
R4962 VGND.n1300 VGND 1.3946
R4963 VGND.n1299 VGND 1.3946
R4964 VGND VGND.n669 1.3946
R4965 VGND.n1115 VGND 1.3946
R4966 VGND VGND.n1116 1.3946
R4967 VGND.n1114 VGND.n1113 1.04507
R4968 VGND.n2708 VGND.n2569 1.00149
R4969 VGND.n2625 VGND.n2624 1.00149
R4970 VGND.n2621 VGND.n192 1.00149
R4971 VGND.n2618 VGND.n193 1.00149
R4972 VGND.n2615 VGND.n198 1.00149
R4973 VGND.n2612 VGND.n199 1.00149
R4974 VGND.n2609 VGND.n204 1.00149
R4975 VGND.n2606 VGND.n205 1.00149
R4976 VGND.n2603 VGND.n210 1.00149
R4977 VGND.n2600 VGND.n211 1.00149
R4978 VGND.n2597 VGND.n216 1.00149
R4979 VGND.n2594 VGND.n217 1.00149
R4980 VGND.n2591 VGND.n222 1.00149
R4981 VGND.n2588 VGND.n223 1.00149
R4982 VGND.n2586 VGND.n30 1.00149
R4983 VGND.n820 VGND.n680 1.00149
R4984 VGND.n817 VGND.n681 1.00149
R4985 VGND.n1138 VGND.n1137 1.00149
R4986 VGND.n1149 VGND.n1148 1.00149
R4987 VGND.n1157 VGND.n1156 1.00149
R4988 VGND.n1153 VGND.n1152 1.00149
R4989 VGND.n1170 VGND.n1169 1.00149
R4990 VGND.n1181 VGND.n1180 1.00149
R4991 VGND.n1189 VGND.n1188 1.00149
R4992 VGND.n1185 VGND.n1184 1.00149
R4993 VGND.n1202 VGND.n1201 1.00149
R4994 VGND.n1213 VGND.n1212 1.00149
R4995 VGND.n1221 VGND.n1219 1.00149
R4996 VGND.n1216 VGND.n784 1.00149
R4997 VGND.n1233 VGND.n786 1.00149
R4998 VGND.n1120 VGND.n823 1.00149
R4999 VGND.n2583 VGND.n2567 0.973133
R5000 VGND.n2834 VGND.n2 0.9305
R5001 VGND.n97 VGND.n93 0.929432
R5002 VGND.n2856 VGND.n2852 0.929432
R5003 VGND.n2888 VGND.n2884 0.929432
R5004 VGND.n70 VGND.n68 0.929432
R5005 VGND.n59 VGND.n1 0.916608
R5006 VGND VGND.n2523 0.839786
R5007 VGND VGND.n2526 0.839786
R5008 VGND VGND.n2529 0.839786
R5009 VGND VGND.n2532 0.839786
R5010 VGND VGND.n2535 0.839786
R5011 VGND VGND.n2538 0.839786
R5012 VGND VGND.n2541 0.839786
R5013 VGND VGND.n2544 0.839786
R5014 VGND VGND.n2547 0.839786
R5015 VGND VGND.n2550 0.839786
R5016 VGND VGND.n2553 0.839786
R5017 VGND VGND.n2556 0.839786
R5018 VGND VGND.n2559 0.839786
R5019 VGND VGND.n2562 0.839786
R5020 VGND VGND.n2565 0.839786
R5021 VGND.n3021 VGND.n3020 0.7755
R5022 VGND.n3022 VGND.n3021 0.774207
R5023 VGND.n117 VGND.n115 0.753441
R5024 VGND.n16 VGND.n14 0.753441
R5025 VGND.n45 VGND.n43 0.753441
R5026 VGND.n2868 VGND.n2845 0.753441
R5027 VGND.n2931 VGND.n2928 0.753441
R5028 VGND.n2973 VGND.n2971 0.753441
R5029 VGND.n3024 VGND.n3023 0.573119
R5030 VGND VGND.n0 0.542567
R5031 VGND.n3024 VGND.n1 0.507317
R5032 VGND.n3005 VGND.n3004 0.404308
R5033 VGND.n1096 VGND.n1093 0.376971
R5034 VGND.n1068 VGND.n1064 0.376971
R5035 VGND.n992 VGND.n991 0.376971
R5036 VGND.n1006 VGND.n1002 0.376971
R5037 VGND.n1037 VGND.n1033 0.376971
R5038 VGND.n84 VGND.n83 0.376971
R5039 VGND.n2914 VGND.n61 0.376971
R5040 VGND VGND.n3024 0.37415
R5041 VGND.n277 VGND.n274 0.362676
R5042 VGND.n1602 VGND.n277 0.362676
R5043 VGND.n1602 VGND.n288 0.362676
R5044 VGND.n508 VGND.n288 0.362676
R5045 VGND.n508 VGND.n507 0.362676
R5046 VGND.n507 VGND.n301 0.362676
R5047 VGND.n452 VGND.n301 0.362676
R5048 VGND.n452 VGND.n451 0.362676
R5049 VGND.n451 VGND.n313 0.362676
R5050 VGND.n396 VGND.n313 0.362676
R5051 VGND.n396 VGND.n395 0.362676
R5052 VGND.n395 VGND.n325 0.362676
R5053 VGND.n325 VGND.n260 0.362676
R5054 VGND.n260 VGND.n31 0.362676
R5055 VGND.n3002 VGND.n31 0.362676
R5056 VGND.n1118 VGND.n897 0.362676
R5057 VGND.n897 VGND.n569 0.362676
R5058 VGND.n1530 VGND.n569 0.362676
R5059 VGND.n1530 VGND.n1529 0.362676
R5060 VGND.n1529 VGND.n570 0.362676
R5061 VGND.n1385 VGND.n570 0.362676
R5062 VGND.n1385 VGND.n657 0.362676
R5063 VGND.n1410 VGND.n657 0.362676
R5064 VGND.n1411 VGND.n1410 0.362676
R5065 VGND.n1411 VGND.n638 0.362676
R5066 VGND.n1435 VGND.n638 0.362676
R5067 VGND.n1435 VGND.n1434 0.362676
R5068 VGND.n1434 VGND.n640 0.362676
R5069 VGND.n640 VGND.n236 0.362676
R5070 VGND.n2711 VGND.n236 0.362676
R5071 VGND.n1280 VGND.n548 0.362676
R5072 VGND.n1628 VGND.n548 0.362676
R5073 VGND.n1629 VGND.n1628 0.362676
R5074 VGND.n1629 VGND.n492 0.362676
R5075 VGND.n1802 VGND.n492 0.362676
R5076 VGND.n1803 VGND.n1802 0.362676
R5077 VGND.n1803 VGND.n436 0.362676
R5078 VGND.n1976 VGND.n436 0.362676
R5079 VGND.n1977 VGND.n1976 0.362676
R5080 VGND.n1977 VGND.n380 0.362676
R5081 VGND.n2150 VGND.n380 0.362676
R5082 VGND.n2151 VGND.n2150 0.362676
R5083 VGND.n2151 VGND.n187 0.362676
R5084 VGND.n2821 VGND.n187 0.362676
R5085 VGND.n2821 VGND.n2820 0.362676
R5086 VGND.n1277 VGND.n1276 0.362676
R5087 VGND.n1276 VGND.n544 0.362676
R5088 VGND.n1641 VGND.n544 0.362676
R5089 VGND.n1642 VGND.n1641 0.362676
R5090 VGND.n1642 VGND.n488 0.362676
R5091 VGND.n1815 VGND.n488 0.362676
R5092 VGND.n1816 VGND.n1815 0.362676
R5093 VGND.n1816 VGND.n432 0.362676
R5094 VGND.n1989 VGND.n432 0.362676
R5095 VGND.n1990 VGND.n1989 0.362676
R5096 VGND.n1990 VGND.n376 0.362676
R5097 VGND.n2163 VGND.n376 0.362676
R5098 VGND.n2164 VGND.n2163 0.362676
R5099 VGND.n2164 VGND.n191 0.362676
R5100 VGND.n2817 VGND.n191 0.362676
R5101 VGND.n1273 VGND.n1272 0.362676
R5102 VGND.n1273 VGND.n540 0.362676
R5103 VGND.n1655 VGND.n540 0.362676
R5104 VGND.n1655 VGND.n1654 0.362676
R5105 VGND.n1654 VGND.n484 0.362676
R5106 VGND.n1829 VGND.n484 0.362676
R5107 VGND.n1829 VGND.n1828 0.362676
R5108 VGND.n1828 VGND.n428 0.362676
R5109 VGND.n2003 VGND.n428 0.362676
R5110 VGND.n2003 VGND.n2002 0.362676
R5111 VGND.n2002 VGND.n361 0.362676
R5112 VGND.n2177 VGND.n361 0.362676
R5113 VGND.n2177 VGND.n2176 0.362676
R5114 VGND.n2176 VGND.n194 0.362676
R5115 VGND.n2814 VGND.n194 0.362676
R5116 VGND.n1269 VGND.n1268 0.362676
R5117 VGND.n1268 VGND.n536 0.362676
R5118 VGND.n1667 VGND.n536 0.362676
R5119 VGND.n1668 VGND.n1667 0.362676
R5120 VGND.n1668 VGND.n480 0.362676
R5121 VGND.n1841 VGND.n480 0.362676
R5122 VGND.n1842 VGND.n1841 0.362676
R5123 VGND.n1842 VGND.n424 0.362676
R5124 VGND.n2015 VGND.n424 0.362676
R5125 VGND.n2016 VGND.n2015 0.362676
R5126 VGND.n2016 VGND.n357 0.362676
R5127 VGND.n2189 VGND.n357 0.362676
R5128 VGND.n2190 VGND.n2189 0.362676
R5129 VGND.n2190 VGND.n197 0.362676
R5130 VGND.n2811 VGND.n197 0.362676
R5131 VGND.n1265 VGND.n1264 0.362676
R5132 VGND.n1265 VGND.n532 0.362676
R5133 VGND.n1681 VGND.n532 0.362676
R5134 VGND.n1681 VGND.n1680 0.362676
R5135 VGND.n1680 VGND.n476 0.362676
R5136 VGND.n1855 VGND.n476 0.362676
R5137 VGND.n1855 VGND.n1854 0.362676
R5138 VGND.n1854 VGND.n420 0.362676
R5139 VGND.n2029 VGND.n420 0.362676
R5140 VGND.n2029 VGND.n2028 0.362676
R5141 VGND.n2028 VGND.n353 0.362676
R5142 VGND.n2203 VGND.n353 0.362676
R5143 VGND.n2203 VGND.n2202 0.362676
R5144 VGND.n2202 VGND.n200 0.362676
R5145 VGND.n2808 VGND.n200 0.362676
R5146 VGND.n1261 VGND.n1260 0.362676
R5147 VGND.n1260 VGND.n528 0.362676
R5148 VGND.n1693 VGND.n528 0.362676
R5149 VGND.n1694 VGND.n1693 0.362676
R5150 VGND.n1694 VGND.n472 0.362676
R5151 VGND.n1867 VGND.n472 0.362676
R5152 VGND.n1868 VGND.n1867 0.362676
R5153 VGND.n1868 VGND.n416 0.362676
R5154 VGND.n2041 VGND.n416 0.362676
R5155 VGND.n2042 VGND.n2041 0.362676
R5156 VGND.n2042 VGND.n349 0.362676
R5157 VGND.n2215 VGND.n349 0.362676
R5158 VGND.n2216 VGND.n2215 0.362676
R5159 VGND.n2216 VGND.n203 0.362676
R5160 VGND.n2805 VGND.n203 0.362676
R5161 VGND.n1257 VGND.n1256 0.362676
R5162 VGND.n1257 VGND.n524 0.362676
R5163 VGND.n1707 VGND.n524 0.362676
R5164 VGND.n1707 VGND.n1706 0.362676
R5165 VGND.n1706 VGND.n468 0.362676
R5166 VGND.n1881 VGND.n468 0.362676
R5167 VGND.n1881 VGND.n1880 0.362676
R5168 VGND.n1880 VGND.n412 0.362676
R5169 VGND.n2055 VGND.n412 0.362676
R5170 VGND.n2055 VGND.n2054 0.362676
R5171 VGND.n2054 VGND.n345 0.362676
R5172 VGND.n2229 VGND.n345 0.362676
R5173 VGND.n2229 VGND.n2228 0.362676
R5174 VGND.n2228 VGND.n206 0.362676
R5175 VGND.n2802 VGND.n206 0.362676
R5176 VGND.n1253 VGND.n1252 0.362676
R5177 VGND.n1252 VGND.n520 0.362676
R5178 VGND.n1719 VGND.n520 0.362676
R5179 VGND.n1720 VGND.n1719 0.362676
R5180 VGND.n1720 VGND.n464 0.362676
R5181 VGND.n1893 VGND.n464 0.362676
R5182 VGND.n1894 VGND.n1893 0.362676
R5183 VGND.n1894 VGND.n408 0.362676
R5184 VGND.n2067 VGND.n408 0.362676
R5185 VGND.n2068 VGND.n2067 0.362676
R5186 VGND.n2068 VGND.n341 0.362676
R5187 VGND.n2241 VGND.n341 0.362676
R5188 VGND.n2242 VGND.n2241 0.362676
R5189 VGND.n2242 VGND.n209 0.362676
R5190 VGND.n2799 VGND.n209 0.362676
R5191 VGND.n1249 VGND.n1248 0.362676
R5192 VGND.n1249 VGND.n516 0.362676
R5193 VGND.n1733 VGND.n516 0.362676
R5194 VGND.n1733 VGND.n1732 0.362676
R5195 VGND.n1732 VGND.n460 0.362676
R5196 VGND.n1907 VGND.n460 0.362676
R5197 VGND.n1907 VGND.n1906 0.362676
R5198 VGND.n1906 VGND.n404 0.362676
R5199 VGND.n2081 VGND.n404 0.362676
R5200 VGND.n2081 VGND.n2080 0.362676
R5201 VGND.n2080 VGND.n337 0.362676
R5202 VGND.n2255 VGND.n337 0.362676
R5203 VGND.n2255 VGND.n2254 0.362676
R5204 VGND.n2254 VGND.n212 0.362676
R5205 VGND.n2796 VGND.n212 0.362676
R5206 VGND.n1245 VGND.n1244 0.362676
R5207 VGND.n1244 VGND.n512 0.362676
R5208 VGND.n1750 VGND.n512 0.362676
R5209 VGND.n1751 VGND.n1750 0.362676
R5210 VGND.n1751 VGND.n456 0.362676
R5211 VGND.n1924 VGND.n456 0.362676
R5212 VGND.n1925 VGND.n1924 0.362676
R5213 VGND.n1925 VGND.n400 0.362676
R5214 VGND.n2098 VGND.n400 0.362676
R5215 VGND.n2099 VGND.n2098 0.362676
R5216 VGND.n2099 VGND.n333 0.362676
R5217 VGND.n2272 VGND.n333 0.362676
R5218 VGND.n2273 VGND.n2272 0.362676
R5219 VGND.n2273 VGND.n215 0.362676
R5220 VGND.n2793 VGND.n215 0.362676
R5221 VGND.n1241 VGND.n1240 0.362676
R5222 VGND.n1241 VGND.n292 0.362676
R5223 VGND.n2374 VGND.n292 0.362676
R5224 VGND.n2374 VGND.n2373 0.362676
R5225 VGND.n2373 VGND.n293 0.362676
R5226 VGND.n2349 VGND.n293 0.362676
R5227 VGND.n2349 VGND.n2348 0.362676
R5228 VGND.n2348 VGND.n305 0.362676
R5229 VGND.n2324 VGND.n305 0.362676
R5230 VGND.n2324 VGND.n2323 0.362676
R5231 VGND.n2323 VGND.n317 0.362676
R5232 VGND.n2299 VGND.n317 0.362676
R5233 VGND.n2299 VGND.n2298 0.362676
R5234 VGND.n2298 VGND.n218 0.362676
R5235 VGND.n2790 VGND.n218 0.362676
R5236 VGND.n2395 VGND.n280 0.362676
R5237 VGND.n2395 VGND.n2394 0.362676
R5238 VGND.n2394 VGND.n281 0.362676
R5239 VGND.n2370 VGND.n281 0.362676
R5240 VGND.n2370 VGND.n2369 0.362676
R5241 VGND.n2369 VGND.n296 0.362676
R5242 VGND.n2345 VGND.n296 0.362676
R5243 VGND.n2345 VGND.n2344 0.362676
R5244 VGND.n2344 VGND.n308 0.362676
R5245 VGND.n2320 VGND.n308 0.362676
R5246 VGND.n2320 VGND.n2319 0.362676
R5247 VGND.n2319 VGND.n320 0.362676
R5248 VGND.n2295 VGND.n320 0.362676
R5249 VGND.n2295 VGND.n221 0.362676
R5250 VGND.n2787 VGND.n221 0.362676
R5251 VGND.n1236 VGND.n285 0.362676
R5252 VGND.n2391 VGND.n285 0.362676
R5253 VGND.n2391 VGND.n2390 0.362676
R5254 VGND.n2390 VGND.n286 0.362676
R5255 VGND.n2366 VGND.n286 0.362676
R5256 VGND.n2366 VGND.n2365 0.362676
R5257 VGND.n2365 VGND.n299 0.362676
R5258 VGND.n2341 VGND.n299 0.362676
R5259 VGND.n2341 VGND.n2340 0.362676
R5260 VGND.n2340 VGND.n311 0.362676
R5261 VGND.n2316 VGND.n311 0.362676
R5262 VGND.n2316 VGND.n2315 0.362676
R5263 VGND.n2315 VGND.n323 0.362676
R5264 VGND.n323 VGND.n224 0.362676
R5265 VGND.n2784 VGND.n224 0.362676
R5266 VGND.n1283 VGND.n562 0.362676
R5267 VGND.n1543 VGND.n562 0.362676
R5268 VGND.n1543 VGND.n1542 0.362676
R5269 VGND.n1542 VGND.n563 0.362676
R5270 VGND.n1366 VGND.n563 0.362676
R5271 VGND.n1366 VGND.n662 0.362676
R5272 VGND.n1406 VGND.n662 0.362676
R5273 VGND.n1407 VGND.n1406 0.362676
R5274 VGND.n1407 VGND.n631 0.362676
R5275 VGND.n1498 VGND.n631 0.362676
R5276 VGND.n1498 VGND.n1497 0.362676
R5277 VGND.n1497 VGND.n183 0.362676
R5278 VGND.n2825 VGND.n183 0.362676
R5279 VGND.n2825 VGND.n2824 0.362676
R5280 VGND.n2824 VGND.n184 0.362676
R5281 VGND.n2623 VGND.n2584 0.349144
R5282 VGND.n2623 VGND.n2622 0.349144
R5283 VGND.n2622 VGND.n2619 0.349144
R5284 VGND.n2619 VGND.n2616 0.349144
R5285 VGND.n2616 VGND.n2613 0.349144
R5286 VGND.n2613 VGND.n2610 0.349144
R5287 VGND.n2610 VGND.n2607 0.349144
R5288 VGND.n2607 VGND.n2604 0.349144
R5289 VGND.n2604 VGND.n2601 0.349144
R5290 VGND.n2601 VGND.n2598 0.349144
R5291 VGND.n2598 VGND.n2595 0.349144
R5292 VGND.n2595 VGND.n2592 0.349144
R5293 VGND.n2592 VGND.n2589 0.349144
R5294 VGND.n1218 VGND.n1217 0.349144
R5295 VGND.n1218 VGND.n1214 0.349144
R5296 VGND.n1214 VGND.n790 0.349144
R5297 VGND.n1186 VGND.n790 0.349144
R5298 VGND.n1187 VGND.n1186 0.349144
R5299 VGND.n1187 VGND.n1182 0.349144
R5300 VGND.n1182 VGND.n798 0.349144
R5301 VGND.n1154 VGND.n798 0.349144
R5302 VGND.n1155 VGND.n1154 0.349144
R5303 VGND.n1155 VGND.n1150 0.349144
R5304 VGND.n1150 VGND.n806 0.349144
R5305 VGND.n818 VGND.n806 0.349144
R5306 VGND.n821 VGND.n818 0.349144
R5307 VGND.n2655 VGND.n2650 0.327628
R5308 VGND.n2659 VGND.n2658 0.327628
R5309 VGND.n2663 VGND.n2646 0.327628
R5310 VGND.n2667 VGND.n2666 0.327628
R5311 VGND.n2671 VGND.n2642 0.327628
R5312 VGND.n2675 VGND.n2674 0.327628
R5313 VGND.n2679 VGND.n2638 0.327628
R5314 VGND.n2683 VGND.n2682 0.327628
R5315 VGND.n2687 VGND.n2634 0.327628
R5316 VGND.n2691 VGND.n2690 0.327628
R5317 VGND.n2695 VGND.n2630 0.327628
R5318 VGND.n2699 VGND.n2698 0.327628
R5319 VGND.n2703 VGND.n2626 0.327628
R5320 VGND.n2707 VGND.n2706 0.327628
R5321 VGND.n2577 VGND.n2575 0.327628
R5322 VGND.n2782 VGND.n2781 0.327628
R5323 VGND.n2778 VGND.n220 0.327628
R5324 VGND.n2773 VGND.n219 0.327628
R5325 VGND.n2768 VGND.n214 0.327628
R5326 VGND.n2763 VGND.n213 0.327628
R5327 VGND.n2758 VGND.n208 0.327628
R5328 VGND.n2753 VGND.n207 0.327628
R5329 VGND.n2748 VGND.n202 0.327628
R5330 VGND.n2743 VGND.n201 0.327628
R5331 VGND.n2738 VGND.n196 0.327628
R5332 VGND.n2733 VGND.n195 0.327628
R5333 VGND.n2728 VGND.n190 0.327628
R5334 VGND.n2723 VGND.n189 0.327628
R5335 VGND.n2718 VGND.n2714 0.327628
R5336 VGND.n235 VGND.n234 0.327628
R5337 VGND.n2487 VGND.n258 0.327628
R5338 VGND.n2482 VGND.n257 0.327628
R5339 VGND.n2477 VGND.n256 0.327628
R5340 VGND.n2472 VGND.n255 0.327628
R5341 VGND.n2467 VGND.n254 0.327628
R5342 VGND.n2462 VGND.n253 0.327628
R5343 VGND.n2457 VGND.n252 0.327628
R5344 VGND.n2452 VGND.n251 0.327628
R5345 VGND.n2447 VGND.n250 0.327628
R5346 VGND.n2442 VGND.n249 0.327628
R5347 VGND.n2437 VGND.n248 0.327628
R5348 VGND.n2504 VGND.n244 0.327628
R5349 VGND.n2507 VGND.n186 0.327628
R5350 VGND.n2512 VGND.n185 0.327628
R5351 VGND.n2516 VGND.n2515 0.327628
R5352 VGND.n2293 VGND.n2292 0.327628
R5353 VGND.n2289 VGND.n329 0.327628
R5354 VGND.n2284 VGND.n328 0.327628
R5355 VGND.n2279 VGND.n2275 0.327628
R5356 VGND.n2252 VGND.n2251 0.327628
R5357 VGND.n2248 VGND.n2244 0.327628
R5358 VGND.n2226 VGND.n2225 0.327628
R5359 VGND.n2222 VGND.n2218 0.327628
R5360 VGND.n2200 VGND.n2199 0.327628
R5361 VGND.n2196 VGND.n2192 0.327628
R5362 VGND.n2174 VGND.n2173 0.327628
R5363 VGND.n2170 VGND.n2166 0.327628
R5364 VGND.n374 VGND.n373 0.327628
R5365 VGND.n2827 VGND.n182 0.327628
R5366 VGND.n2830 VGND.n180 0.327628
R5367 VGND.n2309 VGND.n324 0.327628
R5368 VGND.n2306 VGND.n2302 0.327628
R5369 VGND.n2266 VGND.n327 0.327628
R5370 VGND.n2270 VGND.n2269 0.327628
R5371 VGND.n2261 VGND.n2257 0.327628
R5372 VGND.n2239 VGND.n2238 0.327628
R5373 VGND.n2235 VGND.n2231 0.327628
R5374 VGND.n2213 VGND.n2212 0.327628
R5375 VGND.n2209 VGND.n2205 0.327628
R5376 VGND.n2187 VGND.n2186 0.327628
R5377 VGND.n2183 VGND.n2179 0.327628
R5378 VGND.n2161 VGND.n2160 0.327628
R5379 VGND.n2157 VGND.n2153 0.327628
R5380 VGND.n1431 VGND.n1430 0.327628
R5381 VGND.n1427 VGND.n1420 0.327628
R5382 VGND.n2129 VGND.n322 0.327628
R5383 VGND.n2134 VGND.n321 0.327628
R5384 VGND.n2138 VGND.n2137 0.327628
R5385 VGND.n1446 VGND.n390 0.327628
R5386 VGND.n1451 VGND.n389 0.327628
R5387 VGND.n1456 VGND.n388 0.327628
R5388 VGND.n1461 VGND.n387 0.327628
R5389 VGND.n1466 VGND.n386 0.327628
R5390 VGND.n1471 VGND.n385 0.327628
R5391 VGND.n1476 VGND.n384 0.327628
R5392 VGND.n1481 VGND.n383 0.327628
R5393 VGND.n1486 VGND.n382 0.327628
R5394 VGND.n1491 VGND.n381 0.327628
R5395 VGND.n1495 VGND.n1494 0.327628
R5396 VGND.n1441 VGND.n1437 0.327628
R5397 VGND.n2118 VGND.n399 0.327628
R5398 VGND.n2115 VGND.n319 0.327628
R5399 VGND.n2110 VGND.n318 0.327628
R5400 VGND.n2105 VGND.n2101 0.327628
R5401 VGND.n2078 VGND.n2077 0.327628
R5402 VGND.n2074 VGND.n2070 0.327628
R5403 VGND.n2052 VGND.n2051 0.327628
R5404 VGND.n2048 VGND.n2044 0.327628
R5405 VGND.n2026 VGND.n2025 0.327628
R5406 VGND.n2022 VGND.n2018 0.327628
R5407 VGND.n2000 VGND.n1999 0.327628
R5408 VGND.n1996 VGND.n1992 0.327628
R5409 VGND.n629 VGND.n628 0.327628
R5410 VGND.n1500 VGND.n619 0.327628
R5411 VGND.n1503 VGND.n617 0.327628
R5412 VGND.n2334 VGND.n312 0.327628
R5413 VGND.n2331 VGND.n2327 0.327628
R5414 VGND.n2092 VGND.n316 0.327628
R5415 VGND.n2096 VGND.n2095 0.327628
R5416 VGND.n2087 VGND.n2083 0.327628
R5417 VGND.n2065 VGND.n2064 0.327628
R5418 VGND.n2061 VGND.n2057 0.327628
R5419 VGND.n2039 VGND.n2038 0.327628
R5420 VGND.n2035 VGND.n2031 0.327628
R5421 VGND.n2013 VGND.n2012 0.327628
R5422 VGND.n2009 VGND.n2005 0.327628
R5423 VGND.n1987 VGND.n1986 0.327628
R5424 VGND.n1983 VGND.n1979 0.327628
R5425 VGND.n655 VGND.n654 0.327628
R5426 VGND.n651 VGND.n644 0.327628
R5427 VGND.n1955 VGND.n310 0.327628
R5428 VGND.n1960 VGND.n309 0.327628
R5429 VGND.n1964 VGND.n1963 0.327628
R5430 VGND.n903 VGND.n446 0.327628
R5431 VGND.n908 VGND.n445 0.327628
R5432 VGND.n913 VGND.n444 0.327628
R5433 VGND.n918 VGND.n443 0.327628
R5434 VGND.n923 VGND.n442 0.327628
R5435 VGND.n928 VGND.n441 0.327628
R5436 VGND.n933 VGND.n440 0.327628
R5437 VGND.n938 VGND.n439 0.327628
R5438 VGND.n943 VGND.n438 0.327628
R5439 VGND.n948 VGND.n437 0.327628
R5440 VGND.n953 VGND.n661 0.327628
R5441 VGND.n958 VGND.n660 0.327628
R5442 VGND.n1944 VGND.n455 0.327628
R5443 VGND.n1941 VGND.n307 0.327628
R5444 VGND.n1936 VGND.n306 0.327628
R5445 VGND.n1931 VGND.n1927 0.327628
R5446 VGND.n1904 VGND.n1903 0.327628
R5447 VGND.n1900 VGND.n1896 0.327628
R5448 VGND.n1878 VGND.n1877 0.327628
R5449 VGND.n1874 VGND.n1870 0.327628
R5450 VGND.n1852 VGND.n1851 0.327628
R5451 VGND.n1848 VGND.n1844 0.327628
R5452 VGND.n1826 VGND.n1825 0.327628
R5453 VGND.n1822 VGND.n1818 0.327628
R5454 VGND.n1403 VGND.n1402 0.327628
R5455 VGND.n1399 VGND.n663 0.327628
R5456 VGND.n1394 VGND.n1390 0.327628
R5457 VGND.n2359 VGND.n300 0.327628
R5458 VGND.n2356 VGND.n2352 0.327628
R5459 VGND.n1918 VGND.n304 0.327628
R5460 VGND.n1922 VGND.n1921 0.327628
R5461 VGND.n1913 VGND.n1909 0.327628
R5462 VGND.n1891 VGND.n1890 0.327628
R5463 VGND.n1887 VGND.n1883 0.327628
R5464 VGND.n1865 VGND.n1864 0.327628
R5465 VGND.n1861 VGND.n1857 0.327628
R5466 VGND.n1839 VGND.n1838 0.327628
R5467 VGND.n1835 VGND.n1831 0.327628
R5468 VGND.n1813 VGND.n1812 0.327628
R5469 VGND.n1809 VGND.n1805 0.327628
R5470 VGND.n1383 VGND.n1382 0.327628
R5471 VGND.n1379 VGND.n1372 0.327628
R5472 VGND.n1781 VGND.n298 0.327628
R5473 VGND.n1786 VGND.n297 0.327628
R5474 VGND.n1790 VGND.n1789 0.327628
R5475 VGND.n1316 VGND.n502 0.327628
R5476 VGND.n1321 VGND.n501 0.327628
R5477 VGND.n1326 VGND.n500 0.327628
R5478 VGND.n1331 VGND.n499 0.327628
R5479 VGND.n1336 VGND.n498 0.327628
R5480 VGND.n1341 VGND.n497 0.327628
R5481 VGND.n1346 VGND.n496 0.327628
R5482 VGND.n1351 VGND.n495 0.327628
R5483 VGND.n1356 VGND.n494 0.327628
R5484 VGND.n1361 VGND.n493 0.327628
R5485 VGND.n1365 VGND.n1364 0.327628
R5486 VGND.n1311 VGND.n1304 0.327628
R5487 VGND.n1770 VGND.n511 0.327628
R5488 VGND.n1767 VGND.n295 0.327628
R5489 VGND.n1762 VGND.n294 0.327628
R5490 VGND.n1757 VGND.n1753 0.327628
R5491 VGND.n1730 VGND.n1729 0.327628
R5492 VGND.n1726 VGND.n1722 0.327628
R5493 VGND.n1704 VGND.n1703 0.327628
R5494 VGND.n1700 VGND.n1696 0.327628
R5495 VGND.n1678 VGND.n1677 0.327628
R5496 VGND.n1674 VGND.n1670 0.327628
R5497 VGND.n1652 VGND.n1651 0.327628
R5498 VGND.n1648 VGND.n1644 0.327628
R5499 VGND.n1525 VGND.n1524 0.327628
R5500 VGND.n1521 VGND.n574 0.327628
R5501 VGND.n1516 VGND.n573 0.327628
R5502 VGND.n2384 VGND.n287 0.327628
R5503 VGND.n2381 VGND.n2377 0.327628
R5504 VGND.n1744 VGND.n291 0.327628
R5505 VGND.n1748 VGND.n1747 0.327628
R5506 VGND.n1739 VGND.n1735 0.327628
R5507 VGND.n1717 VGND.n1716 0.327628
R5508 VGND.n1713 VGND.n1709 0.327628
R5509 VGND.n1691 VGND.n1690 0.327628
R5510 VGND.n1687 VGND.n1683 0.327628
R5511 VGND.n1665 VGND.n1664 0.327628
R5512 VGND.n1661 VGND.n1657 0.327628
R5513 VGND.n1639 VGND.n1638 0.327628
R5514 VGND.n1635 VGND.n1631 0.327628
R5515 VGND.n1540 VGND.n1539 0.327628
R5516 VGND.n1536 VGND.n1532 0.327628
R5517 VGND.n1607 VGND.n283 0.327628
R5518 VGND.n1612 VGND.n282 0.327628
R5519 VGND.n1616 VGND.n1615 0.327628
R5520 VGND.n1599 VGND.n558 0.327628
R5521 VGND.n1594 VGND.n557 0.327628
R5522 VGND.n1589 VGND.n556 0.327628
R5523 VGND.n1584 VGND.n555 0.327628
R5524 VGND.n1579 VGND.n554 0.327628
R5525 VGND.n1574 VGND.n553 0.327628
R5526 VGND.n1569 VGND.n552 0.327628
R5527 VGND.n1564 VGND.n551 0.327628
R5528 VGND.n1559 VGND.n550 0.327628
R5529 VGND.n1554 VGND.n549 0.327628
R5530 VGND.n1549 VGND.n1545 0.327628
R5531 VGND.n1297 VGND.n1296 0.327628
R5532 VGND.n2404 VGND.n279 0.327628
R5533 VGND.n2401 VGND.n2397 0.327628
R5534 VGND.n844 VGND.n713 0.327628
R5535 VGND.n849 VGND.n712 0.327628
R5536 VGND.n854 VGND.n707 0.327628
R5537 VGND.n859 VGND.n706 0.327628
R5538 VGND.n864 VGND.n701 0.327628
R5539 VGND.n869 VGND.n700 0.327628
R5540 VGND.n874 VGND.n695 0.327628
R5541 VGND.n879 VGND.n694 0.327628
R5542 VGND.n884 VGND.n689 0.327628
R5543 VGND.n889 VGND.n688 0.327628
R5544 VGND.n893 VGND.n892 0.327628
R5545 VGND.n839 VGND.n827 0.327628
R5546 VGND.n834 VGND.n826 0.327628
R5547 VGND.n1123 VGND.n1121 0.327628
R5548 VGND.n1130 VGND.n1126 0.327628
R5549 VGND.n1133 VGND.n812 0.327628
R5550 VGND.n1143 VGND.n1139 0.327628
R5551 VGND.n1147 VGND.n1146 0.327628
R5552 VGND.n1162 VGND.n1158 0.327628
R5553 VGND.n1165 VGND.n804 0.327628
R5554 VGND.n1175 VGND.n1171 0.327628
R5555 VGND.n1179 VGND.n1178 0.327628
R5556 VGND.n1194 VGND.n1190 0.327628
R5557 VGND.n1197 VGND.n796 0.327628
R5558 VGND.n1207 VGND.n1203 0.327628
R5559 VGND.n1211 VGND.n1210 0.327628
R5560 VGND.n1226 VGND.n1222 0.327628
R5561 VGND.n1229 VGND.n788 0.327628
R5562 VGND.n783 VGND.n782 0.327628
R5563 VGND.n779 VGND.n716 0.327628
R5564 VGND.n774 VGND.n715 0.327628
R5565 VGND.n769 VGND.n710 0.327628
R5566 VGND.n764 VGND.n709 0.327628
R5567 VGND.n759 VGND.n704 0.327628
R5568 VGND.n754 VGND.n703 0.327628
R5569 VGND.n749 VGND.n698 0.327628
R5570 VGND.n744 VGND.n697 0.327628
R5571 VGND.n739 VGND.n692 0.327628
R5572 VGND.n734 VGND.n691 0.327628
R5573 VGND.n729 VGND.n686 0.327628
R5574 VGND.n724 VGND.n685 0.327628
R5575 VGND.n1285 VGND.n679 0.327628
R5576 VGND.n1288 VGND.n677 0.327628
R5577 VGND.n3023 VGND.n2 0.247202
R5578 VGND.n2919 VGND.n59 0.213567
R5579 VGND.n2952 VGND.n2919 0.213567
R5580 VGND.n2953 VGND.n2952 0.213567
R5581 VGND.n2953 VGND.n28 0.213567
R5582 VGND.n1113 VGND.n1090 0.213567
R5583 VGND.n1090 VGND.n1060 0.213567
R5584 VGND.n1060 VGND.n1029 0.213567
R5585 VGND.n1029 VGND.n998 0.213567
R5586 VGND.n998 VGND.n0 0.213567
R5587 VGND.n3005 VGND.n28 0.2073
R5588 VGND.n1115 VGND.n1114 0.17205
R5589 VGND.n2710 VGND 0.169807
R5590 VGND.n2709 VGND 0.169807
R5591 VGND VGND.n188 0.169807
R5592 VGND.n2816 VGND 0.169807
R5593 VGND.n2815 VGND 0.169807
R5594 VGND.n2810 VGND 0.169807
R5595 VGND.n2809 VGND 0.169807
R5596 VGND.n2804 VGND 0.169807
R5597 VGND.n2803 VGND 0.169807
R5598 VGND.n2798 VGND 0.169807
R5599 VGND.n2797 VGND 0.169807
R5600 VGND.n2792 VGND 0.169807
R5601 VGND.n2791 VGND 0.169807
R5602 VGND.n2786 VGND 0.169807
R5603 VGND.n2785 VGND 0.169807
R5604 VGND VGND.n2712 0.169807
R5605 VGND.n2713 VGND 0.169807
R5606 VGND.n2819 VGND 0.169807
R5607 VGND.n2818 VGND 0.169807
R5608 VGND.n2813 VGND 0.169807
R5609 VGND.n2812 VGND 0.169807
R5610 VGND.n2807 VGND 0.169807
R5611 VGND.n2806 VGND 0.169807
R5612 VGND.n2801 VGND 0.169807
R5613 VGND.n2800 VGND 0.169807
R5614 VGND.n2795 VGND 0.169807
R5615 VGND.n2794 VGND 0.169807
R5616 VGND.n2789 VGND 0.169807
R5617 VGND.n2788 VGND 0.169807
R5618 VGND.n2783 VGND 0.169807
R5619 VGND.n2517 VGND 0.169807
R5620 VGND.n2823 VGND 0.169807
R5621 VGND.n2822 VGND 0.169807
R5622 VGND.n2503 VGND 0.169807
R5623 VGND.n2502 VGND 0.169807
R5624 VGND.n2501 VGND 0.169807
R5625 VGND.n2500 VGND 0.169807
R5626 VGND.n2499 VGND 0.169807
R5627 VGND.n2498 VGND 0.169807
R5628 VGND.n2497 VGND 0.169807
R5629 VGND.n2496 VGND 0.169807
R5630 VGND.n2495 VGND 0.169807
R5631 VGND.n2494 VGND 0.169807
R5632 VGND.n2493 VGND 0.169807
R5633 VGND.n2492 VGND 0.169807
R5634 VGND.n639 VGND 0.169807
R5635 VGND.n2826 VGND 0.169807
R5636 VGND VGND.n375 0.169807
R5637 VGND.n2165 VGND 0.169807
R5638 VGND.n2175 VGND 0.169807
R5639 VGND.n2191 VGND 0.169807
R5640 VGND.n2201 VGND 0.169807
R5641 VGND.n2217 VGND 0.169807
R5642 VGND.n2227 VGND 0.169807
R5643 VGND.n2243 VGND 0.169807
R5644 VGND.n2253 VGND 0.169807
R5645 VGND.n2274 VGND 0.169807
R5646 VGND.n2297 VGND 0.169807
R5647 VGND.n2296 VGND 0.169807
R5648 VGND.n2294 VGND 0.169807
R5649 VGND.n1433 VGND 0.169807
R5650 VGND.n1432 VGND 0.169807
R5651 VGND.n2152 VGND 0.169807
R5652 VGND.n2162 VGND 0.169807
R5653 VGND.n2178 VGND 0.169807
R5654 VGND.n2188 VGND 0.169807
R5655 VGND.n2204 VGND 0.169807
R5656 VGND.n2214 VGND 0.169807
R5657 VGND.n2230 VGND 0.169807
R5658 VGND.n2240 VGND 0.169807
R5659 VGND.n2256 VGND 0.169807
R5660 VGND.n2271 VGND 0.169807
R5661 VGND VGND.n2300 0.169807
R5662 VGND.n2301 VGND 0.169807
R5663 VGND.n2314 VGND 0.169807
R5664 VGND.n1436 VGND 0.169807
R5665 VGND.n1496 VGND 0.169807
R5666 VGND.n2149 VGND 0.169807
R5667 VGND.n2148 VGND 0.169807
R5668 VGND.n2147 VGND 0.169807
R5669 VGND.n2146 VGND 0.169807
R5670 VGND.n2145 VGND 0.169807
R5671 VGND.n2144 VGND 0.169807
R5672 VGND.n2143 VGND 0.169807
R5673 VGND.n2142 VGND 0.169807
R5674 VGND.n2141 VGND 0.169807
R5675 VGND.n2140 VGND 0.169807
R5676 VGND.n2139 VGND 0.169807
R5677 VGND.n2318 VGND 0.169807
R5678 VGND.n2317 VGND 0.169807
R5679 VGND.n1414 VGND 0.169807
R5680 VGND.n1499 VGND 0.169807
R5681 VGND.n630 VGND 0.169807
R5682 VGND.n1991 VGND 0.169807
R5683 VGND.n2001 VGND 0.169807
R5684 VGND.n2017 VGND 0.169807
R5685 VGND.n2027 VGND 0.169807
R5686 VGND.n2043 VGND 0.169807
R5687 VGND.n2053 VGND 0.169807
R5688 VGND.n2069 VGND 0.169807
R5689 VGND.n2079 VGND 0.169807
R5690 VGND.n2100 VGND 0.169807
R5691 VGND.n2322 VGND 0.169807
R5692 VGND.n2321 VGND 0.169807
R5693 VGND.n398 VGND 0.169807
R5694 VGND.n1412 VGND 0.169807
R5695 VGND.n656 VGND 0.169807
R5696 VGND.n1978 VGND 0.169807
R5697 VGND.n1988 VGND 0.169807
R5698 VGND.n2004 VGND 0.169807
R5699 VGND.n2014 VGND 0.169807
R5700 VGND.n2030 VGND 0.169807
R5701 VGND.n2040 VGND 0.169807
R5702 VGND.n2056 VGND 0.169807
R5703 VGND.n2066 VGND 0.169807
R5704 VGND.n2082 VGND 0.169807
R5705 VGND.n2097 VGND 0.169807
R5706 VGND VGND.n2325 0.169807
R5707 VGND.n2326 VGND 0.169807
R5708 VGND.n2339 VGND 0.169807
R5709 VGND.n1409 VGND 0.169807
R5710 VGND.n1408 VGND 0.169807
R5711 VGND.n1975 VGND 0.169807
R5712 VGND.n1974 VGND 0.169807
R5713 VGND.n1973 VGND 0.169807
R5714 VGND.n1972 VGND 0.169807
R5715 VGND.n1971 VGND 0.169807
R5716 VGND.n1970 VGND 0.169807
R5717 VGND.n1969 VGND 0.169807
R5718 VGND.n1968 VGND 0.169807
R5719 VGND.n1967 VGND 0.169807
R5720 VGND.n1966 VGND 0.169807
R5721 VGND.n1965 VGND 0.169807
R5722 VGND.n2343 VGND 0.169807
R5723 VGND.n2342 VGND 0.169807
R5724 VGND.n1389 VGND 0.169807
R5725 VGND.n1405 VGND 0.169807
R5726 VGND.n1404 VGND 0.169807
R5727 VGND.n1817 VGND 0.169807
R5728 VGND.n1827 VGND 0.169807
R5729 VGND.n1843 VGND 0.169807
R5730 VGND.n1853 VGND 0.169807
R5731 VGND.n1869 VGND 0.169807
R5732 VGND.n1879 VGND 0.169807
R5733 VGND.n1895 VGND 0.169807
R5734 VGND.n1905 VGND 0.169807
R5735 VGND.n1926 VGND 0.169807
R5736 VGND.n2347 VGND 0.169807
R5737 VGND.n2346 VGND 0.169807
R5738 VGND.n454 VGND 0.169807
R5739 VGND.n1386 VGND 0.169807
R5740 VGND.n1384 VGND 0.169807
R5741 VGND.n1804 VGND 0.169807
R5742 VGND.n1814 VGND 0.169807
R5743 VGND.n1830 VGND 0.169807
R5744 VGND.n1840 VGND 0.169807
R5745 VGND.n1856 VGND 0.169807
R5746 VGND.n1866 VGND 0.169807
R5747 VGND.n1882 VGND 0.169807
R5748 VGND.n1892 VGND 0.169807
R5749 VGND.n1908 VGND 0.169807
R5750 VGND.n1923 VGND 0.169807
R5751 VGND VGND.n2350 0.169807
R5752 VGND.n2351 VGND 0.169807
R5753 VGND.n2364 VGND 0.169807
R5754 VGND.n1368 VGND 0.169807
R5755 VGND.n1367 VGND 0.169807
R5756 VGND.n1801 VGND 0.169807
R5757 VGND.n1800 VGND 0.169807
R5758 VGND.n1799 VGND 0.169807
R5759 VGND.n1798 VGND 0.169807
R5760 VGND.n1797 VGND 0.169807
R5761 VGND.n1796 VGND 0.169807
R5762 VGND.n1795 VGND 0.169807
R5763 VGND.n1794 VGND 0.169807
R5764 VGND.n1793 VGND 0.169807
R5765 VGND.n1792 VGND 0.169807
R5766 VGND.n1791 VGND 0.169807
R5767 VGND.n2368 VGND 0.169807
R5768 VGND.n2367 VGND 0.169807
R5769 VGND.n1528 VGND 0.169807
R5770 VGND.n1527 VGND 0.169807
R5771 VGND.n1526 VGND 0.169807
R5772 VGND.n1643 VGND 0.169807
R5773 VGND.n1653 VGND 0.169807
R5774 VGND.n1669 VGND 0.169807
R5775 VGND.n1679 VGND 0.169807
R5776 VGND.n1695 VGND 0.169807
R5777 VGND.n1705 VGND 0.169807
R5778 VGND.n1721 VGND 0.169807
R5779 VGND.n1731 VGND 0.169807
R5780 VGND.n1752 VGND 0.169807
R5781 VGND.n2372 VGND 0.169807
R5782 VGND.n2371 VGND 0.169807
R5783 VGND.n510 VGND 0.169807
R5784 VGND.n1531 VGND 0.169807
R5785 VGND.n1541 VGND 0.169807
R5786 VGND.n1630 VGND 0.169807
R5787 VGND.n1640 VGND 0.169807
R5788 VGND.n1656 VGND 0.169807
R5789 VGND.n1666 VGND 0.169807
R5790 VGND.n1682 VGND 0.169807
R5791 VGND.n1692 VGND 0.169807
R5792 VGND.n1708 VGND 0.169807
R5793 VGND.n1718 VGND 0.169807
R5794 VGND.n1734 VGND 0.169807
R5795 VGND.n1749 VGND 0.169807
R5796 VGND VGND.n2375 0.169807
R5797 VGND.n2376 VGND 0.169807
R5798 VGND.n2389 VGND 0.169807
R5799 VGND.n1298 VGND 0.169807
R5800 VGND.n1544 VGND 0.169807
R5801 VGND.n1627 VGND 0.169807
R5802 VGND.n1626 VGND 0.169807
R5803 VGND.n1625 VGND 0.169807
R5804 VGND.n1624 VGND 0.169807
R5805 VGND.n1623 VGND 0.169807
R5806 VGND.n1622 VGND 0.169807
R5807 VGND.n1621 VGND 0.169807
R5808 VGND.n1620 VGND 0.169807
R5809 VGND.n1619 VGND 0.169807
R5810 VGND.n1618 VGND 0.169807
R5811 VGND.n1617 VGND 0.169807
R5812 VGND.n2393 VGND 0.169807
R5813 VGND.n2392 VGND 0.169807
R5814 VGND.n896 VGND 0.169807
R5815 VGND.n895 VGND 0.169807
R5816 VGND.n894 VGND 0.169807
R5817 VGND.n1275 VGND 0.169807
R5818 VGND.n1274 VGND 0.169807
R5819 VGND.n1267 VGND 0.169807
R5820 VGND.n1266 VGND 0.169807
R5821 VGND.n1259 VGND 0.169807
R5822 VGND.n1258 VGND 0.169807
R5823 VGND.n1251 VGND 0.169807
R5824 VGND.n1250 VGND 0.169807
R5825 VGND.n1243 VGND 0.169807
R5826 VGND.n1242 VGND 0.169807
R5827 VGND.n2396 VGND 0.169807
R5828 VGND.n284 VGND 0.169807
R5829 VGND.n1119 VGND 0.169807
R5830 VGND.n1282 VGND 0.169807
R5831 VGND.n1281 VGND 0.169807
R5832 VGND VGND.n687 0.169807
R5833 VGND VGND.n690 0.169807
R5834 VGND VGND.n693 0.169807
R5835 VGND VGND.n696 0.169807
R5836 VGND VGND.n699 0.169807
R5837 VGND VGND.n702 0.169807
R5838 VGND VGND.n705 0.169807
R5839 VGND VGND.n708 0.169807
R5840 VGND VGND.n711 0.169807
R5841 VGND VGND.n714 0.169807
R5842 VGND.n1220 VGND 0.169807
R5843 VGND.n1235 VGND 0.169807
R5844 VGND.n1117 VGND 0.169807
R5845 VGND.n1284 VGND 0.169807
R5846 VGND.n1279 VGND 0.169807
R5847 VGND.n1278 VGND 0.169807
R5848 VGND.n1271 VGND 0.169807
R5849 VGND.n1270 VGND 0.169807
R5850 VGND.n1263 VGND 0.169807
R5851 VGND.n1262 VGND 0.169807
R5852 VGND.n1255 VGND 0.169807
R5853 VGND.n1254 VGND 0.169807
R5854 VGND.n1247 VGND 0.169807
R5855 VGND.n1246 VGND 0.169807
R5856 VGND.n1239 VGND 0.169807
R5857 VGND.n1238 VGND 0.169807
R5858 VGND.n1237 VGND 0.169807
R5859 VGND.n109 VGND 0.159538
R5860 VGND.n2870 VGND 0.159538
R5861 VGND.n2410 VGND.n275 0.154425
R5862 VGND.n2410 VGND.n2409 0.154425
R5863 VGND.n2409 VGND.n276 0.154425
R5864 VGND.n289 VGND.n276 0.154425
R5865 VGND.n1775 VGND.n289 0.154425
R5866 VGND.n1776 VGND.n1775 0.154425
R5867 VGND.n1776 VGND.n302 0.154425
R5868 VGND.n1949 VGND.n302 0.154425
R5869 VGND.n1950 VGND.n1949 0.154425
R5870 VGND.n1950 VGND.n314 0.154425
R5871 VGND.n2123 VGND.n314 0.154425
R5872 VGND.n2124 VGND.n2123 0.154425
R5873 VGND.n2124 VGND.n259 0.154425
R5874 VGND.n2431 VGND.n259 0.154425
R5875 VGND.n2432 VGND.n2431 0.154425
R5876 VGND.n2432 VGND.n29 0.154425
R5877 VGND.n3004 VGND.n29 0.154425
R5878 VGND.n1116 VGND.n1115 0.154425
R5879 VGND.n1116 VGND.n669 0.154425
R5880 VGND.n1299 VGND.n669 0.154425
R5881 VGND.n1300 VGND.n1299 0.154425
R5882 VGND.n1301 VGND.n1300 0.154425
R5883 VGND.n1369 VGND.n1301 0.154425
R5884 VGND.n1387 VGND.n1369 0.154425
R5885 VGND.n1388 VGND.n1387 0.154425
R5886 VGND.n1388 VGND.n641 0.154425
R5887 VGND.n1413 VGND.n641 0.154425
R5888 VGND.n1415 VGND.n1413 0.154425
R5889 VGND.n1416 VGND.n1415 0.154425
R5890 VGND.n1417 VGND.n1416 0.154425
R5891 VGND.n1417 VGND.n237 0.154425
R5892 VGND.n2518 VGND.n237 0.154425
R5893 VGND.n2519 VGND.n2518 0.154425
R5894 VGND.n2520 VGND.n2519 0.154425
R5895 VGND.n1100 VGND.n1094 0.144904
R5896 VGND.n1073 VGND.n1065 0.144904
R5897 VGND.n1011 VGND.n1003 0.144904
R5898 VGND.n1042 VGND.n1034 0.144904
R5899 VGND.n2567 VGND.n2566 0.138284
R5900 VGND.n2655 VGND.n2654 0.13638
R5901 VGND.n2658 VGND.n2647 0.13638
R5902 VGND.n2663 VGND.n2662 0.13638
R5903 VGND.n2666 VGND.n2643 0.13638
R5904 VGND.n2671 VGND.n2670 0.13638
R5905 VGND.n2674 VGND.n2639 0.13638
R5906 VGND.n2679 VGND.n2678 0.13638
R5907 VGND.n2682 VGND.n2635 0.13638
R5908 VGND.n2687 VGND.n2686 0.13638
R5909 VGND.n2690 VGND.n2631 0.13638
R5910 VGND.n2695 VGND.n2694 0.13638
R5911 VGND.n2698 VGND.n2627 0.13638
R5912 VGND.n2703 VGND.n2702 0.13638
R5913 VGND.n2706 VGND.n2572 0.13638
R5914 VGND.n2577 VGND.n2576 0.13638
R5915 VGND.n2781 VGND.n227 0.13638
R5916 VGND.n2778 VGND.n2777 0.13638
R5917 VGND.n2773 VGND.n2772 0.13638
R5918 VGND.n2768 VGND.n2767 0.13638
R5919 VGND.n2763 VGND.n2762 0.13638
R5920 VGND.n2758 VGND.n2757 0.13638
R5921 VGND.n2753 VGND.n2752 0.13638
R5922 VGND.n2748 VGND.n2747 0.13638
R5923 VGND.n2743 VGND.n2742 0.13638
R5924 VGND.n2738 VGND.n2737 0.13638
R5925 VGND.n2733 VGND.n2732 0.13638
R5926 VGND.n2728 VGND.n2727 0.13638
R5927 VGND.n2723 VGND.n2722 0.13638
R5928 VGND.n2718 VGND.n2717 0.13638
R5929 VGND.n234 VGND.n232 0.13638
R5930 VGND.n2487 VGND.n2486 0.13638
R5931 VGND.n2482 VGND.n2481 0.13638
R5932 VGND.n2477 VGND.n2476 0.13638
R5933 VGND.n2472 VGND.n2471 0.13638
R5934 VGND.n2467 VGND.n2466 0.13638
R5935 VGND.n2462 VGND.n2461 0.13638
R5936 VGND.n2457 VGND.n2456 0.13638
R5937 VGND.n2452 VGND.n2451 0.13638
R5938 VGND.n2447 VGND.n2446 0.13638
R5939 VGND.n2442 VGND.n2441 0.13638
R5940 VGND.n2437 VGND.n2436 0.13638
R5941 VGND.n246 VGND.n244 0.13638
R5942 VGND.n2507 VGND.n2506 0.13638
R5943 VGND.n2512 VGND.n2511 0.13638
R5944 VGND.n2515 VGND.n242 0.13638
R5945 VGND.n2292 VGND.n332 0.13638
R5946 VGND.n2289 VGND.n2288 0.13638
R5947 VGND.n2284 VGND.n2283 0.13638
R5948 VGND.n2279 VGND.n2278 0.13638
R5949 VGND.n2251 VGND.n340 0.13638
R5950 VGND.n2248 VGND.n2247 0.13638
R5951 VGND.n2225 VGND.n348 0.13638
R5952 VGND.n2222 VGND.n2221 0.13638
R5953 VGND.n2199 VGND.n356 0.13638
R5954 VGND.n2196 VGND.n2195 0.13638
R5955 VGND.n2173 VGND.n364 0.13638
R5956 VGND.n2170 VGND.n2169 0.13638
R5957 VGND.n373 VGND.n370 0.13638
R5958 VGND.n366 VGND.n182 0.13638
R5959 VGND.n2830 VGND.n2829 0.13638
R5960 VGND.n2310 VGND.n2309 0.13638
R5961 VGND.n2306 VGND.n2305 0.13638
R5962 VGND.n2266 VGND.n2265 0.13638
R5963 VGND.n2269 VGND.n336 0.13638
R5964 VGND.n2261 VGND.n2260 0.13638
R5965 VGND.n2238 VGND.n344 0.13638
R5966 VGND.n2235 VGND.n2234 0.13638
R5967 VGND.n2212 VGND.n352 0.13638
R5968 VGND.n2209 VGND.n2208 0.13638
R5969 VGND.n2186 VGND.n360 0.13638
R5970 VGND.n2183 VGND.n2182 0.13638
R5971 VGND.n2160 VGND.n379 0.13638
R5972 VGND.n2157 VGND.n2156 0.13638
R5973 VGND.n1430 VGND.n1423 0.13638
R5974 VGND.n1427 VGND.n1426 0.13638
R5975 VGND.n2129 VGND.n2128 0.13638
R5976 VGND.n2134 VGND.n2133 0.13638
R5977 VGND.n2137 VGND.n393 0.13638
R5978 VGND.n1446 VGND.n1445 0.13638
R5979 VGND.n1451 VGND.n1450 0.13638
R5980 VGND.n1456 VGND.n1455 0.13638
R5981 VGND.n1461 VGND.n1460 0.13638
R5982 VGND.n1466 VGND.n1465 0.13638
R5983 VGND.n1471 VGND.n1470 0.13638
R5984 VGND.n1476 VGND.n1475 0.13638
R5985 VGND.n1481 VGND.n1480 0.13638
R5986 VGND.n1486 VGND.n1485 0.13638
R5987 VGND.n1491 VGND.n1490 0.13638
R5988 VGND.n1494 VGND.n634 0.13638
R5989 VGND.n1441 VGND.n1440 0.13638
R5990 VGND.n2119 VGND.n2118 0.13638
R5991 VGND.n2115 VGND.n2114 0.13638
R5992 VGND.n2110 VGND.n2109 0.13638
R5993 VGND.n2105 VGND.n2104 0.13638
R5994 VGND.n2077 VGND.n407 0.13638
R5995 VGND.n2074 VGND.n2073 0.13638
R5996 VGND.n2051 VGND.n415 0.13638
R5997 VGND.n2048 VGND.n2047 0.13638
R5998 VGND.n2025 VGND.n423 0.13638
R5999 VGND.n2022 VGND.n2021 0.13638
R6000 VGND.n1999 VGND.n431 0.13638
R6001 VGND.n1996 VGND.n1995 0.13638
R6002 VGND.n628 VGND.n625 0.13638
R6003 VGND.n621 VGND.n619 0.13638
R6004 VGND.n1503 VGND.n1502 0.13638
R6005 VGND.n2335 VGND.n2334 0.13638
R6006 VGND.n2331 VGND.n2330 0.13638
R6007 VGND.n2092 VGND.n2091 0.13638
R6008 VGND.n2095 VGND.n403 0.13638
R6009 VGND.n2087 VGND.n2086 0.13638
R6010 VGND.n2064 VGND.n411 0.13638
R6011 VGND.n2061 VGND.n2060 0.13638
R6012 VGND.n2038 VGND.n419 0.13638
R6013 VGND.n2035 VGND.n2034 0.13638
R6014 VGND.n2012 VGND.n427 0.13638
R6015 VGND.n2009 VGND.n2008 0.13638
R6016 VGND.n1986 VGND.n435 0.13638
R6017 VGND.n1983 VGND.n1982 0.13638
R6018 VGND.n654 VGND.n647 0.13638
R6019 VGND.n651 VGND.n650 0.13638
R6020 VGND.n1955 VGND.n1954 0.13638
R6021 VGND.n1960 VGND.n1959 0.13638
R6022 VGND.n1963 VGND.n449 0.13638
R6023 VGND.n903 VGND.n902 0.13638
R6024 VGND.n908 VGND.n907 0.13638
R6025 VGND.n913 VGND.n912 0.13638
R6026 VGND.n918 VGND.n917 0.13638
R6027 VGND.n923 VGND.n922 0.13638
R6028 VGND.n928 VGND.n927 0.13638
R6029 VGND.n933 VGND.n932 0.13638
R6030 VGND.n938 VGND.n937 0.13638
R6031 VGND.n943 VGND.n942 0.13638
R6032 VGND.n948 VGND.n947 0.13638
R6033 VGND.n953 VGND.n952 0.13638
R6034 VGND.n958 VGND.n957 0.13638
R6035 VGND.n1945 VGND.n1944 0.13638
R6036 VGND.n1941 VGND.n1940 0.13638
R6037 VGND.n1936 VGND.n1935 0.13638
R6038 VGND.n1931 VGND.n1930 0.13638
R6039 VGND.n1903 VGND.n463 0.13638
R6040 VGND.n1900 VGND.n1899 0.13638
R6041 VGND.n1877 VGND.n471 0.13638
R6042 VGND.n1874 VGND.n1873 0.13638
R6043 VGND.n1851 VGND.n479 0.13638
R6044 VGND.n1848 VGND.n1847 0.13638
R6045 VGND.n1825 VGND.n487 0.13638
R6046 VGND.n1822 VGND.n1821 0.13638
R6047 VGND.n1402 VGND.n666 0.13638
R6048 VGND.n1399 VGND.n1398 0.13638
R6049 VGND.n1394 VGND.n1393 0.13638
R6050 VGND.n2360 VGND.n2359 0.13638
R6051 VGND.n2356 VGND.n2355 0.13638
R6052 VGND.n1918 VGND.n1917 0.13638
R6053 VGND.n1921 VGND.n459 0.13638
R6054 VGND.n1913 VGND.n1912 0.13638
R6055 VGND.n1890 VGND.n467 0.13638
R6056 VGND.n1887 VGND.n1886 0.13638
R6057 VGND.n1864 VGND.n475 0.13638
R6058 VGND.n1861 VGND.n1860 0.13638
R6059 VGND.n1838 VGND.n483 0.13638
R6060 VGND.n1835 VGND.n1834 0.13638
R6061 VGND.n1812 VGND.n491 0.13638
R6062 VGND.n1809 VGND.n1808 0.13638
R6063 VGND.n1382 VGND.n1375 0.13638
R6064 VGND.n1379 VGND.n1378 0.13638
R6065 VGND.n1781 VGND.n1780 0.13638
R6066 VGND.n1786 VGND.n1785 0.13638
R6067 VGND.n1789 VGND.n505 0.13638
R6068 VGND.n1316 VGND.n1315 0.13638
R6069 VGND.n1321 VGND.n1320 0.13638
R6070 VGND.n1326 VGND.n1325 0.13638
R6071 VGND.n1331 VGND.n1330 0.13638
R6072 VGND.n1336 VGND.n1335 0.13638
R6073 VGND.n1341 VGND.n1340 0.13638
R6074 VGND.n1346 VGND.n1345 0.13638
R6075 VGND.n1351 VGND.n1350 0.13638
R6076 VGND.n1356 VGND.n1355 0.13638
R6077 VGND.n1361 VGND.n1360 0.13638
R6078 VGND.n1364 VGND.n1307 0.13638
R6079 VGND.n1311 VGND.n1310 0.13638
R6080 VGND.n1771 VGND.n1770 0.13638
R6081 VGND.n1767 VGND.n1766 0.13638
R6082 VGND.n1762 VGND.n1761 0.13638
R6083 VGND.n1757 VGND.n1756 0.13638
R6084 VGND.n1729 VGND.n519 0.13638
R6085 VGND.n1726 VGND.n1725 0.13638
R6086 VGND.n1703 VGND.n527 0.13638
R6087 VGND.n1700 VGND.n1699 0.13638
R6088 VGND.n1677 VGND.n535 0.13638
R6089 VGND.n1674 VGND.n1673 0.13638
R6090 VGND.n1651 VGND.n543 0.13638
R6091 VGND.n1648 VGND.n1647 0.13638
R6092 VGND.n1524 VGND.n577 0.13638
R6093 VGND.n1521 VGND.n1520 0.13638
R6094 VGND.n1516 VGND.n1515 0.13638
R6095 VGND.n2385 VGND.n2384 0.13638
R6096 VGND.n2381 VGND.n2380 0.13638
R6097 VGND.n1744 VGND.n1743 0.13638
R6098 VGND.n1747 VGND.n515 0.13638
R6099 VGND.n1739 VGND.n1738 0.13638
R6100 VGND.n1716 VGND.n523 0.13638
R6101 VGND.n1713 VGND.n1712 0.13638
R6102 VGND.n1690 VGND.n531 0.13638
R6103 VGND.n1687 VGND.n1686 0.13638
R6104 VGND.n1664 VGND.n539 0.13638
R6105 VGND.n1661 VGND.n1660 0.13638
R6106 VGND.n1638 VGND.n547 0.13638
R6107 VGND.n1635 VGND.n1634 0.13638
R6108 VGND.n1539 VGND.n566 0.13638
R6109 VGND.n1536 VGND.n1535 0.13638
R6110 VGND.n1607 VGND.n1606 0.13638
R6111 VGND.n1612 VGND.n1611 0.13638
R6112 VGND.n1615 VGND.n561 0.13638
R6113 VGND.n1599 VGND.n1598 0.13638
R6114 VGND.n1594 VGND.n1593 0.13638
R6115 VGND.n1589 VGND.n1588 0.13638
R6116 VGND.n1584 VGND.n1583 0.13638
R6117 VGND.n1579 VGND.n1578 0.13638
R6118 VGND.n1574 VGND.n1573 0.13638
R6119 VGND.n1569 VGND.n1568 0.13638
R6120 VGND.n1564 VGND.n1563 0.13638
R6121 VGND.n1559 VGND.n1558 0.13638
R6122 VGND.n1554 VGND.n1553 0.13638
R6123 VGND.n1549 VGND.n1548 0.13638
R6124 VGND.n1296 VGND.n674 0.13638
R6125 VGND.n2405 VGND.n2404 0.13638
R6126 VGND.n2401 VGND.n2400 0.13638
R6127 VGND.n844 VGND.n843 0.13638
R6128 VGND.n849 VGND.n848 0.13638
R6129 VGND.n854 VGND.n853 0.13638
R6130 VGND.n859 VGND.n858 0.13638
R6131 VGND.n864 VGND.n863 0.13638
R6132 VGND.n869 VGND.n868 0.13638
R6133 VGND.n874 VGND.n873 0.13638
R6134 VGND.n879 VGND.n878 0.13638
R6135 VGND.n884 VGND.n883 0.13638
R6136 VGND.n889 VGND.n888 0.13638
R6137 VGND.n892 VGND.n830 0.13638
R6138 VGND.n839 VGND.n838 0.13638
R6139 VGND.n834 VGND.n833 0.13638
R6140 VGND.n1124 VGND.n1123 0.13638
R6141 VGND.n1130 VGND.n1129 0.13638
R6142 VGND.n1134 VGND.n1133 0.13638
R6143 VGND.n1143 VGND.n1142 0.13638
R6144 VGND.n1146 VGND.n810 0.13638
R6145 VGND.n1162 VGND.n1161 0.13638
R6146 VGND.n1166 VGND.n1165 0.13638
R6147 VGND.n1175 VGND.n1174 0.13638
R6148 VGND.n1178 VGND.n802 0.13638
R6149 VGND.n1194 VGND.n1193 0.13638
R6150 VGND.n1198 VGND.n1197 0.13638
R6151 VGND.n1207 VGND.n1206 0.13638
R6152 VGND.n1210 VGND.n794 0.13638
R6153 VGND.n1226 VGND.n1225 0.13638
R6154 VGND.n1230 VGND.n1229 0.13638
R6155 VGND.n782 VGND.n719 0.13638
R6156 VGND.n779 VGND.n778 0.13638
R6157 VGND.n774 VGND.n773 0.13638
R6158 VGND.n769 VGND.n768 0.13638
R6159 VGND.n764 VGND.n763 0.13638
R6160 VGND.n759 VGND.n758 0.13638
R6161 VGND.n754 VGND.n753 0.13638
R6162 VGND.n749 VGND.n748 0.13638
R6163 VGND.n744 VGND.n743 0.13638
R6164 VGND.n739 VGND.n738 0.13638
R6165 VGND.n734 VGND.n733 0.13638
R6166 VGND.n729 VGND.n728 0.13638
R6167 VGND.n724 VGND.n723 0.13638
R6168 VGND.n683 VGND.n679 0.13638
R6169 VGND.n1288 VGND.n1287 0.13638
R6170 VGND VGND.n109 0.120838
R6171 VGND.n1108 VGND.n1107 0.120292
R6172 VGND.n1107 VGND.n1106 0.120292
R6173 VGND.n1106 VGND.n1092 0.120292
R6174 VGND.n1102 VGND.n1092 0.120292
R6175 VGND.n1102 VGND.n1101 0.120292
R6176 VGND.n1101 VGND.n1100 0.120292
R6177 VGND.n1086 VGND.n1085 0.120292
R6178 VGND.n1081 VGND.n1080 0.120292
R6179 VGND.n1080 VGND.n1079 0.120292
R6180 VGND.n1079 VGND.n1063 0.120292
R6181 VGND.n1075 VGND.n1063 0.120292
R6182 VGND.n1075 VGND.n1074 0.120292
R6183 VGND.n1074 VGND.n1073 0.120292
R6184 VGND.n143 VGND.n120 0.120292
R6185 VGND.n137 VGND.n120 0.120292
R6186 VGND.n137 VGND.n136 0.120292
R6187 VGND.n136 VGND.n124 0.120292
R6188 VGND.n129 VGND.n124 0.120292
R6189 VGND.n129 VGND.n128 0.120292
R6190 VGND.n128 VGND.n127 0.120292
R6191 VGND.n586 VGND.n583 0.120292
R6192 VGND.n587 VGND.n586 0.120292
R6193 VGND.n611 VGND.n588 0.120292
R6194 VGND.n605 VGND.n588 0.120292
R6195 VGND.n605 VGND.n604 0.120292
R6196 VGND.n604 VGND.n592 0.120292
R6197 VGND.n597 VGND.n592 0.120292
R6198 VGND.n597 VGND.n596 0.120292
R6199 VGND.n596 VGND.n595 0.120292
R6200 VGND.n994 VGND.n993 0.120292
R6201 VGND.n987 VGND.n963 0.120292
R6202 VGND.n982 VGND.n963 0.120292
R6203 VGND.n982 VGND.n981 0.120292
R6204 VGND.n978 VGND.n977 0.120292
R6205 VGND.n977 VGND.n972 0.120292
R6206 VGND.n973 VGND.n972 0.120292
R6207 VGND.n1024 VGND.n1023 0.120292
R6208 VGND.n1019 VGND.n1018 0.120292
R6209 VGND.n1018 VGND.n1017 0.120292
R6210 VGND.n1017 VGND.n1001 0.120292
R6211 VGND.n1013 VGND.n1001 0.120292
R6212 VGND.n1013 VGND.n1012 0.120292
R6213 VGND.n1012 VGND.n1011 0.120292
R6214 VGND.n1055 VGND.n1054 0.120292
R6215 VGND.n1050 VGND.n1049 0.120292
R6216 VGND.n1049 VGND.n1048 0.120292
R6217 VGND.n1048 VGND.n1032 0.120292
R6218 VGND.n1044 VGND.n1032 0.120292
R6219 VGND.n1044 VGND.n1043 0.120292
R6220 VGND.n1043 VGND.n1042 0.120292
R6221 VGND.n173 VGND.n150 0.120292
R6222 VGND.n167 VGND.n150 0.120292
R6223 VGND.n167 VGND.n166 0.120292
R6224 VGND.n166 VGND.n154 0.120292
R6225 VGND.n159 VGND.n154 0.120292
R6226 VGND.n159 VGND.n158 0.120292
R6227 VGND.n158 VGND.n157 0.120292
R6228 VGND.n15 VGND.n11 0.120292
R6229 VGND.n20 VGND.n11 0.120292
R6230 VGND.n21 VGND.n20 0.120292
R6231 VGND.n22 VGND.n21 0.120292
R6232 VGND.n22 VGND.n9 0.120292
R6233 VGND.n26 VGND.n9 0.120292
R6234 VGND.n27 VGND.n26 0.120292
R6235 VGND.n101 VGND.n93 0.120292
R6236 VGND.n102 VGND.n101 0.120292
R6237 VGND.n102 VGND.n87 0.120292
R6238 VGND.n107 VGND.n87 0.120292
R6239 VGND.n108 VGND.n107 0.120292
R6240 VGND.n2860 VGND.n2852 0.120292
R6241 VGND.n2861 VGND.n2860 0.120292
R6242 VGND.n2861 VGND.n2846 0.120292
R6243 VGND.n2866 VGND.n2846 0.120292
R6244 VGND.n2867 VGND.n2866 0.120292
R6245 VGND.n2892 VGND.n2884 0.120292
R6246 VGND.n2893 VGND.n2892 0.120292
R6247 VGND.n2893 VGND.n2878 0.120292
R6248 VGND.n2898 VGND.n2878 0.120292
R6249 VGND.n2899 VGND.n2898 0.120292
R6250 VGND.n2903 VGND.n2900 0.120292
R6251 VGND.n75 VGND.n68 0.120292
R6252 VGND.n76 VGND.n75 0.120292
R6253 VGND.n76 VGND.n63 0.120292
R6254 VGND.n81 VGND.n63 0.120292
R6255 VGND.n82 VGND.n81 0.120292
R6256 VGND.n2918 VGND.n60 0.120292
R6257 VGND.n2933 VGND.n2932 0.120292
R6258 VGND.n2933 VGND.n2925 0.120292
R6259 VGND.n2938 VGND.n2925 0.120292
R6260 VGND.n2939 VGND.n2938 0.120292
R6261 VGND.n2940 VGND.n2939 0.120292
R6262 VGND.n2940 VGND.n2923 0.120292
R6263 VGND.n2944 VGND.n2923 0.120292
R6264 VGND.n2946 VGND.n2920 0.120292
R6265 VGND.n2951 VGND.n2920 0.120292
R6266 VGND.n44 VGND.n38 0.120292
R6267 VGND.n49 VGND.n38 0.120292
R6268 VGND.n50 VGND.n49 0.120292
R6269 VGND.n51 VGND.n50 0.120292
R6270 VGND.n51 VGND.n36 0.120292
R6271 VGND.n55 VGND.n36 0.120292
R6272 VGND.n56 VGND.n55 0.120292
R6273 VGND.n2958 VGND.n2957 0.120292
R6274 VGND.n2957 VGND.n2956 0.120292
R6275 VGND.n2972 VGND.n2966 0.120292
R6276 VGND.n2977 VGND.n2966 0.120292
R6277 VGND.n2978 VGND.n2977 0.120292
R6278 VGND.n2979 VGND.n2978 0.120292
R6279 VGND.n2979 VGND.n2964 0.120292
R6280 VGND.n2983 VGND.n2964 0.120292
R6281 VGND.n2984 VGND.n2983 0.120292
R6282 VGND.n2990 VGND.n2989 0.120292
R6283 VGND.n2989 VGND.n2988 0.120292
R6284 VGND VGND.n2870 0.119536
R6285 VGND.n1094 VGND 0.117202
R6286 VGND.n1065 VGND 0.117202
R6287 VGND.n1003 VGND 0.117202
R6288 VGND.n1034 VGND 0.117202
R6289 VGND.n227 VGND.n226 0.110872
R6290 VGND.n2777 VGND.n2776 0.110872
R6291 VGND.n2772 VGND.n2771 0.110872
R6292 VGND.n2767 VGND.n2766 0.110872
R6293 VGND.n2762 VGND.n2761 0.110872
R6294 VGND.n2757 VGND.n2756 0.110872
R6295 VGND.n2752 VGND.n2751 0.110872
R6296 VGND.n2747 VGND.n2746 0.110872
R6297 VGND.n2742 VGND.n2741 0.110872
R6298 VGND.n2737 VGND.n2736 0.110872
R6299 VGND.n2732 VGND.n2731 0.110872
R6300 VGND.n2727 VGND.n2726 0.110872
R6301 VGND.n2722 VGND.n2721 0.110872
R6302 VGND.n2717 VGND.n2716 0.110872
R6303 VGND.n232 VGND.n231 0.110872
R6304 VGND.n2486 VGND.n2485 0.110872
R6305 VGND.n2481 VGND.n2480 0.110872
R6306 VGND.n2476 VGND.n2475 0.110872
R6307 VGND.n2471 VGND.n2470 0.110872
R6308 VGND.n2466 VGND.n2465 0.110872
R6309 VGND.n2461 VGND.n2460 0.110872
R6310 VGND.n2456 VGND.n2455 0.110872
R6311 VGND.n2451 VGND.n2450 0.110872
R6312 VGND.n2446 VGND.n2445 0.110872
R6313 VGND.n2441 VGND.n2440 0.110872
R6314 VGND.n2436 VGND.n2435 0.110872
R6315 VGND.n247 VGND.n246 0.110872
R6316 VGND.n2506 VGND.n2505 0.110872
R6317 VGND.n2511 VGND.n2510 0.110872
R6318 VGND.n242 VGND.n241 0.110872
R6319 VGND.n332 VGND.n331 0.110872
R6320 VGND.n2288 VGND.n2287 0.110872
R6321 VGND.n2283 VGND.n2282 0.110872
R6322 VGND.n2278 VGND.n2277 0.110872
R6323 VGND.n340 VGND.n339 0.110872
R6324 VGND.n2247 VGND.n2246 0.110872
R6325 VGND.n348 VGND.n347 0.110872
R6326 VGND.n2221 VGND.n2220 0.110872
R6327 VGND.n356 VGND.n355 0.110872
R6328 VGND.n2195 VGND.n2194 0.110872
R6329 VGND.n364 VGND.n363 0.110872
R6330 VGND.n2169 VGND.n2168 0.110872
R6331 VGND.n370 VGND.n369 0.110872
R6332 VGND.n367 VGND.n366 0.110872
R6333 VGND.n2829 VGND.n2828 0.110872
R6334 VGND.n2311 VGND.n2310 0.110872
R6335 VGND.n2305 VGND.n2304 0.110872
R6336 VGND.n2265 VGND.n2264 0.110872
R6337 VGND.n336 VGND.n335 0.110872
R6338 VGND.n2260 VGND.n2259 0.110872
R6339 VGND.n344 VGND.n343 0.110872
R6340 VGND.n2234 VGND.n2233 0.110872
R6341 VGND.n352 VGND.n351 0.110872
R6342 VGND.n2208 VGND.n2207 0.110872
R6343 VGND.n360 VGND.n359 0.110872
R6344 VGND.n2182 VGND.n2181 0.110872
R6345 VGND.n379 VGND.n378 0.110872
R6346 VGND.n2156 VGND.n2155 0.110872
R6347 VGND.n1423 VGND.n1422 0.110872
R6348 VGND.n1426 VGND.n1425 0.110872
R6349 VGND.n2128 VGND.n2127 0.110872
R6350 VGND.n2133 VGND.n2132 0.110872
R6351 VGND.n393 VGND.n392 0.110872
R6352 VGND.n1445 VGND.n1444 0.110872
R6353 VGND.n1450 VGND.n1449 0.110872
R6354 VGND.n1455 VGND.n1454 0.110872
R6355 VGND.n1460 VGND.n1459 0.110872
R6356 VGND.n1465 VGND.n1464 0.110872
R6357 VGND.n1470 VGND.n1469 0.110872
R6358 VGND.n1475 VGND.n1474 0.110872
R6359 VGND.n1480 VGND.n1479 0.110872
R6360 VGND.n1485 VGND.n1484 0.110872
R6361 VGND.n1490 VGND.n1489 0.110872
R6362 VGND.n634 VGND.n633 0.110872
R6363 VGND.n1440 VGND.n1439 0.110872
R6364 VGND.n2120 VGND.n2119 0.110872
R6365 VGND.n2114 VGND.n2113 0.110872
R6366 VGND.n2109 VGND.n2108 0.110872
R6367 VGND.n2104 VGND.n2103 0.110872
R6368 VGND.n407 VGND.n406 0.110872
R6369 VGND.n2073 VGND.n2072 0.110872
R6370 VGND.n415 VGND.n414 0.110872
R6371 VGND.n2047 VGND.n2046 0.110872
R6372 VGND.n423 VGND.n422 0.110872
R6373 VGND.n2021 VGND.n2020 0.110872
R6374 VGND.n431 VGND.n430 0.110872
R6375 VGND.n1995 VGND.n1994 0.110872
R6376 VGND.n625 VGND.n624 0.110872
R6377 VGND.n622 VGND.n621 0.110872
R6378 VGND.n1502 VGND.n1501 0.110872
R6379 VGND.n2336 VGND.n2335 0.110872
R6380 VGND.n2330 VGND.n2329 0.110872
R6381 VGND.n2091 VGND.n2090 0.110872
R6382 VGND.n403 VGND.n402 0.110872
R6383 VGND.n2086 VGND.n2085 0.110872
R6384 VGND.n411 VGND.n410 0.110872
R6385 VGND.n2060 VGND.n2059 0.110872
R6386 VGND.n419 VGND.n418 0.110872
R6387 VGND.n2034 VGND.n2033 0.110872
R6388 VGND.n427 VGND.n426 0.110872
R6389 VGND.n2008 VGND.n2007 0.110872
R6390 VGND.n435 VGND.n434 0.110872
R6391 VGND.n1982 VGND.n1981 0.110872
R6392 VGND.n647 VGND.n646 0.110872
R6393 VGND.n650 VGND.n649 0.110872
R6394 VGND.n1954 VGND.n1953 0.110872
R6395 VGND.n1959 VGND.n1958 0.110872
R6396 VGND.n449 VGND.n448 0.110872
R6397 VGND.n902 VGND.n901 0.110872
R6398 VGND.n907 VGND.n906 0.110872
R6399 VGND.n912 VGND.n911 0.110872
R6400 VGND.n917 VGND.n916 0.110872
R6401 VGND.n922 VGND.n921 0.110872
R6402 VGND.n927 VGND.n926 0.110872
R6403 VGND.n932 VGND.n931 0.110872
R6404 VGND.n937 VGND.n936 0.110872
R6405 VGND.n942 VGND.n941 0.110872
R6406 VGND.n947 VGND.n946 0.110872
R6407 VGND.n952 VGND.n951 0.110872
R6408 VGND.n957 VGND.n956 0.110872
R6409 VGND.n1946 VGND.n1945 0.110872
R6410 VGND.n1940 VGND.n1939 0.110872
R6411 VGND.n1935 VGND.n1934 0.110872
R6412 VGND.n1930 VGND.n1929 0.110872
R6413 VGND.n463 VGND.n462 0.110872
R6414 VGND.n1899 VGND.n1898 0.110872
R6415 VGND.n471 VGND.n470 0.110872
R6416 VGND.n1873 VGND.n1872 0.110872
R6417 VGND.n479 VGND.n478 0.110872
R6418 VGND.n1847 VGND.n1846 0.110872
R6419 VGND.n487 VGND.n486 0.110872
R6420 VGND.n1821 VGND.n1820 0.110872
R6421 VGND.n666 VGND.n665 0.110872
R6422 VGND.n1398 VGND.n1397 0.110872
R6423 VGND.n1393 VGND.n1392 0.110872
R6424 VGND.n2361 VGND.n2360 0.110872
R6425 VGND.n2355 VGND.n2354 0.110872
R6426 VGND.n1917 VGND.n1916 0.110872
R6427 VGND.n459 VGND.n458 0.110872
R6428 VGND.n1912 VGND.n1911 0.110872
R6429 VGND.n467 VGND.n466 0.110872
R6430 VGND.n1886 VGND.n1885 0.110872
R6431 VGND.n475 VGND.n474 0.110872
R6432 VGND.n1860 VGND.n1859 0.110872
R6433 VGND.n483 VGND.n482 0.110872
R6434 VGND.n1834 VGND.n1833 0.110872
R6435 VGND.n491 VGND.n490 0.110872
R6436 VGND.n1808 VGND.n1807 0.110872
R6437 VGND.n1375 VGND.n1374 0.110872
R6438 VGND.n1378 VGND.n1377 0.110872
R6439 VGND.n1780 VGND.n1779 0.110872
R6440 VGND.n1785 VGND.n1784 0.110872
R6441 VGND.n505 VGND.n504 0.110872
R6442 VGND.n1315 VGND.n1314 0.110872
R6443 VGND.n1320 VGND.n1319 0.110872
R6444 VGND.n1325 VGND.n1324 0.110872
R6445 VGND.n1330 VGND.n1329 0.110872
R6446 VGND.n1335 VGND.n1334 0.110872
R6447 VGND.n1340 VGND.n1339 0.110872
R6448 VGND.n1345 VGND.n1344 0.110872
R6449 VGND.n1350 VGND.n1349 0.110872
R6450 VGND.n1355 VGND.n1354 0.110872
R6451 VGND.n1360 VGND.n1359 0.110872
R6452 VGND.n1307 VGND.n1306 0.110872
R6453 VGND.n1310 VGND.n1309 0.110872
R6454 VGND.n1772 VGND.n1771 0.110872
R6455 VGND.n1766 VGND.n1765 0.110872
R6456 VGND.n1761 VGND.n1760 0.110872
R6457 VGND.n1756 VGND.n1755 0.110872
R6458 VGND.n519 VGND.n518 0.110872
R6459 VGND.n1725 VGND.n1724 0.110872
R6460 VGND.n527 VGND.n526 0.110872
R6461 VGND.n1699 VGND.n1698 0.110872
R6462 VGND.n535 VGND.n534 0.110872
R6463 VGND.n1673 VGND.n1672 0.110872
R6464 VGND.n543 VGND.n542 0.110872
R6465 VGND.n1647 VGND.n1646 0.110872
R6466 VGND.n577 VGND.n576 0.110872
R6467 VGND.n1520 VGND.n1519 0.110872
R6468 VGND.n1515 VGND.n1514 0.110872
R6469 VGND.n2386 VGND.n2385 0.110872
R6470 VGND.n2380 VGND.n2379 0.110872
R6471 VGND.n1743 VGND.n1742 0.110872
R6472 VGND.n515 VGND.n514 0.110872
R6473 VGND.n1738 VGND.n1737 0.110872
R6474 VGND.n523 VGND.n522 0.110872
R6475 VGND.n1712 VGND.n1711 0.110872
R6476 VGND.n531 VGND.n530 0.110872
R6477 VGND.n1686 VGND.n1685 0.110872
R6478 VGND.n539 VGND.n538 0.110872
R6479 VGND.n1660 VGND.n1659 0.110872
R6480 VGND.n547 VGND.n546 0.110872
R6481 VGND.n1634 VGND.n1633 0.110872
R6482 VGND.n566 VGND.n565 0.110872
R6483 VGND.n1535 VGND.n1534 0.110872
R6484 VGND.n1606 VGND.n1605 0.110872
R6485 VGND.n1611 VGND.n1610 0.110872
R6486 VGND.n561 VGND.n560 0.110872
R6487 VGND.n1598 VGND.n1597 0.110872
R6488 VGND.n1593 VGND.n1592 0.110872
R6489 VGND.n1588 VGND.n1587 0.110872
R6490 VGND.n1583 VGND.n1582 0.110872
R6491 VGND.n1578 VGND.n1577 0.110872
R6492 VGND.n1573 VGND.n1572 0.110872
R6493 VGND.n1568 VGND.n1567 0.110872
R6494 VGND.n1563 VGND.n1562 0.110872
R6495 VGND.n1558 VGND.n1557 0.110872
R6496 VGND.n1553 VGND.n1552 0.110872
R6497 VGND.n1548 VGND.n1547 0.110872
R6498 VGND.n674 VGND.n673 0.110872
R6499 VGND.n2406 VGND.n2405 0.110872
R6500 VGND.n2400 VGND.n2399 0.110872
R6501 VGND.n843 VGND.n842 0.110872
R6502 VGND.n848 VGND.n847 0.110872
R6503 VGND.n853 VGND.n852 0.110872
R6504 VGND.n858 VGND.n857 0.110872
R6505 VGND.n863 VGND.n862 0.110872
R6506 VGND.n868 VGND.n867 0.110872
R6507 VGND.n873 VGND.n872 0.110872
R6508 VGND.n878 VGND.n877 0.110872
R6509 VGND.n883 VGND.n882 0.110872
R6510 VGND.n888 VGND.n887 0.110872
R6511 VGND.n830 VGND.n829 0.110872
R6512 VGND.n838 VGND.n837 0.110872
R6513 VGND.n833 VGND.n832 0.110872
R6514 VGND.n1125 VGND.n1124 0.110872
R6515 VGND.n1129 VGND.n1128 0.110872
R6516 VGND.n1135 VGND.n1134 0.110872
R6517 VGND.n1142 VGND.n1141 0.110872
R6518 VGND.n810 VGND.n809 0.110872
R6519 VGND.n1161 VGND.n1160 0.110872
R6520 VGND.n1167 VGND.n1166 0.110872
R6521 VGND.n1174 VGND.n1173 0.110872
R6522 VGND.n802 VGND.n801 0.110872
R6523 VGND.n1193 VGND.n1192 0.110872
R6524 VGND.n1199 VGND.n1198 0.110872
R6525 VGND.n1206 VGND.n1205 0.110872
R6526 VGND.n794 VGND.n793 0.110872
R6527 VGND.n1225 VGND.n1224 0.110872
R6528 VGND.n1231 VGND.n1230 0.110872
R6529 VGND.n719 VGND.n718 0.110872
R6530 VGND.n778 VGND.n777 0.110872
R6531 VGND.n773 VGND.n772 0.110872
R6532 VGND.n768 VGND.n767 0.110872
R6533 VGND.n763 VGND.n762 0.110872
R6534 VGND.n758 VGND.n757 0.110872
R6535 VGND.n753 VGND.n752 0.110872
R6536 VGND.n748 VGND.n747 0.110872
R6537 VGND.n743 VGND.n742 0.110872
R6538 VGND.n738 VGND.n737 0.110872
R6539 VGND.n733 VGND.n732 0.110872
R6540 VGND.n728 VGND.n727 0.110872
R6541 VGND.n723 VGND.n722 0.110872
R6542 VGND.n684 VGND.n683 0.110872
R6543 VGND.n1287 VGND.n1286 0.110872
R6544 VGND.n1086 VGND 0.0981562
R6545 VGND.n994 VGND 0.0981562
R6546 VGND.n1055 VGND 0.0981562
R6547 VGND VGND.n143 0.0968542
R6548 VGND VGND.n611 0.0968542
R6549 VGND VGND.n987 0.0968542
R6550 VGND.n1024 VGND 0.0968542
R6551 VGND VGND.n173 0.0968542
R6552 VGND.n15 VGND 0.0968542
R6553 VGND VGND.n2903 0.0968542
R6554 VGND VGND.n60 0.0968542
R6555 VGND.n2932 VGND 0.0968542
R6556 VGND.n44 VGND 0.0968542
R6557 VGND.n2972 VGND 0.0968542
R6558 VGND.n2520 VGND 0.088625
R6559 VGND.n2710 VGND 0.0790114
R6560 VGND VGND.n2709 0.0790114
R6561 VGND VGND.n188 0.0790114
R6562 VGND.n2816 VGND 0.0790114
R6563 VGND VGND.n2815 0.0790114
R6564 VGND.n2810 VGND 0.0790114
R6565 VGND VGND.n2809 0.0790114
R6566 VGND.n2804 VGND 0.0790114
R6567 VGND VGND.n2803 0.0790114
R6568 VGND.n2798 VGND 0.0790114
R6569 VGND VGND.n2797 0.0790114
R6570 VGND.n2792 VGND 0.0790114
R6571 VGND VGND.n2791 0.0790114
R6572 VGND.n2786 VGND 0.0790114
R6573 VGND VGND.n2785 0.0790114
R6574 VGND.n3003 VGND 0.0790114
R6575 VGND.n2712 VGND 0.0790114
R6576 VGND.n2713 VGND 0.0790114
R6577 VGND.n2819 VGND 0.0790114
R6578 VGND VGND.n2818 0.0790114
R6579 VGND.n2813 VGND 0.0790114
R6580 VGND VGND.n2812 0.0790114
R6581 VGND.n2807 VGND 0.0790114
R6582 VGND VGND.n2806 0.0790114
R6583 VGND.n2801 VGND 0.0790114
R6584 VGND VGND.n2800 0.0790114
R6585 VGND.n2795 VGND 0.0790114
R6586 VGND VGND.n2794 0.0790114
R6587 VGND.n2789 VGND 0.0790114
R6588 VGND VGND.n2788 0.0790114
R6589 VGND.n2783 VGND 0.0790114
R6590 VGND.n3001 VGND 0.0790114
R6591 VGND VGND.n2517 0.0790114
R6592 VGND.n2823 VGND 0.0790114
R6593 VGND VGND.n2822 0.0790114
R6594 VGND.n2503 VGND 0.0790114
R6595 VGND VGND.n2502 0.0790114
R6596 VGND VGND.n2501 0.0790114
R6597 VGND VGND.n2500 0.0790114
R6598 VGND VGND.n2499 0.0790114
R6599 VGND VGND.n2498 0.0790114
R6600 VGND VGND.n2497 0.0790114
R6601 VGND VGND.n2496 0.0790114
R6602 VGND VGND.n2495 0.0790114
R6603 VGND VGND.n2494 0.0790114
R6604 VGND VGND.n2493 0.0790114
R6605 VGND VGND.n2492 0.0790114
R6606 VGND VGND.n2491 0.0790114
R6607 VGND.n639 VGND 0.0790114
R6608 VGND.n2826 VGND 0.0790114
R6609 VGND.n375 VGND 0.0790114
R6610 VGND.n2165 VGND 0.0790114
R6611 VGND.n2175 VGND 0.0790114
R6612 VGND.n2191 VGND 0.0790114
R6613 VGND.n2201 VGND 0.0790114
R6614 VGND.n2217 VGND 0.0790114
R6615 VGND.n2227 VGND 0.0790114
R6616 VGND.n2243 VGND 0.0790114
R6617 VGND.n2253 VGND 0.0790114
R6618 VGND.n2274 VGND 0.0790114
R6619 VGND.n2297 VGND 0.0790114
R6620 VGND VGND.n2296 0.0790114
R6621 VGND VGND.n2294 0.0790114
R6622 VGND.n2430 VGND 0.0790114
R6623 VGND.n1433 VGND 0.0790114
R6624 VGND VGND.n1432 0.0790114
R6625 VGND.n2152 VGND 0.0790114
R6626 VGND.n2162 VGND 0.0790114
R6627 VGND.n2178 VGND 0.0790114
R6628 VGND.n2188 VGND 0.0790114
R6629 VGND.n2204 VGND 0.0790114
R6630 VGND.n2214 VGND 0.0790114
R6631 VGND.n2230 VGND 0.0790114
R6632 VGND.n2240 VGND 0.0790114
R6633 VGND.n2256 VGND 0.0790114
R6634 VGND.n2271 VGND 0.0790114
R6635 VGND.n2300 VGND 0.0790114
R6636 VGND.n2301 VGND 0.0790114
R6637 VGND.n2314 VGND 0.0790114
R6638 VGND VGND.n2313 0.0790114
R6639 VGND.n1436 VGND 0.0790114
R6640 VGND.n1496 VGND 0.0790114
R6641 VGND.n2149 VGND 0.0790114
R6642 VGND VGND.n2148 0.0790114
R6643 VGND VGND.n2147 0.0790114
R6644 VGND VGND.n2146 0.0790114
R6645 VGND VGND.n2145 0.0790114
R6646 VGND VGND.n2144 0.0790114
R6647 VGND VGND.n2143 0.0790114
R6648 VGND VGND.n2142 0.0790114
R6649 VGND VGND.n2141 0.0790114
R6650 VGND VGND.n2140 0.0790114
R6651 VGND VGND.n2139 0.0790114
R6652 VGND.n2318 VGND 0.0790114
R6653 VGND VGND.n2317 0.0790114
R6654 VGND.n2125 VGND 0.0790114
R6655 VGND VGND.n1414 0.0790114
R6656 VGND.n1499 VGND 0.0790114
R6657 VGND VGND.n630 0.0790114
R6658 VGND.n1991 VGND 0.0790114
R6659 VGND.n2001 VGND 0.0790114
R6660 VGND.n2017 VGND 0.0790114
R6661 VGND.n2027 VGND 0.0790114
R6662 VGND.n2043 VGND 0.0790114
R6663 VGND.n2053 VGND 0.0790114
R6664 VGND.n2069 VGND 0.0790114
R6665 VGND.n2079 VGND 0.0790114
R6666 VGND.n2100 VGND 0.0790114
R6667 VGND.n2322 VGND 0.0790114
R6668 VGND VGND.n2321 0.0790114
R6669 VGND.n398 VGND 0.0790114
R6670 VGND.n2122 VGND 0.0790114
R6671 VGND VGND.n1412 0.0790114
R6672 VGND VGND.n656 0.0790114
R6673 VGND.n1978 VGND 0.0790114
R6674 VGND.n1988 VGND 0.0790114
R6675 VGND.n2004 VGND 0.0790114
R6676 VGND.n2014 VGND 0.0790114
R6677 VGND.n2030 VGND 0.0790114
R6678 VGND.n2040 VGND 0.0790114
R6679 VGND.n2056 VGND 0.0790114
R6680 VGND.n2066 VGND 0.0790114
R6681 VGND.n2082 VGND 0.0790114
R6682 VGND.n2097 VGND 0.0790114
R6683 VGND.n2325 VGND 0.0790114
R6684 VGND.n2326 VGND 0.0790114
R6685 VGND.n2339 VGND 0.0790114
R6686 VGND VGND.n2338 0.0790114
R6687 VGND.n1409 VGND 0.0790114
R6688 VGND VGND.n1408 0.0790114
R6689 VGND.n1975 VGND 0.0790114
R6690 VGND VGND.n1974 0.0790114
R6691 VGND VGND.n1973 0.0790114
R6692 VGND VGND.n1972 0.0790114
R6693 VGND VGND.n1971 0.0790114
R6694 VGND VGND.n1970 0.0790114
R6695 VGND VGND.n1969 0.0790114
R6696 VGND VGND.n1968 0.0790114
R6697 VGND VGND.n1967 0.0790114
R6698 VGND VGND.n1966 0.0790114
R6699 VGND VGND.n1965 0.0790114
R6700 VGND.n2343 VGND 0.0790114
R6701 VGND VGND.n2342 0.0790114
R6702 VGND.n1951 VGND 0.0790114
R6703 VGND.n1389 VGND 0.0790114
R6704 VGND.n1405 VGND 0.0790114
R6705 VGND VGND.n1404 0.0790114
R6706 VGND.n1817 VGND 0.0790114
R6707 VGND.n1827 VGND 0.0790114
R6708 VGND.n1843 VGND 0.0790114
R6709 VGND.n1853 VGND 0.0790114
R6710 VGND.n1869 VGND 0.0790114
R6711 VGND.n1879 VGND 0.0790114
R6712 VGND.n1895 VGND 0.0790114
R6713 VGND.n1905 VGND 0.0790114
R6714 VGND.n1926 VGND 0.0790114
R6715 VGND.n2347 VGND 0.0790114
R6716 VGND VGND.n2346 0.0790114
R6717 VGND.n454 VGND 0.0790114
R6718 VGND.n1948 VGND 0.0790114
R6719 VGND VGND.n1386 0.0790114
R6720 VGND VGND.n1384 0.0790114
R6721 VGND.n1804 VGND 0.0790114
R6722 VGND.n1814 VGND 0.0790114
R6723 VGND.n1830 VGND 0.0790114
R6724 VGND.n1840 VGND 0.0790114
R6725 VGND.n1856 VGND 0.0790114
R6726 VGND.n1866 VGND 0.0790114
R6727 VGND.n1882 VGND 0.0790114
R6728 VGND.n1892 VGND 0.0790114
R6729 VGND.n1908 VGND 0.0790114
R6730 VGND.n1923 VGND 0.0790114
R6731 VGND.n2350 VGND 0.0790114
R6732 VGND.n2351 VGND 0.0790114
R6733 VGND.n2364 VGND 0.0790114
R6734 VGND VGND.n2363 0.0790114
R6735 VGND VGND.n1368 0.0790114
R6736 VGND VGND.n1367 0.0790114
R6737 VGND.n1801 VGND 0.0790114
R6738 VGND VGND.n1800 0.0790114
R6739 VGND VGND.n1799 0.0790114
R6740 VGND VGND.n1798 0.0790114
R6741 VGND VGND.n1797 0.0790114
R6742 VGND VGND.n1796 0.0790114
R6743 VGND VGND.n1795 0.0790114
R6744 VGND VGND.n1794 0.0790114
R6745 VGND VGND.n1793 0.0790114
R6746 VGND VGND.n1792 0.0790114
R6747 VGND VGND.n1791 0.0790114
R6748 VGND.n2368 VGND 0.0790114
R6749 VGND VGND.n2367 0.0790114
R6750 VGND.n1777 VGND 0.0790114
R6751 VGND.n1528 VGND 0.0790114
R6752 VGND VGND.n1527 0.0790114
R6753 VGND VGND.n1526 0.0790114
R6754 VGND.n1643 VGND 0.0790114
R6755 VGND.n1653 VGND 0.0790114
R6756 VGND.n1669 VGND 0.0790114
R6757 VGND.n1679 VGND 0.0790114
R6758 VGND.n1695 VGND 0.0790114
R6759 VGND.n1705 VGND 0.0790114
R6760 VGND.n1721 VGND 0.0790114
R6761 VGND.n1731 VGND 0.0790114
R6762 VGND.n1752 VGND 0.0790114
R6763 VGND.n2372 VGND 0.0790114
R6764 VGND VGND.n2371 0.0790114
R6765 VGND.n510 VGND 0.0790114
R6766 VGND.n1774 VGND 0.0790114
R6767 VGND.n1531 VGND 0.0790114
R6768 VGND.n1541 VGND 0.0790114
R6769 VGND.n1630 VGND 0.0790114
R6770 VGND.n1640 VGND 0.0790114
R6771 VGND.n1656 VGND 0.0790114
R6772 VGND.n1666 VGND 0.0790114
R6773 VGND.n1682 VGND 0.0790114
R6774 VGND.n1692 VGND 0.0790114
R6775 VGND.n1708 VGND 0.0790114
R6776 VGND.n1718 VGND 0.0790114
R6777 VGND.n1734 VGND 0.0790114
R6778 VGND.n1749 VGND 0.0790114
R6779 VGND.n2375 VGND 0.0790114
R6780 VGND.n2376 VGND 0.0790114
R6781 VGND.n2389 VGND 0.0790114
R6782 VGND VGND.n2388 0.0790114
R6783 VGND VGND.n1298 0.0790114
R6784 VGND.n1544 VGND 0.0790114
R6785 VGND.n1627 VGND 0.0790114
R6786 VGND VGND.n1626 0.0790114
R6787 VGND VGND.n1625 0.0790114
R6788 VGND VGND.n1624 0.0790114
R6789 VGND VGND.n1623 0.0790114
R6790 VGND VGND.n1622 0.0790114
R6791 VGND VGND.n1621 0.0790114
R6792 VGND VGND.n1620 0.0790114
R6793 VGND VGND.n1619 0.0790114
R6794 VGND VGND.n1618 0.0790114
R6795 VGND VGND.n1617 0.0790114
R6796 VGND.n2393 VGND 0.0790114
R6797 VGND VGND.n2392 0.0790114
R6798 VGND.n1603 VGND 0.0790114
R6799 VGND.n896 VGND 0.0790114
R6800 VGND VGND.n895 0.0790114
R6801 VGND VGND.n894 0.0790114
R6802 VGND.n1275 VGND 0.0790114
R6803 VGND VGND.n1274 0.0790114
R6804 VGND.n1267 VGND 0.0790114
R6805 VGND VGND.n1266 0.0790114
R6806 VGND.n1259 VGND 0.0790114
R6807 VGND VGND.n1258 0.0790114
R6808 VGND.n1251 VGND 0.0790114
R6809 VGND VGND.n1250 0.0790114
R6810 VGND.n1243 VGND 0.0790114
R6811 VGND VGND.n1242 0.0790114
R6812 VGND.n2396 VGND 0.0790114
R6813 VGND.n284 VGND 0.0790114
R6814 VGND.n2408 VGND 0.0790114
R6815 VGND.n1119 VGND 0.0790114
R6816 VGND.n1282 VGND 0.0790114
R6817 VGND VGND.n1281 0.0790114
R6818 VGND.n687 VGND 0.0790114
R6819 VGND.n690 VGND 0.0790114
R6820 VGND.n693 VGND 0.0790114
R6821 VGND.n696 VGND 0.0790114
R6822 VGND.n699 VGND 0.0790114
R6823 VGND.n702 VGND 0.0790114
R6824 VGND.n705 VGND 0.0790114
R6825 VGND.n708 VGND 0.0790114
R6826 VGND.n711 VGND 0.0790114
R6827 VGND.n714 VGND 0.0790114
R6828 VGND.n1220 VGND 0.0790114
R6829 VGND.n1235 VGND 0.0790114
R6830 VGND VGND.n1234 0.0790114
R6831 VGND.n1117 VGND 0.0790114
R6832 VGND.n1284 VGND 0.0790114
R6833 VGND.n1279 VGND 0.0790114
R6834 VGND VGND.n1278 0.0790114
R6835 VGND.n1271 VGND 0.0790114
R6836 VGND VGND.n1270 0.0790114
R6837 VGND.n1263 VGND 0.0790114
R6838 VGND VGND.n1262 0.0790114
R6839 VGND.n1255 VGND 0.0790114
R6840 VGND VGND.n1254 0.0790114
R6841 VGND.n1247 VGND 0.0790114
R6842 VGND VGND.n1246 0.0790114
R6843 VGND.n1239 VGND 0.0790114
R6844 VGND VGND.n1238 0.0790114
R6845 VGND VGND.n1237 0.0790114
R6846 VGND.n2411 VGND 0.0790114
R6847 VGND.n3023 VGND.n3022 0.0732323
R6848 VGND.n2654 VGND.n2653 0.0656596
R6849 VGND.n2649 VGND.n2647 0.0656596
R6850 VGND.n2662 VGND.n2661 0.0656596
R6851 VGND.n2645 VGND.n2643 0.0656596
R6852 VGND.n2670 VGND.n2669 0.0656596
R6853 VGND.n2641 VGND.n2639 0.0656596
R6854 VGND.n2678 VGND.n2677 0.0656596
R6855 VGND.n2637 VGND.n2635 0.0656596
R6856 VGND.n2686 VGND.n2685 0.0656596
R6857 VGND.n2633 VGND.n2631 0.0656596
R6858 VGND.n2694 VGND.n2693 0.0656596
R6859 VGND.n2629 VGND.n2627 0.0656596
R6860 VGND.n2702 VGND.n2701 0.0656596
R6861 VGND.n2580 VGND.n2572 0.0656596
R6862 VGND.n2576 VGND.n2571 0.0656596
R6863 VGND.n2564 VGND 0.063
R6864 VGND.n2561 VGND 0.063
R6865 VGND.n2558 VGND 0.063
R6866 VGND.n2555 VGND 0.063
R6867 VGND.n2552 VGND 0.063
R6868 VGND.n2549 VGND 0.063
R6869 VGND.n2546 VGND 0.063
R6870 VGND.n2543 VGND 0.063
R6871 VGND.n2540 VGND 0.063
R6872 VGND.n2537 VGND 0.063
R6873 VGND.n2534 VGND 0.063
R6874 VGND.n2531 VGND 0.063
R6875 VGND.n2528 VGND 0.063
R6876 VGND.n2525 VGND 0.063
R6877 VGND.n2522 VGND 0.063
R6878 VGND.n1108 VGND 0.0603958
R6879 VGND.n1085 VGND 0.0603958
R6880 VGND VGND.n1084 0.0603958
R6881 VGND.n1081 VGND 0.0603958
R6882 VGND.n145 VGND 0.0603958
R6883 VGND VGND.n144 0.0603958
R6884 VGND.n127 VGND 0.0603958
R6885 VGND.n613 VGND 0.0603958
R6886 VGND VGND.n612 0.0603958
R6887 VGND.n595 VGND 0.0603958
R6888 VGND.n989 VGND 0.0603958
R6889 VGND VGND.n988 0.0603958
R6890 VGND.n981 VGND 0.0603958
R6891 VGND.n978 VGND 0.0603958
R6892 VGND.n973 VGND 0.0603958
R6893 VGND.n1023 VGND 0.0603958
R6894 VGND VGND.n1022 0.0603958
R6895 VGND.n1019 VGND 0.0603958
R6896 VGND.n1054 VGND 0.0603958
R6897 VGND VGND.n1053 0.0603958
R6898 VGND.n1050 VGND 0.0603958
R6899 VGND.n175 VGND 0.0603958
R6900 VGND VGND.n174 0.0603958
R6901 VGND.n157 VGND 0.0603958
R6902 VGND VGND.n27 0.0603958
R6903 VGND.n3006 VGND 0.0603958
R6904 VGND.n111 VGND 0.0603958
R6905 VGND VGND.n110 0.0603958
R6906 VGND.n2872 VGND 0.0603958
R6907 VGND VGND.n2871 0.0603958
R6908 VGND.n2905 VGND 0.0603958
R6909 VGND VGND.n2904 0.0603958
R6910 VGND.n2900 VGND 0.0603958
R6911 VGND.n2912 VGND 0.0603958
R6912 VGND.n2913 VGND 0.0603958
R6913 VGND VGND.n2944 0.0603958
R6914 VGND.n2945 VGND 0.0603958
R6915 VGND.n2946 VGND 0.0603958
R6916 VGND VGND.n56 0.0603958
R6917 VGND.n57 VGND 0.0603958
R6918 VGND.n2958 VGND 0.0603958
R6919 VGND VGND.n2984 0.0603958
R6920 VGND.n2985 VGND 0.0603958
R6921 VGND.n2990 VGND 0.0603958
R6922 VGND.n2653 VGND 0.0574853
R6923 VGND.n2649 VGND 0.0574853
R6924 VGND.n2661 VGND 0.0574853
R6925 VGND.n2645 VGND 0.0574853
R6926 VGND.n2669 VGND 0.0574853
R6927 VGND.n2641 VGND 0.0574853
R6928 VGND.n2677 VGND 0.0574853
R6929 VGND.n2637 VGND 0.0574853
R6930 VGND.n2685 VGND 0.0574853
R6931 VGND.n2633 VGND 0.0574853
R6932 VGND.n2693 VGND 0.0574853
R6933 VGND.n2629 VGND 0.0574853
R6934 VGND.n2701 VGND 0.0574853
R6935 VGND.n2580 VGND 0.0574853
R6936 VGND.n2571 VGND 0.0574853
R6937 VGND.n822 VGND 0.0489375
R6938 VGND.n785 VGND 0.0489375
R6939 VGND.n2585 VGND 0.0489375
R6940 VGND.n2582 VGND 0.0489375
R6941 VGND.n2568 VGND 0.0489375
R6942 VGND.n2581 VGND 0.0489375
R6943 VGND.n2620 VGND 0.0489375
R6944 VGND.n2617 VGND 0.0489375
R6945 VGND.n2614 VGND 0.0489375
R6946 VGND.n2611 VGND 0.0489375
R6947 VGND.n2608 VGND 0.0489375
R6948 VGND.n2605 VGND 0.0489375
R6949 VGND.n2602 VGND 0.0489375
R6950 VGND.n2599 VGND 0.0489375
R6951 VGND.n2596 VGND 0.0489375
R6952 VGND.n2593 VGND 0.0489375
R6953 VGND.n2590 VGND 0.0489375
R6954 VGND.n2587 VGND 0.0489375
R6955 VGND.n819 VGND 0.0489375
R6956 VGND.n816 VGND 0.0489375
R6957 VGND.n1136 VGND 0.0489375
R6958 VGND.n807 VGND 0.0489375
R6959 VGND.n805 VGND 0.0489375
R6960 VGND.n1151 VGND 0.0489375
R6961 VGND.n1168 VGND 0.0489375
R6962 VGND.n799 VGND 0.0489375
R6963 VGND.n797 VGND 0.0489375
R6964 VGND.n1183 VGND 0.0489375
R6965 VGND.n1200 VGND 0.0489375
R6966 VGND.n791 VGND 0.0489375
R6967 VGND.n789 VGND 0.0489375
R6968 VGND.n1215 VGND 0.0489375
R6969 VGND VGND.n2574 0.037734
R6970 VGND.n226 VGND 0.037734
R6971 VGND.n2776 VGND 0.037734
R6972 VGND.n2771 VGND 0.037734
R6973 VGND.n2766 VGND 0.037734
R6974 VGND.n2761 VGND 0.037734
R6975 VGND.n2756 VGND 0.037734
R6976 VGND.n2751 VGND 0.037734
R6977 VGND.n2746 VGND 0.037734
R6978 VGND.n2741 VGND 0.037734
R6979 VGND.n2736 VGND 0.037734
R6980 VGND.n2731 VGND 0.037734
R6981 VGND.n2726 VGND 0.037734
R6982 VGND.n2721 VGND 0.037734
R6983 VGND.n2716 VGND 0.037734
R6984 VGND.n231 VGND 0.037734
R6985 VGND VGND.n229 0.037734
R6986 VGND.n2485 VGND 0.037734
R6987 VGND.n2480 VGND 0.037734
R6988 VGND.n2475 VGND 0.037734
R6989 VGND.n2470 VGND 0.037734
R6990 VGND.n2465 VGND 0.037734
R6991 VGND.n2460 VGND 0.037734
R6992 VGND.n2455 VGND 0.037734
R6993 VGND.n2450 VGND 0.037734
R6994 VGND.n2445 VGND 0.037734
R6995 VGND.n2440 VGND 0.037734
R6996 VGND.n2435 VGND 0.037734
R6997 VGND VGND.n247 0.037734
R6998 VGND.n2505 VGND 0.037734
R6999 VGND.n2510 VGND 0.037734
R7000 VGND.n241 VGND 0.037734
R7001 VGND VGND.n239 0.037734
R7002 VGND.n331 VGND 0.037734
R7003 VGND.n2287 VGND 0.037734
R7004 VGND.n2282 VGND 0.037734
R7005 VGND.n2277 VGND 0.037734
R7006 VGND.n339 VGND 0.037734
R7007 VGND.n2246 VGND 0.037734
R7008 VGND.n347 VGND 0.037734
R7009 VGND.n2220 VGND 0.037734
R7010 VGND.n355 VGND 0.037734
R7011 VGND.n2194 VGND 0.037734
R7012 VGND.n363 VGND 0.037734
R7013 VGND.n2168 VGND 0.037734
R7014 VGND.n369 VGND 0.037734
R7015 VGND VGND.n367 0.037734
R7016 VGND.n2828 VGND 0.037734
R7017 VGND VGND.n179 0.037734
R7018 VGND VGND.n2311 0.037734
R7019 VGND.n2304 VGND 0.037734
R7020 VGND.n2264 VGND 0.037734
R7021 VGND.n335 VGND 0.037734
R7022 VGND.n2259 VGND 0.037734
R7023 VGND.n343 VGND 0.037734
R7024 VGND.n2233 VGND 0.037734
R7025 VGND.n351 VGND 0.037734
R7026 VGND.n2207 VGND 0.037734
R7027 VGND.n359 VGND 0.037734
R7028 VGND.n2181 VGND 0.037734
R7029 VGND.n378 VGND 0.037734
R7030 VGND.n2155 VGND 0.037734
R7031 VGND.n1422 VGND 0.037734
R7032 VGND.n1425 VGND 0.037734
R7033 VGND VGND.n1419 0.037734
R7034 VGND.n2127 VGND 0.037734
R7035 VGND.n2132 VGND 0.037734
R7036 VGND.n392 VGND 0.037734
R7037 VGND.n1444 VGND 0.037734
R7038 VGND.n1449 VGND 0.037734
R7039 VGND.n1454 VGND 0.037734
R7040 VGND.n1459 VGND 0.037734
R7041 VGND.n1464 VGND 0.037734
R7042 VGND.n1469 VGND 0.037734
R7043 VGND.n1474 VGND 0.037734
R7044 VGND.n1479 VGND 0.037734
R7045 VGND.n1484 VGND 0.037734
R7046 VGND.n1489 VGND 0.037734
R7047 VGND.n633 VGND 0.037734
R7048 VGND.n1439 VGND 0.037734
R7049 VGND VGND.n637 0.037734
R7050 VGND VGND.n2120 0.037734
R7051 VGND.n2113 VGND 0.037734
R7052 VGND.n2108 VGND 0.037734
R7053 VGND.n2103 VGND 0.037734
R7054 VGND.n406 VGND 0.037734
R7055 VGND.n2072 VGND 0.037734
R7056 VGND.n414 VGND 0.037734
R7057 VGND.n2046 VGND 0.037734
R7058 VGND.n422 VGND 0.037734
R7059 VGND.n2020 VGND 0.037734
R7060 VGND.n430 VGND 0.037734
R7061 VGND.n1994 VGND 0.037734
R7062 VGND.n624 VGND 0.037734
R7063 VGND VGND.n622 0.037734
R7064 VGND.n1501 VGND 0.037734
R7065 VGND VGND.n616 0.037734
R7066 VGND VGND.n2336 0.037734
R7067 VGND.n2329 VGND 0.037734
R7068 VGND.n2090 VGND 0.037734
R7069 VGND.n402 VGND 0.037734
R7070 VGND.n2085 VGND 0.037734
R7071 VGND.n410 VGND 0.037734
R7072 VGND.n2059 VGND 0.037734
R7073 VGND.n418 VGND 0.037734
R7074 VGND.n2033 VGND 0.037734
R7075 VGND.n426 VGND 0.037734
R7076 VGND.n2007 VGND 0.037734
R7077 VGND.n434 VGND 0.037734
R7078 VGND.n1981 VGND 0.037734
R7079 VGND.n646 VGND 0.037734
R7080 VGND.n649 VGND 0.037734
R7081 VGND VGND.n643 0.037734
R7082 VGND.n1953 VGND 0.037734
R7083 VGND.n1958 VGND 0.037734
R7084 VGND.n448 VGND 0.037734
R7085 VGND.n901 VGND 0.037734
R7086 VGND.n906 VGND 0.037734
R7087 VGND.n911 VGND 0.037734
R7088 VGND.n916 VGND 0.037734
R7089 VGND.n921 VGND 0.037734
R7090 VGND.n926 VGND 0.037734
R7091 VGND.n931 VGND 0.037734
R7092 VGND.n936 VGND 0.037734
R7093 VGND.n941 VGND 0.037734
R7094 VGND.n946 VGND 0.037734
R7095 VGND.n951 VGND 0.037734
R7096 VGND.n956 VGND 0.037734
R7097 VGND VGND.n659 0.037734
R7098 VGND VGND.n1946 0.037734
R7099 VGND.n1939 VGND 0.037734
R7100 VGND.n1934 VGND 0.037734
R7101 VGND.n1929 VGND 0.037734
R7102 VGND.n462 VGND 0.037734
R7103 VGND.n1898 VGND 0.037734
R7104 VGND.n470 VGND 0.037734
R7105 VGND.n1872 VGND 0.037734
R7106 VGND.n478 VGND 0.037734
R7107 VGND.n1846 VGND 0.037734
R7108 VGND.n486 VGND 0.037734
R7109 VGND.n1820 VGND 0.037734
R7110 VGND.n665 VGND 0.037734
R7111 VGND.n1397 VGND 0.037734
R7112 VGND.n1392 VGND 0.037734
R7113 VGND VGND.n668 0.037734
R7114 VGND VGND.n2361 0.037734
R7115 VGND.n2354 VGND 0.037734
R7116 VGND.n1916 VGND 0.037734
R7117 VGND.n458 VGND 0.037734
R7118 VGND.n1911 VGND 0.037734
R7119 VGND.n466 VGND 0.037734
R7120 VGND.n1885 VGND 0.037734
R7121 VGND.n474 VGND 0.037734
R7122 VGND.n1859 VGND 0.037734
R7123 VGND.n482 VGND 0.037734
R7124 VGND.n1833 VGND 0.037734
R7125 VGND.n490 VGND 0.037734
R7126 VGND.n1807 VGND 0.037734
R7127 VGND.n1374 VGND 0.037734
R7128 VGND.n1377 VGND 0.037734
R7129 VGND VGND.n1371 0.037734
R7130 VGND.n1779 VGND 0.037734
R7131 VGND.n1784 VGND 0.037734
R7132 VGND.n504 VGND 0.037734
R7133 VGND.n1314 VGND 0.037734
R7134 VGND.n1319 VGND 0.037734
R7135 VGND.n1324 VGND 0.037734
R7136 VGND.n1329 VGND 0.037734
R7137 VGND.n1334 VGND 0.037734
R7138 VGND.n1339 VGND 0.037734
R7139 VGND.n1344 VGND 0.037734
R7140 VGND.n1349 VGND 0.037734
R7141 VGND.n1354 VGND 0.037734
R7142 VGND.n1359 VGND 0.037734
R7143 VGND.n1306 VGND 0.037734
R7144 VGND.n1309 VGND 0.037734
R7145 VGND VGND.n1303 0.037734
R7146 VGND VGND.n1772 0.037734
R7147 VGND.n1765 VGND 0.037734
R7148 VGND.n1760 VGND 0.037734
R7149 VGND.n1755 VGND 0.037734
R7150 VGND.n518 VGND 0.037734
R7151 VGND.n1724 VGND 0.037734
R7152 VGND.n526 VGND 0.037734
R7153 VGND.n1698 VGND 0.037734
R7154 VGND.n534 VGND 0.037734
R7155 VGND.n1672 VGND 0.037734
R7156 VGND.n542 VGND 0.037734
R7157 VGND.n1646 VGND 0.037734
R7158 VGND.n576 VGND 0.037734
R7159 VGND.n1519 VGND 0.037734
R7160 VGND.n1514 VGND 0.037734
R7161 VGND VGND.n572 0.037734
R7162 VGND VGND.n2386 0.037734
R7163 VGND.n2379 VGND 0.037734
R7164 VGND.n1742 VGND 0.037734
R7165 VGND.n514 VGND 0.037734
R7166 VGND.n1737 VGND 0.037734
R7167 VGND.n522 VGND 0.037734
R7168 VGND.n1711 VGND 0.037734
R7169 VGND.n530 VGND 0.037734
R7170 VGND.n1685 VGND 0.037734
R7171 VGND.n538 VGND 0.037734
R7172 VGND.n1659 VGND 0.037734
R7173 VGND.n546 VGND 0.037734
R7174 VGND.n1633 VGND 0.037734
R7175 VGND.n565 VGND 0.037734
R7176 VGND.n1534 VGND 0.037734
R7177 VGND VGND.n568 0.037734
R7178 VGND.n1605 VGND 0.037734
R7179 VGND.n1610 VGND 0.037734
R7180 VGND.n560 VGND 0.037734
R7181 VGND.n1597 VGND 0.037734
R7182 VGND.n1592 VGND 0.037734
R7183 VGND.n1587 VGND 0.037734
R7184 VGND.n1582 VGND 0.037734
R7185 VGND.n1577 VGND 0.037734
R7186 VGND.n1572 VGND 0.037734
R7187 VGND.n1567 VGND 0.037734
R7188 VGND.n1562 VGND 0.037734
R7189 VGND.n1557 VGND 0.037734
R7190 VGND.n1552 VGND 0.037734
R7191 VGND.n1547 VGND 0.037734
R7192 VGND.n673 VGND 0.037734
R7193 VGND VGND.n671 0.037734
R7194 VGND VGND.n2406 0.037734
R7195 VGND.n2399 VGND 0.037734
R7196 VGND.n842 VGND 0.037734
R7197 VGND.n847 VGND 0.037734
R7198 VGND.n852 VGND 0.037734
R7199 VGND.n857 VGND 0.037734
R7200 VGND.n862 VGND 0.037734
R7201 VGND.n867 VGND 0.037734
R7202 VGND.n872 VGND 0.037734
R7203 VGND.n877 VGND 0.037734
R7204 VGND.n882 VGND 0.037734
R7205 VGND.n887 VGND 0.037734
R7206 VGND.n829 VGND 0.037734
R7207 VGND.n837 VGND 0.037734
R7208 VGND.n832 VGND 0.037734
R7209 VGND VGND.n825 0.037734
R7210 VGND VGND.n815 0.037734
R7211 VGND VGND.n1125 0.037734
R7212 VGND.n1128 VGND 0.037734
R7213 VGND VGND.n1135 0.037734
R7214 VGND.n1141 VGND 0.037734
R7215 VGND.n809 VGND 0.037734
R7216 VGND.n1160 VGND 0.037734
R7217 VGND VGND.n1167 0.037734
R7218 VGND.n1173 VGND 0.037734
R7219 VGND.n801 VGND 0.037734
R7220 VGND.n1192 VGND 0.037734
R7221 VGND VGND.n1199 0.037734
R7222 VGND.n1205 VGND 0.037734
R7223 VGND.n793 VGND 0.037734
R7224 VGND.n1224 VGND 0.037734
R7225 VGND VGND.n1231 0.037734
R7226 VGND.n718 VGND 0.037734
R7227 VGND.n777 VGND 0.037734
R7228 VGND.n772 VGND 0.037734
R7229 VGND.n767 VGND 0.037734
R7230 VGND.n762 VGND 0.037734
R7231 VGND.n757 VGND 0.037734
R7232 VGND.n752 VGND 0.037734
R7233 VGND.n747 VGND 0.037734
R7234 VGND.n742 VGND 0.037734
R7235 VGND.n737 VGND 0.037734
R7236 VGND.n732 VGND 0.037734
R7237 VGND.n727 VGND 0.037734
R7238 VGND.n722 VGND 0.037734
R7239 VGND VGND.n684 0.037734
R7240 VGND.n1286 VGND 0.037734
R7241 VGND VGND.n676 0.037734
R7242 VGND.n1112 VGND 0.0343542
R7243 VGND.n1084 VGND 0.0343542
R7244 VGND.n145 VGND 0.0343542
R7245 VGND.n613 VGND 0.0343542
R7246 VGND.n989 VGND 0.0343542
R7247 VGND.n1022 VGND 0.0343542
R7248 VGND.n1053 VGND 0.0343542
R7249 VGND.n175 VGND 0.0343542
R7250 VGND.n3006 VGND 0.0330521
R7251 VGND.n111 VGND 0.0330521
R7252 VGND.n2872 VGND 0.0330521
R7253 VGND.n2905 VGND 0.0330521
R7254 VGND VGND.n2912 0.0330521
R7255 VGND VGND.n2945 0.0330521
R7256 VGND VGND.n57 0.0330521
R7257 VGND VGND.n2985 0.0330521
R7258 VGND.n3005 VGND 0.024
R7259 VGND.n1 VGND 0.024
R7260 VGND.n144 VGND 0.0239375
R7261 VGND.n612 VGND 0.0239375
R7262 VGND.n174 VGND 0.0239375
R7263 VGND.n2904 VGND 0.0239375
R7264 VGND.n2913 VGND 0.0239375
R7265 VGND.n1089 VGND 0.0226354
R7266 VGND VGND.n119 0.0226354
R7267 VGND.n997 VGND 0.0226354
R7268 VGND.n988 VGND 0.0226354
R7269 VGND.n1028 VGND 0.0226354
R7270 VGND VGND.n2918 0.0226354
R7271 VGND.n2956 VGND 0.0226354
R7272 VGND.n2988 VGND 0.0226354
R7273 VGND VGND.n587 0.0213333
R7274 VGND.n993 VGND 0.0213333
R7275 VGND.n1059 VGND 0.0213333
R7276 VGND VGND.n108 0.0213333
R7277 VGND.n110 VGND 0.0213333
R7278 VGND VGND.n2867 0.0213333
R7279 VGND.n2871 VGND 0.0213333
R7280 VGND VGND.n2899 0.0213333
R7281 VGND.n82 VGND 0.0213333
R7282 VGND VGND.n2951 0.0213333
R7283 VGND.n3005 VGND 0.0161667
R7284 VGND.n2575 VGND 0.00980851
R7285 VGND.n3000 VGND 0.00980851
R7286 VGND.n2782 VGND 0.00980851
R7287 VGND VGND.n220 0.00980851
R7288 VGND VGND.n219 0.00980851
R7289 VGND VGND.n214 0.00980851
R7290 VGND VGND.n213 0.00980851
R7291 VGND VGND.n208 0.00980851
R7292 VGND VGND.n207 0.00980851
R7293 VGND VGND.n202 0.00980851
R7294 VGND VGND.n201 0.00980851
R7295 VGND VGND.n196 0.00980851
R7296 VGND VGND.n195 0.00980851
R7297 VGND VGND.n190 0.00980851
R7298 VGND VGND.n189 0.00980851
R7299 VGND.n2714 VGND 0.00980851
R7300 VGND.n235 VGND 0.00980851
R7301 VGND.n2490 VGND 0.00980851
R7302 VGND VGND.n258 0.00980851
R7303 VGND VGND.n257 0.00980851
R7304 VGND VGND.n256 0.00980851
R7305 VGND VGND.n255 0.00980851
R7306 VGND VGND.n254 0.00980851
R7307 VGND VGND.n253 0.00980851
R7308 VGND VGND.n252 0.00980851
R7309 VGND VGND.n251 0.00980851
R7310 VGND VGND.n250 0.00980851
R7311 VGND VGND.n249 0.00980851
R7312 VGND.n248 VGND 0.00980851
R7313 VGND VGND.n2504 0.00980851
R7314 VGND VGND.n186 0.00980851
R7315 VGND VGND.n185 0.00980851
R7316 VGND.n2516 VGND 0.00980851
R7317 VGND.n2429 VGND 0.00980851
R7318 VGND.n2293 VGND 0.00980851
R7319 VGND VGND.n329 0.00980851
R7320 VGND VGND.n328 0.00980851
R7321 VGND.n2275 VGND 0.00980851
R7322 VGND.n2252 VGND 0.00980851
R7323 VGND.n2244 VGND 0.00980851
R7324 VGND.n2226 VGND 0.00980851
R7325 VGND.n2218 VGND 0.00980851
R7326 VGND.n2200 VGND 0.00980851
R7327 VGND.n2192 VGND 0.00980851
R7328 VGND.n2174 VGND 0.00980851
R7329 VGND.n2166 VGND 0.00980851
R7330 VGND.n374 VGND 0.00980851
R7331 VGND VGND.n2827 0.00980851
R7332 VGND.n180 VGND 0.00980851
R7333 VGND.n2312 VGND 0.00980851
R7334 VGND VGND.n324 0.00980851
R7335 VGND.n2302 VGND 0.00980851
R7336 VGND VGND.n327 0.00980851
R7337 VGND.n2270 VGND 0.00980851
R7338 VGND.n2257 VGND 0.00980851
R7339 VGND.n2239 VGND 0.00980851
R7340 VGND.n2231 VGND 0.00980851
R7341 VGND.n2213 VGND 0.00980851
R7342 VGND.n2205 VGND 0.00980851
R7343 VGND.n2187 VGND 0.00980851
R7344 VGND.n2179 VGND 0.00980851
R7345 VGND.n2161 VGND 0.00980851
R7346 VGND.n2153 VGND 0.00980851
R7347 VGND.n1431 VGND 0.00980851
R7348 VGND.n1420 VGND 0.00980851
R7349 VGND VGND.n2126 0.00980851
R7350 VGND VGND.n322 0.00980851
R7351 VGND VGND.n321 0.00980851
R7352 VGND.n2138 VGND 0.00980851
R7353 VGND VGND.n390 0.00980851
R7354 VGND VGND.n389 0.00980851
R7355 VGND VGND.n388 0.00980851
R7356 VGND VGND.n387 0.00980851
R7357 VGND VGND.n386 0.00980851
R7358 VGND VGND.n385 0.00980851
R7359 VGND VGND.n384 0.00980851
R7360 VGND VGND.n383 0.00980851
R7361 VGND VGND.n382 0.00980851
R7362 VGND VGND.n381 0.00980851
R7363 VGND.n1495 VGND 0.00980851
R7364 VGND.n1437 VGND 0.00980851
R7365 VGND.n2121 VGND 0.00980851
R7366 VGND VGND.n399 0.00980851
R7367 VGND VGND.n319 0.00980851
R7368 VGND VGND.n318 0.00980851
R7369 VGND.n2101 VGND 0.00980851
R7370 VGND.n2078 VGND 0.00980851
R7371 VGND.n2070 VGND 0.00980851
R7372 VGND.n2052 VGND 0.00980851
R7373 VGND.n2044 VGND 0.00980851
R7374 VGND.n2026 VGND 0.00980851
R7375 VGND.n2018 VGND 0.00980851
R7376 VGND.n2000 VGND 0.00980851
R7377 VGND.n1992 VGND 0.00980851
R7378 VGND.n629 VGND 0.00980851
R7379 VGND VGND.n1500 0.00980851
R7380 VGND.n617 VGND 0.00980851
R7381 VGND.n2337 VGND 0.00980851
R7382 VGND VGND.n312 0.00980851
R7383 VGND.n2327 VGND 0.00980851
R7384 VGND VGND.n316 0.00980851
R7385 VGND.n2096 VGND 0.00980851
R7386 VGND.n2083 VGND 0.00980851
R7387 VGND.n2065 VGND 0.00980851
R7388 VGND.n2057 VGND 0.00980851
R7389 VGND.n2039 VGND 0.00980851
R7390 VGND.n2031 VGND 0.00980851
R7391 VGND.n2013 VGND 0.00980851
R7392 VGND.n2005 VGND 0.00980851
R7393 VGND.n1987 VGND 0.00980851
R7394 VGND.n1979 VGND 0.00980851
R7395 VGND.n655 VGND 0.00980851
R7396 VGND.n644 VGND 0.00980851
R7397 VGND VGND.n1952 0.00980851
R7398 VGND VGND.n310 0.00980851
R7399 VGND VGND.n309 0.00980851
R7400 VGND.n1964 VGND 0.00980851
R7401 VGND VGND.n446 0.00980851
R7402 VGND VGND.n445 0.00980851
R7403 VGND VGND.n444 0.00980851
R7404 VGND VGND.n443 0.00980851
R7405 VGND VGND.n442 0.00980851
R7406 VGND VGND.n441 0.00980851
R7407 VGND VGND.n440 0.00980851
R7408 VGND VGND.n439 0.00980851
R7409 VGND VGND.n438 0.00980851
R7410 VGND VGND.n437 0.00980851
R7411 VGND VGND.n661 0.00980851
R7412 VGND.n660 VGND 0.00980851
R7413 VGND.n1947 VGND 0.00980851
R7414 VGND VGND.n455 0.00980851
R7415 VGND VGND.n307 0.00980851
R7416 VGND VGND.n306 0.00980851
R7417 VGND.n1927 VGND 0.00980851
R7418 VGND.n1904 VGND 0.00980851
R7419 VGND.n1896 VGND 0.00980851
R7420 VGND.n1878 VGND 0.00980851
R7421 VGND.n1870 VGND 0.00980851
R7422 VGND.n1852 VGND 0.00980851
R7423 VGND.n1844 VGND 0.00980851
R7424 VGND.n1826 VGND 0.00980851
R7425 VGND.n1818 VGND 0.00980851
R7426 VGND.n1403 VGND 0.00980851
R7427 VGND VGND.n663 0.00980851
R7428 VGND.n1390 VGND 0.00980851
R7429 VGND.n2362 VGND 0.00980851
R7430 VGND VGND.n300 0.00980851
R7431 VGND.n2352 VGND 0.00980851
R7432 VGND VGND.n304 0.00980851
R7433 VGND.n1922 VGND 0.00980851
R7434 VGND.n1909 VGND 0.00980851
R7435 VGND.n1891 VGND 0.00980851
R7436 VGND.n1883 VGND 0.00980851
R7437 VGND.n1865 VGND 0.00980851
R7438 VGND.n1857 VGND 0.00980851
R7439 VGND.n1839 VGND 0.00980851
R7440 VGND.n1831 VGND 0.00980851
R7441 VGND.n1813 VGND 0.00980851
R7442 VGND.n1805 VGND 0.00980851
R7443 VGND.n1383 VGND 0.00980851
R7444 VGND.n1372 VGND 0.00980851
R7445 VGND VGND.n1778 0.00980851
R7446 VGND VGND.n298 0.00980851
R7447 VGND VGND.n297 0.00980851
R7448 VGND.n1790 VGND 0.00980851
R7449 VGND VGND.n502 0.00980851
R7450 VGND VGND.n501 0.00980851
R7451 VGND VGND.n500 0.00980851
R7452 VGND VGND.n499 0.00980851
R7453 VGND VGND.n498 0.00980851
R7454 VGND VGND.n497 0.00980851
R7455 VGND VGND.n496 0.00980851
R7456 VGND VGND.n495 0.00980851
R7457 VGND VGND.n494 0.00980851
R7458 VGND VGND.n493 0.00980851
R7459 VGND.n1365 VGND 0.00980851
R7460 VGND.n1304 VGND 0.00980851
R7461 VGND.n1773 VGND 0.00980851
R7462 VGND VGND.n511 0.00980851
R7463 VGND VGND.n295 0.00980851
R7464 VGND VGND.n294 0.00980851
R7465 VGND.n1753 VGND 0.00980851
R7466 VGND.n1730 VGND 0.00980851
R7467 VGND.n1722 VGND 0.00980851
R7468 VGND.n1704 VGND 0.00980851
R7469 VGND.n1696 VGND 0.00980851
R7470 VGND.n1678 VGND 0.00980851
R7471 VGND.n1670 VGND 0.00980851
R7472 VGND.n1652 VGND 0.00980851
R7473 VGND.n1644 VGND 0.00980851
R7474 VGND.n1525 VGND 0.00980851
R7475 VGND VGND.n574 0.00980851
R7476 VGND.n573 VGND 0.00980851
R7477 VGND.n2387 VGND 0.00980851
R7478 VGND VGND.n287 0.00980851
R7479 VGND.n2377 VGND 0.00980851
R7480 VGND VGND.n291 0.00980851
R7481 VGND.n1748 VGND 0.00980851
R7482 VGND.n1735 VGND 0.00980851
R7483 VGND.n1717 VGND 0.00980851
R7484 VGND.n1709 VGND 0.00980851
R7485 VGND.n1691 VGND 0.00980851
R7486 VGND.n1683 VGND 0.00980851
R7487 VGND.n1665 VGND 0.00980851
R7488 VGND.n1657 VGND 0.00980851
R7489 VGND.n1639 VGND 0.00980851
R7490 VGND.n1631 VGND 0.00980851
R7491 VGND.n1540 VGND 0.00980851
R7492 VGND.n1532 VGND 0.00980851
R7493 VGND VGND.n1604 0.00980851
R7494 VGND VGND.n283 0.00980851
R7495 VGND VGND.n282 0.00980851
R7496 VGND.n1616 VGND 0.00980851
R7497 VGND VGND.n558 0.00980851
R7498 VGND VGND.n557 0.00980851
R7499 VGND VGND.n556 0.00980851
R7500 VGND VGND.n555 0.00980851
R7501 VGND VGND.n554 0.00980851
R7502 VGND VGND.n553 0.00980851
R7503 VGND VGND.n552 0.00980851
R7504 VGND VGND.n551 0.00980851
R7505 VGND VGND.n550 0.00980851
R7506 VGND VGND.n549 0.00980851
R7507 VGND.n1545 VGND 0.00980851
R7508 VGND.n1297 VGND 0.00980851
R7509 VGND.n2407 VGND 0.00980851
R7510 VGND VGND.n279 0.00980851
R7511 VGND.n2397 VGND 0.00980851
R7512 VGND VGND.n713 0.00980851
R7513 VGND VGND.n712 0.00980851
R7514 VGND VGND.n707 0.00980851
R7515 VGND VGND.n706 0.00980851
R7516 VGND VGND.n701 0.00980851
R7517 VGND VGND.n700 0.00980851
R7518 VGND VGND.n695 0.00980851
R7519 VGND VGND.n694 0.00980851
R7520 VGND VGND.n689 0.00980851
R7521 VGND VGND.n688 0.00980851
R7522 VGND.n893 VGND 0.00980851
R7523 VGND VGND.n827 0.00980851
R7524 VGND.n826 VGND 0.00980851
R7525 VGND.n1121 VGND 0.00980851
R7526 VGND.n1126 VGND 0.00980851
R7527 VGND VGND.n812 0.00980851
R7528 VGND.n1139 VGND 0.00980851
R7529 VGND.n1147 VGND 0.00980851
R7530 VGND.n1158 VGND 0.00980851
R7531 VGND VGND.n804 0.00980851
R7532 VGND.n1171 VGND 0.00980851
R7533 VGND.n1179 VGND 0.00980851
R7534 VGND.n1190 VGND 0.00980851
R7535 VGND VGND.n796 0.00980851
R7536 VGND.n1203 VGND 0.00980851
R7537 VGND.n1211 VGND 0.00980851
R7538 VGND.n1222 VGND 0.00980851
R7539 VGND VGND.n788 0.00980851
R7540 VGND.n1232 VGND 0.00980851
R7541 VGND.n2412 VGND 0.00980851
R7542 VGND.n783 VGND 0.00980851
R7543 VGND VGND.n716 0.00980851
R7544 VGND VGND.n715 0.00980851
R7545 VGND VGND.n710 0.00980851
R7546 VGND VGND.n709 0.00980851
R7547 VGND VGND.n704 0.00980851
R7548 VGND VGND.n703 0.00980851
R7549 VGND VGND.n698 0.00980851
R7550 VGND VGND.n697 0.00980851
R7551 VGND VGND.n692 0.00980851
R7552 VGND VGND.n691 0.00980851
R7553 VGND VGND.n686 0.00980851
R7554 VGND.n685 VGND 0.00980851
R7555 VGND VGND.n1285 0.00980851
R7556 VGND.n677 VGND 0.00980851
R7557 VGND.n3022 VGND 0.00851991
R7558 VGND.n2653 VGND.n2651 0.00182979
R7559 VGND.n2650 VGND.n2649 0.00182979
R7560 VGND.n2661 VGND.n2659 0.00182979
R7561 VGND.n2646 VGND.n2645 0.00182979
R7562 VGND.n2669 VGND.n2667 0.00182979
R7563 VGND.n2642 VGND.n2641 0.00182979
R7564 VGND.n2677 VGND.n2675 0.00182979
R7565 VGND.n2638 VGND.n2637 0.00182979
R7566 VGND.n2685 VGND.n2683 0.00182979
R7567 VGND.n2634 VGND.n2633 0.00182979
R7568 VGND.n2693 VGND.n2691 0.00182979
R7569 VGND.n2630 VGND.n2629 0.00182979
R7570 VGND.n2701 VGND.n2699 0.00182979
R7571 VGND.n2626 VGND.n2580 0.00182979
R7572 VGND.n2707 VGND.n2571 0.00182979
R7573 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7574 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7575 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7576 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7577 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7578 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7579 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7580 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7581 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7582 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7583 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7584 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7585 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7586 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7587 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7588 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7589 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7590 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7591 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7592 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7593 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7594 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7595 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7596 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7597 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7598 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7599 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7600 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7601 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7602 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7603 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7604 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7605 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7606 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7607 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7608 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7609 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7610 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7611 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7612 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7613 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7614 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7615 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7616 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7617 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7618 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7619 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7620 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7621 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7622 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7623 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7624 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7625 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7626 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7627 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7628 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7629 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7630 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7631 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7632 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7633 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7634 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7635 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7636 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7637 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7638 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7639 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7640 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7641 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7642 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7643 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7644 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7645 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7646 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7647 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7648 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7649 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7650 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7651 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7652 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7653 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7654 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7655 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7656 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7657 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7658 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7659 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7660 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7661 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7662 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7663 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7664 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7665 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7666 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7667 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7668 XThR.Tn[2].n7 XThR.Tn[2].n5 135.249
R7669 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R7670 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R7671 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R7672 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R7673 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R7674 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7675 XThR.Tn[2].n1 XThR.Tn[2].t6 26.5955
R7676 XThR.Tn[2].n1 XThR.Tn[2].t5 26.5955
R7677 XThR.Tn[2].n0 XThR.Tn[2].t7 26.5955
R7678 XThR.Tn[2].n0 XThR.Tn[2].t4 26.5955
R7679 XThR.Tn[2].n3 XThR.Tn[2].t10 24.9236
R7680 XThR.Tn[2].n3 XThR.Tn[2].t11 24.9236
R7681 XThR.Tn[2].n4 XThR.Tn[2].t9 24.9236
R7682 XThR.Tn[2].n4 XThR.Tn[2].t8 24.9236
R7683 XThR.Tn[2].n5 XThR.Tn[2].t1 24.9236
R7684 XThR.Tn[2].n5 XThR.Tn[2].t2 24.9236
R7685 XThR.Tn[2].n6 XThR.Tn[2].t3 24.9236
R7686 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R7687 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7688 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7689 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7690 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7691 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7692 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7693 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7694 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7695 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7696 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7697 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7698 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7699 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7700 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7701 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7702 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7703 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7704 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7705 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7706 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7707 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7708 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7709 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7710 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7711 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7712 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7713 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7714 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7715 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7716 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7717 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7718 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7719 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7720 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7721 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7722 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7723 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7724 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7725 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7726 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7727 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7728 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7729 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7730 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7731 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7732 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7733 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7734 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7735 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7736 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7737 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7738 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7739 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7740 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7741 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7742 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7743 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7744 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7745 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7746 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7747 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7748 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7749 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7750 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7751 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7752 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7753 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7754 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7755 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7756 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7757 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7758 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7759 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7760 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7761 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7762 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7763 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7764 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7765 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7766 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7767 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7768 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7769 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7770 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7771 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7772 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7773 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7774 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7775 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7776 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7777 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7778 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7779 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7780 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7781 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7782 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7783 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7784 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7785 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7786 VPWR.n2837 VPWR.n2823 2618.82
R7787 VPWR.n2835 VPWR.n2829 2618.82
R7788 VPWR.n2853 VPWR.n2823 1916.47
R7789 VPWR.n2828 VPWR.n2827 1916.47
R7790 VPWR.n2827 VPWR.n2821 1916.47
R7791 VPWR.n2829 VPWR.n2822 1916.47
R7792 VPWR.n2852 VPWR.n2824 1912.94
R7793 VPWR.n2849 VPWR.n2843 1560
R7794 VPWR.n2850 VPWR.n2824 1408.24
R7795 VPWR.n2853 VPWR.n2852 1210.59
R7796 VPWR.n2851 VPWR.n2821 1210.59
R7797 VPWR.n2380 VPWR.t148 1005.7
R7798 VPWR.t366 VPWR.n485 1005.7
R7799 VPWR.t215 VPWR.n2210 1005.7
R7800 VPWR.n639 VPWR.t323 1005.7
R7801 VPWR.n2184 VPWR.t49 1005.7
R7802 VPWR.t156 VPWR.n677 1005.7
R7803 VPWR.t116 VPWR.n2014 1005.7
R7804 VPWR.n831 VPWR.t221 1005.7
R7805 VPWR.n1988 VPWR.t41 1005.7
R7806 VPWR.t228 VPWR.n869 1005.7
R7807 VPWR.n447 VPWR.t33 1005.7
R7808 VPWR.t336 VPWR.n1818 1005.7
R7809 VPWR.t318 VPWR.n2406 1005.7
R7810 VPWR.n1023 VPWR.t188 1005.7
R7811 VPWR.t358 VPWR.n293 1005.7
R7812 VPWR.n1792 VPWR.t299 1005.7
R7813 VPWR.n2591 VPWR.t250 1005.7
R7814 VPWR.n1062 VPWR.t134 1005.7
R7815 VPWR.t710 VPWR.n2309 983.14
R7816 VPWR.n2310 VPWR.t841 983.14
R7817 VPWR.t1406 VPWR.n2319 983.14
R7818 VPWR.n2320 VPWR.t1027 983.14
R7819 VPWR.t1567 VPWR.n2329 983.14
R7820 VPWR.n2330 VPWR.t963 983.14
R7821 VPWR.t736 VPWR.n2339 983.14
R7822 VPWR.n2340 VPWR.t858 983.14
R7823 VPWR.t479 VPWR.n2349 983.14
R7824 VPWR.n2350 VPWR.t664 983.14
R7825 VPWR.t1577 VPWR.n2359 983.14
R7826 VPWR.n2360 VPWR.t471 983.14
R7827 VPWR.t453 VPWR.n2369 983.14
R7828 VPWR.n2370 VPWR.t1491 983.14
R7829 VPWR.t694 VPWR.n2379 983.14
R7830 VPWR.n542 VPWR.t1126 983.14
R7831 VPWR.n541 VPWR.t419 983.14
R7832 VPWR.n537 VPWR.t1382 983.14
R7833 VPWR.n533 VPWR.t1057 983.14
R7834 VPWR.n529 VPWR.t827 983.14
R7835 VPWR.n525 VPWR.t708 983.14
R7836 VPWR.n521 VPWR.t716 983.14
R7837 VPWR.n517 VPWR.t1108 983.14
R7838 VPWR.n513 VPWR.t1012 983.14
R7839 VPWR.n509 VPWR.t1832 983.14
R7840 VPWR.n505 VPWR.t1045 983.14
R7841 VPWR.n501 VPWR.t1195 983.14
R7842 VPWR.n497 VPWR.t815 983.14
R7843 VPWR.n493 VPWR.t1466 983.14
R7844 VPWR.n489 VPWR.t622 983.14
R7845 VPWR.n2281 VPWR.t533 983.14
R7846 VPWR.n2280 VPWR.t1597 983.14
R7847 VPWR.n2271 VPWR.t1360 983.14
R7848 VPWR.n2270 VPWR.t1632 983.14
R7849 VPWR.n2261 VPWR.t1513 983.14
R7850 VPWR.n2260 VPWR.t559 983.14
R7851 VPWR.n2251 VPWR.t1800 983.14
R7852 VPWR.n2250 VPWR.t905 983.14
R7853 VPWR.n2241 VPWR.t951 983.14
R7854 VPWR.n2240 VPWR.t612 983.14
R7855 VPWR.n2231 VPWR.t1680 983.14
R7856 VPWR.n2230 VPWR.t1762 983.14
R7857 VPWR.n2221 VPWR.t1700 983.14
R7858 VPWR.n2220 VPWR.t939 983.14
R7859 VPWR.n2211 VPWR.t756 983.14
R7860 VPWR.t1152 VPWR.n582 983.14
R7861 VPWR.t1609 VPWR.n586 983.14
R7862 VPWR.t1374 VPWR.n590 983.14
R7863 VPWR.t1063 VPWR.n594 983.14
R7864 VPWR.t1544 VPWR.n598 983.14
R7865 VPWR.t543 VPWR.n602 983.14
R7866 VPWR.t726 VPWR.n606 983.14
R7867 VPWR.t1018 VPWR.n610 983.14
R7868 VPWR.t1918 VPWR.n614 983.14
R7869 VPWR.t640 VPWR.n618 983.14
R7870 VPWR.t1055 VPWR.n622 983.14
R7871 VPWR.t1181 VPWR.n626 983.14
R7872 VPWR.t922 VPWR.n630 983.14
R7873 VPWR.t680 VPWR.n634 983.14
R7874 VPWR.t628 VPWR.n638 983.14
R7875 VPWR.t1724 VPWR.n2113 983.14
R7876 VPWR.n2114 VPWR.t1583 983.14
R7877 VPWR.t1394 VPWR.n2123 983.14
R7878 VPWR.n2124 VPWR.t802 983.14
R7879 VPWR.t1666 VPWR.n2133 983.14
R7880 VPWR.n2134 VPWR.t591 983.14
R7881 VPWR.t1898 VPWR.n2143 983.14
R7882 VPWR.n2144 VPWR.t577 983.14
R7883 VPWR.t1599 VPWR.n2153 983.14
R7884 VPWR.n2154 VPWR.t1820 983.14
R7885 VPWR.t553 VPWR.n2163 983.14
R7886 VPWR.n2164 VPWR.t1205 983.14
R7887 VPWR.t805 VPWR.n2173 983.14
R7888 VPWR.n2174 VPWR.t997 983.14
R7889 VPWR.t1808 VPWR.n2183 983.14
R7890 VPWR.n734 VPWR.t901 983.14
R7891 VPWR.n733 VPWR.t839 983.14
R7892 VPWR.n729 VPWR.t1408 983.14
R7893 VPWR.n725 VPWR.t1025 983.14
R7894 VPWR.n721 VPWR.t521 983.14
R7895 VPWR.n717 VPWR.t961 983.14
R7896 VPWR.n713 VPWR.t734 983.14
R7897 VPWR.n709 VPWR.t856 983.14
R7898 VPWR.n705 VPWR.t477 983.14
R7899 VPWR.n701 VPWR.t662 983.14
R7900 VPWR.n697 VPWR.t1575 983.14
R7901 VPWR.n693 VPWR.t469 983.14
R7902 VPWR.n689 VPWR.t451 983.14
R7903 VPWR.n685 VPWR.t1784 983.14
R7904 VPWR.n681 VPWR.t692 983.14
R7905 VPWR.n2085 VPWR.t829 983.14
R7906 VPWR.n2084 VPWR.t1521 983.14
R7907 VPWR.n2075 VPWR.t1402 983.14
R7908 VPWR.n2074 VPWR.t1029 983.14
R7909 VPWR.n2065 VPWR.t1573 983.14
R7910 VPWR.n2064 VPWR.t969 983.14
R7911 VPWR.n2055 VPWR.t1894 983.14
R7912 VPWR.n2054 VPWR.t981 983.14
R7913 VPWR.n2045 VPWR.t1118 983.14
R7914 VPWR.n2044 VPWR.t670 983.14
R7915 VPWR.n2035 VPWR.t549 983.14
R7916 VPWR.n2034 VPWR.t1756 983.14
R7917 VPWR.n2025 VPWR.t455 983.14
R7918 VPWR.n2024 VPWR.t1615 983.14
R7919 VPWR.n2015 VPWR.t696 983.14
R7920 VPWR.t531 VPWR.n774 983.14
R7921 VPWR.t1595 VPWR.n778 983.14
R7922 VPWR.t1362 VPWR.n782 983.14
R7923 VPWR.t1628 VPWR.n786 983.14
R7924 VPWR.t1511 VPWR.n790 983.14
R7925 VPWR.t557 VPWR.n794 983.14
R7926 VPWR.t1798 VPWR.n798 983.14
R7927 VPWR.t919 VPWR.n802 983.14
R7928 VPWR.t847 VPWR.n806 983.14
R7929 VPWR.t610 VPWR.n810 983.14
R7930 VPWR.t1213 VPWR.n814 983.14
R7931 VPWR.t1760 VPWR.n818 983.14
R7932 VPWR.t1696 VPWR.n822 983.14
R7933 VPWR.t937 VPWR.n826 983.14
R7934 VPWR.t752 VPWR.n830 983.14
R7935 VPWR.t1726 VPWR.n1917 983.14
R7936 VPWR.n1918 VPWR.t1585 983.14
R7937 VPWR.t1392 VPWR.n1927 983.14
R7938 VPWR.n1928 VPWR.t1851 983.14
R7939 VPWR.t1534 VPWR.n1937 983.14
R7940 VPWR.n1938 VPWR.t593 983.14
R7941 VPWR.t1900 VPWR.n1947 983.14
R7942 VPWR.n1948 VPWR.t864 983.14
R7943 VPWR.t1601 VPWR.n1957 983.14
R7944 VPWR.n1958 VPWR.t1822 983.14
R7945 VPWR.t1471 VPWR.n1967 983.14
R7946 VPWR.n1968 VPWR.t1207 983.14
R7947 VPWR.t807 VPWR.n1977 983.14
R7948 VPWR.n1978 VPWR.t999 983.14
R7949 VPWR.t1810 VPWR.n1987 983.14
R7950 VPWR.n926 VPWR.t529 983.14
R7951 VPWR.n925 VPWR.t1593 983.14
R7952 VPWR.n921 VPWR.t1364 983.14
R7953 VPWR.n917 VPWR.t1626 983.14
R7954 VPWR.n913 VPWR.t1509 983.14
R7955 VPWR.n909 VPWR.t555 983.14
R7956 VPWR.n905 VPWR.t1796 983.14
R7957 VPWR.n901 VPWR.t915 983.14
R7958 VPWR.n897 VPWR.t845 983.14
R7959 VPWR.n893 VPWR.t608 983.14
R7960 VPWR.n889 VPWR.t1211 983.14
R7961 VPWR.n885 VPWR.t1172 983.14
R7962 VPWR.n881 VPWR.t1692 983.14
R7963 VPWR.n877 VPWR.t935 983.14
R7964 VPWR.n873 VPWR.t750 983.14
R7965 VPWR.t1728 VPWR.n390 983.14
R7966 VPWR.t1587 VPWR.n394 983.14
R7967 VPWR.t1390 VPWR.n398 983.14
R7968 VPWR.t1855 VPWR.n402 983.14
R7969 VPWR.t1536 VPWR.n406 983.14
R7970 VPWR.t595 VPWR.n410 983.14
R7971 VPWR.t1902 VPWR.n414 983.14
R7972 VPWR.t866 VPWR.n418 983.14
R7973 VPWR.t1603 VPWR.n422 983.14
R7974 VPWR.t1824 VPWR.n426 983.14
R7975 VPWR.t1473 VPWR.n430 983.14
R7976 VPWR.t1239 VPWR.n434 983.14
R7977 VPWR.t809 VPWR.n438 983.14
R7978 VPWR.t1001 VPWR.n442 983.14
R7979 VPWR.t1814 VPWR.n446 983.14
R7980 VPWR.n1889 VPWR.t1739 983.14
R7981 VPWR.n1888 VPWR.t425 983.14
R7982 VPWR.n1879 VPWR.t1376 983.14
R7983 VPWR.n1878 VPWR.t1061 983.14
R7984 VPWR.n1869 VPWR.t1717 983.14
R7985 VPWR.n1868 VPWR.t539 983.14
R7986 VPWR.n1859 VPWR.t722 983.14
R7987 VPWR.n1858 VPWR.t1016 983.14
R7988 VPWR.n1849 VPWR.t1914 983.14
R7989 VPWR.n1848 VPWR.t638 983.14
R7990 VPWR.n1839 VPWR.t1051 983.14
R7991 VPWR.n1838 VPWR.t1179 983.14
R7992 VPWR.n1829 VPWR.t821 983.14
R7993 VPWR.n1828 VPWR.t678 983.14
R7994 VPWR.n1819 VPWR.t626 983.14
R7995 VPWR.n2477 VPWR.t1154 983.14
R7996 VPWR.n2476 VPWR.t1611 983.14
R7997 VPWR.n2467 VPWR.t1372 983.14
R7998 VPWR.n2466 VPWR.t1067 983.14
R7999 VPWR.n2457 VPWR.t1546 983.14
R8000 VPWR.n2456 VPWR.t545 983.14
R8001 VPWR.n2447 VPWR.t728 983.14
R8002 VPWR.n2446 VPWR.t1020 983.14
R8003 VPWR.n2437 VPWR.t1920 983.14
R8004 VPWR.n2436 VPWR.t642 983.14
R8005 VPWR.n2427 VPWR.t1098 983.14
R8006 VPWR.n2426 VPWR.t1183 983.14
R8007 VPWR.n2417 VPWR.t924 983.14
R8008 VPWR.n2416 VPWR.t682 983.14
R8009 VPWR.n2407 VPWR.t632 983.14
R8010 VPWR.t893 VPWR.n966 983.14
R8011 VPWR.t1084 VPWR.n970 983.14
R8012 VPWR.t1354 VPWR.n974 983.14
R8013 VPWR.t1638 VPWR.n978 983.14
R8014 VPWR.t515 VPWR.n982 983.14
R8015 VPWR.t565 VPWR.n986 983.14
R8016 VPWR.t740 VPWR.n990 983.14
R8017 VPWR.t909 VPWR.n994 983.14
R8018 VPWR.t957 VPWR.n998 983.14
R8019 VPWR.t614 VPWR.n1002 983.14
R8020 VPWR.t1686 VPWR.n1006 983.14
R8021 VPWR.t1764 VPWR.n1010 983.14
R8022 VPWR.t1704 VPWR.n1014 983.14
R8023 VPWR.t1174 VPWR.n1018 983.14
R8024 VPWR.t762 VPWR.n1022 983.14
R8025 VPWR.n350 VPWR.t1128 983.14
R8026 VPWR.n349 VPWR.t421 983.14
R8027 VPWR.n345 VPWR.t1380 983.14
R8028 VPWR.n341 VPWR.t1059 983.14
R8029 VPWR.n337 VPWR.t1713 983.14
R8030 VPWR.n333 VPWR.t535 983.14
R8031 VPWR.n329 VPWR.t718 983.14
R8032 VPWR.n325 VPWR.t1112 983.14
R8033 VPWR.n321 VPWR.t1014 983.14
R8034 VPWR.n317 VPWR.t1834 983.14
R8035 VPWR.n313 VPWR.t1047 983.14
R8036 VPWR.n309 VPWR.t1197 983.14
R8037 VPWR.n305 VPWR.t819 983.14
R8038 VPWR.n301 VPWR.t1468 983.14
R8039 VPWR.n297 VPWR.t624 983.14
R8040 VPWR.t269 VPWR.n1468 983.14
R8041 VPWR.t371 VPWR.n1475 983.14
R8042 VPWR.t142 VPWR.n1481 983.14
R8043 VPWR.t244 VPWR.n1492 983.14
R8044 VPWR.n1493 VPWR.t266 983.14
R8045 VPWR.t17 VPWR.n1506 983.14
R8046 VPWR.n1507 VPWR.t139 983.14
R8047 VPWR.t280 VPWR.n1520 983.14
R8048 VPWR.n1521 VPWR.t296 983.14
R8049 VPWR.n1536 VPWR.t36 983.14
R8050 VPWR.n1535 VPWR.t169 983.14
R8051 VPWR.n1761 VPWR.t210 983.14
R8052 VPWR.n1760 VPWR.t46 983.14
R8053 VPWR.n1749 VPWR.t83 983.14
R8054 VPWR.t191 VPWR.n1791 983.14
R8055 VPWR.t197 VPWR.n2506 983.14
R8056 VPWR.n2507 VPWR.t309 983.14
R8057 VPWR.t74 VPWR.n2518 983.14
R8058 VPWR.n2519 VPWR.t182 983.14
R8059 VPWR.t194 VPWR.n2530 983.14
R8060 VPWR.n2531 VPWR.t350 983.14
R8061 VPWR.t71 VPWR.n2542 983.14
R8062 VPWR.n2543 VPWR.t231 983.14
R8063 VPWR.t247 VPWR.n2554 983.14
R8064 VPWR.n2555 VPWR.t377 983.14
R8065 VPWR.t121 VPWR.n2566 983.14
R8066 VPWR.n2567 VPWR.t151 983.14
R8067 VPWR.t1 VPWR.n2578 983.14
R8068 VPWR.n2579 VPWR.t20 983.14
R8069 VPWR.t145 VPWR.n2590 983.14
R8070 VPWR.n1594 VPWR.t80 983.14
R8071 VPWR.n1593 VPWR.t185 983.14
R8072 VPWR.t347 VPWR.n1182 983.14
R8073 VPWR.t65 VPWR.n1185 983.14
R8074 VPWR.n1220 VPWR.t77 983.14
R8075 VPWR.n1219 VPWR.t236 983.14
R8076 VPWR.n1216 VPWR.t344 983.14
R8077 VPWR.n1213 VPWR.t105 983.14
R8078 VPWR.n1205 VPWR.t131 983.14
R8079 VPWR.n1202 VPWR.t258 983.14
R8080 VPWR.n1199 VPWR.t4 983.14
R8081 VPWR.n1191 VPWR.t25 983.14
R8082 VPWR.n1188 VPWR.t263 983.14
R8083 VPWR.n1740 VPWR.t291 983.14
R8084 VPWR.n1739 VPWR.t11 983.14
R8085 VPWR.n1308 VPWR.t415 877.144
R8086 VPWR.n2723 VPWR.t1319 877.144
R8087 VPWR.n2843 VPWR.n2822 857.648
R8088 VPWR.n1122 VPWR.t313 738.074
R8089 VPWR.n99 VPWR.t53 738.074
R8090 VPWR.n290 VPWR.t1426 738.074
R8091 VPWR.n68 VPWR.t122 738.074
R8092 VPWR.n346 VPWR.t1129 738.074
R8093 VPWR.n98 VPWR.t198 738.074
R8094 VPWR.n963 VPWR.t1411 738.074
R8095 VPWR.n356 VPWR.t1419 738.074
R8096 VPWR.n357 VPWR.t1155 738.074
R8097 VPWR.n318 VPWR.t1113 738.074
R8098 VPWR.n75 VPWR.t232 738.074
R8099 VPWR.n971 VPWR.t1085 738.074
R8100 VPWR.n369 VPWR.t729 738.074
R8101 VPWR.n322 VPWR.t719 738.074
R8102 VPWR.n80 VPWR.t72 738.074
R8103 VPWR.n932 VPWR.t1423 738.074
R8104 VPWR.n933 VPWR.t1740 738.074
R8105 VPWR.n936 VPWR.t426 738.074
R8106 VPWR.n387 VPWR.t1430 738.074
R8107 VPWR.n391 VPWR.t1729 738.074
R8108 VPWR.n395 VPWR.t1588 738.074
R8109 VPWR.n365 VPWR.t1547 738.074
R8110 VPWR.n330 VPWR.t1714 738.074
R8111 VPWR.n86 VPWR.t195 738.074
R8112 VPWR.n937 VPWR.t1377 738.074
R8113 VPWR.n403 VPWR.t1856 738.074
R8114 VPWR.n364 VPWR.t1068 738.074
R8115 VPWR.n334 VPWR.t1060 738.074
R8116 VPWR.n87 VPWR.t183 738.074
R8117 VPWR.n481 VPWR.t1438 738.074
R8118 VPWR.n480 VPWR.t711 738.074
R8119 VPWR.n477 VPWR.t842 738.074
R8120 VPWR.n476 VPWR.t1407 738.074
R8121 VPWR.n472 VPWR.t1568 738.074
R8122 VPWR.n469 VPWR.t964 738.074
R8123 VPWR.n468 VPWR.t737 738.074
R8124 VPWR.n465 VPWR.t859 738.074
R8125 VPWR.n464 VPWR.t480 738.074
R8126 VPWR.n461 VPWR.t665 738.074
R8127 VPWR.n460 VPWR.t1578 738.074
R8128 VPWR.n457 VPWR.t472 738.074
R8129 VPWR.n456 VPWR.t454 738.074
R8130 VPWR.n453 VPWR.t1492 738.074
R8131 VPWR.n452 VPWR.t695 738.074
R8132 VPWR.n473 VPWR.t1028 738.074
R8133 VPWR.n482 VPWR.t1428 738.074
R8134 VPWR.n538 VPWR.t1127 738.074
R8135 VPWR.n534 VPWR.t420 738.074
R8136 VPWR.n530 VPWR.t1383 738.074
R8137 VPWR.n522 VPWR.t828 738.074
R8138 VPWR.n518 VPWR.t709 738.074
R8139 VPWR.n514 VPWR.t717 738.074
R8140 VPWR.n510 VPWR.t1109 738.074
R8141 VPWR.n506 VPWR.t1013 738.074
R8142 VPWR.n502 VPWR.t1833 738.074
R8143 VPWR.n498 VPWR.t1046 738.074
R8144 VPWR.n494 VPWR.t1196 738.074
R8145 VPWR.n490 VPWR.t816 738.074
R8146 VPWR.n486 VPWR.t1467 738.074
R8147 VPWR.n483 VPWR.t623 738.074
R8148 VPWR.n526 VPWR.t1058 738.074
R8149 VPWR.n548 VPWR.t1413 738.074
R8150 VPWR.n549 VPWR.t534 738.074
R8151 VPWR.n552 VPWR.t1598 738.074
R8152 VPWR.n553 VPWR.t1361 738.074
R8153 VPWR.n557 VPWR.t1514 738.074
R8154 VPWR.n560 VPWR.t560 738.074
R8155 VPWR.n561 VPWR.t1801 738.074
R8156 VPWR.n564 VPWR.t906 738.074
R8157 VPWR.n565 VPWR.t952 738.074
R8158 VPWR.n568 VPWR.t613 738.074
R8159 VPWR.n569 VPWR.t1681 738.074
R8160 VPWR.n572 VPWR.t1763 738.074
R8161 VPWR.n573 VPWR.t1701 738.074
R8162 VPWR.n576 VPWR.t940 738.074
R8163 VPWR.n577 VPWR.t757 738.074
R8164 VPWR.n556 VPWR.t1633 738.074
R8165 VPWR.n579 VPWR.t1421 738.074
R8166 VPWR.n583 VPWR.t1153 738.074
R8167 VPWR.n587 VPWR.t1610 738.074
R8168 VPWR.n591 VPWR.t1375 738.074
R8169 VPWR.n599 VPWR.t1545 738.074
R8170 VPWR.n603 VPWR.t544 738.074
R8171 VPWR.n607 VPWR.t727 738.074
R8172 VPWR.n611 VPWR.t1019 738.074
R8173 VPWR.n615 VPWR.t1919 738.074
R8174 VPWR.n619 VPWR.t641 738.074
R8175 VPWR.n623 VPWR.t1056 738.074
R8176 VPWR.n627 VPWR.t1182 738.074
R8177 VPWR.n631 VPWR.t923 738.074
R8178 VPWR.n635 VPWR.t681 738.074
R8179 VPWR.n578 VPWR.t629 738.074
R8180 VPWR.n595 VPWR.t1064 738.074
R8181 VPWR.n673 VPWR.t1434 738.074
R8182 VPWR.n672 VPWR.t1725 738.074
R8183 VPWR.n669 VPWR.t1584 738.074
R8184 VPWR.n668 VPWR.t1395 738.074
R8185 VPWR.n664 VPWR.t1667 738.074
R8186 VPWR.n661 VPWR.t592 738.074
R8187 VPWR.n660 VPWR.t1899 738.074
R8188 VPWR.n657 VPWR.t578 738.074
R8189 VPWR.n656 VPWR.t1600 738.074
R8190 VPWR.n653 VPWR.t1821 738.074
R8191 VPWR.n652 VPWR.t554 738.074
R8192 VPWR.n649 VPWR.t1206 738.074
R8193 VPWR.n648 VPWR.t806 738.074
R8194 VPWR.n645 VPWR.t998 738.074
R8195 VPWR.n644 VPWR.t1809 738.074
R8196 VPWR.n665 VPWR.t803 738.074
R8197 VPWR.n674 VPWR.t1440 738.074
R8198 VPWR.n730 VPWR.t902 738.074
R8199 VPWR.n726 VPWR.t840 738.074
R8200 VPWR.n722 VPWR.t1409 738.074
R8201 VPWR.n714 VPWR.t522 738.074
R8202 VPWR.n710 VPWR.t962 738.074
R8203 VPWR.n706 VPWR.t735 738.074
R8204 VPWR.n702 VPWR.t857 738.074
R8205 VPWR.n698 VPWR.t478 738.074
R8206 VPWR.n694 VPWR.t663 738.074
R8207 VPWR.n690 VPWR.t1576 738.074
R8208 VPWR.n686 VPWR.t470 738.074
R8209 VPWR.n682 VPWR.t452 738.074
R8210 VPWR.n678 VPWR.t1785 738.074
R8211 VPWR.n675 VPWR.t693 738.074
R8212 VPWR.n718 VPWR.t1026 738.074
R8213 VPWR.n740 VPWR.t1436 738.074
R8214 VPWR.n741 VPWR.t830 738.074
R8215 VPWR.n744 VPWR.t1522 738.074
R8216 VPWR.n745 VPWR.t1403 738.074
R8217 VPWR.n749 VPWR.t1574 738.074
R8218 VPWR.n752 VPWR.t970 738.074
R8219 VPWR.n753 VPWR.t1895 738.074
R8220 VPWR.n756 VPWR.t982 738.074
R8221 VPWR.n757 VPWR.t1119 738.074
R8222 VPWR.n760 VPWR.t671 738.074
R8223 VPWR.n761 VPWR.t550 738.074
R8224 VPWR.n764 VPWR.t1757 738.074
R8225 VPWR.n765 VPWR.t456 738.074
R8226 VPWR.n768 VPWR.t1616 738.074
R8227 VPWR.n769 VPWR.t697 738.074
R8228 VPWR.n748 VPWR.t1030 738.074
R8229 VPWR.n771 VPWR.t1415 738.074
R8230 VPWR.n775 VPWR.t532 738.074
R8231 VPWR.n779 VPWR.t1596 738.074
R8232 VPWR.n783 VPWR.t1363 738.074
R8233 VPWR.n791 VPWR.t1512 738.074
R8234 VPWR.n795 VPWR.t558 738.074
R8235 VPWR.n799 VPWR.t1799 738.074
R8236 VPWR.n803 VPWR.t920 738.074
R8237 VPWR.n807 VPWR.t848 738.074
R8238 VPWR.n811 VPWR.t611 738.074
R8239 VPWR.n815 VPWR.t1214 738.074
R8240 VPWR.n819 VPWR.t1761 738.074
R8241 VPWR.n823 VPWR.t1697 738.074
R8242 VPWR.n827 VPWR.t938 738.074
R8243 VPWR.n770 VPWR.t753 738.074
R8244 VPWR.n787 VPWR.t1629 738.074
R8245 VPWR.n865 VPWR.t1432 738.074
R8246 VPWR.n864 VPWR.t1727 738.074
R8247 VPWR.n861 VPWR.t1586 738.074
R8248 VPWR.n860 VPWR.t1393 738.074
R8249 VPWR.n856 VPWR.t1535 738.074
R8250 VPWR.n853 VPWR.t594 738.074
R8251 VPWR.n852 VPWR.t1901 738.074
R8252 VPWR.n849 VPWR.t865 738.074
R8253 VPWR.n848 VPWR.t1602 738.074
R8254 VPWR.n845 VPWR.t1823 738.074
R8255 VPWR.n844 VPWR.t1472 738.074
R8256 VPWR.n841 VPWR.t1208 738.074
R8257 VPWR.n840 VPWR.t808 738.074
R8258 VPWR.n837 VPWR.t1000 738.074
R8259 VPWR.n836 VPWR.t1811 738.074
R8260 VPWR.n857 VPWR.t1852 738.074
R8261 VPWR.n866 VPWR.t1417 738.074
R8262 VPWR.n922 VPWR.t530 738.074
R8263 VPWR.n918 VPWR.t1594 738.074
R8264 VPWR.n914 VPWR.t1365 738.074
R8265 VPWR.n906 VPWR.t1510 738.074
R8266 VPWR.n902 VPWR.t556 738.074
R8267 VPWR.n898 VPWR.t1797 738.074
R8268 VPWR.n894 VPWR.t916 738.074
R8269 VPWR.n890 VPWR.t846 738.074
R8270 VPWR.n886 VPWR.t609 738.074
R8271 VPWR.n882 VPWR.t1212 738.074
R8272 VPWR.n878 VPWR.t1173 738.074
R8273 VPWR.n874 VPWR.t1693 738.074
R8274 VPWR.n870 VPWR.t936 738.074
R8275 VPWR.n867 VPWR.t751 738.074
R8276 VPWR.n910 VPWR.t1627 738.074
R8277 VPWR.n940 VPWR.t1062 738.074
R8278 VPWR.n979 VPWR.t1639 738.074
R8279 VPWR.n1179 VPWR.t66 738.074
R8280 VPWR.n399 VPWR.t1391 738.074
R8281 VPWR.n361 VPWR.t1373 738.074
R8282 VPWR.n338 VPWR.t1381 738.074
R8283 VPWR.n92 VPWR.t75 738.074
R8284 VPWR.n975 VPWR.t1355 738.074
R8285 VPWR.n1183 VPWR.t348 738.074
R8286 VPWR.n941 VPWR.t1718 738.074
R8287 VPWR.n983 VPWR.t516 738.074
R8288 VPWR.n1217 VPWR.t78 738.074
R8289 VPWR.n407 VPWR.t1537 738.074
R8290 VPWR.n415 VPWR.t1903 738.074
R8291 VPWR.n419 VPWR.t867 738.074
R8292 VPWR.n423 VPWR.t1604 738.074
R8293 VPWR.n427 VPWR.t1825 738.074
R8294 VPWR.n431 VPWR.t1474 738.074
R8295 VPWR.n435 VPWR.t1240 738.074
R8296 VPWR.n439 VPWR.t810 738.074
R8297 VPWR.n443 VPWR.t1002 738.074
R8298 VPWR.n386 VPWR.t1815 738.074
R8299 VPWR.n411 VPWR.t596 738.074
R8300 VPWR.n368 VPWR.t546 738.074
R8301 VPWR.n326 VPWR.t536 738.074
R8302 VPWR.n81 VPWR.t351 738.074
R8303 VPWR.n987 VPWR.t566 738.074
R8304 VPWR.n1214 VPWR.t237 738.074
R8305 VPWR.n944 VPWR.t540 738.074
R8306 VPWR.n948 VPWR.t1017 738.074
R8307 VPWR.n949 VPWR.t1915 738.074
R8308 VPWR.n952 VPWR.t639 738.074
R8309 VPWR.n953 VPWR.t1052 738.074
R8310 VPWR.n956 VPWR.t1180 738.074
R8311 VPWR.n957 VPWR.t822 738.074
R8312 VPWR.n960 VPWR.t679 738.074
R8313 VPWR.n961 VPWR.t627 738.074
R8314 VPWR.n945 VPWR.t723 738.074
R8315 VPWR.n991 VPWR.t741 738.074
R8316 VPWR.n1206 VPWR.t345 738.074
R8317 VPWR.n360 VPWR.t1612 738.074
R8318 VPWR.n342 VPWR.t422 738.074
R8319 VPWR.n93 VPWR.t310 738.074
R8320 VPWR.n1180 VPWR.t186 738.074
R8321 VPWR.n995 VPWR.t910 738.074
R8322 VPWR.n1203 VPWR.t106 738.074
R8323 VPWR.n372 VPWR.t1021 738.074
R8324 VPWR.n376 VPWR.t643 738.074
R8325 VPWR.n377 VPWR.t1099 738.074
R8326 VPWR.n380 VPWR.t1184 738.074
R8327 VPWR.n381 VPWR.t925 738.074
R8328 VPWR.n384 VPWR.t683 738.074
R8329 VPWR.n385 VPWR.t633 738.074
R8330 VPWR.n373 VPWR.t1921 738.074
R8331 VPWR.n314 VPWR.t1015 738.074
R8332 VPWR.n74 VPWR.t248 738.074
R8333 VPWR.n1200 VPWR.t132 738.074
R8334 VPWR.n999 VPWR.t958 738.074
R8335 VPWR.n1003 VPWR.t615 738.074
R8336 VPWR.n1007 VPWR.t1687 738.074
R8337 VPWR.n1011 VPWR.t1765 738.074
R8338 VPWR.n1015 VPWR.t1705 738.074
R8339 VPWR.n1019 VPWR.t1175 738.074
R8340 VPWR.n962 VPWR.t763 738.074
R8341 VPWR.n967 VPWR.t894 738.074
R8342 VPWR.n1123 VPWR.t81 738.074
R8343 VPWR.n310 VPWR.t1835 738.074
R8344 VPWR.n69 VPWR.t378 738.074
R8345 VPWR.n1192 VPWR.t259 738.074
R8346 VPWR.n1189 VPWR.t5 738.074
R8347 VPWR.n306 VPWR.t1048 738.074
R8348 VPWR.n302 VPWR.t1198 738.074
R8349 VPWR.n294 VPWR.t1469 738.074
R8350 VPWR.n291 VPWR.t625 738.074
R8351 VPWR.n298 VPWR.t820 738.074
R8352 VPWR.n1058 VPWR.t264 738.074
R8353 VPWR.n1186 VPWR.t26 738.074
R8354 VPWR.n63 VPWR.t152 738.074
R8355 VPWR.n62 VPWR.t2 738.074
R8356 VPWR.n57 VPWR.t21 738.074
R8357 VPWR.n56 VPWR.t146 738.074
R8358 VPWR.n1059 VPWR.t292 738.074
R8359 VPWR.n1061 VPWR.t12 738.074
R8360 VPWR.n2856 VPWR.n2821 702.354
R8361 VPWR.n2856 VPWR.n2822 702.354
R8362 VPWR.n2854 VPWR.n2853 702.354
R8363 VPWR.n2854 VPWR.n2821 702.354
R8364 VPWR.n2837 VPWR.n2828 702.354
R8365 VPWR.n2850 VPWR.n2849 702.354
R8366 VPWR.n2835 VPWR.n2828 702.354
R8367 VPWR.n2815 VPWR.t978 651.634
R8368 VPWR.n2831 VPWR.t1424 651.505
R8369 VPWR.n2825 VPWR.t1265 651.505
R8370 VPWR.n2862 VPWR.t1131 651.431
R8371 VPWR.n1061 VPWR.t135 646.071
R8372 VPWR.n1122 VPWR.t31 646.071
R8373 VPWR.n1059 VPWR.t284 646.071
R8374 VPWR.n56 VPWR.t251 646.071
R8375 VPWR.n62 VPWR.t375 646.071
R8376 VPWR.n99 VPWR.t160 646.071
R8377 VPWR.n1053 VPWR.t450 646.071
R8378 VPWR.n1231 VPWR.t975 646.071
R8379 VPWR.n298 VPWR.t485 646.071
R8380 VPWR.n290 VPWR.t1159 646.071
R8381 VPWR.n306 VPWR.t1188 646.071
R8382 VPWR.n68 VPWR.t114 646.071
R8383 VPWR.n1153 VPWR.t1107 646.071
R8384 VPWR.n346 VPWR.t1608 646.071
R8385 VPWR.n98 VPWR.t289 646.071
R8386 VPWR.n967 VPWR.t1089 646.071
R8387 VPWR.n963 VPWR.t713 646.071
R8388 VPWR.n999 VPWR.t667 646.071
R8389 VPWR.n373 VPWR.t653 646.071
R8390 VPWR.n356 VPWR.t973 646.071
R8391 VPWR.n357 VPWR.t836 646.071
R8392 VPWR.n372 VPWR.t1482 646.071
R8393 VPWR.n318 VPWR.t1917 646.071
R8394 VPWR.n75 VPWR.t219 646.071
R8395 VPWR.n971 VPWR.t1389 646.071
R8396 VPWR.n369 VPWR.t914 646.071
R8397 VPWR.n322 VPWR.t904 646.071
R8398 VPWR.n80 VPWR.t91 646.071
R8399 VPWR.n945 VPWR.t908 646.071
R8400 VPWR.n932 VPWR.t1161 646.071
R8401 VPWR.n933 VPWR.t1614 646.071
R8402 VPWR.n936 VPWR.t1353 646.071
R8403 VPWR.n944 VPWR.t731 646.071
R8404 VPWR.n411 VPWR.t1909 646.071
R8405 VPWR.n387 VPWR.t1125 646.071
R8406 VPWR.n391 VPWR.t1007 646.071
R8407 VPWR.n395 VPWR.t1367 646.071
R8408 VPWR.n407 VPWR.t707 646.071
R8409 VPWR.n365 VPWR.t689 646.071
R8410 VPWR.n330 VPWR.t542 646.071
R8411 VPWR.n86 VPWR.t332 646.071
R8412 VPWR.n937 VPWR.t1631 646.071
R8413 VPWR.n403 VPWR.t1564 646.071
R8414 VPWR.n364 VPWR.t1553 646.071
R8415 VPWR.n334 VPWR.t1720 646.071
R8416 VPWR.n87 VPWR.t177 646.071
R8417 VPWR.n473 VPWR.t1572 646.071
R8418 VPWR.n481 VPWR.t832 646.071
R8419 VPWR.n480 VPWR.t1520 646.071
R8420 VPWR.n477 VPWR.t1385 646.071
R8421 VPWR.n476 VPWR.t1858 646.071
R8422 VPWR.n472 VPWR.t968 646.071
R8423 VPWR.n469 VPWR.t1893 646.071
R8424 VPWR.n468 VPWR.t871 646.071
R8425 VPWR.n465 VPWR.t1117 646.071
R8426 VPWR.n464 VPWR.t673 646.071
R8427 VPWR.n461 VPWR.t1582 646.071
R8428 VPWR.n460 VPWR.t1759 646.071
R8429 VPWR.n457 VPWR.t814 646.071
R8430 VPWR.n456 VPWR.t1618 646.071
R8431 VPWR.n453 VPWR.t1817 646.071
R8432 VPWR.n452 VPWR.t149 646.071
R8433 VPWR.n526 VPWR.t1716 646.071
R8434 VPWR.n482 VPWR.t1157 646.071
R8435 VPWR.n538 VPWR.t424 646.071
R8436 VPWR.n534 VPWR.t1359 646.071
R8437 VPWR.n530 VPWR.t1190 646.071
R8438 VPWR.n522 VPWR.t538 646.071
R8439 VPWR.n518 VPWR.t721 646.071
R8440 VPWR.n514 VPWR.t918 646.071
R8441 VPWR.n510 VPWR.t1913 646.071
R8442 VPWR.n506 VPWR.t645 646.071
R8443 VPWR.n502 VPWR.t1050 646.071
R8444 VPWR.n498 VPWR.t1186 646.071
R8445 VPWR.n494 VPWR.t1695 646.071
R8446 VPWR.n490 VPWR.t685 646.071
R8447 VPWR.n486 VPWR.t747 646.071
R8448 VPWR.n483 VPWR.t367 646.071
R8449 VPWR.n556 VPWR.t518 646.071
R8450 VPWR.n548 VPWR.t900 646.071
R8451 VPWR.n549 VPWR.t1087 646.071
R8452 VPWR.n552 VPWR.t1397 646.071
R8453 VPWR.n553 VPWR.t1036 646.071
R8454 VPWR.n557 VPWR.t568 646.071
R8455 VPWR.n560 VPWR.t743 646.071
R8456 VPWR.n561 VPWR.t574 646.071
R8457 VPWR.n564 VPWR.t960 646.071
R8458 VPWR.n565 VPWR.t621 646.071
R8459 VPWR.n568 VPWR.t1689 646.071
R8460 VPWR.n569 VPWR.t468 646.071
R8461 VPWR.n572 VPWR.t462 646.071
R8462 VPWR.n573 VPWR.t1783 646.071
R8463 VPWR.n576 VPWR.t1805 646.071
R8464 VPWR.n577 VPWR.t216 646.071
R8465 VPWR.n595 VPWR.t1551 646.071
R8466 VPWR.n579 VPWR.t1163 646.071
R8467 VPWR.n583 VPWR.t1911 646.071
R8468 VPWR.n587 VPWR.t1351 646.071
R8469 VPWR.n591 VPWR.t1635 646.071
R8470 VPWR.n599 VPWR.t687 646.071
R8471 VPWR.n603 VPWR.t1791 646.071
R8472 VPWR.n607 VPWR.t912 646.071
R8473 VPWR.n611 VPWR.t1925 646.071
R8474 VPWR.n615 VPWR.t651 646.071
R8475 VPWR.n619 VPWR.t1103 646.071
R8476 VPWR.n623 VPWR.t1460 646.071
R8477 VPWR.n627 VPWR.t1707 646.071
R8478 VPWR.n631 VPWR.t489 646.071
R8479 VPWR.n635 VPWR.t759 646.071
R8480 VPWR.n578 VPWR.t324 646.071
R8481 VPWR.n665 VPWR.t1560 646.071
R8482 VPWR.n673 VPWR.t980 646.071
R8483 VPWR.n672 VPWR.t1590 646.071
R8484 VPWR.n669 VPWR.t1371 646.071
R8485 VPWR.n668 VPWR.t1066 646.071
R8486 VPWR.n664 VPWR.t703 646.071
R8487 VPWR.n661 VPWR.t1905 646.071
R8488 VPWR.n660 VPWR.t1023 646.071
R8489 VPWR.n657 VPWR.t1606 646.071
R8490 VPWR.n656 VPWR.t1827 646.071
R8491 VPWR.n653 VPWR.t1476 646.071
R8492 VPWR.n652 VPWR.t1242 646.071
R8493 VPWR.n649 VPWR.t927 646.071
R8494 VPWR.n648 VPWR.t510 646.071
R8495 VPWR.n645 VPWR.t631 646.071
R8496 VPWR.n644 VPWR.t50 646.071
R8497 VPWR.n718 VPWR.t1570 646.071
R8498 VPWR.n674 VPWR.t715 646.071
R8499 VPWR.n730 VPWR.t844 646.071
R8500 VPWR.n726 VPWR.t1387 646.071
R8501 VPWR.n722 VPWR.t1854 646.071
R8502 VPWR.n714 VPWR.t966 646.071
R8503 VPWR.n710 VPWR.t1891 646.071
R8504 VPWR.n706 VPWR.t869 646.071
R8505 VPWR.n702 VPWR.t1115 646.071
R8506 VPWR.n698 VPWR.t669 646.071
R8507 VPWR.n694 VPWR.t1580 646.071
R8508 VPWR.n690 VPWR.t1755 646.071
R8509 VPWR.n686 VPWR.t812 646.071
R8510 VPWR.n682 VPWR.t1496 646.071
R8511 VPWR.n678 VPWR.t1813 646.071
R8512 VPWR.n675 VPWR.t157 646.071
R8513 VPWR.n748 VPWR.t1665 646.071
R8514 VPWR.n740 VPWR.t834 646.071
R8515 VPWR.n741 VPWR.t1524 646.071
R8516 VPWR.n744 VPWR.t1379 646.071
R8517 VPWR.n745 VPWR.t1860 646.071
R8518 VPWR.n749 VPWR.t590 646.071
R8519 VPWR.n752 VPWR.t1897 646.071
R8520 VPWR.n753 VPWR.t1111 646.071
R8521 VPWR.n756 VPWR.t1121 646.071
R8522 VPWR.n757 VPWR.t675 646.071
R8523 VPWR.n760 VPWR.t552 646.071
R8524 VPWR.n761 VPWR.t1204 646.071
R8525 VPWR.n764 VPWR.t818 646.071
R8526 VPWR.n765 VPWR.t1620 646.071
R8527 VPWR.n768 VPWR.t1819 646.071
R8528 VPWR.n769 VPWR.t117 646.071
R8529 VPWR.n787 VPWR.t1518 646.071
R8530 VPWR.n771 VPWR.t898 646.071
R8531 VPWR.n775 VPWR.t1083 646.071
R8532 VPWR.n779 VPWR.t1399 646.071
R8533 VPWR.n783 VPWR.t1034 646.071
R8534 VPWR.n791 VPWR.t564 646.071
R8535 VPWR.n795 VPWR.t739 646.071
R8536 VPWR.n799 VPWR.t572 646.071
R8537 VPWR.n803 VPWR.t956 646.071
R8538 VPWR.n807 VPWR.t619 646.071
R8539 VPWR.n811 VPWR.t1685 646.071
R8540 VPWR.n815 VPWR.t466 646.071
R8541 VPWR.n819 VPWR.t460 646.071
R8542 VPWR.n823 VPWR.t1781 646.071
R8543 VPWR.n827 VPWR.t701 646.071
R8544 VPWR.n770 VPWR.t222 646.071
R8545 VPWR.n857 VPWR.t1562 646.071
R8546 VPWR.n865 VPWR.t1123 646.071
R8547 VPWR.n864 VPWR.t1592 646.071
R8548 VPWR.n861 VPWR.t1369 646.071
R8549 VPWR.n860 VPWR.t1070 646.071
R8550 VPWR.n856 VPWR.t705 646.071
R8551 VPWR.n853 VPWR.t1907 646.071
R8552 VPWR.n852 VPWR.t385 646.071
R8553 VPWR.n849 VPWR.t1009 646.071
R8554 VPWR.n848 VPWR.t1829 646.071
R8555 VPWR.n845 VPWR.t1478 646.071
R8556 VPWR.n844 VPWR.t1244 646.071
R8557 VPWR.n841 VPWR.t929 646.071
R8558 VPWR.n840 VPWR.t512 646.071
R8559 VPWR.n837 VPWR.t635 646.071
R8560 VPWR.n836 VPWR.t42 646.071
R8561 VPWR.n910 VPWR.t1516 646.071
R8562 VPWR.n866 VPWR.t896 646.071
R8563 VPWR.n922 VPWR.t1081 646.071
R8564 VPWR.n918 VPWR.t1401 646.071
R8565 VPWR.n914 VPWR.t1032 646.071
R8566 VPWR.n906 VPWR.t562 646.071
R8567 VPWR.n902 VPWR.t1803 646.071
R8568 VPWR.n898 VPWR.t984 646.071
R8569 VPWR.n894 VPWR.t954 646.071
R8570 VPWR.n890 VPWR.t617 646.071
R8571 VPWR.n886 VPWR.t1683 646.071
R8572 VPWR.n882 VPWR.t1767 646.071
R8573 VPWR.n878 VPWR.t458 646.071
R8574 VPWR.n874 VPWR.t1779 646.071
R8575 VPWR.n870 VPWR.t699 646.071
R8576 VPWR.n867 VPWR.t229 646.071
R8577 VPWR.n940 VPWR.t1549 646.071
R8578 VPWR.n979 VPWR.t520 646.071
R8579 VPWR.n1227 VPWR.t1224 646.071
R8580 VPWR.n1179 VPWR.t61 646.071
R8581 VPWR.n399 VPWR.t1072 646.071
R8582 VPWR.n361 VPWR.t1637 646.071
R8583 VPWR.n338 VPWR.t1192 646.071
R8584 VPWR.n92 VPWR.t69 646.071
R8585 VPWR.n975 VPWR.t1038 646.071
R8586 VPWR.n1485 VPWR.t1641 646.071
R8587 VPWR.n1183 VPWR.t340 646.071
R8588 VPWR.n941 VPWR.t548 646.071
R8589 VPWR.n983 VPWR.t570 646.071
R8590 VPWR.n1173 VPWR.t691 646.071
R8591 VPWR.n1217 VPWR.t208 646.071
R8592 VPWR.n415 VPWR.t387 646.071
R8593 VPWR.n419 VPWR.t1011 646.071
R8594 VPWR.n423 VPWR.t1831 646.071
R8595 VPWR.n427 VPWR.t1480 646.071
R8596 VPWR.n431 VPWR.t1246 646.071
R8597 VPWR.n435 VPWR.t931 646.071
R8598 VPWR.n439 VPWR.t514 646.071
R8599 VPWR.n443 VPWR.t637 646.071
R8600 VPWR.n386 VPWR.t34 646.071
R8601 VPWR.n368 VPWR.t1793 646.071
R8602 VPWR.n326 VPWR.t725 646.071
R8603 VPWR.n81 VPWR.t56 646.071
R8604 VPWR.n987 VPWR.t745 646.071
R8605 VPWR.n1169 VPWR.t1795 646.071
R8606 VPWR.n1214 VPWR.t316 646.071
R8607 VPWR.n948 VPWR.t1923 646.071
R8608 VPWR.n949 VPWR.t649 646.071
R8609 VPWR.n952 VPWR.t1101 646.071
R8610 VPWR.n953 VPWR.t1458 646.071
R8611 VPWR.n956 VPWR.t1703 646.071
R8612 VPWR.n957 VPWR.t487 646.071
R8613 VPWR.n960 VPWR.t755 646.071
R8614 VPWR.n961 VPWR.t337 646.071
R8615 VPWR.n991 VPWR.t576 646.071
R8616 VPWR.n1163 VPWR.t855 646.071
R8617 VPWR.n1206 VPWR.t356 646.071
R8618 VPWR.n360 VPWR.t1349 646.071
R8619 VPWR.n342 VPWR.t1357 646.071
R8620 VPWR.n93 VPWR.t307 646.071
R8621 VPWR.n1479 VPWR.t1405 646.071
R8622 VPWR.n1180 VPWR.t180 646.071
R8623 VPWR.n995 VPWR.t476 646.071
R8624 VPWR.n1159 VPWR.t1484 646.071
R8625 VPWR.n1203 VPWR.t101 646.071
R8626 VPWR.n376 VPWR.t1105 646.071
R8627 VPWR.n377 VPWR.t1462 646.071
R8628 VPWR.n380 VPWR.t1709 646.071
R8629 VPWR.n381 VPWR.t861 646.071
R8630 VPWR.n384 VPWR.t761 646.071
R8631 VPWR.n385 VPWR.t319 646.071
R8632 VPWR.n314 VPWR.t647 646.071
R8633 VPWR.n74 VPWR.t329 646.071
R8634 VPWR.n1149 VPWR.t1789 646.071
R8635 VPWR.n1200 VPWR.t205 646.071
R8636 VPWR.n1003 VPWR.t1691 646.071
R8637 VPWR.n1007 VPWR.t474 646.071
R8638 VPWR.n1011 VPWR.t464 646.071
R8639 VPWR.n1015 VPWR.t1494 646.071
R8640 VPWR.n1019 VPWR.t1807 646.071
R8641 VPWR.n962 VPWR.t189 646.071
R8642 VPWR.n1472 VPWR.t838 646.071
R8643 VPWR.n1123 VPWR.t167 646.071
R8644 VPWR.n310 VPWR.t1054 646.071
R8645 VPWR.n69 VPWR.t96 646.071
R8646 VPWR.n1192 VPWR.t364 646.071
R8647 VPWR.n1049 VPWR.t1171 646.071
R8648 VPWR.n1189 VPWR.t383 646.071
R8649 VPWR.n302 VPWR.t1699 646.071
R8650 VPWR.n294 VPWR.t749 646.071
R8651 VPWR.n291 VPWR.t359 646.071
R8652 VPWR.n1058 VPWR.t256 646.071
R8653 VPWR.n1748 VPWR.t863 646.071
R8654 VPWR.n1036 VPWR.t765 646.071
R8655 VPWR.n1032 VPWR.t300 646.071
R8656 VPWR.n1186 VPWR.t127 646.071
R8657 VPWR.n63 VPWR.t242 646.071
R8658 VPWR.n57 VPWR.t15 646.071
R8659 VPWR.n1230 VPWR.t109 642.13
R8660 VPWR.n1152 VPWR.t37 642.13
R8661 VPWR.n1226 VPWR.t245 642.13
R8662 VPWR.n1484 VPWR.t143 642.13
R8663 VPWR.n1172 VPWR.t267 642.13
R8664 VPWR.n1168 VPWR.t18 642.13
R8665 VPWR.n1162 VPWR.t140 642.13
R8666 VPWR.n1478 VPWR.t372 642.13
R8667 VPWR.n1158 VPWR.t281 642.13
R8668 VPWR.n1148 VPWR.t297 642.13
R8669 VPWR.n1471 VPWR.t270 642.13
R8670 VPWR.n1048 VPWR.t170 642.13
R8671 VPWR.n1747 VPWR.t47 642.13
R8672 VPWR.n1035 VPWR.t84 642.13
R8673 VPWR.n1031 VPWR.t192 642.13
R8674 VPWR.n1052 VPWR.t211 642.13
R8675 VPWR.n2309 VPWR.t831 629.652
R8676 VPWR.n2310 VPWR.t1519 629.652
R8677 VPWR.n2319 VPWR.t1384 629.652
R8678 VPWR.n2320 VPWR.t1857 629.652
R8679 VPWR.n2329 VPWR.t1571 629.652
R8680 VPWR.n2330 VPWR.t967 629.652
R8681 VPWR.n2339 VPWR.t1892 629.652
R8682 VPWR.n2340 VPWR.t870 629.652
R8683 VPWR.n2349 VPWR.t1116 629.652
R8684 VPWR.n2350 VPWR.t672 629.652
R8685 VPWR.n2359 VPWR.t1581 629.652
R8686 VPWR.n2360 VPWR.t1758 629.652
R8687 VPWR.n2369 VPWR.t813 629.652
R8688 VPWR.n2370 VPWR.t1617 629.652
R8689 VPWR.n2379 VPWR.t1816 629.652
R8690 VPWR.n542 VPWR.t1156 629.652
R8691 VPWR.t423 VPWR.n541 629.652
R8692 VPWR.t1358 VPWR.n537 629.652
R8693 VPWR.t1189 VPWR.n533 629.652
R8694 VPWR.t1715 VPWR.n529 629.652
R8695 VPWR.t537 VPWR.n525 629.652
R8696 VPWR.t720 VPWR.n521 629.652
R8697 VPWR.t917 VPWR.n517 629.652
R8698 VPWR.t1912 VPWR.n513 629.652
R8699 VPWR.t644 VPWR.n509 629.652
R8700 VPWR.t1049 VPWR.n505 629.652
R8701 VPWR.t1185 VPWR.n501 629.652
R8702 VPWR.t1694 VPWR.n497 629.652
R8703 VPWR.t684 VPWR.n493 629.652
R8704 VPWR.t746 VPWR.n489 629.652
R8705 VPWR.n2281 VPWR.t899 629.652
R8706 VPWR.t1086 VPWR.n2280 629.652
R8707 VPWR.n2271 VPWR.t1396 629.652
R8708 VPWR.t1035 VPWR.n2270 629.652
R8709 VPWR.n2261 VPWR.t517 629.652
R8710 VPWR.t567 VPWR.n2260 629.652
R8711 VPWR.n2251 VPWR.t742 629.652
R8712 VPWR.t573 VPWR.n2250 629.652
R8713 VPWR.n2241 VPWR.t959 629.652
R8714 VPWR.t620 VPWR.n2240 629.652
R8715 VPWR.n2231 VPWR.t1688 629.652
R8716 VPWR.t467 VPWR.n2230 629.652
R8717 VPWR.n2221 VPWR.t461 629.652
R8718 VPWR.t1782 VPWR.n2220 629.652
R8719 VPWR.n2211 VPWR.t1804 629.652
R8720 VPWR.n582 VPWR.t1162 629.652
R8721 VPWR.n586 VPWR.t1910 629.652
R8722 VPWR.n590 VPWR.t1350 629.652
R8723 VPWR.n594 VPWR.t1634 629.652
R8724 VPWR.n598 VPWR.t1550 629.652
R8725 VPWR.n602 VPWR.t686 629.652
R8726 VPWR.n606 VPWR.t1790 629.652
R8727 VPWR.n610 VPWR.t911 629.652
R8728 VPWR.n614 VPWR.t1924 629.652
R8729 VPWR.n618 VPWR.t650 629.652
R8730 VPWR.n622 VPWR.t1102 629.652
R8731 VPWR.n626 VPWR.t1459 629.652
R8732 VPWR.n630 VPWR.t1706 629.652
R8733 VPWR.n634 VPWR.t488 629.652
R8734 VPWR.n638 VPWR.t758 629.652
R8735 VPWR.n2113 VPWR.t979 629.652
R8736 VPWR.n2114 VPWR.t1589 629.652
R8737 VPWR.n2123 VPWR.t1370 629.652
R8738 VPWR.n2124 VPWR.t1065 629.652
R8739 VPWR.n2133 VPWR.t1559 629.652
R8740 VPWR.n2134 VPWR.t702 629.652
R8741 VPWR.n2143 VPWR.t1904 629.652
R8742 VPWR.n2144 VPWR.t1022 629.652
R8743 VPWR.n2153 VPWR.t1605 629.652
R8744 VPWR.n2154 VPWR.t1826 629.652
R8745 VPWR.n2163 VPWR.t1475 629.652
R8746 VPWR.n2164 VPWR.t1241 629.652
R8747 VPWR.n2173 VPWR.t926 629.652
R8748 VPWR.n2174 VPWR.t509 629.652
R8749 VPWR.n2183 VPWR.t630 629.652
R8750 VPWR.n734 VPWR.t714 629.652
R8751 VPWR.t843 VPWR.n733 629.652
R8752 VPWR.t1386 VPWR.n729 629.652
R8753 VPWR.t1853 VPWR.n725 629.652
R8754 VPWR.t1569 VPWR.n721 629.652
R8755 VPWR.t965 VPWR.n717 629.652
R8756 VPWR.t1890 VPWR.n713 629.652
R8757 VPWR.t868 VPWR.n709 629.652
R8758 VPWR.t1114 VPWR.n705 629.652
R8759 VPWR.t668 VPWR.n701 629.652
R8760 VPWR.t1579 VPWR.n697 629.652
R8761 VPWR.t1754 VPWR.n693 629.652
R8762 VPWR.t811 VPWR.n689 629.652
R8763 VPWR.t1495 VPWR.n685 629.652
R8764 VPWR.t1812 VPWR.n681 629.652
R8765 VPWR.n2085 VPWR.t833 629.652
R8766 VPWR.t1523 VPWR.n2084 629.652
R8767 VPWR.n2075 VPWR.t1378 629.652
R8768 VPWR.t1859 VPWR.n2074 629.652
R8769 VPWR.n2065 VPWR.t1664 629.652
R8770 VPWR.t589 VPWR.n2064 629.652
R8771 VPWR.n2055 VPWR.t1896 629.652
R8772 VPWR.t1110 VPWR.n2054 629.652
R8773 VPWR.n2045 VPWR.t1120 629.652
R8774 VPWR.t674 VPWR.n2044 629.652
R8775 VPWR.n2035 VPWR.t551 629.652
R8776 VPWR.t1203 VPWR.n2034 629.652
R8777 VPWR.n2025 VPWR.t817 629.652
R8778 VPWR.t1619 VPWR.n2024 629.652
R8779 VPWR.n2015 VPWR.t1818 629.652
R8780 VPWR.n774 VPWR.t897 629.652
R8781 VPWR.n778 VPWR.t1082 629.652
R8782 VPWR.n782 VPWR.t1398 629.652
R8783 VPWR.n786 VPWR.t1033 629.652
R8784 VPWR.n790 VPWR.t1517 629.652
R8785 VPWR.n794 VPWR.t563 629.652
R8786 VPWR.n798 VPWR.t738 629.652
R8787 VPWR.n802 VPWR.t571 629.652
R8788 VPWR.n806 VPWR.t955 629.652
R8789 VPWR.n810 VPWR.t618 629.652
R8790 VPWR.n814 VPWR.t1684 629.652
R8791 VPWR.n818 VPWR.t465 629.652
R8792 VPWR.n822 VPWR.t459 629.652
R8793 VPWR.n826 VPWR.t1780 629.652
R8794 VPWR.n830 VPWR.t700 629.652
R8795 VPWR.n1917 VPWR.t1122 629.652
R8796 VPWR.n1918 VPWR.t1591 629.652
R8797 VPWR.n1927 VPWR.t1368 629.652
R8798 VPWR.n1928 VPWR.t1069 629.652
R8799 VPWR.n1937 VPWR.t1561 629.652
R8800 VPWR.n1938 VPWR.t704 629.652
R8801 VPWR.n1947 VPWR.t1906 629.652
R8802 VPWR.n1948 VPWR.t384 629.652
R8803 VPWR.n1957 VPWR.t1008 629.652
R8804 VPWR.n1958 VPWR.t1828 629.652
R8805 VPWR.n1967 VPWR.t1477 629.652
R8806 VPWR.n1968 VPWR.t1243 629.652
R8807 VPWR.n1977 VPWR.t928 629.652
R8808 VPWR.n1978 VPWR.t511 629.652
R8809 VPWR.n1987 VPWR.t634 629.652
R8810 VPWR.n926 VPWR.t895 629.652
R8811 VPWR.t1080 VPWR.n925 629.652
R8812 VPWR.t1400 VPWR.n921 629.652
R8813 VPWR.t1031 VPWR.n917 629.652
R8814 VPWR.t1515 VPWR.n913 629.652
R8815 VPWR.t561 VPWR.n909 629.652
R8816 VPWR.t1802 VPWR.n905 629.652
R8817 VPWR.t983 VPWR.n901 629.652
R8818 VPWR.t953 VPWR.n897 629.652
R8819 VPWR.t616 VPWR.n893 629.652
R8820 VPWR.t1682 VPWR.n889 629.652
R8821 VPWR.t1766 VPWR.n885 629.652
R8822 VPWR.t457 VPWR.n881 629.652
R8823 VPWR.t1778 VPWR.n877 629.652
R8824 VPWR.t698 VPWR.n873 629.652
R8825 VPWR.n390 VPWR.t1124 629.652
R8826 VPWR.n394 VPWR.t1006 629.652
R8827 VPWR.n398 VPWR.t1366 629.652
R8828 VPWR.n402 VPWR.t1071 629.652
R8829 VPWR.n406 VPWR.t1563 629.652
R8830 VPWR.n410 VPWR.t706 629.652
R8831 VPWR.n414 VPWR.t1908 629.652
R8832 VPWR.n418 VPWR.t386 629.652
R8833 VPWR.n422 VPWR.t1010 629.652
R8834 VPWR.n426 VPWR.t1830 629.652
R8835 VPWR.n430 VPWR.t1479 629.652
R8836 VPWR.n434 VPWR.t1245 629.652
R8837 VPWR.n438 VPWR.t930 629.652
R8838 VPWR.n442 VPWR.t513 629.652
R8839 VPWR.n446 VPWR.t636 629.652
R8840 VPWR.n1889 VPWR.t1160 629.652
R8841 VPWR.t1613 VPWR.n1888 629.652
R8842 VPWR.n1879 VPWR.t1352 629.652
R8843 VPWR.t1630 VPWR.n1878 629.652
R8844 VPWR.n1869 VPWR.t1548 629.652
R8845 VPWR.t547 VPWR.n1868 629.652
R8846 VPWR.n1859 VPWR.t730 629.652
R8847 VPWR.t907 VPWR.n1858 629.652
R8848 VPWR.n1849 VPWR.t1922 629.652
R8849 VPWR.t648 VPWR.n1848 629.652
R8850 VPWR.n1839 VPWR.t1100 629.652
R8851 VPWR.t1457 VPWR.n1838 629.652
R8852 VPWR.n1829 VPWR.t1702 629.652
R8853 VPWR.t486 VPWR.n1828 629.652
R8854 VPWR.n1819 VPWR.t754 629.652
R8855 VPWR.n2477 VPWR.t972 629.652
R8856 VPWR.t835 VPWR.n2476 629.652
R8857 VPWR.n2467 VPWR.t1348 629.652
R8858 VPWR.t1636 VPWR.n2466 629.652
R8859 VPWR.n2457 VPWR.t1552 629.652
R8860 VPWR.t688 VPWR.n2456 629.652
R8861 VPWR.n2447 VPWR.t1792 629.652
R8862 VPWR.t913 VPWR.n2446 629.652
R8863 VPWR.n2437 VPWR.t1481 629.652
R8864 VPWR.t652 VPWR.n2436 629.652
R8865 VPWR.n2427 VPWR.t1104 629.652
R8866 VPWR.t1461 VPWR.n2426 629.652
R8867 VPWR.n2417 VPWR.t1708 629.652
R8868 VPWR.t860 VPWR.n2416 629.652
R8869 VPWR.n2407 VPWR.t760 629.652
R8870 VPWR.n966 VPWR.t712 629.652
R8871 VPWR.n970 VPWR.t1088 629.652
R8872 VPWR.n974 VPWR.t1388 629.652
R8873 VPWR.n978 VPWR.t1037 629.652
R8874 VPWR.n982 VPWR.t519 629.652
R8875 VPWR.n986 VPWR.t569 629.652
R8876 VPWR.n990 VPWR.t744 629.652
R8877 VPWR.n994 VPWR.t575 629.652
R8878 VPWR.n998 VPWR.t475 629.652
R8879 VPWR.n1002 VPWR.t666 629.652
R8880 VPWR.n1006 VPWR.t1690 629.652
R8881 VPWR.n1010 VPWR.t473 629.652
R8882 VPWR.n1014 VPWR.t463 629.652
R8883 VPWR.n1018 VPWR.t1493 629.652
R8884 VPWR.n1022 VPWR.t1806 629.652
R8885 VPWR.n350 VPWR.t1158 629.652
R8886 VPWR.t1607 VPWR.n349 629.652
R8887 VPWR.t1356 VPWR.n345 629.652
R8888 VPWR.t1191 VPWR.n341 629.652
R8889 VPWR.t1719 VPWR.n337 629.652
R8890 VPWR.t541 VPWR.n333 629.652
R8891 VPWR.t724 VPWR.n329 629.652
R8892 VPWR.t903 VPWR.n325 629.652
R8893 VPWR.t1916 VPWR.n321 629.652
R8894 VPWR.t646 VPWR.n317 629.652
R8895 VPWR.t1053 VPWR.n313 629.652
R8896 VPWR.t1187 VPWR.n309 629.652
R8897 VPWR.t1698 VPWR.n305 629.652
R8898 VPWR.t484 VPWR.n301 629.652
R8899 VPWR.t748 VPWR.n297 629.652
R8900 VPWR.n1468 VPWR.t974 629.652
R8901 VPWR.n1475 VPWR.t837 629.652
R8902 VPWR.n1481 VPWR.t1404 629.652
R8903 VPWR.n1492 VPWR.t1640 629.652
R8904 VPWR.n1493 VPWR.t1223 629.652
R8905 VPWR.n1506 VPWR.t690 629.652
R8906 VPWR.n1507 VPWR.t1794 629.652
R8907 VPWR.n1520 VPWR.t854 629.652
R8908 VPWR.n1521 VPWR.t1483 629.652
R8909 VPWR.n1536 VPWR.t1788 629.652
R8910 VPWR.t1106 VPWR.n1535 629.652
R8911 VPWR.n1761 VPWR.t1170 629.652
R8912 VPWR.t449 VPWR.n1760 629.652
R8913 VPWR.n1749 VPWR.t862 629.652
R8914 VPWR.n1791 VPWR.t764 629.652
R8915 VPWR.n2506 VPWR.t159 629.652
R8916 VPWR.n2507 VPWR.t288 629.652
R8917 VPWR.n2518 VPWR.t306 629.652
R8918 VPWR.n2519 VPWR.t68 629.652
R8919 VPWR.n2530 VPWR.t176 629.652
R8920 VPWR.n2531 VPWR.t331 629.652
R8921 VPWR.n2542 VPWR.t55 629.652
R8922 VPWR.n2543 VPWR.t90 629.652
R8923 VPWR.n2554 VPWR.t218 629.652
R8924 VPWR.n2555 VPWR.t328 629.652
R8925 VPWR.n2566 VPWR.t95 629.652
R8926 VPWR.n2567 VPWR.t113 629.652
R8927 VPWR.n2578 VPWR.t241 629.652
R8928 VPWR.n2579 VPWR.t374 629.652
R8929 VPWR.n2590 VPWR.t14 629.652
R8930 VPWR.n1594 VPWR.t30 629.652
R8931 VPWR.t166 VPWR.n1593 629.652
R8932 VPWR.n1182 VPWR.t179 629.652
R8933 VPWR.n1185 VPWR.t339 629.652
R8934 VPWR.n1220 VPWR.t60 629.652
R8935 VPWR.t207 VPWR.n1219 629.652
R8936 VPWR.t315 VPWR.n1216 629.652
R8937 VPWR.t355 VPWR.n1213 629.652
R8938 VPWR.t100 VPWR.n1205 629.652
R8939 VPWR.t204 VPWR.n1202 629.652
R8940 VPWR.t363 VPWR.n1199 629.652
R8941 VPWR.t382 VPWR.n1191 629.652
R8942 VPWR.t126 VPWR.n1188 629.652
R8943 VPWR.n1740 VPWR.t255 629.652
R8944 VPWR.t283 VPWR.n1739 629.652
R8945 VPWR.n2836 VPWR.t1264 531.804
R8946 VPWR.n2855 VPWR.t1264 531.804
R8947 VPWR.n2851 VPWR.n2850 504.707
R8948 VPWR.t831 VPWR.t1097 486.048
R8949 VPWR.t1519 VPWR.t1623 486.048
R8950 VPWR.t1645 VPWR.t1384 486.048
R8951 VPWR.t1857 VPWR.t1644 486.048
R8952 VPWR.t1096 VPWR.t1571 486.048
R8953 VPWR.t967 VPWR.t800 486.048
R8954 VPWR.t799 VPWR.t1892 486.048
R8955 VPWR.t870 VPWR.t1095 486.048
R8956 VPWR.t1625 VPWR.t1116 486.048
R8957 VPWR.t672 VPWR.t801 486.048
R8958 VPWR.t1643 VPWR.t1581 486.048
R8959 VPWR.t1758 VPWR.t1642 486.048
R8960 VPWR.t798 VPWR.t813 486.048
R8961 VPWR.t1617 VPWR.t797 486.048
R8962 VPWR.t1646 VPWR.t1816 486.048
R8963 VPWR.t148 VPWR.t1624 486.048
R8964 VPWR.t1156 VPWR.t1233 486.048
R8965 VPWR.t1554 VPWR.t423 486.048
R8966 VPWR.t1237 VPWR.t1358 486.048
R8967 VPWR.t1236 VPWR.t1189 486.048
R8968 VPWR.t1558 VPWR.t1715 486.048
R8969 VPWR.t1452 VPWR.t537 486.048
R8970 VPWR.t1451 VPWR.t720 486.048
R8971 VPWR.t1557 VPWR.t917 486.048
R8972 VPWR.t1556 VPWR.t1912 486.048
R8973 VPWR.t1453 VPWR.t644 486.048
R8974 VPWR.t1235 VPWR.t1049 486.048
R8975 VPWR.t1234 VPWR.t1185 486.048
R8976 VPWR.t1450 VPWR.t1694 486.048
R8977 VPWR.t1449 VPWR.t684 486.048
R8978 VPWR.t1238 VPWR.t746 486.048
R8979 VPWR.t1555 VPWR.t366 486.048
R8980 VPWR.t899 VPWR.t1274 486.048
R8981 VPWR.t1221 VPWR.t1086 486.048
R8982 VPWR.t1396 VPWR.t430 486.048
R8983 VPWR.t429 VPWR.t1035 486.048
R8984 VPWR.t517 VPWR.t1273 486.048
R8985 VPWR.t1219 VPWR.t567 486.048
R8986 VPWR.t742 VPWR.t1218 486.048
R8987 VPWR.t1272 VPWR.t573 486.048
R8988 VPWR.t959 VPWR.t1271 486.048
R8989 VPWR.t1220 VPWR.t620 486.048
R8990 VPWR.t1688 VPWR.t428 486.048
R8991 VPWR.t427 VPWR.t467 486.048
R8992 VPWR.t461 VPWR.t1217 486.048
R8993 VPWR.t1216 VPWR.t1782 486.048
R8994 VPWR.t1804 VPWR.t1215 486.048
R8995 VPWR.t1222 VPWR.t215 486.048
R8996 VPWR.t1162 VPWR.t1446 486.048
R8997 VPWR.t1910 VPWR.t1441 486.048
R8998 VPWR.t1350 VPWR.t607 486.048
R8999 VPWR.t1634 VPWR.t606 486.048
R9000 VPWR.t1550 VPWR.t1445 486.048
R9001 VPWR.t686 VPWR.t1168 486.048
R9002 VPWR.t1790 VPWR.t1167 486.048
R9003 VPWR.t911 VPWR.t1444 486.048
R9004 VPWR.t1924 VPWR.t1443 486.048
R9005 VPWR.t650 VPWR.t1169 486.048
R9006 VPWR.t1102 VPWR.t1448 486.048
R9007 VPWR.t1459 VPWR.t1447 486.048
R9008 VPWR.t1706 VPWR.t1166 486.048
R9009 VPWR.t488 VPWR.t1165 486.048
R9010 VPWR.t758 VPWR.t1164 486.048
R9011 VPWR.t323 VPWR.t1442 486.048
R9012 VPWR.t979 VPWR.t1506 486.048
R9013 VPWR.t1589 VPWR.t921 486.048
R9014 VPWR.t496 VPWR.t1370 486.048
R9015 VPWR.t1065 VPWR.t495 486.048
R9016 VPWR.t1505 VPWR.t1559 486.048
R9017 VPWR.t702 VPWR.t1565 486.048
R9018 VPWR.t1005 VPWR.t1904 486.048
R9019 VPWR.t1022 VPWR.t826 486.048
R9020 VPWR.t825 VPWR.t1605 486.048
R9021 VPWR.t1826 VPWR.t1566 486.048
R9022 VPWR.t1508 VPWR.t1475 486.048
R9023 VPWR.t1241 VPWR.t1507 486.048
R9024 VPWR.t1004 VPWR.t926 486.048
R9025 VPWR.t509 VPWR.t1003 486.048
R9026 VPWR.t497 VPWR.t630 486.048
R9027 VPWR.t49 VPWR.t824 486.048
R9028 VPWR.t714 VPWR.t600 486.048
R9029 VPWR.t732 VPWR.t843 486.048
R9030 VPWR.t605 VPWR.t1386 486.048
R9031 VPWR.t604 VPWR.t1853 486.048
R9032 VPWR.t599 VPWR.t1569 486.048
R9033 VPWR.t1043 VPWR.t965 486.048
R9034 VPWR.t1042 VPWR.t1890 486.048
R9035 VPWR.t598 VPWR.t868 486.048
R9036 VPWR.t1712 VPWR.t1114 486.048
R9037 VPWR.t1044 VPWR.t668 486.048
R9038 VPWR.t603 VPWR.t1579 486.048
R9039 VPWR.t602 VPWR.t1754 486.048
R9040 VPWR.t1041 VPWR.t811 486.048
R9041 VPWR.t1040 VPWR.t1495 486.048
R9042 VPWR.t1039 VPWR.t1812 486.048
R9043 VPWR.t733 VPWR.t156 486.048
R9044 VPWR.t833 VPWR.t789 486.048
R9045 VPWR.t1078 VPWR.t1523 486.048
R9046 VPWR.t1378 VPWR.t793 486.048
R9047 VPWR.t792 VPWR.t1859 486.048
R9048 VPWR.t1664 VPWR.t788 486.048
R9049 VPWR.t1076 VPWR.t589 486.048
R9050 VPWR.t1896 VPWR.t1075 486.048
R9051 VPWR.t787 VPWR.t1110 486.048
R9052 VPWR.t1120 VPWR.t786 486.048
R9053 VPWR.t1077 VPWR.t674 486.048
R9054 VPWR.t551 VPWR.t791 486.048
R9055 VPWR.t790 VPWR.t1203 486.048
R9056 VPWR.t817 VPWR.t1074 486.048
R9057 VPWR.t1073 VPWR.t1619 486.048
R9058 VPWR.t1818 VPWR.t794 486.048
R9059 VPWR.t785 VPWR.t116 486.048
R9060 VPWR.t897 VPWR.t1753 486.048
R9061 VPWR.t1082 VPWR.t1748 486.048
R9062 VPWR.t1398 VPWR.t1771 486.048
R9063 VPWR.t1033 VPWR.t1770 486.048
R9064 VPWR.t1517 VPWR.t1752 486.048
R9065 VPWR.t563 VPWR.t1776 486.048
R9066 VPWR.t738 VPWR.t1775 486.048
R9067 VPWR.t571 VPWR.t1751 486.048
R9068 VPWR.t955 VPWR.t1750 486.048
R9069 VPWR.t618 VPWR.t1777 486.048
R9070 VPWR.t1684 VPWR.t1769 486.048
R9071 VPWR.t465 VPWR.t1768 486.048
R9072 VPWR.t459 VPWR.t1774 486.048
R9073 VPWR.t1780 VPWR.t1773 486.048
R9074 VPWR.t700 VPWR.t1772 486.048
R9075 VPWR.t221 VPWR.t1749 486.048
R9076 VPWR.t1122 VPWR.t1846 486.048
R9077 VPWR.t1591 VPWR.t852 486.048
R9078 VPWR.t1836 VPWR.t1368 486.048
R9079 VPWR.t1069 VPWR.t1849 486.048
R9080 VPWR.t1845 VPWR.t1561 486.048
R9081 VPWR.t704 VPWR.t1841 486.048
R9082 VPWR.t1840 VPWR.t1906 486.048
R9083 VPWR.t384 VPWR.t1844 486.048
R9084 VPWR.t1843 VPWR.t1008 486.048
R9085 VPWR.t1828 VPWR.t1842 486.048
R9086 VPWR.t1848 VPWR.t1477 486.048
R9087 VPWR.t1243 VPWR.t1847 486.048
R9088 VPWR.t1839 VPWR.t928 486.048
R9089 VPWR.t511 VPWR.t1838 486.048
R9090 VPWR.t1837 VPWR.t634 486.048
R9091 VPWR.t41 VPWR.t853 486.048
R9092 VPWR.t895 VPWR.t1652 486.048
R9093 VPWR.t1647 VPWR.t1080 486.048
R9094 VPWR.t391 VPWR.t1400 486.048
R9095 VPWR.t390 VPWR.t1031 486.048
R9096 VPWR.t1651 VPWR.t1515 486.048
R9097 VPWR.t1529 VPWR.t561 486.048
R9098 VPWR.t1528 VPWR.t1802 486.048
R9099 VPWR.t1650 VPWR.t983 486.048
R9100 VPWR.t1649 VPWR.t953 486.048
R9101 VPWR.t1530 VPWR.t616 486.048
R9102 VPWR.t389 VPWR.t1682 486.048
R9103 VPWR.t388 VPWR.t1766 486.048
R9104 VPWR.t1527 VPWR.t457 486.048
R9105 VPWR.t1526 VPWR.t1778 486.048
R9106 VPWR.t1525 VPWR.t698 486.048
R9107 VPWR.t1648 VPWR.t228 486.048
R9108 VPWR.t1124 VPWR.t1673 486.048
R9109 VPWR.t1006 VPWR.t1225 486.048
R9110 VPWR.t1366 VPWR.t1230 486.048
R9111 VPWR.t1071 VPWR.t1229 486.048
R9112 VPWR.t1563 VPWR.t1672 486.048
R9113 VPWR.t706 VPWR.t1677 486.048
R9114 VPWR.t1908 VPWR.t1676 486.048
R9115 VPWR.t386 VPWR.t1671 486.048
R9116 VPWR.t1010 VPWR.t1227 486.048
R9117 VPWR.t1830 VPWR.t1678 486.048
R9118 VPWR.t1479 VPWR.t1228 486.048
R9119 VPWR.t1245 VPWR.t1674 486.048
R9120 VPWR.t930 VPWR.t1675 486.048
R9121 VPWR.t513 VPWR.t1232 486.048
R9122 VPWR.t636 VPWR.t1231 486.048
R9123 VPWR.t33 VPWR.t1226 486.048
R9124 VPWR.t1160 VPWR.t1487 486.048
R9125 VPWR.t434 VPWR.t1613 486.048
R9126 VPWR.t1352 VPWR.t1202 486.048
R9127 VPWR.t1490 VPWR.t1630 486.048
R9128 VPWR.t1548 VPWR.t1486 486.048
R9129 VPWR.t432 VPWR.t547 486.048
R9130 VPWR.t730 VPWR.t431 486.048
R9131 VPWR.t1485 VPWR.t907 486.048
R9132 VPWR.t1922 VPWR.t436 486.048
R9133 VPWR.t433 VPWR.t648 486.048
R9134 VPWR.t1100 VPWR.t1489 486.048
R9135 VPWR.t1488 VPWR.t1457 486.048
R9136 VPWR.t1702 VPWR.t1456 486.048
R9137 VPWR.t1455 VPWR.t486 486.048
R9138 VPWR.t754 VPWR.t1454 486.048
R9139 VPWR.t435 VPWR.t336 486.048
R9140 VPWR.t972 VPWR.t1279 486.048
R9141 VPWR.t1663 VPWR.t835 486.048
R9142 VPWR.t1348 VPWR.t498 486.048
R9143 VPWR.t1533 VPWR.t1636 486.048
R9144 VPWR.t1552 VPWR.t1278 486.048
R9145 VPWR.t1661 VPWR.t688 486.048
R9146 VPWR.t1792 VPWR.t1660 486.048
R9147 VPWR.t1277 VPWR.t913 486.048
R9148 VPWR.t1481 VPWR.t1276 486.048
R9149 VPWR.t1662 VPWR.t652 486.048
R9150 VPWR.t1104 VPWR.t1532 486.048
R9151 VPWR.t1531 VPWR.t1461 486.048
R9152 VPWR.t1708 VPWR.t501 486.048
R9153 VPWR.t500 VPWR.t860 486.048
R9154 VPWR.t760 VPWR.t499 486.048
R9155 VPWR.t1275 VPWR.t318 486.048
R9156 VPWR.t712 VPWR.t1260 486.048
R9157 VPWR.t1088 VPWR.t481 486.048
R9158 VPWR.t1388 VPWR.t525 486.048
R9159 VPWR.t1037 VPWR.t524 486.048
R9160 VPWR.t519 VPWR.t796 486.048
R9161 VPWR.t569 VPWR.t948 486.048
R9162 VPWR.t744 VPWR.t947 486.048
R9163 VPWR.t575 VPWR.t795 486.048
R9164 VPWR.t475 VPWR.t483 486.048
R9165 VPWR.t666 VPWR.t949 486.048
R9166 VPWR.t1690 VPWR.t523 486.048
R9167 VPWR.t473 VPWR.t1261 486.048
R9168 VPWR.t463 VPWR.t946 486.048
R9169 VPWR.t1493 VPWR.t945 486.048
R9170 VPWR.t1806 VPWR.t526 486.048
R9171 VPWR.t188 VPWR.t482 486.048
R9172 VPWR.t1158 VPWR.t1877 486.048
R9173 VPWR.t1656 VPWR.t1607 486.048
R9174 VPWR.t1881 VPWR.t1356 486.048
R9175 VPWR.t1880 VPWR.t1191 486.048
R9176 VPWR.t1876 VPWR.t1719 486.048
R9177 VPWR.t1654 VPWR.t541 486.048
R9178 VPWR.t1653 VPWR.t724 486.048
R9179 VPWR.t1659 VPWR.t903 486.048
R9180 VPWR.t1658 VPWR.t1916 486.048
R9181 VPWR.t1655 VPWR.t646 486.048
R9182 VPWR.t1879 VPWR.t1053 486.048
R9183 VPWR.t1878 VPWR.t1187 486.048
R9184 VPWR.t1194 VPWR.t1698 486.048
R9185 VPWR.t1193 VPWR.t484 486.048
R9186 VPWR.t804 VPWR.t748 486.048
R9187 VPWR.t1657 VPWR.t358 486.048
R9188 VPWR.t974 VPWR.t93 486.048
R9189 VPWR.t837 VPWR.t224 486.048
R9190 VPWR.t1404 VPWR.t353 486.048
R9191 VPWR.t1640 VPWR.t9 486.048
R9192 VPWR.t1223 VPWR.t119 486.048
R9193 VPWR.t274 VPWR.t690 486.048
R9194 VPWR.t1794 VPWR.t276 486.048
R9195 VPWR.t124 VPWR.t854 486.048
R9196 VPWR.t1483 VPWR.t154 486.048
R9197 VPWR.t272 VPWR.t1788 486.048
R9198 VPWR.t23 VPWR.t1106 486.048
R9199 VPWR.t39 VPWR.t1170 486.048
R9200 VPWR.t286 VPWR.t449 486.048
R9201 VPWR.t862 VPWR.t304 486.048
R9202 VPWR.t342 VPWR.t764 486.048
R9203 VPWR.t299 VPWR.t174 486.048
R9204 VPWR.t159 VPWR.t28 486.048
R9205 VPWR.t288 VPWR.t164 486.048
R9206 VPWR.t294 VPWR.t306 486.048
R9207 VPWR.t68 VPWR.t334 486.048
R9208 VPWR.t58 VPWR.t176 486.048
R9209 VPWR.t331 VPWR.t202 486.048
R9210 VPWR.t226 VPWR.t55 486.048
R9211 VPWR.t90 VPWR.t63 486.048
R9212 VPWR.t98 VPWR.t218 486.048
R9213 VPWR.t328 VPWR.t200 486.048
R9214 VPWR.t361 VPWR.t95 486.048
R9215 VPWR.t113 VPWR.t380 486.048
R9216 VPWR.t234 VPWR.t241 486.048
R9217 VPWR.t374 VPWR.t253 486.048
R9218 VPWR.t278 VPWR.t14 486.048
R9219 VPWR.t250 VPWR.t129 486.048
R9220 VPWR.t30 VPWR.t302 486.048
R9221 VPWR.t44 VPWR.t166 486.048
R9222 VPWR.t179 VPWR.t172 486.048
R9223 VPWR.t339 VPWR.t213 486.048
R9224 VPWR.t60 VPWR.t321 486.048
R9225 VPWR.t88 VPWR.t207 486.048
R9226 VPWR.t103 VPWR.t315 486.048
R9227 VPWR.t326 VPWR.t355 486.048
R9228 VPWR.t369 VPWR.t100 486.048
R9229 VPWR.t86 VPWR.t204 486.048
R9230 VPWR.t239 VPWR.t363 486.048
R9231 VPWR.t261 VPWR.t382 486.048
R9232 VPWR.t111 VPWR.t126 486.048
R9233 VPWR.t137 VPWR.t255 486.048
R9234 VPWR.t162 VPWR.t283 486.048
R9235 VPWR.t134 VPWR.t7 486.048
R9236 VPWR.t1097 VPWR.t1437 463.954
R9237 VPWR.t1623 VPWR.t710 463.954
R9238 VPWR.t841 VPWR.t1645 463.954
R9239 VPWR.t1644 VPWR.t1406 463.954
R9240 VPWR.t1027 VPWR.t1096 463.954
R9241 VPWR.t800 VPWR.t1567 463.954
R9242 VPWR.t963 VPWR.t799 463.954
R9243 VPWR.t1095 VPWR.t736 463.954
R9244 VPWR.t858 VPWR.t1625 463.954
R9245 VPWR.t801 VPWR.t479 463.954
R9246 VPWR.t664 VPWR.t1643 463.954
R9247 VPWR.t1642 VPWR.t1577 463.954
R9248 VPWR.t471 VPWR.t798 463.954
R9249 VPWR.t797 VPWR.t453 463.954
R9250 VPWR.t1491 VPWR.t1646 463.954
R9251 VPWR.t1624 VPWR.t694 463.954
R9252 VPWR.t1233 VPWR.t1427 463.954
R9253 VPWR.t1126 VPWR.t1554 463.954
R9254 VPWR.t419 VPWR.t1237 463.954
R9255 VPWR.t1382 VPWR.t1236 463.954
R9256 VPWR.t1057 VPWR.t1558 463.954
R9257 VPWR.t827 VPWR.t1452 463.954
R9258 VPWR.t708 VPWR.t1451 463.954
R9259 VPWR.t716 VPWR.t1557 463.954
R9260 VPWR.t1108 VPWR.t1556 463.954
R9261 VPWR.t1012 VPWR.t1453 463.954
R9262 VPWR.t1832 VPWR.t1235 463.954
R9263 VPWR.t1045 VPWR.t1234 463.954
R9264 VPWR.t1195 VPWR.t1450 463.954
R9265 VPWR.t815 VPWR.t1449 463.954
R9266 VPWR.t1466 VPWR.t1238 463.954
R9267 VPWR.t622 VPWR.t1555 463.954
R9268 VPWR.t1274 VPWR.t1412 463.954
R9269 VPWR.t533 VPWR.t1221 463.954
R9270 VPWR.t430 VPWR.t1597 463.954
R9271 VPWR.t1360 VPWR.t429 463.954
R9272 VPWR.t1273 VPWR.t1632 463.954
R9273 VPWR.t1513 VPWR.t1219 463.954
R9274 VPWR.t1218 VPWR.t559 463.954
R9275 VPWR.t1800 VPWR.t1272 463.954
R9276 VPWR.t1271 VPWR.t905 463.954
R9277 VPWR.t951 VPWR.t1220 463.954
R9278 VPWR.t428 VPWR.t612 463.954
R9279 VPWR.t1680 VPWR.t427 463.954
R9280 VPWR.t1217 VPWR.t1762 463.954
R9281 VPWR.t1700 VPWR.t1216 463.954
R9282 VPWR.t1215 VPWR.t939 463.954
R9283 VPWR.t756 VPWR.t1222 463.954
R9284 VPWR.t1446 VPWR.t1420 463.954
R9285 VPWR.t1441 VPWR.t1152 463.954
R9286 VPWR.t607 VPWR.t1609 463.954
R9287 VPWR.t606 VPWR.t1374 463.954
R9288 VPWR.t1445 VPWR.t1063 463.954
R9289 VPWR.t1168 VPWR.t1544 463.954
R9290 VPWR.t1167 VPWR.t543 463.954
R9291 VPWR.t1444 VPWR.t726 463.954
R9292 VPWR.t1443 VPWR.t1018 463.954
R9293 VPWR.t1169 VPWR.t1918 463.954
R9294 VPWR.t1448 VPWR.t640 463.954
R9295 VPWR.t1447 VPWR.t1055 463.954
R9296 VPWR.t1166 VPWR.t1181 463.954
R9297 VPWR.t1165 VPWR.t922 463.954
R9298 VPWR.t1164 VPWR.t680 463.954
R9299 VPWR.t1442 VPWR.t628 463.954
R9300 VPWR.t1506 VPWR.t1433 463.954
R9301 VPWR.t921 VPWR.t1724 463.954
R9302 VPWR.t1583 VPWR.t496 463.954
R9303 VPWR.t495 VPWR.t1394 463.954
R9304 VPWR.t802 VPWR.t1505 463.954
R9305 VPWR.t1565 VPWR.t1666 463.954
R9306 VPWR.t591 VPWR.t1005 463.954
R9307 VPWR.t826 VPWR.t1898 463.954
R9308 VPWR.t577 VPWR.t825 463.954
R9309 VPWR.t1566 VPWR.t1599 463.954
R9310 VPWR.t1820 VPWR.t1508 463.954
R9311 VPWR.t1507 VPWR.t553 463.954
R9312 VPWR.t1205 VPWR.t1004 463.954
R9313 VPWR.t1003 VPWR.t805 463.954
R9314 VPWR.t997 VPWR.t497 463.954
R9315 VPWR.t824 VPWR.t1808 463.954
R9316 VPWR.t600 VPWR.t1439 463.954
R9317 VPWR.t901 VPWR.t732 463.954
R9318 VPWR.t839 VPWR.t605 463.954
R9319 VPWR.t1408 VPWR.t604 463.954
R9320 VPWR.t1025 VPWR.t599 463.954
R9321 VPWR.t521 VPWR.t1043 463.954
R9322 VPWR.t961 VPWR.t1042 463.954
R9323 VPWR.t734 VPWR.t598 463.954
R9324 VPWR.t856 VPWR.t1712 463.954
R9325 VPWR.t477 VPWR.t1044 463.954
R9326 VPWR.t662 VPWR.t603 463.954
R9327 VPWR.t1575 VPWR.t602 463.954
R9328 VPWR.t469 VPWR.t1041 463.954
R9329 VPWR.t451 VPWR.t1040 463.954
R9330 VPWR.t1784 VPWR.t1039 463.954
R9331 VPWR.t692 VPWR.t733 463.954
R9332 VPWR.t789 VPWR.t1435 463.954
R9333 VPWR.t829 VPWR.t1078 463.954
R9334 VPWR.t793 VPWR.t1521 463.954
R9335 VPWR.t1402 VPWR.t792 463.954
R9336 VPWR.t788 VPWR.t1029 463.954
R9337 VPWR.t1573 VPWR.t1076 463.954
R9338 VPWR.t1075 VPWR.t969 463.954
R9339 VPWR.t1894 VPWR.t787 463.954
R9340 VPWR.t786 VPWR.t981 463.954
R9341 VPWR.t1118 VPWR.t1077 463.954
R9342 VPWR.t791 VPWR.t670 463.954
R9343 VPWR.t549 VPWR.t790 463.954
R9344 VPWR.t1074 VPWR.t1756 463.954
R9345 VPWR.t455 VPWR.t1073 463.954
R9346 VPWR.t794 VPWR.t1615 463.954
R9347 VPWR.t696 VPWR.t785 463.954
R9348 VPWR.t1753 VPWR.t1414 463.954
R9349 VPWR.t1748 VPWR.t531 463.954
R9350 VPWR.t1771 VPWR.t1595 463.954
R9351 VPWR.t1770 VPWR.t1362 463.954
R9352 VPWR.t1752 VPWR.t1628 463.954
R9353 VPWR.t1776 VPWR.t1511 463.954
R9354 VPWR.t1775 VPWR.t557 463.954
R9355 VPWR.t1751 VPWR.t1798 463.954
R9356 VPWR.t1750 VPWR.t919 463.954
R9357 VPWR.t1777 VPWR.t847 463.954
R9358 VPWR.t1769 VPWR.t610 463.954
R9359 VPWR.t1768 VPWR.t1213 463.954
R9360 VPWR.t1774 VPWR.t1760 463.954
R9361 VPWR.t1773 VPWR.t1696 463.954
R9362 VPWR.t1772 VPWR.t937 463.954
R9363 VPWR.t1749 VPWR.t752 463.954
R9364 VPWR.t1846 VPWR.t1431 463.954
R9365 VPWR.t852 VPWR.t1726 463.954
R9366 VPWR.t1585 VPWR.t1836 463.954
R9367 VPWR.t1849 VPWR.t1392 463.954
R9368 VPWR.t1851 VPWR.t1845 463.954
R9369 VPWR.t1841 VPWR.t1534 463.954
R9370 VPWR.t593 VPWR.t1840 463.954
R9371 VPWR.t1844 VPWR.t1900 463.954
R9372 VPWR.t864 VPWR.t1843 463.954
R9373 VPWR.t1842 VPWR.t1601 463.954
R9374 VPWR.t1822 VPWR.t1848 463.954
R9375 VPWR.t1847 VPWR.t1471 463.954
R9376 VPWR.t1207 VPWR.t1839 463.954
R9377 VPWR.t1838 VPWR.t807 463.954
R9378 VPWR.t999 VPWR.t1837 463.954
R9379 VPWR.t853 VPWR.t1810 463.954
R9380 VPWR.t1652 VPWR.t1416 463.954
R9381 VPWR.t529 VPWR.t1647 463.954
R9382 VPWR.t1593 VPWR.t391 463.954
R9383 VPWR.t1364 VPWR.t390 463.954
R9384 VPWR.t1626 VPWR.t1651 463.954
R9385 VPWR.t1509 VPWR.t1529 463.954
R9386 VPWR.t555 VPWR.t1528 463.954
R9387 VPWR.t1796 VPWR.t1650 463.954
R9388 VPWR.t915 VPWR.t1649 463.954
R9389 VPWR.t845 VPWR.t1530 463.954
R9390 VPWR.t608 VPWR.t389 463.954
R9391 VPWR.t1211 VPWR.t388 463.954
R9392 VPWR.t1172 VPWR.t1527 463.954
R9393 VPWR.t1692 VPWR.t1526 463.954
R9394 VPWR.t935 VPWR.t1525 463.954
R9395 VPWR.t750 VPWR.t1648 463.954
R9396 VPWR.t1673 VPWR.t1429 463.954
R9397 VPWR.t1225 VPWR.t1728 463.954
R9398 VPWR.t1230 VPWR.t1587 463.954
R9399 VPWR.t1229 VPWR.t1390 463.954
R9400 VPWR.t1672 VPWR.t1855 463.954
R9401 VPWR.t1677 VPWR.t1536 463.954
R9402 VPWR.t1676 VPWR.t595 463.954
R9403 VPWR.t1671 VPWR.t1902 463.954
R9404 VPWR.t1227 VPWR.t866 463.954
R9405 VPWR.t1678 VPWR.t1603 463.954
R9406 VPWR.t1228 VPWR.t1824 463.954
R9407 VPWR.t1674 VPWR.t1473 463.954
R9408 VPWR.t1675 VPWR.t1239 463.954
R9409 VPWR.t1232 VPWR.t809 463.954
R9410 VPWR.t1231 VPWR.t1001 463.954
R9411 VPWR.t1226 VPWR.t1814 463.954
R9412 VPWR.t1487 VPWR.t1422 463.954
R9413 VPWR.t1739 VPWR.t434 463.954
R9414 VPWR.t1202 VPWR.t425 463.954
R9415 VPWR.t1376 VPWR.t1490 463.954
R9416 VPWR.t1486 VPWR.t1061 463.954
R9417 VPWR.t1717 VPWR.t432 463.954
R9418 VPWR.t431 VPWR.t539 463.954
R9419 VPWR.t722 VPWR.t1485 463.954
R9420 VPWR.t436 VPWR.t1016 463.954
R9421 VPWR.t1914 VPWR.t433 463.954
R9422 VPWR.t1489 VPWR.t638 463.954
R9423 VPWR.t1051 VPWR.t1488 463.954
R9424 VPWR.t1456 VPWR.t1179 463.954
R9425 VPWR.t821 VPWR.t1455 463.954
R9426 VPWR.t1454 VPWR.t678 463.954
R9427 VPWR.t626 VPWR.t435 463.954
R9428 VPWR.t1279 VPWR.t1418 463.954
R9429 VPWR.t1154 VPWR.t1663 463.954
R9430 VPWR.t498 VPWR.t1611 463.954
R9431 VPWR.t1372 VPWR.t1533 463.954
R9432 VPWR.t1278 VPWR.t1067 463.954
R9433 VPWR.t1546 VPWR.t1661 463.954
R9434 VPWR.t1660 VPWR.t545 463.954
R9435 VPWR.t728 VPWR.t1277 463.954
R9436 VPWR.t1276 VPWR.t1020 463.954
R9437 VPWR.t1920 VPWR.t1662 463.954
R9438 VPWR.t1532 VPWR.t642 463.954
R9439 VPWR.t1098 VPWR.t1531 463.954
R9440 VPWR.t501 VPWR.t1183 463.954
R9441 VPWR.t924 VPWR.t500 463.954
R9442 VPWR.t499 VPWR.t682 463.954
R9443 VPWR.t632 VPWR.t1275 463.954
R9444 VPWR.t1260 VPWR.t1410 463.954
R9445 VPWR.t481 VPWR.t893 463.954
R9446 VPWR.t525 VPWR.t1084 463.954
R9447 VPWR.t524 VPWR.t1354 463.954
R9448 VPWR.t796 VPWR.t1638 463.954
R9449 VPWR.t948 VPWR.t515 463.954
R9450 VPWR.t947 VPWR.t565 463.954
R9451 VPWR.t795 VPWR.t740 463.954
R9452 VPWR.t483 VPWR.t909 463.954
R9453 VPWR.t949 VPWR.t957 463.954
R9454 VPWR.t523 VPWR.t614 463.954
R9455 VPWR.t1261 VPWR.t1686 463.954
R9456 VPWR.t946 VPWR.t1764 463.954
R9457 VPWR.t945 VPWR.t1704 463.954
R9458 VPWR.t526 VPWR.t1174 463.954
R9459 VPWR.t482 VPWR.t762 463.954
R9460 VPWR.t1877 VPWR.t1425 463.954
R9461 VPWR.t1128 VPWR.t1656 463.954
R9462 VPWR.t421 VPWR.t1881 463.954
R9463 VPWR.t1380 VPWR.t1880 463.954
R9464 VPWR.t1059 VPWR.t1876 463.954
R9465 VPWR.t1713 VPWR.t1654 463.954
R9466 VPWR.t535 VPWR.t1653 463.954
R9467 VPWR.t718 VPWR.t1659 463.954
R9468 VPWR.t1112 VPWR.t1658 463.954
R9469 VPWR.t1014 VPWR.t1655 463.954
R9470 VPWR.t1834 VPWR.t1879 463.954
R9471 VPWR.t1047 VPWR.t1878 463.954
R9472 VPWR.t1197 VPWR.t1194 463.954
R9473 VPWR.t819 VPWR.t1193 463.954
R9474 VPWR.t1468 VPWR.t804 463.954
R9475 VPWR.t624 VPWR.t1657 463.954
R9476 VPWR.t93 VPWR.t108 463.954
R9477 VPWR.t224 VPWR.t269 463.954
R9478 VPWR.t353 VPWR.t371 463.954
R9479 VPWR.t9 VPWR.t142 463.954
R9480 VPWR.t119 VPWR.t244 463.954
R9481 VPWR.t266 VPWR.t274 463.954
R9482 VPWR.t276 VPWR.t17 463.954
R9483 VPWR.t139 VPWR.t124 463.954
R9484 VPWR.t154 VPWR.t280 463.954
R9485 VPWR.t296 VPWR.t272 463.954
R9486 VPWR.t36 VPWR.t23 463.954
R9487 VPWR.t169 VPWR.t39 463.954
R9488 VPWR.t210 VPWR.t286 463.954
R9489 VPWR.t304 VPWR.t46 463.954
R9490 VPWR.t83 VPWR.t342 463.954
R9491 VPWR.t174 VPWR.t191 463.954
R9492 VPWR.t28 VPWR.t52 463.954
R9493 VPWR.t164 VPWR.t197 463.954
R9494 VPWR.t309 VPWR.t294 463.954
R9495 VPWR.t334 VPWR.t74 463.954
R9496 VPWR.t182 VPWR.t58 463.954
R9497 VPWR.t202 VPWR.t194 463.954
R9498 VPWR.t350 VPWR.t226 463.954
R9499 VPWR.t63 VPWR.t71 463.954
R9500 VPWR.t231 VPWR.t98 463.954
R9501 VPWR.t200 VPWR.t247 463.954
R9502 VPWR.t377 VPWR.t361 463.954
R9503 VPWR.t380 VPWR.t121 463.954
R9504 VPWR.t151 VPWR.t234 463.954
R9505 VPWR.t253 VPWR.t1 463.954
R9506 VPWR.t20 VPWR.t278 463.954
R9507 VPWR.t129 VPWR.t145 463.954
R9508 VPWR.t302 VPWR.t312 463.954
R9509 VPWR.t80 VPWR.t44 463.954
R9510 VPWR.t172 VPWR.t185 463.954
R9511 VPWR.t213 VPWR.t347 463.954
R9512 VPWR.t321 VPWR.t65 463.954
R9513 VPWR.t77 VPWR.t88 463.954
R9514 VPWR.t236 VPWR.t103 463.954
R9515 VPWR.t344 VPWR.t326 463.954
R9516 VPWR.t105 VPWR.t369 463.954
R9517 VPWR.t131 VPWR.t86 463.954
R9518 VPWR.t258 VPWR.t239 463.954
R9519 VPWR.t4 VPWR.t261 463.954
R9520 VPWR.t25 VPWR.t111 463.954
R9521 VPWR.t263 VPWR.t137 463.954
R9522 VPWR.t291 VPWR.t162 463.954
R9523 VPWR.t7 VPWR.t11 463.954
R9524 VPWR.n2626 VPWR.t1140 428.822
R9525 VPWR.n1595 VPWR.n1594 376.045
R9526 VPWR.n2506 VPWR.n2505 376.045
R9527 VPWR.n1468 VPWR.n1467 376.045
R9528 VPWR.n351 VPWR.n350 376.045
R9529 VPWR.n2568 VPWR.n2567 376.045
R9530 VPWR.n1535 VPWR.n1534 376.045
R9531 VPWR.n349 VPWR.n348 376.045
R9532 VPWR.n2508 VPWR.n2507 376.045
R9533 VPWR.n966 VPWR.n965 376.045
R9534 VPWR.n2478 VPWR.n2477 376.045
R9535 VPWR.n2476 VPWR.n2475 376.045
R9536 VPWR.n321 VPWR.n320 376.045
R9537 VPWR.n2554 VPWR.n2553 376.045
R9538 VPWR.n974 VPWR.n973 376.045
R9539 VPWR.n2446 VPWR.n2445 376.045
R9540 VPWR.n325 VPWR.n324 376.045
R9541 VPWR.n2544 VPWR.n2543 376.045
R9542 VPWR.n1890 VPWR.n1889 376.045
R9543 VPWR.n1888 VPWR.n1887 376.045
R9544 VPWR.n1880 VPWR.n1879 376.045
R9545 VPWR.n390 VPWR.n389 376.045
R9546 VPWR.n394 VPWR.n393 376.045
R9547 VPWR.n398 VPWR.n397 376.045
R9548 VPWR.n2456 VPWR.n2455 376.045
R9549 VPWR.n333 VPWR.n332 376.045
R9550 VPWR.n2532 VPWR.n2531 376.045
R9551 VPWR.n1878 VPWR.n1877 376.045
R9552 VPWR.n406 VPWR.n405 376.045
R9553 VPWR.n2458 VPWR.n2457 376.045
R9554 VPWR.n337 VPWR.n336 376.045
R9555 VPWR.n2530 VPWR.n2529 376.045
R9556 VPWR.n2309 VPWR.n2308 376.045
R9557 VPWR.n2311 VPWR.n2310 376.045
R9558 VPWR.n2319 VPWR.n2318 376.045
R9559 VPWR.n2321 VPWR.n2320 376.045
R9560 VPWR.n2331 VPWR.n2330 376.045
R9561 VPWR.n2339 VPWR.n2338 376.045
R9562 VPWR.n2341 VPWR.n2340 376.045
R9563 VPWR.n2349 VPWR.n2348 376.045
R9564 VPWR.n2351 VPWR.n2350 376.045
R9565 VPWR.n2359 VPWR.n2358 376.045
R9566 VPWR.n2361 VPWR.n2360 376.045
R9567 VPWR.n2369 VPWR.n2368 376.045
R9568 VPWR.n2371 VPWR.n2370 376.045
R9569 VPWR.n2379 VPWR.n2378 376.045
R9570 VPWR.n2329 VPWR.n2328 376.045
R9571 VPWR.n543 VPWR.n542 376.045
R9572 VPWR.n541 VPWR.n540 376.045
R9573 VPWR.n537 VPWR.n536 376.045
R9574 VPWR.n533 VPWR.n532 376.045
R9575 VPWR.n525 VPWR.n524 376.045
R9576 VPWR.n521 VPWR.n520 376.045
R9577 VPWR.n517 VPWR.n516 376.045
R9578 VPWR.n513 VPWR.n512 376.045
R9579 VPWR.n509 VPWR.n508 376.045
R9580 VPWR.n505 VPWR.n504 376.045
R9581 VPWR.n501 VPWR.n500 376.045
R9582 VPWR.n497 VPWR.n496 376.045
R9583 VPWR.n493 VPWR.n492 376.045
R9584 VPWR.n489 VPWR.n488 376.045
R9585 VPWR.n529 VPWR.n528 376.045
R9586 VPWR.n2282 VPWR.n2281 376.045
R9587 VPWR.n2280 VPWR.n2279 376.045
R9588 VPWR.n2272 VPWR.n2271 376.045
R9589 VPWR.n2270 VPWR.n2269 376.045
R9590 VPWR.n2260 VPWR.n2259 376.045
R9591 VPWR.n2252 VPWR.n2251 376.045
R9592 VPWR.n2250 VPWR.n2249 376.045
R9593 VPWR.n2242 VPWR.n2241 376.045
R9594 VPWR.n2240 VPWR.n2239 376.045
R9595 VPWR.n2232 VPWR.n2231 376.045
R9596 VPWR.n2230 VPWR.n2229 376.045
R9597 VPWR.n2222 VPWR.n2221 376.045
R9598 VPWR.n2220 VPWR.n2219 376.045
R9599 VPWR.n2212 VPWR.n2211 376.045
R9600 VPWR.n2262 VPWR.n2261 376.045
R9601 VPWR.n582 VPWR.n581 376.045
R9602 VPWR.n586 VPWR.n585 376.045
R9603 VPWR.n590 VPWR.n589 376.045
R9604 VPWR.n594 VPWR.n593 376.045
R9605 VPWR.n602 VPWR.n601 376.045
R9606 VPWR.n606 VPWR.n605 376.045
R9607 VPWR.n610 VPWR.n609 376.045
R9608 VPWR.n614 VPWR.n613 376.045
R9609 VPWR.n618 VPWR.n617 376.045
R9610 VPWR.n622 VPWR.n621 376.045
R9611 VPWR.n626 VPWR.n625 376.045
R9612 VPWR.n630 VPWR.n629 376.045
R9613 VPWR.n634 VPWR.n633 376.045
R9614 VPWR.n638 VPWR.n637 376.045
R9615 VPWR.n598 VPWR.n597 376.045
R9616 VPWR.n2113 VPWR.n2112 376.045
R9617 VPWR.n2115 VPWR.n2114 376.045
R9618 VPWR.n2123 VPWR.n2122 376.045
R9619 VPWR.n2125 VPWR.n2124 376.045
R9620 VPWR.n2135 VPWR.n2134 376.045
R9621 VPWR.n2143 VPWR.n2142 376.045
R9622 VPWR.n2145 VPWR.n2144 376.045
R9623 VPWR.n2153 VPWR.n2152 376.045
R9624 VPWR.n2155 VPWR.n2154 376.045
R9625 VPWR.n2163 VPWR.n2162 376.045
R9626 VPWR.n2165 VPWR.n2164 376.045
R9627 VPWR.n2173 VPWR.n2172 376.045
R9628 VPWR.n2175 VPWR.n2174 376.045
R9629 VPWR.n2183 VPWR.n2182 376.045
R9630 VPWR.n2133 VPWR.n2132 376.045
R9631 VPWR.n735 VPWR.n734 376.045
R9632 VPWR.n733 VPWR.n732 376.045
R9633 VPWR.n729 VPWR.n728 376.045
R9634 VPWR.n725 VPWR.n724 376.045
R9635 VPWR.n717 VPWR.n716 376.045
R9636 VPWR.n713 VPWR.n712 376.045
R9637 VPWR.n709 VPWR.n708 376.045
R9638 VPWR.n705 VPWR.n704 376.045
R9639 VPWR.n701 VPWR.n700 376.045
R9640 VPWR.n697 VPWR.n696 376.045
R9641 VPWR.n693 VPWR.n692 376.045
R9642 VPWR.n689 VPWR.n688 376.045
R9643 VPWR.n685 VPWR.n684 376.045
R9644 VPWR.n681 VPWR.n680 376.045
R9645 VPWR.n721 VPWR.n720 376.045
R9646 VPWR.n2086 VPWR.n2085 376.045
R9647 VPWR.n2084 VPWR.n2083 376.045
R9648 VPWR.n2076 VPWR.n2075 376.045
R9649 VPWR.n2074 VPWR.n2073 376.045
R9650 VPWR.n2064 VPWR.n2063 376.045
R9651 VPWR.n2056 VPWR.n2055 376.045
R9652 VPWR.n2054 VPWR.n2053 376.045
R9653 VPWR.n2046 VPWR.n2045 376.045
R9654 VPWR.n2044 VPWR.n2043 376.045
R9655 VPWR.n2036 VPWR.n2035 376.045
R9656 VPWR.n2034 VPWR.n2033 376.045
R9657 VPWR.n2026 VPWR.n2025 376.045
R9658 VPWR.n2024 VPWR.n2023 376.045
R9659 VPWR.n2016 VPWR.n2015 376.045
R9660 VPWR.n2066 VPWR.n2065 376.045
R9661 VPWR.n774 VPWR.n773 376.045
R9662 VPWR.n778 VPWR.n777 376.045
R9663 VPWR.n782 VPWR.n781 376.045
R9664 VPWR.n786 VPWR.n785 376.045
R9665 VPWR.n794 VPWR.n793 376.045
R9666 VPWR.n798 VPWR.n797 376.045
R9667 VPWR.n802 VPWR.n801 376.045
R9668 VPWR.n806 VPWR.n805 376.045
R9669 VPWR.n810 VPWR.n809 376.045
R9670 VPWR.n814 VPWR.n813 376.045
R9671 VPWR.n818 VPWR.n817 376.045
R9672 VPWR.n822 VPWR.n821 376.045
R9673 VPWR.n826 VPWR.n825 376.045
R9674 VPWR.n830 VPWR.n829 376.045
R9675 VPWR.n790 VPWR.n789 376.045
R9676 VPWR.n1917 VPWR.n1916 376.045
R9677 VPWR.n1919 VPWR.n1918 376.045
R9678 VPWR.n1927 VPWR.n1926 376.045
R9679 VPWR.n1929 VPWR.n1928 376.045
R9680 VPWR.n1939 VPWR.n1938 376.045
R9681 VPWR.n1947 VPWR.n1946 376.045
R9682 VPWR.n1949 VPWR.n1948 376.045
R9683 VPWR.n1957 VPWR.n1956 376.045
R9684 VPWR.n1959 VPWR.n1958 376.045
R9685 VPWR.n1967 VPWR.n1966 376.045
R9686 VPWR.n1969 VPWR.n1968 376.045
R9687 VPWR.n1977 VPWR.n1976 376.045
R9688 VPWR.n1979 VPWR.n1978 376.045
R9689 VPWR.n1987 VPWR.n1986 376.045
R9690 VPWR.n1937 VPWR.n1936 376.045
R9691 VPWR.n927 VPWR.n926 376.045
R9692 VPWR.n925 VPWR.n924 376.045
R9693 VPWR.n921 VPWR.n920 376.045
R9694 VPWR.n917 VPWR.n916 376.045
R9695 VPWR.n909 VPWR.n908 376.045
R9696 VPWR.n905 VPWR.n904 376.045
R9697 VPWR.n901 VPWR.n900 376.045
R9698 VPWR.n897 VPWR.n896 376.045
R9699 VPWR.n893 VPWR.n892 376.045
R9700 VPWR.n889 VPWR.n888 376.045
R9701 VPWR.n885 VPWR.n884 376.045
R9702 VPWR.n881 VPWR.n880 376.045
R9703 VPWR.n877 VPWR.n876 376.045
R9704 VPWR.n873 VPWR.n872 376.045
R9705 VPWR.n913 VPWR.n912 376.045
R9706 VPWR.n1870 VPWR.n1869 376.045
R9707 VPWR.n982 VPWR.n981 376.045
R9708 VPWR.n1494 VPWR.n1493 376.045
R9709 VPWR.n1221 VPWR.n1220 376.045
R9710 VPWR.n402 VPWR.n401 376.045
R9711 VPWR.n2466 VPWR.n2465 376.045
R9712 VPWR.n341 VPWR.n340 376.045
R9713 VPWR.n2520 VPWR.n2519 376.045
R9714 VPWR.n978 VPWR.n977 376.045
R9715 VPWR.n1492 VPWR.n1491 376.045
R9716 VPWR.n1185 VPWR.n1184 376.045
R9717 VPWR.n1868 VPWR.n1867 376.045
R9718 VPWR.n986 VPWR.n985 376.045
R9719 VPWR.n1506 VPWR.n1505 376.045
R9720 VPWR.n1219 VPWR.n1218 376.045
R9721 VPWR.n410 VPWR.n409 376.045
R9722 VPWR.n418 VPWR.n417 376.045
R9723 VPWR.n422 VPWR.n421 376.045
R9724 VPWR.n426 VPWR.n425 376.045
R9725 VPWR.n430 VPWR.n429 376.045
R9726 VPWR.n434 VPWR.n433 376.045
R9727 VPWR.n438 VPWR.n437 376.045
R9728 VPWR.n442 VPWR.n441 376.045
R9729 VPWR.n446 VPWR.n445 376.045
R9730 VPWR.n414 VPWR.n413 376.045
R9731 VPWR.n2448 VPWR.n2447 376.045
R9732 VPWR.n329 VPWR.n328 376.045
R9733 VPWR.n2542 VPWR.n2541 376.045
R9734 VPWR.n990 VPWR.n989 376.045
R9735 VPWR.n1508 VPWR.n1507 376.045
R9736 VPWR.n1216 VPWR.n1215 376.045
R9737 VPWR.n1860 VPWR.n1859 376.045
R9738 VPWR.n1850 VPWR.n1849 376.045
R9739 VPWR.n1848 VPWR.n1847 376.045
R9740 VPWR.n1840 VPWR.n1839 376.045
R9741 VPWR.n1838 VPWR.n1837 376.045
R9742 VPWR.n1830 VPWR.n1829 376.045
R9743 VPWR.n1828 VPWR.n1827 376.045
R9744 VPWR.n1820 VPWR.n1819 376.045
R9745 VPWR.n1858 VPWR.n1857 376.045
R9746 VPWR.n994 VPWR.n993 376.045
R9747 VPWR.n1520 VPWR.n1519 376.045
R9748 VPWR.n1213 VPWR.n1212 376.045
R9749 VPWR.n2468 VPWR.n2467 376.045
R9750 VPWR.n345 VPWR.n344 376.045
R9751 VPWR.n2518 VPWR.n2517 376.045
R9752 VPWR.n1481 VPWR.n1480 376.045
R9753 VPWR.n1182 VPWR.n1181 376.045
R9754 VPWR.n998 VPWR.n997 376.045
R9755 VPWR.n1522 VPWR.n1521 376.045
R9756 VPWR.n1205 VPWR.n1204 376.045
R9757 VPWR.n2438 VPWR.n2437 376.045
R9758 VPWR.n2428 VPWR.n2427 376.045
R9759 VPWR.n2426 VPWR.n2425 376.045
R9760 VPWR.n2418 VPWR.n2417 376.045
R9761 VPWR.n2416 VPWR.n2415 376.045
R9762 VPWR.n2408 VPWR.n2407 376.045
R9763 VPWR.n2436 VPWR.n2435 376.045
R9764 VPWR.n317 VPWR.n316 376.045
R9765 VPWR.n2556 VPWR.n2555 376.045
R9766 VPWR.n1537 VPWR.n1536 376.045
R9767 VPWR.n1202 VPWR.n1201 376.045
R9768 VPWR.n1002 VPWR.n1001 376.045
R9769 VPWR.n1006 VPWR.n1005 376.045
R9770 VPWR.n1010 VPWR.n1009 376.045
R9771 VPWR.n1014 VPWR.n1013 376.045
R9772 VPWR.n1018 VPWR.n1017 376.045
R9773 VPWR.n1022 VPWR.n1021 376.045
R9774 VPWR.n970 VPWR.n969 376.045
R9775 VPWR.n1475 VPWR.n1474 376.045
R9776 VPWR.n1593 VPWR.n1592 376.045
R9777 VPWR.n313 VPWR.n312 376.045
R9778 VPWR.n2566 VPWR.n2565 376.045
R9779 VPWR.n1199 VPWR.n1198 376.045
R9780 VPWR.n1762 VPWR.n1761 376.045
R9781 VPWR.n1191 VPWR.n1190 376.045
R9782 VPWR.n309 VPWR.n308 376.045
R9783 VPWR.n305 VPWR.n304 376.045
R9784 VPWR.n297 VPWR.n296 376.045
R9785 VPWR.n301 VPWR.n300 376.045
R9786 VPWR.n1741 VPWR.n1740 376.045
R9787 VPWR.n1750 VPWR.n1749 376.045
R9788 VPWR.n1791 VPWR.n1790 376.045
R9789 VPWR.n1760 VPWR.n1759 376.045
R9790 VPWR.n1188 VPWR.n1187 376.045
R9791 VPWR.n2578 VPWR.n2577 376.045
R9792 VPWR.n2580 VPWR.n2579 376.045
R9793 VPWR.n2590 VPWR.n2589 376.045
R9794 VPWR.n1739 VPWR.n1738 376.045
R9795 VPWR.n1339 VPWR.t876 342.841
R9796 VPWR.n1378 VPWR.t778 342.841
R9797 VPWR.n1415 VPWR.t772 342.841
R9798 VPWR.n2693 VPWR.t976 342.841
R9799 VPWR.n2656 VPWR.t884 342.841
R9800 VPWR.n2599 VPWR.t1141 342.841
R9801 VPWR.n1339 VPWR.t1867 342.839
R9802 VPWR.n1378 VPWR.t1178 342.839
R9803 VPWR.n1415 VPWR.t656 342.839
R9804 VPWR.n2693 VPWR.t403 342.839
R9805 VPWR.n2656 VPWR.t1464 342.839
R9806 VPWR.n2599 VPWR.t1248 342.839
R9807 VPWR.n2842 VPWR.n2824 339.212
R9808 VPWR.n1306 VPWR.t873 338.488
R9809 VPWR.n2729 VPWR.t1887 338.488
R9810 VPWR.n1315 VPWR.n1314 327.377
R9811 VPWR.n1308 VPWR.n1307 327.377
R9812 VPWR.n1322 VPWR.n1321 327.377
R9813 VPWR.n1352 VPWR.n1350 327.377
R9814 VPWR.n1345 VPWR.n1343 327.377
R9815 VPWR.n1360 VPWR.n1358 327.377
R9816 VPWR.n1391 VPWR.n1389 327.377
R9817 VPWR.n1384 VPWR.n1382 327.377
R9818 VPWR.n1399 VPWR.n1397 327.377
R9819 VPWR.n1428 VPWR.n1426 327.377
R9820 VPWR.n1421 VPWR.n1419 327.377
R9821 VPWR.n1436 VPWR.n1434 327.377
R9822 VPWR.n1324 VPWR.n1323 327.375
R9823 VPWR.n1352 VPWR.n1351 327.375
R9824 VPWR.n1345 VPWR.n1344 327.375
R9825 VPWR.n1360 VPWR.n1359 327.375
R9826 VPWR.n1391 VPWR.n1390 327.375
R9827 VPWR.n1384 VPWR.n1383 327.375
R9828 VPWR.n1399 VPWR.n1398 327.375
R9829 VPWR.n1428 VPWR.n1427 327.375
R9830 VPWR.n1421 VPWR.n1420 327.375
R9831 VPWR.n1436 VPWR.n1435 327.375
R9832 VPWR.n1 VPWR 325.546
R9833 VPWR.n2667 VPWR.t402 322.262
R9834 VPWR.n2630 VPWR.t883 322.262
R9835 VPWR.n2805 VPWR.n2804 321.642
R9836 VPWR.n2722 VPWR.n2712 320.976
R9837 VPWR.n2716 VPWR.n2715 320.976
R9838 VPWR.n2710 VPWR.n2709 320.976
R9839 VPWR.n2680 VPWR.n2679 320.976
R9840 VPWR.n2686 VPWR.n2675 320.976
R9841 VPWR.n2672 VPWR.n2671 320.976
R9842 VPWR.n2643 VPWR.n2642 320.976
R9843 VPWR.n2649 VPWR.n2638 320.976
R9844 VPWR.n2635 VPWR.n2634 320.976
R9845 VPWR.n2610 VPWR.n2606 320.976
R9846 VPWR.n2614 VPWR.n2613 320.976
R9847 VPWR.n2620 VPWR.n2602 320.976
R9848 VPWR.n2727 VPWR.n2708 320.976
R9849 VPWR.n2680 VPWR.n2678 320.976
R9850 VPWR.n2686 VPWR.n2674 320.976
R9851 VPWR.n2672 VPWR.n2670 320.976
R9852 VPWR.n2643 VPWR.n2641 320.976
R9853 VPWR.n2649 VPWR.n2637 320.976
R9854 VPWR.n2635 VPWR.n2633 320.976
R9855 VPWR.n2610 VPWR.n2605 320.976
R9856 VPWR.n2614 VPWR.n2612 320.976
R9857 VPWR.n2620 VPWR.n2601 320.976
R9858 VPWR.n2801 VPWR 319.627
R9859 VPWR.n6 VPWR.n5 316.245
R9860 VPWR.n1241 VPWR.n1239 316.245
R9861 VPWR.n1264 VPWR.n1262 316.245
R9862 VPWR.n1288 VPWR.n1286 316.245
R9863 VPWR.n2784 VPWR.n2783 316.245
R9864 VPWR.n2764 VPWR.n2763 316.245
R9865 VPWR.n2745 VPWR.n2744 316.245
R9866 VPWR.n1241 VPWR.n1240 316.245
R9867 VPWR.n1264 VPWR.n1263 316.245
R9868 VPWR.n1288 VPWR.n1287 316.245
R9869 VPWR.n2784 VPWR.n2782 316.245
R9870 VPWR.n2764 VPWR.n2762 316.245
R9871 VPWR.n2745 VPWR.n2743 316.245
R9872 VPWR.n2630 VPWR.t527 313.87
R9873 VPWR.n10 VPWR.n4 310.502
R9874 VPWR.n1246 VPWR.n1238 310.502
R9875 VPWR.n1269 VPWR.n1261 310.502
R9876 VPWR.n1293 VPWR.n1285 310.502
R9877 VPWR.n2803 VPWR.n2802 310.502
R9878 VPWR.n2788 VPWR.n2787 310.502
R9879 VPWR.n2768 VPWR.n2767 310.502
R9880 VPWR.n2749 VPWR.n2748 310.502
R9881 VPWR.n1246 VPWR.n1245 310.5
R9882 VPWR.n1269 VPWR.n1268 310.5
R9883 VPWR.n1293 VPWR.n1292 310.5
R9884 VPWR.n2788 VPWR.n2786 310.5
R9885 VPWR.n2768 VPWR.n2766 310.5
R9886 VPWR.n2749 VPWR.n2747 310.5
R9887 VPWR.n2834 VPWR.n2833 279.341
R9888 VPWR.n2839 VPWR.n2838 279.341
R9889 VPWR.n1412 VPWR.t1024 255.905
R9890 VPWR.n2663 VPWR.t1079 255.905
R9891 VPWR.n1275 VPWR.t508 255.904
R9892 VPWR.n1412 VPWR.t1622 255.904
R9893 VPWR.n2774 VPWR.t1735 255.904
R9894 VPWR.n2663 VPWR.t528 255.904
R9895 VPWR.n1303 VPWR.t1747 254.019
R9896 VPWR.n2735 VPWR.t944 254.019
R9897 VPWR.n1335 VPWR.t1745 252.948
R9898 VPWR.n2737 VPWR.t942 252.948
R9899 VPWR.n1373 VPWR.t971 250.722
R9900 VPWR.n2700 VPWR.t996 250.722
R9901 VPWR.n1310 VPWR.t585 249.901
R9902 VPWR.n1346 VPWR.t1869 249.901
R9903 VPWR.n1385 VPWR.t1255 249.901
R9904 VPWR.n1422 VPWR.t1871 249.901
R9905 VPWR.n2714 VPWR.t1331 249.901
R9906 VPWR.n2677 VPWR.t1328 249.901
R9907 VPWR.n2640 VPWR.t1342 249.901
R9908 VPWR.n2607 VPWR.t1296 249.901
R9909 VPWR.n1346 VPWR.t1542 249.901
R9910 VPWR.n1385 VPWR.t445 249.901
R9911 VPWR.n1422 VPWR.t932 249.901
R9912 VPWR.n2677 VPWR.t1341 249.901
R9913 VPWR.n2640 VPWR.t1294 249.901
R9914 VPWR.n2607 VPWR.t1317 249.901
R9915 VPWR.n1253 VPWR.t1093 249.363
R9916 VPWR.n1338 VPWR.t985 249.363
R9917 VPWR.n2811 VPWR.t1133 249.363
R9918 VPWR.n2795 VPWR.t774 249.363
R9919 VPWR.n2698 VPWR.t1270 249.363
R9920 VPWR.n17 VPWR.t1723 249.362
R9921 VPWR.n1253 VPWR.t1262 249.362
R9922 VPWR.n2795 VPWR.t395 249.362
R9923 VPWR.t502 VPWR.t1722 248.599
R9924 VPWR.t992 VPWR.t1497 248.599
R9925 VPWR.t1497 VPWR.t1501 248.599
R9926 VPWR.t1501 VPWR.t988 248.599
R9927 VPWR.t988 VPWR.t412 248.599
R9928 VPWR.t412 VPWR.t416 248.599
R9929 VPWR.t416 VPWR.t448 248.599
R9930 VPWR.t448 VPWR.t1873 248.599
R9931 VPWR.t1538 VPWR.t1540 248.599
R9932 VPWR.t1540 VPWR.t584 248.599
R9933 VPWR.t1344 VPWR.t1320 248.599
R9934 VPWR.t1308 VPWR.t1344 248.599
R9935 VPWR.t1282 VPWR.t1308 248.599
R9936 VPWR.t1884 VPWR.t1282 248.599
R9937 VPWR.t676 VPWR.t1884 248.599
R9938 VPWR.t491 VPWR.t676 248.599
R9939 VPWR.t417 VPWR.t491 248.599
R9940 VPWR.t1736 VPWR.t1132 248.599
R9941 VPWR.t1288 VPWR.t1330 248.599
R9942 VPWR.t1336 VPWR.t1288 248.599
R9943 VPWR.n15 VPWR.t503 247.394
R9944 VPWR.n1251 VPWR.t506 247.394
R9945 VPWR.n2809 VPWR.t1737 247.394
R9946 VPWR.n2793 VPWR.t1731 247.394
R9947 VPWR.n1251 VPWR.t504 247.394
R9948 VPWR.n2793 VPWR.t1733 247.394
R9949 VPWR.n1304 VPWR.t588 244.737
R9950 VPWR.n2730 VPWR.t1346 244.737
R9951 VPWR.n1374 VPWR.t1470 243.886
R9952 VPWR.n2701 VPWR.t850 243.886
R9953 VPWR.n1277 VPWR.t1721 243.512
R9954 VPWR.n1300 VPWR.t1094 243.512
R9955 VPWR.n1303 VPWR.t987 243.512
R9956 VPWR.n2776 VPWR.t1135 243.512
R9957 VPWR.n2756 VPWR.t775 243.512
R9958 VPWR.n2735 VPWR.t1268 243.512
R9959 VPWR.n1300 VPWR.t1263 243.512
R9960 VPWR.n2756 VPWR.t393 243.512
R9961 VPWR.n1329 VPWR.t1746 238.339
R9962 VPWR.n2705 VPWR.t943 238.339
R9963 VPWR.n2855 VPWR.t977 237.99
R9964 VPWR.n2667 VPWR.t1269 234.982
R9965 VPWR.t933 VPWR.t1538 228.101
R9966 VPWR.t1314 VPWR.t1336 228.101
R9967 VPWR.n2801 VPWR 224.923
R9968 VPWR.n1 VPWR 219.004
R9969 VPWR.n1444 VPWR.n1443 214.613
R9970 VPWR.n1444 VPWR.n1442 214.613
R9971 VPWR.n1236 VPWR.n1235 214.326
R9972 VPWR.n1259 VPWR.n1258 214.326
R9973 VPWR.n1283 VPWR.n1282 214.326
R9974 VPWR.n1368 VPWR.n1367 214.326
R9975 VPWR.n1407 VPWR.n1406 214.326
R9976 VPWR.n1236 VPWR.n1234 214.326
R9977 VPWR.n1259 VPWR.n1257 214.326
R9978 VPWR.n1283 VPWR.n1281 214.326
R9979 VPWR.n1368 VPWR.n1366 214.326
R9980 VPWR.n1407 VPWR.n1405 214.326
R9981 VPWR.n2 VPWR.n1 213.119
R9982 VPWR.n2808 VPWR.n2801 213.119
R9983 VPWR VPWR.t502 207.166
R9984 VPWR.n2840 VPWR.n2839 204.424
R9985 VPWR.n2830 VPWR.n2817 204.424
R9986 VPWR.n2833 VPWR.n2820 204.424
R9987 VPWR.n2844 VPWR.n2841 204.048
R9988 VPWR VPWR.t417 201.246
R9989 VPWR.t584 VPWR 189.409
R9990 VPWR.n2741 VPWR 184.63
R9991 VPWR.n1329 VPWR 182.952
R9992 VPWR.n2760 VPWR 182.952
R9993 VPWR.n2780 VPWR 181.273
R9994 VPWR.t527 VPWR 177.916
R9995 VPWR.n2848 VPWR.n2847 166.4
R9996 VPWR.n1770 VPWR.n1768 161.365
R9997 VPWR.n1041 VPWR.n1039 161.365
R9998 VPWR.n1545 VPWR.n1543 161.365
R9999 VPWR.n1550 VPWR.n1548 161.365
R10000 VPWR.n1555 VPWR.n1553 161.365
R10001 VPWR.n1560 VPWR.n1558 161.365
R10002 VPWR.n1565 VPWR.n1563 161.365
R10003 VPWR.n1570 VPWR.n1568 161.365
R10004 VPWR.n1575 VPWR.n1573 161.365
R10005 VPWR.n1580 VPWR.n1578 161.365
R10006 VPWR.n1135 VPWR.n1133 161.365
R10007 VPWR.n1460 VPWR.n1458 161.365
R10008 VPWR.n1455 VPWR.n1453 161.365
R10009 VPWR.n1775 VPWR.n1773 161.365
R10010 VPWR.n1783 VPWR.n1781 161.365
R10011 VPWR.n1779 VPWR.n1777 161.365
R10012 VPWR VPWR.n53 161.363
R10013 VPWR VPWR.n51 161.363
R10014 VPWR VPWR.n49 161.363
R10015 VPWR VPWR.n47 161.363
R10016 VPWR VPWR.n45 161.363
R10017 VPWR VPWR.n43 161.363
R10018 VPWR VPWR.n41 161.363
R10019 VPWR VPWR.n39 161.363
R10020 VPWR VPWR.n37 161.363
R10021 VPWR VPWR.n35 161.363
R10022 VPWR VPWR.n33 161.363
R10023 VPWR VPWR.n31 161.363
R10024 VPWR VPWR.n29 161.363
R10025 VPWR VPWR.n27 161.363
R10026 VPWR VPWR.n25 161.363
R10027 VPWR VPWR.n23 161.363
R10028 VPWR.n1115 VPWR.n1114 161.303
R10029 VPWR.n107 VPWR.n106 161.303
R10030 VPWR.n1120 VPWR.n1119 161.3
R10031 VPWR.n1599 VPWR.n1598 161.3
R10032 VPWR.n1602 VPWR.n1601 161.3
R10033 VPWR.n1111 VPWR.n1110 161.3
R10034 VPWR.n1126 VPWR.n1125 161.3
R10035 VPWR.n1107 VPWR.n1106 161.3
R10036 VPWR.n1612 VPWR.n1611 161.3
R10037 VPWR.n1615 VPWR.n1614 161.3
R10038 VPWR.n1618 VPWR.n1617 161.3
R10039 VPWR.n1623 VPWR.n1622 161.3
R10040 VPWR.n1626 VPWR.n1625 161.3
R10041 VPWR.n1629 VPWR.n1628 161.3
R10042 VPWR.n1101 VPWR.n1100 161.3
R10043 VPWR.n1177 VPWR.n1176 161.3
R10044 VPWR.n1097 VPWR.n1096 161.3
R10045 VPWR.n1639 VPWR.n1638 161.3
R10046 VPWR.n1642 VPWR.n1641 161.3
R10047 VPWR.n1645 VPWR.n1644 161.3
R10048 VPWR.n1650 VPWR.n1649 161.3
R10049 VPWR.n1653 VPWR.n1652 161.3
R10050 VPWR.n1656 VPWR.n1655 161.3
R10051 VPWR.n1091 VPWR.n1090 161.3
R10052 VPWR.n1209 VPWR.n1208 161.3
R10053 VPWR.n1087 VPWR.n1086 161.3
R10054 VPWR.n1666 VPWR.n1665 161.3
R10055 VPWR.n1669 VPWR.n1668 161.3
R10056 VPWR.n1672 VPWR.n1671 161.3
R10057 VPWR.n1677 VPWR.n1676 161.3
R10058 VPWR.n1680 VPWR.n1679 161.3
R10059 VPWR.n1683 VPWR.n1682 161.3
R10060 VPWR.n1081 VPWR.n1080 161.3
R10061 VPWR.n1195 VPWR.n1194 161.3
R10062 VPWR.n1077 VPWR.n1076 161.3
R10063 VPWR.n1693 VPWR.n1692 161.3
R10064 VPWR.n1696 VPWR.n1695 161.3
R10065 VPWR.n1699 VPWR.n1698 161.3
R10066 VPWR.n1704 VPWR.n1703 161.3
R10067 VPWR.n1707 VPWR.n1706 161.3
R10068 VPWR.n1710 VPWR.n1709 161.3
R10069 VPWR.n1070 VPWR.n1069 161.3
R10070 VPWR.n1719 VPWR.n1718 161.3
R10071 VPWR.n1722 VPWR.n1721 161.3
R10072 VPWR.n1717 VPWR.n1716 161.3
R10073 VPWR.n1734 VPWR.n1733 161.3
R10074 VPWR.n1117 VPWR.n1116 161.3
R10075 VPWR.n1731 VPWR.n1730 161.3
R10076 VPWR.n1065 VPWR.n1064 161.3
R10077 VPWR.n126 VPWR.n125 161.3
R10078 VPWR.n117 VPWR.n116 161.3
R10079 VPWR.n120 VPWR.n119 161.3
R10080 VPWR.n115 VPWR.n114 161.3
R10081 VPWR.n138 VPWR.n137 161.3
R10082 VPWR.n128 VPWR.n127 161.3
R10083 VPWR.n109 VPWR.n108 161.3
R10084 VPWR.n105 VPWR.n104 161.3
R10085 VPWR.n288 VPWR.n287 161.3
R10086 VPWR.n285 VPWR.n284 161.3
R10087 VPWR.n101 VPWR.n100 161.3
R10088 VPWR.n272 VPWR.n271 161.3
R10089 VPWR.n275 VPWR.n274 161.3
R10090 VPWR.n270 VPWR.n269 161.3
R10091 VPWR.n260 VPWR.n259 161.3
R10092 VPWR.n263 VPWR.n262 161.3
R10093 VPWR.n258 VPWR.n257 161.3
R10094 VPWR.n248 VPWR.n247 161.3
R10095 VPWR.n251 VPWR.n250 161.3
R10096 VPWR.n246 VPWR.n245 161.3
R10097 VPWR.n236 VPWR.n235 161.3
R10098 VPWR.n239 VPWR.n238 161.3
R10099 VPWR.n234 VPWR.n233 161.3
R10100 VPWR.n224 VPWR.n223 161.3
R10101 VPWR.n227 VPWR.n226 161.3
R10102 VPWR.n222 VPWR.n221 161.3
R10103 VPWR.n212 VPWR.n211 161.3
R10104 VPWR.n215 VPWR.n214 161.3
R10105 VPWR.n210 VPWR.n209 161.3
R10106 VPWR.n200 VPWR.n199 161.3
R10107 VPWR.n203 VPWR.n202 161.3
R10108 VPWR.n198 VPWR.n197 161.3
R10109 VPWR.n188 VPWR.n187 161.3
R10110 VPWR.n191 VPWR.n190 161.3
R10111 VPWR.n186 VPWR.n185 161.3
R10112 VPWR.n176 VPWR.n175 161.3
R10113 VPWR.n179 VPWR.n178 161.3
R10114 VPWR.n174 VPWR.n173 161.3
R10115 VPWR.n164 VPWR.n163 161.3
R10116 VPWR.n167 VPWR.n166 161.3
R10117 VPWR.n162 VPWR.n161 161.3
R10118 VPWR.n152 VPWR.n151 161.3
R10119 VPWR.n155 VPWR.n154 161.3
R10120 VPWR.n150 VPWR.n149 161.3
R10121 VPWR.n140 VPWR.n139 161.3
R10122 VPWR.n143 VPWR.n142 161.3
R10123 VPWR.n131 VPWR.n130 161.3
R10124 VPWR.n1601 VPWR.t43 161.202
R10125 VPWR.n1106 VPWR.t171 161.202
R10126 VPWR.n1617 VPWR.t212 161.202
R10127 VPWR.n1628 VPWR.t320 161.202
R10128 VPWR.n1096 VPWR.t87 161.202
R10129 VPWR.n1644 VPWR.t102 161.202
R10130 VPWR.n1655 VPWR.t325 161.202
R10131 VPWR.n1086 VPWR.t368 161.202
R10132 VPWR.n1671 VPWR.t85 161.202
R10133 VPWR.n1682 VPWR.t238 161.202
R10134 VPWR.n1076 VPWR.t260 161.202
R10135 VPWR.n1698 VPWR.t110 161.202
R10136 VPWR.n1709 VPWR.t136 161.202
R10137 VPWR.n1721 VPWR.t161 161.202
R10138 VPWR.n1116 VPWR.t301 161.202
R10139 VPWR.n1730 VPWR.t6 161.202
R10140 VPWR.n119 VPWR.t128 161.202
R10141 VPWR.n108 VPWR.t27 161.202
R10142 VPWR.n284 VPWR.t163 161.202
R10143 VPWR.n274 VPWR.t293 161.202
R10144 VPWR.n262 VPWR.t333 161.202
R10145 VPWR.n250 VPWR.t57 161.202
R10146 VPWR.n238 VPWR.t201 161.202
R10147 VPWR.n226 VPWR.t225 161.202
R10148 VPWR.n214 VPWR.t62 161.202
R10149 VPWR.n202 VPWR.t97 161.202
R10150 VPWR.n190 VPWR.t199 161.202
R10151 VPWR.n178 VPWR.t360 161.202
R10152 VPWR.n166 VPWR.t379 161.202
R10153 VPWR.n154 VPWR.t233 161.202
R10154 VPWR.n1768 VPWR.t285 161.202
R10155 VPWR.n1039 VPWR.t38 161.202
R10156 VPWR.n1543 VPWR.t22 161.202
R10157 VPWR.n1548 VPWR.t271 161.202
R10158 VPWR.n1553 VPWR.t153 161.202
R10159 VPWR.n1558 VPWR.t123 161.202
R10160 VPWR.n1563 VPWR.t275 161.202
R10161 VPWR.n1568 VPWR.t273 161.202
R10162 VPWR.n1573 VPWR.t118 161.202
R10163 VPWR.n1578 VPWR.t8 161.202
R10164 VPWR.n1133 VPWR.t352 161.202
R10165 VPWR.n1458 VPWR.t223 161.202
R10166 VPWR.n1453 VPWR.t92 161.202
R10167 VPWR.n1773 VPWR.t303 161.202
R10168 VPWR.n1781 VPWR.t341 161.202
R10169 VPWR.n1777 VPWR.t173 161.202
R10170 VPWR.n142 VPWR.t252 161.202
R10171 VPWR.n130 VPWR.t277 161.202
R10172 VPWR.n1119 VPWR.t29 161.106
R10173 VPWR.n1110 VPWR.t165 161.106
R10174 VPWR.n1611 VPWR.t178 161.106
R10175 VPWR.n1622 VPWR.t338 161.106
R10176 VPWR.n1100 VPWR.t59 161.106
R10177 VPWR.n1638 VPWR.t206 161.106
R10178 VPWR.n1649 VPWR.t314 161.106
R10179 VPWR.n1090 VPWR.t354 161.106
R10180 VPWR.n1665 VPWR.t99 161.106
R10181 VPWR.n1676 VPWR.t203 161.106
R10182 VPWR.n1080 VPWR.t362 161.106
R10183 VPWR.n1692 VPWR.t381 161.106
R10184 VPWR.n1703 VPWR.t125 161.106
R10185 VPWR.n1069 VPWR.t254 161.106
R10186 VPWR.n1716 VPWR.t282 161.106
R10187 VPWR.n1064 VPWR.t133 161.106
R10188 VPWR.n125 VPWR.t13 161.106
R10189 VPWR.n114 VPWR.t249 161.106
R10190 VPWR.n137 VPWR.t373 161.106
R10191 VPWR.n104 VPWR.t158 161.106
R10192 VPWR.n100 VPWR.t287 161.106
R10193 VPWR.n269 VPWR.t305 161.106
R10194 VPWR.n257 VPWR.t67 161.106
R10195 VPWR.n245 VPWR.t175 161.106
R10196 VPWR.n233 VPWR.t330 161.106
R10197 VPWR.n221 VPWR.t54 161.106
R10198 VPWR.n209 VPWR.t89 161.106
R10199 VPWR.n197 VPWR.t217 161.106
R10200 VPWR.n185 VPWR.t327 161.106
R10201 VPWR.n173 VPWR.t94 161.106
R10202 VPWR.n161 VPWR.t112 161.106
R10203 VPWR.n149 VPWR.t240 161.106
R10204 VPWR.n53 VPWR.t357 161.106
R10205 VPWR.n51 VPWR.t317 161.106
R10206 VPWR.n49 VPWR.t32 161.106
R10207 VPWR.n47 VPWR.t147 161.106
R10208 VPWR.n45 VPWR.t365 161.106
R10209 VPWR.n43 VPWR.t214 161.106
R10210 VPWR.n41 VPWR.t322 161.106
R10211 VPWR.n39 VPWR.t48 161.106
R10212 VPWR.n37 VPWR.t155 161.106
R10213 VPWR.n35 VPWR.t115 161.106
R10214 VPWR.n33 VPWR.t220 161.106
R10215 VPWR.n31 VPWR.t40 161.106
R10216 VPWR.n29 VPWR.t227 161.106
R10217 VPWR.n27 VPWR.t335 161.106
R10218 VPWR.n25 VPWR.t187 161.106
R10219 VPWR.n23 VPWR.t298 161.106
R10220 VPWR.n1598 VPWR.t79 159.978
R10221 VPWR.n1125 VPWR.t184 159.978
R10222 VPWR.n1614 VPWR.t346 159.978
R10223 VPWR.n1625 VPWR.t64 159.978
R10224 VPWR.n1176 VPWR.t76 159.978
R10225 VPWR.n1641 VPWR.t235 159.978
R10226 VPWR.n1652 VPWR.t343 159.978
R10227 VPWR.n1208 VPWR.t104 159.978
R10228 VPWR.n1668 VPWR.t130 159.978
R10229 VPWR.n1679 VPWR.t257 159.978
R10230 VPWR.n1194 VPWR.t3 159.978
R10231 VPWR.n1695 VPWR.t24 159.978
R10232 VPWR.n1706 VPWR.t262 159.978
R10233 VPWR.n1718 VPWR.t290 159.978
R10234 VPWR.n1733 VPWR.t10 159.978
R10235 VPWR.n1114 VPWR.t311 159.978
R10236 VPWR.n116 VPWR.t144 159.978
R10237 VPWR.n127 VPWR.t19 159.978
R10238 VPWR.n106 VPWR.t51 159.978
R10239 VPWR.n287 VPWR.t196 159.978
R10240 VPWR.n271 VPWR.t308 159.978
R10241 VPWR.n259 VPWR.t73 159.978
R10242 VPWR.n247 VPWR.t181 159.978
R10243 VPWR.n235 VPWR.t193 159.978
R10244 VPWR.n223 VPWR.t349 159.978
R10245 VPWR.n211 VPWR.t70 159.978
R10246 VPWR.n199 VPWR.t230 159.978
R10247 VPWR.n187 VPWR.t246 159.978
R10248 VPWR.n175 VPWR.t376 159.978
R10249 VPWR.n163 VPWR.t120 159.978
R10250 VPWR.n151 VPWR.t150 159.978
R10251 VPWR.n1228 VPWR.t107 159.978
R10252 VPWR.n1150 VPWR.t35 159.978
R10253 VPWR.n1224 VPWR.t243 159.978
R10254 VPWR.n1482 VPWR.t141 159.978
R10255 VPWR.n1170 VPWR.t265 159.978
R10256 VPWR.n1166 VPWR.t16 159.978
R10257 VPWR.n1160 VPWR.t138 159.978
R10258 VPWR.n1476 VPWR.t370 159.978
R10259 VPWR.n1156 VPWR.t279 159.978
R10260 VPWR.n1146 VPWR.t295 159.978
R10261 VPWR.n1469 VPWR.t268 159.978
R10262 VPWR.n1046 VPWR.t168 159.978
R10263 VPWR.n1745 VPWR.t45 159.978
R10264 VPWR.n1033 VPWR.t82 159.978
R10265 VPWR.n1029 VPWR.t190 159.978
R10266 VPWR.n1050 VPWR.t209 159.978
R10267 VPWR.n139 VPWR.t0 159.978
R10268 VPWR.n1229 VPWR.n1228 152
R10269 VPWR.n1151 VPWR.n1150 152
R10270 VPWR.n1225 VPWR.n1224 152
R10271 VPWR.n1483 VPWR.n1482 152
R10272 VPWR.n1171 VPWR.n1170 152
R10273 VPWR.n1167 VPWR.n1166 152
R10274 VPWR.n1161 VPWR.n1160 152
R10275 VPWR.n1477 VPWR.n1476 152
R10276 VPWR.n1157 VPWR.n1156 152
R10277 VPWR.n1147 VPWR.n1146 152
R10278 VPWR.n1470 VPWR.n1469 152
R10279 VPWR.n1047 VPWR.n1046 152
R10280 VPWR.n1746 VPWR.n1745 152
R10281 VPWR.n1034 VPWR.n1033 152
R10282 VPWR.n1030 VPWR.n1029 152
R10283 VPWR.n1051 VPWR.n1050 152
R10284 VPWR.n2845 VPWR.n2844 150.213
R10285 VPWR.n1601 VPWR.t2063 145.137
R10286 VPWR.n1106 VPWR.t2014 145.137
R10287 VPWR.n1617 VPWR.t2000 145.137
R10288 VPWR.n1628 VPWR.t1962 145.137
R10289 VPWR.n1096 VPWR.t2049 145.137
R10290 VPWR.n1644 VPWR.t2042 145.137
R10291 VPWR.n1655 VPWR.t1959 145.137
R10292 VPWR.n1086 VPWR.t1945 145.137
R10293 VPWR.n1671 VPWR.t2050 145.137
R10294 VPWR.n1682 VPWR.t1993 145.137
R10295 VPWR.n1076 VPWR.t1988 145.137
R10296 VPWR.n1698 VPWR.t2040 145.137
R10297 VPWR.n1709 VPWR.t2033 145.137
R10298 VPWR.n1721 VPWR.t2019 145.137
R10299 VPWR.n1116 VPWR.t1969 145.137
R10300 VPWR.n1730 VPWR.t1937 145.137
R10301 VPWR.n119 VPWR.t2048 145.137
R10302 VPWR.n108 VPWR.t1934 145.137
R10303 VPWR.n284 VPWR.t2030 145.137
R10304 VPWR.n274 VPWR.t1983 145.137
R10305 VPWR.n262 VPWR.t1971 145.137
R10306 VPWR.n250 VPWR.t1930 145.137
R10307 VPWR.n238 VPWR.t2016 145.137
R10308 VPWR.n226 VPWR.t2008 145.137
R10309 VPWR.n214 VPWR.t1928 145.137
R10310 VPWR.n202 VPWR.t2057 145.137
R10311 VPWR.n190 VPWR.t2017 145.137
R10312 VPWR.n178 VPWR.t1961 145.137
R10313 VPWR.n166 VPWR.t1952 145.137
R10314 VPWR.n154 VPWR.t2007 145.137
R10315 VPWR.n1768 VPWR.t1976 145.137
R10316 VPWR.n1039 VPWR.t2065 145.137
R10317 VPWR.n1543 VPWR.t1929 145.137
R10318 VPWR.n1548 VPWR.t1986 145.137
R10319 VPWR.n1553 VPWR.t2025 145.137
R10320 VPWR.n1558 VPWR.t2037 145.137
R10321 VPWR.n1563 VPWR.t1979 145.137
R10322 VPWR.n1568 VPWR.t1985 145.137
R10323 VPWR.n1573 VPWR.t2039 145.137
R10324 VPWR.n1578 VPWR.t1936 145.137
R10325 VPWR.n1133 VPWR.t1950 145.137
R10326 VPWR.n1458 VPWR.t1996 145.137
R10327 VPWR.n1453 VPWR.t2045 145.137
R10328 VPWR.n1773 VPWR.t1968 145.137
R10329 VPWR.n1781 VPWR.t1953 145.137
R10330 VPWR.n1777 VPWR.t2013 145.137
R10331 VPWR.n142 VPWR.t1999 145.137
R10332 VPWR.n130 VPWR.t1990 145.137
R10333 VPWR.n1119 VPWR.t2067 145.038
R10334 VPWR.n1110 VPWR.t2018 145.038
R10335 VPWR.n1611 VPWR.t2010 145.038
R10336 VPWR.n1622 VPWR.t1955 145.038
R10337 VPWR.n1100 VPWR.t2059 145.038
R10338 VPWR.n1638 VPWR.t2002 145.038
R10339 VPWR.n1649 VPWR.t1964 145.038
R10340 VPWR.n1090 VPWR.t1949 145.038
R10341 VPWR.n1665 VPWR.t2043 145.038
R10342 VPWR.n1676 VPWR.t2003 145.038
R10343 VPWR.n1080 VPWR.t1947 145.038
R10344 VPWR.n1692 VPWR.t1939 145.038
R10345 VPWR.n1703 VPWR.t2036 145.038
R10346 VPWR.n1069 VPWR.t1989 145.038
R10347 VPWR.n1716 VPWR.t1977 145.038
R10348 VPWR.n1064 VPWR.t2034 145.038
R10349 VPWR.n125 VPWR.t1940 145.038
R10350 VPWR.n114 VPWR.t2001 145.038
R10351 VPWR.n137 VPWR.t1954 145.038
R10352 VPWR.n104 VPWR.t2032 145.038
R10353 VPWR.n100 VPWR.t1987 145.038
R10354 VPWR.n269 VPWR.t1980 145.038
R10355 VPWR.n257 VPWR.t2068 145.038
R10356 VPWR.n245 VPWR.t2027 145.038
R10357 VPWR.n233 VPWR.t1972 145.038
R10358 VPWR.n221 VPWR.t1931 145.038
R10359 VPWR.n209 VPWR.t2060 145.038
R10360 VPWR.n197 VPWR.t2009 145.038
R10361 VPWR.n185 VPWR.t1973 145.038
R10362 VPWR.n173 VPWR.t2058 145.038
R10363 VPWR.n161 VPWR.t2052 145.038
R10364 VPWR.n149 VPWR.t2004 145.038
R10365 VPWR.n53 VPWR.t2053 145.038
R10366 VPWR.n51 VPWR.t1963 145.038
R10367 VPWR.n49 VPWR.t2066 145.038
R10368 VPWR.n47 VPWR.t2026 145.038
R10369 VPWR.n45 VPWR.t1946 145.038
R10370 VPWR.n43 VPWR.t2051 145.038
R10371 VPWR.n41 VPWR.t2069 145.038
R10372 VPWR.n39 VPWR.t2028 145.038
R10373 VPWR.n37 VPWR.t2022 145.038
R10374 VPWR.n35 VPWR.t1943 145.038
R10375 VPWR.n33 VPWR.t1997 145.038
R10376 VPWR.n31 VPWR.t2064 145.038
R10377 VPWR.n29 VPWR.t1995 145.038
R10378 VPWR.n27 VPWR.t1956 145.038
R10379 VPWR.n25 VPWR.t2021 145.038
R10380 VPWR.n23 VPWR.t1970 145.038
R10381 VPWR.n1598 VPWR.t1966 143.911
R10382 VPWR.n1125 VPWR.t2062 143.911
R10383 VPWR.n1614 VPWR.t2047 143.911
R10384 VPWR.n1625 VPWR.t1965 143.911
R10385 VPWR.n1176 VPWR.t1958 143.911
R10386 VPWR.n1641 VPWR.t1944 143.911
R10387 VPWR.n1652 VPWR.t2005 143.911
R10388 VPWR.n1208 VPWR.t1992 143.911
R10389 VPWR.n1668 VPWR.t1941 143.911
R10390 VPWR.n1679 VPWR.t2038 143.911
R10391 VPWR.n1194 VPWR.t2031 143.911
R10392 VPWR.n1695 VPWR.t1978 143.911
R10393 VPWR.n1706 VPWR.t1935 143.911
R10394 VPWR.n1718 VPWR.t2024 143.911
R10395 VPWR.n1733 VPWR.t1984 143.911
R10396 VPWR.n1114 VPWR.t2012 143.911
R10397 VPWR.n116 VPWR.t1951 143.911
R10398 VPWR.n127 VPWR.t1991 143.911
R10399 VPWR.n106 VPWR.t1981 143.911
R10400 VPWR.n287 VPWR.t1933 143.911
R10401 VPWR.n271 VPWR.t2029 143.911
R10402 VPWR.n259 VPWR.t2015 143.911
R10403 VPWR.n247 VPWR.t1932 143.911
R10404 VPWR.n235 VPWR.t1926 143.911
R10405 VPWR.n223 VPWR.t2056 143.911
R10406 VPWR.n211 VPWR.t1974 143.911
R10407 VPWR.n199 VPWR.t1960 143.911
R10408 VPWR.n187 VPWR.t2054 143.911
R10409 VPWR.n175 VPWR.t2006 143.911
R10410 VPWR.n163 VPWR.t1998 143.911
R10411 VPWR.n151 VPWR.t1942 143.911
R10412 VPWR.n1228 VPWR.t1948 143.911
R10413 VPWR.n1150 VPWR.t1975 143.911
R10414 VPWR.n1224 VPWR.t2041 143.911
R10415 VPWR.n1482 VPWR.t1982 143.911
R10416 VPWR.n1170 VPWR.t2035 143.911
R10417 VPWR.n1166 VPWR.t2023 143.911
R10418 VPWR.n1160 VPWR.t1938 143.911
R10419 VPWR.n1476 VPWR.t1994 143.911
R10420 VPWR.n1156 VPWR.t1927 143.911
R10421 VPWR.n1146 VPWR.t2020 143.911
R10422 VPWR.n1469 VPWR.t2044 143.911
R10423 VPWR.n1046 VPWR.t1967 143.911
R10424 VPWR.n1745 VPWR.t2011 143.911
R10425 VPWR.n1033 VPWR.t1957 143.911
R10426 VPWR.n1029 VPWR.t2061 143.911
R10427 VPWR.n1050 VPWR.t2055 143.911
R10428 VPWR.n139 VPWR.t2046 143.911
R10429 VPWR.t1503 VPWR.t933 140.989
R10430 VPWR.t1299 VPWR.t1286 140.989
R10431 VPWR.t1326 VPWR.t1299 140.989
R10432 VPWR.t1302 VPWR.t1326 140.989
R10433 VPWR.t410 VPWR.t1302 140.989
R10434 VPWR.t404 VPWR.t410 140.989
R10435 VPWR.t396 VPWR.t404 140.989
R10436 VPWR.t398 VPWR.t396 140.989
R10437 VPWR.t1730 VPWR.t394 140.989
R10438 VPWR.t1338 VPWR.t1305 140.989
R10439 VPWR.t1292 VPWR.t1338 140.989
R10440 VPWR.t1339 VPWR.t1292 140.989
R10441 VPWR.t877 VPWR.t1339 140.989
R10442 VPWR.t889 VPWR.t877 140.989
R10443 VPWR.t881 VPWR.t889 140.989
R10444 VPWR.t885 VPWR.t881 140.989
R10445 VPWR.t1283 VPWR.t1324 140.989
R10446 VPWR.t1313 VPWR.t1283 140.989
R10447 VPWR.t1287 VPWR.t1313 140.989
R10448 VPWR.t1144 VPWR.t1287 140.989
R10449 VPWR.t1142 VPWR.t1144 140.989
R10450 VPWR.t1148 VPWR.t1142 140.989
R10451 VPWR.t1136 VPWR.t1148 140.989
R10452 VPWR.t1882 VPWR.t1314 140.989
R10453 VPWR.t1284 VPWR.t1327 140.989
R10454 VPWR.t1334 VPWR.t1284 140.989
R10455 VPWR.t1311 VPWR.t1334 140.989
R10456 VPWR.t406 VPWR.t1311 140.989
R10457 VPWR.t400 VPWR.t406 140.989
R10458 VPWR.t408 VPWR.t400 140.989
R10459 VPWR.t402 VPWR.t408 140.989
R10460 VPWR.t1306 VPWR.t1293 140.989
R10461 VPWR.t1280 VPWR.t1306 140.989
R10462 VPWR.t1332 VPWR.t1280 140.989
R10463 VPWR.t887 VPWR.t1332 140.989
R10464 VPWR.t879 VPWR.t887 140.989
R10465 VPWR.t891 VPWR.t879 140.989
R10466 VPWR.t883 VPWR.t891 140.989
R10467 VPWR.t1303 VPWR.t1295 140.989
R10468 VPWR.t1309 VPWR.t1303 140.989
R10469 VPWR.t1297 VPWR.t1309 140.989
R10470 VPWR.t1146 VPWR.t1297 140.989
R10471 VPWR.t1150 VPWR.t1146 140.989
R10472 VPWR.t1138 VPWR.t1150 140.989
R10473 VPWR.t1140 VPWR.t1138 140.989
R10474 VPWR VPWR.n1442 133.312
R10475 VPWR.n2841 VPWR.n2840 129.13
R10476 VPWR.n2858 VPWR.n2819 129.13
R10477 VPWR.n2780 VPWR 127.562
R10478 VPWR.n2760 VPWR 127.562
R10479 VPWR.n2741 VPWR 127.562
R10480 VPWR VPWR.t1345 125.883
R10481 VPWR.n2705 VPWR 125.883
R10482 VPWR.t1732 VPWR.t392 120.849
R10483 VPWR.t986 VPWR.t1744 117.492
R10484 VPWR.t1267 VPWR.t941 117.492
R10485 VPWR.t849 VPWR 115.814
R10486 VPWR VPWR.t398 114.135
R10487 VPWR VPWR.t885 114.135
R10488 VPWR VPWR.t1136 114.135
R10489 VPWR.n2859 VPWR.n2817 111.059
R10490 VPWR.t1266 VPWR 107.421
R10491 VPWR.n1330 VPWR.n1329 106.561
R10492 VPWR.n2781 VPWR.n2780 106.561
R10493 VPWR.n2761 VPWR.n2760 106.561
R10494 VPWR.n2742 VPWR.n2741 106.561
R10495 VPWR.n2706 VPWR.n2705 106.561
R10496 VPWR.n2668 VPWR.n2667 106.561
R10497 VPWR.n2631 VPWR.n2630 106.561
R10498 VPWR VPWR.t1736 106.543
R10499 VPWR VPWR.n1234 104.8
R10500 VPWR VPWR.n1257 104.8
R10501 VPWR VPWR.n1281 104.8
R10502 VPWR VPWR.n1366 104.8
R10503 VPWR VPWR.n1405 104.8
R10504 VPWR.n1443 VPWR 100.883
R10505 VPWR VPWR.t992 100.624
R10506 VPWR.t1130 VPWR.t977 97.9386
R10507 VPWR.n2859 VPWR.n2858 93.3652
R10508 VPWR.n1231 VPWR.n1230 91.8492
R10509 VPWR.n1153 VPWR.n1152 91.8492
R10510 VPWR.n1227 VPWR.n1226 91.8492
R10511 VPWR.n1485 VPWR.n1484 91.8492
R10512 VPWR.n1173 VPWR.n1172 91.8492
R10513 VPWR.n1169 VPWR.n1168 91.8492
R10514 VPWR.n1163 VPWR.n1162 91.8492
R10515 VPWR.n1479 VPWR.n1478 91.8492
R10516 VPWR.n1159 VPWR.n1158 91.8492
R10517 VPWR.n1149 VPWR.n1148 91.8492
R10518 VPWR.n1472 VPWR.n1471 91.8492
R10519 VPWR.n1049 VPWR.n1048 91.8492
R10520 VPWR.n1748 VPWR.n1747 91.8492
R10521 VPWR.n1036 VPWR.n1035 91.8492
R10522 VPWR.n1032 VPWR.n1031 91.8492
R10523 VPWR.n1053 VPWR.n1052 91.8492
R10524 VPWR.n2847 VPWR.n2820 91.4829
R10525 VPWR.t1130 VPWR.n2842 90.0872
R10526 VPWR.t1330 VPWR 88.7855
R10527 VPWR.n1235 VPWR 79.407
R10528 VPWR.n1258 VPWR 79.407
R10529 VPWR.n1282 VPWR 79.407
R10530 VPWR.n1367 VPWR 79.407
R10531 VPWR.n1406 VPWR 79.407
R10532 VPWR.t1269 VPWR.t995 78.8874
R10533 VPWR.n2840 VPWR.n2818 74.9181
R10534 VPWR.n2858 VPWR.n2818 74.9181
R10535 VPWR.n2858 VPWR.n2857 74.9181
R10536 VPWR.n2857 VPWR.n2820 74.9181
R10537 VPWR.t587 VPWR.t872 70.4952
R10538 VPWR.t872 VPWR.t438 70.4952
R10539 VPWR.t438 VPWR.t1499 70.4952
R10540 VPWR.t1499 VPWR.t1742 70.4952
R10541 VPWR.t1742 VPWR.t990 70.4952
R10542 VPWR.t990 VPWR.t414 70.4952
R10543 VPWR.t414 VPWR.t1503 70.4952
R10544 VPWR.t1318 VPWR.t1882 70.4952
R10545 VPWR.t1888 VPWR.t1318 70.4952
R10546 VPWR.t1290 VPWR.t1888 70.4952
R10547 VPWR.t493 VPWR.t1290 70.4952
R10548 VPWR.t1322 VPWR.t493 70.4952
R10549 VPWR.t1886 VPWR.t1322 70.4952
R10550 VPWR.t1345 VPWR.t1886 70.4952
R10551 VPWR VPWR.t587 68.8168
R10552 VPWR.t1738 VPWR.t1734 68.8168
R10553 VPWR.t995 VPWR.t849 62.103
R10554 VPWR VPWR.t1730 60.4245
R10555 VPWR.n2849 VPWR.n2842 59.762
R10556 VPWR.n2845 VPWR.n2819 53.8358
R10557 VPWR.t1734 VPWR.t1134 52.0323
R10558 VPWR.t950 VPWR 50.3539
R10559 VPWR VPWR.t1738 50.3539
R10560 VPWR VPWR.t1732 50.3539
R10561 VPWR.t1327 VPWR 50.3539
R10562 VPWR.t1293 VPWR 50.3539
R10563 VPWR.t1295 VPWR 50.3539
R10564 VPWR.n2854 VPWR.n2818 46.2505
R10565 VPWR.n2855 VPWR.n2854 46.2505
R10566 VPWR.n2835 VPWR.n2834 46.2505
R10567 VPWR.n2836 VPWR.n2835 46.2505
R10568 VPWR.n2838 VPWR.n2837 46.2505
R10569 VPWR.n2837 VPWR.n2836 46.2505
R10570 VPWR.n2844 VPWR.n2824 46.2505
R10571 VPWR.n2857 VPWR.n2856 46.2505
R10572 VPWR.n2856 VPWR.n2855 46.2505
R10573 VPWR.n2849 VPWR.n2848 46.2505
R10574 VPWR.n2846 VPWR.n2845 45.9299
R10575 VPWR.n2832 VPWR.n2830 44.8005
R10576 VPWR.n2830 VPWR.n2826 44.8005
R10577 VPWR.n2847 VPWR.n2843 37.0005
R10578 VPWR.n2843 VPWR.t977 37.0005
R10579 VPWR.n1230 VPWR.n1229 34.7473
R10580 VPWR.n1152 VPWR.n1151 34.7473
R10581 VPWR.n1226 VPWR.n1225 34.7473
R10582 VPWR.n1484 VPWR.n1483 34.7473
R10583 VPWR.n1172 VPWR.n1171 34.7473
R10584 VPWR.n1168 VPWR.n1167 34.7473
R10585 VPWR.n1162 VPWR.n1161 34.7473
R10586 VPWR.n1478 VPWR.n1477 34.7473
R10587 VPWR.n1158 VPWR.n1157 34.7473
R10588 VPWR.n1148 VPWR.n1147 34.7473
R10589 VPWR.n1471 VPWR.n1470 34.7473
R10590 VPWR.n1048 VPWR.n1047 34.7473
R10591 VPWR.n1747 VPWR.n1746 34.7473
R10592 VPWR.n1035 VPWR.n1034 34.7473
R10593 VPWR.n1031 VPWR.n1030 34.7473
R10594 VPWR.n1052 VPWR.n1051 34.7473
R10595 VPWR.n1299 VPWR.n1298 34.6358
R10596 VPWR.n1357 VPWR.n1341 34.6358
R10597 VPWR.n1362 VPWR.n1361 34.6358
R10598 VPWR.n1396 VPWR.n1380 34.6358
R10599 VPWR.n1401 VPWR.n1400 34.6358
R10600 VPWR.n1411 VPWR.n1377 34.6358
R10601 VPWR.n1433 VPWR.n1417 34.6358
R10602 VPWR.n1438 VPWR.n1437 34.6358
R10603 VPWR.n2755 VPWR.n2754 34.6358
R10604 VPWR.n2721 VPWR.n2713 34.6358
R10605 VPWR.n2728 VPWR.n2727 34.6358
R10606 VPWR.n2685 VPWR.n2676 34.6358
R10607 VPWR.n2688 VPWR.n2687 34.6358
R10608 VPWR.n2692 VPWR.n2691 34.6358
R10609 VPWR.n2648 VPWR.n2639 34.6358
R10610 VPWR.n2651 VPWR.n2650 34.6358
R10611 VPWR.n2655 VPWR.n2654 34.6358
R10612 VPWR.n2662 VPWR.n2661 34.6358
R10613 VPWR.n2615 VPWR.n2611 34.6358
R10614 VPWR.n2619 VPWR.n2603 34.6358
R10615 VPWR.n2622 VPWR.n2621 34.6358
R10616 VPWR.n1316 VPWR.n1315 32.0005
R10617 VPWR.n1353 VPWR.n1352 32.0005
R10618 VPWR.n1392 VPWR.n1391 32.0005
R10619 VPWR.n1429 VPWR.n1428 32.0005
R10620 VPWR.n2717 VPWR.n2716 30.8711
R10621 VPWR.n2681 VPWR.n2680 30.8711
R10622 VPWR.n2644 VPWR.n2643 30.8711
R10623 VPWR.n2610 VPWR.n2609 30.8711
R10624 VPWR.n2834 VPWR.n2832 30.1181
R10625 VPWR.n2838 VPWR.n2826 30.1181
R10626 VPWR.n2848 VPWR.n2846 28.9887
R10627 VPWR.n1325 VPWR.n1324 28.2358
R10628 VPWR.n5 VPWR.t1502 26.5955
R10629 VPWR.n5 VPWR.t989 26.5955
R10630 VPWR.n4 VPWR.t993 26.5955
R10631 VPWR.n4 VPWR.t1498 26.5955
R10632 VPWR.n1240 VPWR.t1865 26.5955
R10633 VPWR.n1240 VPWR.t1864 26.5955
R10634 VPWR.n1239 VPWR.t875 26.5955
R10635 VPWR.n1239 VPWR.t1710 26.5955
R10636 VPWR.n1245 VPWR.t1861 26.5955
R10637 VPWR.n1245 VPWR.t1866 26.5955
R10638 VPWR.n1238 VPWR.t1090 26.5955
R10639 VPWR.n1238 VPWR.t874 26.5955
R10640 VPWR.n1263 VPWR.t1668 26.5955
R10641 VPWR.n1263 VPWR.t1669 26.5955
R10642 VPWR.n1262 VPWR.t779 26.5955
R10643 VPWR.n1262 VPWR.t776 26.5955
R10644 VPWR.n1268 VPWR.t1177 26.5955
R10645 VPWR.n1268 VPWR.t1679 26.5955
R10646 VPWR.n1261 VPWR.t782 26.5955
R10647 VPWR.n1261 VPWR.t780 26.5955
R10648 VPWR.n1287 VPWR.t654 26.5955
R10649 VPWR.n1287 VPWR.t661 26.5955
R10650 VPWR.n1286 VPWR.t770 26.5955
R10651 VPWR.n1286 VPWR.t769 26.5955
R10652 VPWR.n1292 VPWR.t658 26.5955
R10653 VPWR.n1292 VPWR.t655 26.5955
R10654 VPWR.n1285 VPWR.t773 26.5955
R10655 VPWR.n1285 VPWR.t771 26.5955
R10656 VPWR.n1314 VPWR.t1539 26.5955
R10657 VPWR.n1314 VPWR.t1541 26.5955
R10658 VPWR.n1307 VPWR.t1504 26.5955
R10659 VPWR.n1307 VPWR.t934 26.5955
R10660 VPWR.n1321 VPWR.t1500 26.5955
R10661 VPWR.n1321 VPWR.t991 26.5955
R10662 VPWR.n1323 VPWR.t439 26.5955
R10663 VPWR.n1323 VPWR.t1743 26.5955
R10664 VPWR.n1351 VPWR.t1872 26.5955
R10665 VPWR.n1351 VPWR.t1875 26.5955
R10666 VPWR.n1350 VPWR.t1259 26.5955
R10667 VPWR.n1350 VPWR.t580 26.5955
R10668 VPWR.n1344 VPWR.t1868 26.5955
R10669 VPWR.n1344 VPWR.t447 26.5955
R10670 VPWR.n1343 VPWR.t1091 26.5955
R10671 VPWR.n1343 VPWR.t1257 26.5955
R10672 VPWR.n1359 VPWR.t1863 26.5955
R10673 VPWR.n1359 VPWR.t1862 26.5955
R10674 VPWR.n1358 VPWR.t1711 26.5955
R10675 VPWR.n1358 VPWR.t1092 26.5955
R10676 VPWR.n1390 VPWR.t1256 26.5955
R10677 VPWR.n1390 VPWR.t1787 26.5955
R10678 VPWR.n1389 VPWR.t1874 26.5955
R10679 VPWR.n1389 VPWR.t1741 26.5955
R10680 VPWR.n1383 VPWR.t1850 26.5955
R10681 VPWR.n1383 VPWR.t1543 26.5955
R10682 VPWR.n1382 VPWR.t783 26.5955
R10683 VPWR.n1382 VPWR.t1870 26.5955
R10684 VPWR.n1398 VPWR.t1670 26.5955
R10685 VPWR.n1398 VPWR.t1176 26.5955
R10686 VPWR.n1397 VPWR.t784 26.5955
R10687 VPWR.n1397 VPWR.t781 26.5955
R10688 VPWR.n1427 VPWR.t586 26.5955
R10689 VPWR.n1427 VPWR.t441 26.5955
R10690 VPWR.n1426 VPWR.t1786 26.5955
R10691 VPWR.n1426 VPWR.t582 26.5955
R10692 VPWR.n1420 VPWR.t657 26.5955
R10693 VPWR.n1420 VPWR.t583 26.5955
R10694 VPWR.n1419 VPWR.t767 26.5955
R10695 VPWR.n1419 VPWR.t1258 26.5955
R10696 VPWR.n1435 VPWR.t660 26.5955
R10697 VPWR.n1435 VPWR.t659 26.5955
R10698 VPWR.n1434 VPWR.t768 26.5955
R10699 VPWR.n1434 VPWR.t766 26.5955
R10700 VPWR.n2802 VPWR.t492 26.5955
R10701 VPWR.n2802 VPWR.t418 26.5955
R10702 VPWR.n2804 VPWR.t1885 26.5955
R10703 VPWR.n2804 VPWR.t677 26.5955
R10704 VPWR.n2782 VPWR.t411 26.5955
R10705 VPWR.n2782 VPWR.t405 26.5955
R10706 VPWR.n2783 VPWR.t851 26.5955
R10707 VPWR.n2783 VPWR.t1621 26.5955
R10708 VPWR.n2786 VPWR.t397 26.5955
R10709 VPWR.n2786 VPWR.t399 26.5955
R10710 VPWR.n2787 VPWR.t994 26.5955
R10711 VPWR.n2787 VPWR.t601 26.5955
R10712 VPWR.n2762 VPWR.t1199 26.5955
R10713 VPWR.n2762 VPWR.t1463 26.5955
R10714 VPWR.n2763 VPWR.t878 26.5955
R10715 VPWR.n2763 VPWR.t890 26.5955
R10716 VPWR.n2766 VPWR.t1210 26.5955
R10717 VPWR.n2766 VPWR.t1209 26.5955
R10718 VPWR.n2767 VPWR.t882 26.5955
R10719 VPWR.n2767 VPWR.t886 26.5955
R10720 VPWR.n2743 VPWR.t1252 26.5955
R10721 VPWR.n2743 VPWR.t1249 26.5955
R10722 VPWR.n2744 VPWR.t1145 26.5955
R10723 VPWR.n2744 VPWR.t1143 26.5955
R10724 VPWR.n2747 VPWR.t1253 26.5955
R10725 VPWR.n2747 VPWR.t1254 26.5955
R10726 VPWR.n2748 VPWR.t1149 26.5955
R10727 VPWR.n2748 VPWR.t1137 26.5955
R10728 VPWR.n2708 VPWR.t1291 26.5955
R10729 VPWR.n2708 VPWR.t1323 26.5955
R10730 VPWR.n2712 VPWR.t1315 26.5955
R10731 VPWR.n2712 VPWR.t1883 26.5955
R10732 VPWR.n2715 VPWR.t1289 26.5955
R10733 VPWR.n2715 VPWR.t1337 26.5955
R10734 VPWR.n2709 VPWR.t1889 26.5955
R10735 VPWR.n2709 VPWR.t494 26.5955
R10736 VPWR.n2679 VPWR.t1285 26.5955
R10737 VPWR.n2679 VPWR.t1335 26.5955
R10738 VPWR.n2678 VPWR.t1301 26.5955
R10739 VPWR.n2678 VPWR.t1347 26.5955
R10740 VPWR.n2675 VPWR.t1312 26.5955
R10741 VPWR.n2675 VPWR.t823 26.5955
R10742 VPWR.n2674 VPWR.t1329 26.5955
R10743 VPWR.n2674 VPWR.t407 26.5955
R10744 VPWR.n2671 VPWR.t490 26.5955
R10745 VPWR.n2671 VPWR.t597 26.5955
R10746 VPWR.n2670 VPWR.t401 26.5955
R10747 VPWR.n2670 VPWR.t409 26.5955
R10748 VPWR.n2642 VPWR.t1307 26.5955
R10749 VPWR.n2642 VPWR.t1281 26.5955
R10750 VPWR.n2641 VPWR.t1325 26.5955
R10751 VPWR.n2641 VPWR.t1300 26.5955
R10752 VPWR.n2638 VPWR.t1333 26.5955
R10753 VPWR.n2638 VPWR.t888 26.5955
R10754 VPWR.n2637 VPWR.t1343 26.5955
R10755 VPWR.n2637 VPWR.t1201 26.5955
R10756 VPWR.n2634 VPWR.t880 26.5955
R10757 VPWR.n2634 VPWR.t892 26.5955
R10758 VPWR.n2633 VPWR.t1465 26.5955
R10759 VPWR.n2633 VPWR.t1200 26.5955
R10760 VPWR.n2606 VPWR.t1304 26.5955
R10761 VPWR.n2606 VPWR.t1310 26.5955
R10762 VPWR.n2605 VPWR.t1340 26.5955
R10763 VPWR.n2605 VPWR.t1321 26.5955
R10764 VPWR.n2613 VPWR.t1316 26.5955
R10765 VPWR.n2613 VPWR.t1147 26.5955
R10766 VPWR.n2612 VPWR.t1298 26.5955
R10767 VPWR.n2612 VPWR.t1250 26.5955
R10768 VPWR.n2602 VPWR.t1151 26.5955
R10769 VPWR.n2602 VPWR.t1139 26.5955
R10770 VPWR.n2601 VPWR.t1247 26.5955
R10771 VPWR.n2601 VPWR.t1251 26.5955
R10772 VPWR.n17 VPWR.n16 25.977
R10773 VPWR.n1253 VPWR.n1252 25.977
R10774 VPWR.n1313 VPWR.n1310 25.977
R10775 VPWR.n1349 VPWR.n1346 25.977
R10776 VPWR.n1372 VPWR.n1338 25.977
R10777 VPWR.n1388 VPWR.n1385 25.977
R10778 VPWR.n1425 VPWR.n1422 25.977
R10779 VPWR.n2811 VPWR.n2810 25.977
R10780 VPWR.n2795 VPWR.n2794 25.977
R10781 VPWR.n2717 VPWR.n2714 25.977
R10782 VPWR.n2681 VPWR.n2677 25.977
R10783 VPWR.n2699 VPWR.n2698 25.977
R10784 VPWR.n2644 VPWR.n2640 25.977
R10785 VPWR.n2609 VPWR.n2607 25.977
R10786 VPWR.n1335 VPWR.n1334 25.224
R10787 VPWR.n2737 VPWR.n2736 25.224
R10788 VPWR.n2722 VPWR.n2721 24.8476
R10789 VPWR.n2686 VPWR.n2685 24.8476
R10790 VPWR.n2649 VPWR.n2648 24.8476
R10791 VPWR.n2615 VPWR.n2614 24.8476
R10792 VPWR.n16 VPWR.n15 24.4711
R10793 VPWR.n1252 VPWR.n1251 24.4711
R10794 VPWR.n1315 VPWR.n1313 24.4711
R10795 VPWR.n1352 VPWR.n1349 24.4711
R10796 VPWR.n1391 VPWR.n1388 24.4711
R10797 VPWR.n1428 VPWR.n1425 24.4711
R10798 VPWR.n2810 VPWR.n2809 24.4711
R10799 VPWR.n2794 VPWR.n2793 24.4711
R10800 VPWR.n11 VPWR.n2 23.7181
R10801 VPWR.n1247 VPWR.n1236 23.7181
R10802 VPWR.n1270 VPWR.n1259 23.7181
R10803 VPWR.n1274 VPWR.n1259 23.7181
R10804 VPWR.n1294 VPWR.n1283 23.7181
R10805 VPWR.n1298 VPWR.n1283 23.7181
R10806 VPWR.n1330 VPWR.n1328 23.7181
R10807 VPWR.n1368 VPWR.n1365 23.7181
R10808 VPWR.n1407 VPWR.n1404 23.7181
R10809 VPWR.n1407 VPWR.n1377 23.7181
R10810 VPWR.n1444 VPWR.n1441 23.7181
R10811 VPWR.n2808 VPWR.n2807 23.7181
R10812 VPWR.n2789 VPWR.n2781 23.7181
R10813 VPWR.n2769 VPWR.n2761 23.7181
R10814 VPWR.n2773 VPWR.n2761 23.7181
R10815 VPWR.n2750 VPWR.n2742 23.7181
R10816 VPWR.n2754 VPWR.n2742 23.7181
R10817 VPWR.n2731 VPWR.n2706 23.7181
R10818 VPWR.n2694 VPWR.n2668 23.7181
R10819 VPWR.n2657 VPWR.n2631 23.7181
R10820 VPWR.n2661 VPWR.n2631 23.7181
R10821 VPWR.n2626 VPWR.n2625 23.7181
R10822 VPWR.t1746 VPWR.t986 23.4987
R10823 VPWR.t943 VPWR.t1267 23.4987
R10824 VPWR.n2852 VPWR.n2841 23.1255
R10825 VPWR.n2852 VPWR.t1130 23.1255
R10826 VPWR.n2851 VPWR.n2819 23.1255
R10827 VPWR.t1130 VPWR.n2851 23.1255
R10828 VPWR.n11 VPWR.n10 22.9652
R10829 VPWR.n1247 VPWR.n1246 22.9652
R10830 VPWR.n1270 VPWR.n1269 22.9652
R10831 VPWR.n1294 VPWR.n1293 22.9652
R10832 VPWR.n2807 VPWR.n2803 22.9652
R10833 VPWR.n2789 VPWR.n2788 22.9652
R10834 VPWR.n2769 VPWR.n2768 22.9652
R10835 VPWR.n2750 VPWR.n2749 22.9652
R10836 VPWR.n1320 VPWR.n1308 22.2123
R10837 VPWR.n2724 VPWR.n2723 22.2123
R10838 VPWR.n10 VPWR.n3 21.4593
R10839 VPWR.n1246 VPWR.n1237 21.4593
R10840 VPWR.n1269 VPWR.n1260 21.4593
R10841 VPWR.n1293 VPWR.n1284 21.4593
R10842 VPWR.n1442 VPWR.t581 20.5957
R10843 VPWR.n1443 VPWR.t440 20.5957
R10844 VPWR.n1277 VPWR.n1276 19.9534
R10845 VPWR.n1300 VPWR.n1299 19.9534
R10846 VPWR.n1334 VPWR.n1303 19.9534
R10847 VPWR.n2776 VPWR.n2775 19.9534
R10848 VPWR.n2756 VPWR.n2755 19.9534
R10849 VPWR.n2736 VPWR.n2735 19.9534
R10850 VPWR.n2724 VPWR.n2710 18.824
R10851 VPWR.n2688 VPWR.n2672 18.824
R10852 VPWR.n2651 VPWR.n2635 18.824
R10853 VPWR.n2620 VPWR.n2619 18.824
R10854 VPWR.n1316 VPWR.n1308 18.4476
R10855 VPWR.n1353 VPWR.n1345 18.4476
R10856 VPWR.n1373 VPWR.n1372 18.4476
R10857 VPWR.n1392 VPWR.n1384 18.4476
R10858 VPWR.n1429 VPWR.n1421 18.4476
R10859 VPWR.n2700 VPWR.n2699 18.4476
R10860 VPWR.n1413 VPWR.n1412 17.5829
R10861 VPWR.n2664 VPWR.n2663 17.5829
R10862 VPWR.n6 VPWR.n3 16.9417
R10863 VPWR.n1241 VPWR.n1237 16.9417
R10864 VPWR.n1264 VPWR.n1260 16.9417
R10865 VPWR.n1288 VPWR.n1284 16.9417
R10866 VPWR.n2730 VPWR.n2729 16.5652
R10867 VPWR.n1306 VPWR.n1304 16.1887
R10868 VPWR.n1374 VPWR.n1373 16.1887
R10869 VPWR.n2701 VPWR.n2700 16.1887
R10870 VPWR.n1235 VPWR.t443 16.0935
R10871 VPWR.n1258 VPWR.t507 16.0935
R10872 VPWR.n1282 VPWR.t413 16.0935
R10873 VPWR.n1367 VPWR.t446 16.0935
R10874 VPWR.n1406 VPWR.t444 16.0935
R10875 VPWR.n1234 VPWR.t437 16.0935
R10876 VPWR.n1257 VPWR.t442 16.0935
R10877 VPWR.n1281 VPWR.t505 16.0935
R10878 VPWR.n1366 VPWR.t579 16.0935
R10879 VPWR.n1405 VPWR.t777 16.0935
R10880 VPWR.n1325 VPWR.n1306 15.8123
R10881 VPWR.n2727 VPWR.n2710 15.8123
R10882 VPWR.n2729 VPWR.n2728 15.8123
R10883 VPWR.n2691 VPWR.n2672 15.8123
R10884 VPWR.n2654 VPWR.n2635 15.8123
R10885 VPWR.n2621 VPWR.n2620 15.8123
R10886 VPWR.n1330 VPWR.n1303 13.5534
R10887 VPWR.n2735 VPWR.n2706 13.5534
R10888 VPWR.n2839 VPWR.n2823 13.2148
R10889 VPWR.n2823 VPWR.t1264 13.2148
R10890 VPWR.n2827 VPWR.n2817 13.2148
R10891 VPWR.n2827 VPWR.t1264 13.2148
R10892 VPWR.n2833 VPWR.n2829 13.2148
R10893 VPWR.n2829 VPWR.t1264 13.2148
R10894 VPWR.n15 VPWR.n2 12.8005
R10895 VPWR.n1251 VPWR.n1236 12.8005
R10896 VPWR.n1368 VPWR.n1338 12.8005
R10897 VPWR.n2809 VPWR.n2808 12.8005
R10898 VPWR.n2793 VPWR.n2781 12.8005
R10899 VPWR.n2698 VPWR.n2668 12.8005
R10900 VPWR.n1322 VPWR.n1320 12.424
R10901 VPWR.n1360 VPWR.n1357 12.424
R10902 VPWR.n1399 VPWR.n1396 12.424
R10903 VPWR.n1436 VPWR.n1433 12.424
R10904 VPWR.n1276 VPWR.n1275 10.5417
R10905 VPWR.n1412 VPWR.n1411 10.5417
R10906 VPWR.n2775 VPWR.n2774 10.5417
R10907 VPWR.n2663 VPWR.n2662 10.5417
R10908 VPWR.n2687 VPWR.n2686 9.78874
R10909 VPWR.n2650 VPWR.n2649 9.78874
R10910 VPWR.n2614 VPWR.n2603 9.78874
R10911 VPWR.n1361 VPWR.n1360 9.41227
R10912 VPWR.n1365 VPWR.n1339 9.41227
R10913 VPWR.n1400 VPWR.n1399 9.41227
R10914 VPWR.n1404 VPWR.n1378 9.41227
R10915 VPWR.n1437 VPWR.n1436 9.41227
R10916 VPWR.n1441 VPWR.n1415 9.41227
R10917 VPWR.n2694 VPWR.n2693 9.41227
R10918 VPWR.n2657 VPWR.n2656 9.41227
R10919 VPWR.n2625 VPWR.n2599 9.41227
R10920 VPWR.n1229 VPWR 9.37021
R10921 VPWR.n1151 VPWR 9.37021
R10922 VPWR.n1225 VPWR 9.37021
R10923 VPWR.n1483 VPWR 9.37021
R10924 VPWR.n1171 VPWR 9.37021
R10925 VPWR.n1167 VPWR 9.37021
R10926 VPWR.n1161 VPWR 9.37021
R10927 VPWR.n1477 VPWR 9.37021
R10928 VPWR.n1157 VPWR 9.37021
R10929 VPWR.n1147 VPWR 9.37021
R10930 VPWR.n1470 VPWR 9.37021
R10931 VPWR.n1047 VPWR 9.37021
R10932 VPWR.n1746 VPWR 9.37021
R10933 VPWR.n1034 VPWR 9.37021
R10934 VPWR.n1030 VPWR 9.37021
R10935 VPWR.n1051 VPWR 9.37021
R10936 VPWR.n1467 VPWR.n1466 9.33404
R10937 VPWR.n352 VPWR.n351 9.33404
R10938 VPWR.n1534 VPWR.n1533 9.33404
R10939 VPWR.n348 VPWR.n347 9.33404
R10940 VPWR.n965 VPWR.n964 9.33404
R10941 VPWR.n2479 VPWR.n2478 9.33404
R10942 VPWR.n2475 VPWR.n2474 9.33404
R10943 VPWR.n320 VPWR.n319 9.33404
R10944 VPWR.n973 VPWR.n972 9.33404
R10945 VPWR.n2445 VPWR.n2444 9.33404
R10946 VPWR.n324 VPWR.n323 9.33404
R10947 VPWR.n1891 VPWR.n1890 9.33404
R10948 VPWR.n1887 VPWR.n1886 9.33404
R10949 VPWR.n1881 VPWR.n1880 9.33404
R10950 VPWR.n389 VPWR.n388 9.33404
R10951 VPWR.n393 VPWR.n392 9.33404
R10952 VPWR.n397 VPWR.n396 9.33404
R10953 VPWR.n2455 VPWR.n2454 9.33404
R10954 VPWR.n332 VPWR.n331 9.33404
R10955 VPWR.n1877 VPWR.n1876 9.33404
R10956 VPWR.n405 VPWR.n404 9.33404
R10957 VPWR.n2459 VPWR.n2458 9.33404
R10958 VPWR.n336 VPWR.n335 9.33404
R10959 VPWR.n2308 VPWR.n2307 9.33404
R10960 VPWR.n2312 VPWR.n2311 9.33404
R10961 VPWR.n2318 VPWR.n2317 9.33404
R10962 VPWR.n2322 VPWR.n2321 9.33404
R10963 VPWR.n2332 VPWR.n2331 9.33404
R10964 VPWR.n2338 VPWR.n2337 9.33404
R10965 VPWR.n2342 VPWR.n2341 9.33404
R10966 VPWR.n2348 VPWR.n2347 9.33404
R10967 VPWR.n2352 VPWR.n2351 9.33404
R10968 VPWR.n2358 VPWR.n2357 9.33404
R10969 VPWR.n2362 VPWR.n2361 9.33404
R10970 VPWR.n2368 VPWR.n2367 9.33404
R10971 VPWR.n2372 VPWR.n2371 9.33404
R10972 VPWR.n2378 VPWR.n2377 9.33404
R10973 VPWR.n2381 VPWR.n2380 9.33404
R10974 VPWR.n2328 VPWR.n2327 9.33404
R10975 VPWR.n544 VPWR.n543 9.33404
R10976 VPWR.n540 VPWR.n539 9.33404
R10977 VPWR.n536 VPWR.n535 9.33404
R10978 VPWR.n532 VPWR.n531 9.33404
R10979 VPWR.n524 VPWR.n523 9.33404
R10980 VPWR.n520 VPWR.n519 9.33404
R10981 VPWR.n516 VPWR.n515 9.33404
R10982 VPWR.n512 VPWR.n511 9.33404
R10983 VPWR.n508 VPWR.n507 9.33404
R10984 VPWR.n504 VPWR.n503 9.33404
R10985 VPWR.n500 VPWR.n499 9.33404
R10986 VPWR.n496 VPWR.n495 9.33404
R10987 VPWR.n492 VPWR.n491 9.33404
R10988 VPWR.n488 VPWR.n487 9.33404
R10989 VPWR.n485 VPWR.n484 9.33404
R10990 VPWR.n528 VPWR.n527 9.33404
R10991 VPWR.n2283 VPWR.n2282 9.33404
R10992 VPWR.n2279 VPWR.n2278 9.33404
R10993 VPWR.n2273 VPWR.n2272 9.33404
R10994 VPWR.n2269 VPWR.n2268 9.33404
R10995 VPWR.n2259 VPWR.n2258 9.33404
R10996 VPWR.n2253 VPWR.n2252 9.33404
R10997 VPWR.n2249 VPWR.n2248 9.33404
R10998 VPWR.n2243 VPWR.n2242 9.33404
R10999 VPWR.n2239 VPWR.n2238 9.33404
R11000 VPWR.n2233 VPWR.n2232 9.33404
R11001 VPWR.n2229 VPWR.n2228 9.33404
R11002 VPWR.n2223 VPWR.n2222 9.33404
R11003 VPWR.n2219 VPWR.n2218 9.33404
R11004 VPWR.n2213 VPWR.n2212 9.33404
R11005 VPWR.n2210 VPWR.n2209 9.33404
R11006 VPWR.n2263 VPWR.n2262 9.33404
R11007 VPWR.n581 VPWR.n580 9.33404
R11008 VPWR.n585 VPWR.n584 9.33404
R11009 VPWR.n589 VPWR.n588 9.33404
R11010 VPWR.n593 VPWR.n592 9.33404
R11011 VPWR.n601 VPWR.n600 9.33404
R11012 VPWR.n605 VPWR.n604 9.33404
R11013 VPWR.n609 VPWR.n608 9.33404
R11014 VPWR.n613 VPWR.n612 9.33404
R11015 VPWR.n617 VPWR.n616 9.33404
R11016 VPWR.n621 VPWR.n620 9.33404
R11017 VPWR.n625 VPWR.n624 9.33404
R11018 VPWR.n629 VPWR.n628 9.33404
R11019 VPWR.n633 VPWR.n632 9.33404
R11020 VPWR.n637 VPWR.n636 9.33404
R11021 VPWR.n640 VPWR.n639 9.33404
R11022 VPWR.n597 VPWR.n596 9.33404
R11023 VPWR.n2112 VPWR.n2111 9.33404
R11024 VPWR.n2116 VPWR.n2115 9.33404
R11025 VPWR.n2122 VPWR.n2121 9.33404
R11026 VPWR.n2126 VPWR.n2125 9.33404
R11027 VPWR.n2136 VPWR.n2135 9.33404
R11028 VPWR.n2142 VPWR.n2141 9.33404
R11029 VPWR.n2146 VPWR.n2145 9.33404
R11030 VPWR.n2152 VPWR.n2151 9.33404
R11031 VPWR.n2156 VPWR.n2155 9.33404
R11032 VPWR.n2162 VPWR.n2161 9.33404
R11033 VPWR.n2166 VPWR.n2165 9.33404
R11034 VPWR.n2172 VPWR.n2171 9.33404
R11035 VPWR.n2176 VPWR.n2175 9.33404
R11036 VPWR.n2182 VPWR.n2181 9.33404
R11037 VPWR.n2185 VPWR.n2184 9.33404
R11038 VPWR.n2132 VPWR.n2131 9.33404
R11039 VPWR.n736 VPWR.n735 9.33404
R11040 VPWR.n732 VPWR.n731 9.33404
R11041 VPWR.n728 VPWR.n727 9.33404
R11042 VPWR.n724 VPWR.n723 9.33404
R11043 VPWR.n716 VPWR.n715 9.33404
R11044 VPWR.n712 VPWR.n711 9.33404
R11045 VPWR.n708 VPWR.n707 9.33404
R11046 VPWR.n704 VPWR.n703 9.33404
R11047 VPWR.n700 VPWR.n699 9.33404
R11048 VPWR.n696 VPWR.n695 9.33404
R11049 VPWR.n692 VPWR.n691 9.33404
R11050 VPWR.n688 VPWR.n687 9.33404
R11051 VPWR.n684 VPWR.n683 9.33404
R11052 VPWR.n680 VPWR.n679 9.33404
R11053 VPWR.n677 VPWR.n676 9.33404
R11054 VPWR.n720 VPWR.n719 9.33404
R11055 VPWR.n2087 VPWR.n2086 9.33404
R11056 VPWR.n2083 VPWR.n2082 9.33404
R11057 VPWR.n2077 VPWR.n2076 9.33404
R11058 VPWR.n2073 VPWR.n2072 9.33404
R11059 VPWR.n2063 VPWR.n2062 9.33404
R11060 VPWR.n2057 VPWR.n2056 9.33404
R11061 VPWR.n2053 VPWR.n2052 9.33404
R11062 VPWR.n2047 VPWR.n2046 9.33404
R11063 VPWR.n2043 VPWR.n2042 9.33404
R11064 VPWR.n2037 VPWR.n2036 9.33404
R11065 VPWR.n2033 VPWR.n2032 9.33404
R11066 VPWR.n2027 VPWR.n2026 9.33404
R11067 VPWR.n2023 VPWR.n2022 9.33404
R11068 VPWR.n2017 VPWR.n2016 9.33404
R11069 VPWR.n2014 VPWR.n2013 9.33404
R11070 VPWR.n2067 VPWR.n2066 9.33404
R11071 VPWR.n773 VPWR.n772 9.33404
R11072 VPWR.n777 VPWR.n776 9.33404
R11073 VPWR.n781 VPWR.n780 9.33404
R11074 VPWR.n785 VPWR.n784 9.33404
R11075 VPWR.n793 VPWR.n792 9.33404
R11076 VPWR.n797 VPWR.n796 9.33404
R11077 VPWR.n801 VPWR.n800 9.33404
R11078 VPWR.n805 VPWR.n804 9.33404
R11079 VPWR.n809 VPWR.n808 9.33404
R11080 VPWR.n813 VPWR.n812 9.33404
R11081 VPWR.n817 VPWR.n816 9.33404
R11082 VPWR.n821 VPWR.n820 9.33404
R11083 VPWR.n825 VPWR.n824 9.33404
R11084 VPWR.n829 VPWR.n828 9.33404
R11085 VPWR.n832 VPWR.n831 9.33404
R11086 VPWR.n789 VPWR.n788 9.33404
R11087 VPWR.n1916 VPWR.n1915 9.33404
R11088 VPWR.n1920 VPWR.n1919 9.33404
R11089 VPWR.n1926 VPWR.n1925 9.33404
R11090 VPWR.n1930 VPWR.n1929 9.33404
R11091 VPWR.n1940 VPWR.n1939 9.33404
R11092 VPWR.n1946 VPWR.n1945 9.33404
R11093 VPWR.n1950 VPWR.n1949 9.33404
R11094 VPWR.n1956 VPWR.n1955 9.33404
R11095 VPWR.n1960 VPWR.n1959 9.33404
R11096 VPWR.n1966 VPWR.n1965 9.33404
R11097 VPWR.n1970 VPWR.n1969 9.33404
R11098 VPWR.n1976 VPWR.n1975 9.33404
R11099 VPWR.n1980 VPWR.n1979 9.33404
R11100 VPWR.n1986 VPWR.n1985 9.33404
R11101 VPWR.n1989 VPWR.n1988 9.33404
R11102 VPWR.n1936 VPWR.n1935 9.33404
R11103 VPWR.n928 VPWR.n927 9.33404
R11104 VPWR.n924 VPWR.n923 9.33404
R11105 VPWR.n920 VPWR.n919 9.33404
R11106 VPWR.n916 VPWR.n915 9.33404
R11107 VPWR.n908 VPWR.n907 9.33404
R11108 VPWR.n904 VPWR.n903 9.33404
R11109 VPWR.n900 VPWR.n899 9.33404
R11110 VPWR.n896 VPWR.n895 9.33404
R11111 VPWR.n892 VPWR.n891 9.33404
R11112 VPWR.n888 VPWR.n887 9.33404
R11113 VPWR.n884 VPWR.n883 9.33404
R11114 VPWR.n880 VPWR.n879 9.33404
R11115 VPWR.n876 VPWR.n875 9.33404
R11116 VPWR.n872 VPWR.n871 9.33404
R11117 VPWR.n869 VPWR.n868 9.33404
R11118 VPWR.n912 VPWR.n911 9.33404
R11119 VPWR.n1871 VPWR.n1870 9.33404
R11120 VPWR.n981 VPWR.n980 9.33404
R11121 VPWR.n1495 VPWR.n1494 9.33404
R11122 VPWR.n401 VPWR.n400 9.33404
R11123 VPWR.n2465 VPWR.n2464 9.33404
R11124 VPWR.n340 VPWR.n339 9.33404
R11125 VPWR.n977 VPWR.n976 9.33404
R11126 VPWR.n1491 VPWR.n1490 9.33404
R11127 VPWR.n1867 VPWR.n1866 9.33404
R11128 VPWR.n985 VPWR.n984 9.33404
R11129 VPWR.n1505 VPWR.n1504 9.33404
R11130 VPWR.n409 VPWR.n408 9.33404
R11131 VPWR.n417 VPWR.n416 9.33404
R11132 VPWR.n421 VPWR.n420 9.33404
R11133 VPWR.n425 VPWR.n424 9.33404
R11134 VPWR.n429 VPWR.n428 9.33404
R11135 VPWR.n433 VPWR.n432 9.33404
R11136 VPWR.n437 VPWR.n436 9.33404
R11137 VPWR.n441 VPWR.n440 9.33404
R11138 VPWR.n445 VPWR.n444 9.33404
R11139 VPWR.n448 VPWR.n447 9.33404
R11140 VPWR.n413 VPWR.n412 9.33404
R11141 VPWR.n2449 VPWR.n2448 9.33404
R11142 VPWR.n328 VPWR.n327 9.33404
R11143 VPWR.n989 VPWR.n988 9.33404
R11144 VPWR.n1509 VPWR.n1508 9.33404
R11145 VPWR.n1861 VPWR.n1860 9.33404
R11146 VPWR.n1851 VPWR.n1850 9.33404
R11147 VPWR.n1847 VPWR.n1846 9.33404
R11148 VPWR.n1841 VPWR.n1840 9.33404
R11149 VPWR.n1837 VPWR.n1836 9.33404
R11150 VPWR.n1831 VPWR.n1830 9.33404
R11151 VPWR.n1827 VPWR.n1826 9.33404
R11152 VPWR.n1821 VPWR.n1820 9.33404
R11153 VPWR.n1818 VPWR.n1817 9.33404
R11154 VPWR.n1857 VPWR.n1856 9.33404
R11155 VPWR.n993 VPWR.n992 9.33404
R11156 VPWR.n1519 VPWR.n1518 9.33404
R11157 VPWR.n2469 VPWR.n2468 9.33404
R11158 VPWR.n344 VPWR.n343 9.33404
R11159 VPWR.n1480 VPWR.n1130 9.33404
R11160 VPWR.n997 VPWR.n996 9.33404
R11161 VPWR.n1523 VPWR.n1522 9.33404
R11162 VPWR.n2439 VPWR.n2438 9.33404
R11163 VPWR.n2429 VPWR.n2428 9.33404
R11164 VPWR.n2425 VPWR.n2424 9.33404
R11165 VPWR.n2419 VPWR.n2418 9.33404
R11166 VPWR.n2415 VPWR.n2414 9.33404
R11167 VPWR.n2409 VPWR.n2408 9.33404
R11168 VPWR.n2406 VPWR.n2405 9.33404
R11169 VPWR.n2435 VPWR.n2434 9.33404
R11170 VPWR.n316 VPWR.n315 9.33404
R11171 VPWR.n1538 VPWR.n1537 9.33404
R11172 VPWR.n1001 VPWR.n1000 9.33404
R11173 VPWR.n1005 VPWR.n1004 9.33404
R11174 VPWR.n1009 VPWR.n1008 9.33404
R11175 VPWR.n1013 VPWR.n1012 9.33404
R11176 VPWR.n1017 VPWR.n1016 9.33404
R11177 VPWR.n1021 VPWR.n1020 9.33404
R11178 VPWR.n1024 VPWR.n1023 9.33404
R11179 VPWR.n969 VPWR.n968 9.33404
R11180 VPWR.n1474 VPWR.n1473 9.33404
R11181 VPWR.n312 VPWR.n311 9.33404
R11182 VPWR.n1763 VPWR.n1762 9.33404
R11183 VPWR.n308 VPWR.n307 9.33404
R11184 VPWR.n304 VPWR.n303 9.33404
R11185 VPWR.n296 VPWR.n295 9.33404
R11186 VPWR.n293 VPWR.n292 9.33404
R11187 VPWR.n300 VPWR.n299 9.33404
R11188 VPWR.n1751 VPWR.n1750 9.33404
R11189 VPWR.n1790 VPWR.n1789 9.33404
R11190 VPWR.n1793 VPWR.n1792 9.33404
R11191 VPWR.n1759 VPWR.n1758 9.33404
R11192 VPWR.n2714 VPWR 9.32394
R11193 VPWR.n2677 VPWR 9.32394
R11194 VPWR.n2640 VPWR 9.32394
R11195 VPWR VPWR.n2607 9.32394
R11196 VPWR.n18 VPWR.n17 9.3005
R11197 VPWR.n15 VPWR.n14 9.3005
R11198 VPWR.n13 VPWR.n2 9.3005
R11199 VPWR.n10 VPWR.n9 9.3005
R11200 VPWR.n8 VPWR.n3 9.3005
R11201 VPWR.n12 VPWR.n11 9.3005
R11202 VPWR.n16 VPWR.n0 9.3005
R11203 VPWR.n1254 VPWR.n1253 9.3005
R11204 VPWR.n1251 VPWR.n1250 9.3005
R11205 VPWR.n1249 VPWR.n1236 9.3005
R11206 VPWR.n1246 VPWR.n1244 9.3005
R11207 VPWR.n1243 VPWR.n1237 9.3005
R11208 VPWR.n1248 VPWR.n1247 9.3005
R11209 VPWR.n1252 VPWR.n1233 9.3005
R11210 VPWR.n1278 VPWR.n1277 9.3005
R11211 VPWR.n1272 VPWR.n1259 9.3005
R11212 VPWR.n1269 VPWR.n1267 9.3005
R11213 VPWR.n1266 VPWR.n1260 9.3005
R11214 VPWR.n1271 VPWR.n1270 9.3005
R11215 VPWR.n1274 VPWR.n1273 9.3005
R11216 VPWR.n1276 VPWR.n1256 9.3005
R11217 VPWR.n1301 VPWR.n1300 9.3005
R11218 VPWR.n1296 VPWR.n1283 9.3005
R11219 VPWR.n1293 VPWR.n1291 9.3005
R11220 VPWR.n1290 VPWR.n1284 9.3005
R11221 VPWR.n1295 VPWR.n1294 9.3005
R11222 VPWR.n1298 VPWR.n1297 9.3005
R11223 VPWR.n1299 VPWR.n1280 9.3005
R11224 VPWR.n1332 VPWR.n1303 9.3005
R11225 VPWR.n1331 VPWR.n1330 9.3005
R11226 VPWR.n1311 VPWR.n1310 9.3005
R11227 VPWR.n1313 VPWR.n1312 9.3005
R11228 VPWR.n1315 VPWR.n1309 9.3005
R11229 VPWR.n1317 VPWR.n1316 9.3005
R11230 VPWR.n1318 VPWR.n1308 9.3005
R11231 VPWR.n1320 VPWR.n1319 9.3005
R11232 VPWR.n1324 VPWR.n1305 9.3005
R11233 VPWR.n1326 VPWR.n1325 9.3005
R11234 VPWR.n1328 VPWR.n1327 9.3005
R11235 VPWR.n1334 VPWR.n1333 9.3005
R11236 VPWR.n1336 VPWR.n1335 9.3005
R11237 VPWR.n1375 VPWR.n1374 9.3005
R11238 VPWR.n1370 VPWR.n1338 9.3005
R11239 VPWR.n1369 VPWR.n1368 9.3005
R11240 VPWR.n1347 VPWR.n1346 9.3005
R11241 VPWR.n1349 VPWR.n1348 9.3005
R11242 VPWR.n1352 VPWR.n1342 9.3005
R11243 VPWR.n1354 VPWR.n1353 9.3005
R11244 VPWR.n1355 VPWR.n1341 9.3005
R11245 VPWR.n1357 VPWR.n1356 9.3005
R11246 VPWR.n1361 VPWR.n1340 9.3005
R11247 VPWR.n1363 VPWR.n1362 9.3005
R11248 VPWR.n1365 VPWR.n1364 9.3005
R11249 VPWR.n1372 VPWR.n1371 9.3005
R11250 VPWR.n1408 VPWR.n1407 9.3005
R11251 VPWR.n1386 VPWR.n1385 9.3005
R11252 VPWR.n1388 VPWR.n1387 9.3005
R11253 VPWR.n1391 VPWR.n1381 9.3005
R11254 VPWR.n1393 VPWR.n1392 9.3005
R11255 VPWR.n1394 VPWR.n1380 9.3005
R11256 VPWR.n1396 VPWR.n1395 9.3005
R11257 VPWR.n1400 VPWR.n1379 9.3005
R11258 VPWR.n1402 VPWR.n1401 9.3005
R11259 VPWR.n1404 VPWR.n1403 9.3005
R11260 VPWR.n1409 VPWR.n1377 9.3005
R11261 VPWR.n1411 VPWR.n1410 9.3005
R11262 VPWR.n1445 VPWR.n1444 9.3005
R11263 VPWR.n1423 VPWR.n1422 9.3005
R11264 VPWR.n1425 VPWR.n1424 9.3005
R11265 VPWR.n1428 VPWR.n1418 9.3005
R11266 VPWR.n1430 VPWR.n1429 9.3005
R11267 VPWR.n1431 VPWR.n1417 9.3005
R11268 VPWR.n1433 VPWR.n1432 9.3005
R11269 VPWR.n1437 VPWR.n1416 9.3005
R11270 VPWR.n1439 VPWR.n1438 9.3005
R11271 VPWR.n1441 VPWR.n1440 9.3005
R11272 VPWR.n2807 VPWR.n2806 9.3005
R11273 VPWR.n2808 VPWR.n2800 9.3005
R11274 VPWR.n2809 VPWR.n2799 9.3005
R11275 VPWR.n2810 VPWR.n2798 9.3005
R11276 VPWR.n2812 VPWR.n2811 9.3005
R11277 VPWR.n2796 VPWR.n2795 9.3005
R11278 VPWR.n2790 VPWR.n2789 9.3005
R11279 VPWR.n2791 VPWR.n2781 9.3005
R11280 VPWR.n2793 VPWR.n2792 9.3005
R11281 VPWR.n2794 VPWR.n2779 9.3005
R11282 VPWR.n2777 VPWR.n2776 9.3005
R11283 VPWR.n2775 VPWR.n2759 9.3005
R11284 VPWR.n2770 VPWR.n2769 9.3005
R11285 VPWR.n2771 VPWR.n2761 9.3005
R11286 VPWR.n2773 VPWR.n2772 9.3005
R11287 VPWR.n2757 VPWR.n2756 9.3005
R11288 VPWR.n2751 VPWR.n2750 9.3005
R11289 VPWR.n2752 VPWR.n2742 9.3005
R11290 VPWR.n2754 VPWR.n2753 9.3005
R11291 VPWR.n2755 VPWR.n2740 9.3005
R11292 VPWR.n2738 VPWR.n2737 9.3005
R11293 VPWR.n2718 VPWR.n2717 9.3005
R11294 VPWR.n2719 VPWR.n2713 9.3005
R11295 VPWR.n2721 VPWR.n2720 9.3005
R11296 VPWR.n2723 VPWR.n2711 9.3005
R11297 VPWR.n2725 VPWR.n2724 9.3005
R11298 VPWR.n2727 VPWR.n2726 9.3005
R11299 VPWR.n2728 VPWR.n2707 9.3005
R11300 VPWR.n2732 VPWR.n2731 9.3005
R11301 VPWR.n2733 VPWR.n2706 9.3005
R11302 VPWR.n2735 VPWR.n2734 9.3005
R11303 VPWR.n2736 VPWR.n2704 9.3005
R11304 VPWR.n2702 VPWR.n2701 9.3005
R11305 VPWR.n2682 VPWR.n2681 9.3005
R11306 VPWR.n2683 VPWR.n2676 9.3005
R11307 VPWR.n2685 VPWR.n2684 9.3005
R11308 VPWR.n2687 VPWR.n2673 9.3005
R11309 VPWR.n2689 VPWR.n2688 9.3005
R11310 VPWR.n2691 VPWR.n2690 9.3005
R11311 VPWR.n2692 VPWR.n2669 9.3005
R11312 VPWR.n2695 VPWR.n2694 9.3005
R11313 VPWR.n2696 VPWR.n2668 9.3005
R11314 VPWR.n2698 VPWR.n2697 9.3005
R11315 VPWR.n2699 VPWR.n2666 9.3005
R11316 VPWR.n2645 VPWR.n2644 9.3005
R11317 VPWR.n2646 VPWR.n2639 9.3005
R11318 VPWR.n2648 VPWR.n2647 9.3005
R11319 VPWR.n2650 VPWR.n2636 9.3005
R11320 VPWR.n2652 VPWR.n2651 9.3005
R11321 VPWR.n2654 VPWR.n2653 9.3005
R11322 VPWR.n2655 VPWR.n2632 9.3005
R11323 VPWR.n2658 VPWR.n2657 9.3005
R11324 VPWR.n2659 VPWR.n2631 9.3005
R11325 VPWR.n2661 VPWR.n2660 9.3005
R11326 VPWR.n2662 VPWR.n2629 9.3005
R11327 VPWR.n2627 VPWR.n2626 9.3005
R11328 VPWR.n2609 VPWR.n2608 9.3005
R11329 VPWR.n2611 VPWR.n2604 9.3005
R11330 VPWR.n2616 VPWR.n2615 9.3005
R11331 VPWR.n2617 VPWR.n2603 9.3005
R11332 VPWR.n2619 VPWR.n2618 9.3005
R11333 VPWR.n2621 VPWR.n2600 9.3005
R11334 VPWR.n2623 VPWR.n2622 9.3005
R11335 VPWR.n2625 VPWR.n2624 9.3005
R11336 VPWR.n2505 VPWR.n2504 9.3005
R11337 VPWR.n2569 VPWR.n2568 9.3005
R11338 VPWR.n2509 VPWR.n2508 9.3005
R11339 VPWR.n2553 VPWR.n2552 9.3005
R11340 VPWR.n2545 VPWR.n2544 9.3005
R11341 VPWR.n2533 VPWR.n2532 9.3005
R11342 VPWR.n2529 VPWR.n2528 9.3005
R11343 VPWR.n1222 VPWR.n1221 9.3005
R11344 VPWR.n2521 VPWR.n2520 9.3005
R11345 VPWR.n1184 VPWR.n1102 9.3005
R11346 VPWR.n1218 VPWR.n1094 9.3005
R11347 VPWR.n2541 VPWR.n2540 9.3005
R11348 VPWR.n1215 VPWR.n1092 9.3005
R11349 VPWR.n1212 VPWR.n1211 9.3005
R11350 VPWR.n2517 VPWR.n2516 9.3005
R11351 VPWR.n1181 VPWR.n1104 9.3005
R11352 VPWR.n1204 VPWR.n1084 9.3005
R11353 VPWR.n2557 VPWR.n2556 9.3005
R11354 VPWR.n1201 VPWR.n1082 9.3005
R11355 VPWR.n1592 VPWR.n1591 9.3005
R11356 VPWR.n2565 VPWR.n2564 9.3005
R11357 VPWR.n1198 VPWR.n1197 9.3005
R11358 VPWR.n1190 VPWR.n1074 9.3005
R11359 VPWR.n1742 VPWR.n1741 9.3005
R11360 VPWR.n1187 VPWR.n1071 9.3005
R11361 VPWR.n2577 VPWR.n2576 9.3005
R11362 VPWR.n2581 VPWR.n2580 9.3005
R11363 VPWR.n2592 VPWR.n2591 9.3005
R11364 VPWR.n2589 VPWR.n2588 9.3005
R11365 VPWR.n1738 VPWR.n1737 9.3005
R11366 VPWR.n1063 VPWR.n1062 9.3005
R11367 VPWR.n1596 VPWR.n1595 9.3005
R11368 VPWR.n1275 VPWR.n1274 8.28285
R11369 VPWR.n2774 VPWR.n2773 8.28285
R11370 VPWR.n1607 VPWR.n1109 8.25914
R11371 VPWR.n1728 VPWR.n1727 8.25914
R11372 VPWR.n281 VPWR.n113 8.25914
R11373 VPWR.n136 VPWR.n124 8.25914
R11374 VPWR.n1780 VPWR.n1779 7.91351
R11375 VPWR.n1771 VPWR.n1770 7.9105
R11376 VPWR.n1042 VPWR.n1041 7.9105
R11377 VPWR.n1546 VPWR.n1545 7.9105
R11378 VPWR.n1551 VPWR.n1550 7.9105
R11379 VPWR.n1556 VPWR.n1555 7.9105
R11380 VPWR.n1561 VPWR.n1560 7.9105
R11381 VPWR.n1566 VPWR.n1565 7.9105
R11382 VPWR.n1571 VPWR.n1570 7.9105
R11383 VPWR.n1576 VPWR.n1575 7.9105
R11384 VPWR.n1581 VPWR.n1580 7.9105
R11385 VPWR.n1136 VPWR.n1135 7.9105
R11386 VPWR.n1461 VPWR.n1460 7.9105
R11387 VPWR.n1456 VPWR.n1455 7.9105
R11388 VPWR.n1776 VPWR.n1775 7.9105
R11389 VPWR.n1784 VPWR.n1783 7.9105
R11390 VPWR.n282 VPWR.n281 7.9105
R11391 VPWR.n280 VPWR.n279 7.9105
R11392 VPWR.n268 VPWR.n267 7.9105
R11393 VPWR.n256 VPWR.n255 7.9105
R11394 VPWR.n244 VPWR.n243 7.9105
R11395 VPWR.n232 VPWR.n231 7.9105
R11396 VPWR.n220 VPWR.n219 7.9105
R11397 VPWR.n208 VPWR.n207 7.9105
R11398 VPWR.n196 VPWR.n195 7.9105
R11399 VPWR.n184 VPWR.n183 7.9105
R11400 VPWR.n172 VPWR.n171 7.9105
R11401 VPWR.n160 VPWR.n159 7.9105
R11402 VPWR.n148 VPWR.n147 7.9105
R11403 VPWR.n136 VPWR.n135 7.9105
R11404 VPWR.n1727 VPWR.n1726 7.9105
R11405 VPWR.n1715 VPWR.n1714 7.9105
R11406 VPWR.n1701 VPWR.n1068 7.9105
R11407 VPWR.n1690 VPWR.n1689 7.9105
R11408 VPWR.n1688 VPWR.n1687 7.9105
R11409 VPWR.n1674 VPWR.n1079 7.9105
R11410 VPWR.n1663 VPWR.n1662 7.9105
R11411 VPWR.n1661 VPWR.n1660 7.9105
R11412 VPWR.n1647 VPWR.n1089 7.9105
R11413 VPWR.n1636 VPWR.n1635 7.9105
R11414 VPWR.n1634 VPWR.n1633 7.9105
R11415 VPWR.n1620 VPWR.n1099 7.9105
R11416 VPWR.n1609 VPWR.n1608 7.9105
R11417 VPWR.n1607 VPWR.n1606 7.9105
R11418 VPWR.n26 VPWR.n24 7.8627
R11419 VPWR.n7 VPWR.n6 7.56315
R11420 VPWR.n1242 VPWR.n1241 7.56315
R11421 VPWR.n1265 VPWR.n1264 7.56315
R11422 VPWR.n1289 VPWR.n1288 7.56315
R11423 VPWR.n2805 VPWR.n2803 6.4511
R11424 VPWR.n2788 VPWR.n2785 6.4511
R11425 VPWR.n2768 VPWR.n2765 6.4511
R11426 VPWR.n2749 VPWR.n2746 6.4511
R11427 VPWR.n1362 VPWR.n1339 6.4005
R11428 VPWR.n1401 VPWR.n1378 6.4005
R11429 VPWR.n1438 VPWR.n1415 6.4005
R11430 VPWR.n2723 VPWR.n2722 6.4005
R11431 VPWR.n2693 VPWR.n2692 6.4005
R11432 VPWR.n2656 VPWR.n2655 6.4005
R11433 VPWR.n2622 VPWR.n2599 6.4005
R11434 VPWR.n1595 VPWR.n1122 6.04494
R11435 VPWR.n2505 VPWR.n99 6.04494
R11436 VPWR.n1467 VPWR.n1231 6.04494
R11437 VPWR.n351 VPWR.n290 6.04494
R11438 VPWR.n2568 VPWR.n68 6.04494
R11439 VPWR.n1534 VPWR.n1153 6.04494
R11440 VPWR.n348 VPWR.n346 6.04494
R11441 VPWR.n2508 VPWR.n98 6.04494
R11442 VPWR.n965 VPWR.n963 6.04494
R11443 VPWR.n2478 VPWR.n356 6.04494
R11444 VPWR.n2475 VPWR.n357 6.04494
R11445 VPWR.n320 VPWR.n318 6.04494
R11446 VPWR.n2553 VPWR.n75 6.04494
R11447 VPWR.n973 VPWR.n971 6.04494
R11448 VPWR.n2445 VPWR.n369 6.04494
R11449 VPWR.n324 VPWR.n322 6.04494
R11450 VPWR.n2544 VPWR.n80 6.04494
R11451 VPWR.n1890 VPWR.n932 6.04494
R11452 VPWR.n1887 VPWR.n933 6.04494
R11453 VPWR.n1880 VPWR.n936 6.04494
R11454 VPWR.n389 VPWR.n387 6.04494
R11455 VPWR.n393 VPWR.n391 6.04494
R11456 VPWR.n397 VPWR.n395 6.04494
R11457 VPWR.n2455 VPWR.n365 6.04494
R11458 VPWR.n332 VPWR.n330 6.04494
R11459 VPWR.n2532 VPWR.n86 6.04494
R11460 VPWR.n1877 VPWR.n937 6.04494
R11461 VPWR.n405 VPWR.n403 6.04494
R11462 VPWR.n2458 VPWR.n364 6.04494
R11463 VPWR.n336 VPWR.n334 6.04494
R11464 VPWR.n2529 VPWR.n87 6.04494
R11465 VPWR.n2308 VPWR.n481 6.04494
R11466 VPWR.n2311 VPWR.n480 6.04494
R11467 VPWR.n2318 VPWR.n477 6.04494
R11468 VPWR.n2321 VPWR.n476 6.04494
R11469 VPWR.n2331 VPWR.n472 6.04494
R11470 VPWR.n2338 VPWR.n469 6.04494
R11471 VPWR.n2341 VPWR.n468 6.04494
R11472 VPWR.n2348 VPWR.n465 6.04494
R11473 VPWR.n2351 VPWR.n464 6.04494
R11474 VPWR.n2358 VPWR.n461 6.04494
R11475 VPWR.n2361 VPWR.n460 6.04494
R11476 VPWR.n2368 VPWR.n457 6.04494
R11477 VPWR.n2371 VPWR.n456 6.04494
R11478 VPWR.n2378 VPWR.n453 6.04494
R11479 VPWR.n2380 VPWR.n452 6.04494
R11480 VPWR.n2328 VPWR.n473 6.04494
R11481 VPWR.n543 VPWR.n482 6.04494
R11482 VPWR.n540 VPWR.n538 6.04494
R11483 VPWR.n536 VPWR.n534 6.04494
R11484 VPWR.n532 VPWR.n530 6.04494
R11485 VPWR.n524 VPWR.n522 6.04494
R11486 VPWR.n520 VPWR.n518 6.04494
R11487 VPWR.n516 VPWR.n514 6.04494
R11488 VPWR.n512 VPWR.n510 6.04494
R11489 VPWR.n508 VPWR.n506 6.04494
R11490 VPWR.n504 VPWR.n502 6.04494
R11491 VPWR.n500 VPWR.n498 6.04494
R11492 VPWR.n496 VPWR.n494 6.04494
R11493 VPWR.n492 VPWR.n490 6.04494
R11494 VPWR.n488 VPWR.n486 6.04494
R11495 VPWR.n485 VPWR.n483 6.04494
R11496 VPWR.n528 VPWR.n526 6.04494
R11497 VPWR.n2282 VPWR.n548 6.04494
R11498 VPWR.n2279 VPWR.n549 6.04494
R11499 VPWR.n2272 VPWR.n552 6.04494
R11500 VPWR.n2269 VPWR.n553 6.04494
R11501 VPWR.n2259 VPWR.n557 6.04494
R11502 VPWR.n2252 VPWR.n560 6.04494
R11503 VPWR.n2249 VPWR.n561 6.04494
R11504 VPWR.n2242 VPWR.n564 6.04494
R11505 VPWR.n2239 VPWR.n565 6.04494
R11506 VPWR.n2232 VPWR.n568 6.04494
R11507 VPWR.n2229 VPWR.n569 6.04494
R11508 VPWR.n2222 VPWR.n572 6.04494
R11509 VPWR.n2219 VPWR.n573 6.04494
R11510 VPWR.n2212 VPWR.n576 6.04494
R11511 VPWR.n2210 VPWR.n577 6.04494
R11512 VPWR.n2262 VPWR.n556 6.04494
R11513 VPWR.n581 VPWR.n579 6.04494
R11514 VPWR.n585 VPWR.n583 6.04494
R11515 VPWR.n589 VPWR.n587 6.04494
R11516 VPWR.n593 VPWR.n591 6.04494
R11517 VPWR.n601 VPWR.n599 6.04494
R11518 VPWR.n605 VPWR.n603 6.04494
R11519 VPWR.n609 VPWR.n607 6.04494
R11520 VPWR.n613 VPWR.n611 6.04494
R11521 VPWR.n617 VPWR.n615 6.04494
R11522 VPWR.n621 VPWR.n619 6.04494
R11523 VPWR.n625 VPWR.n623 6.04494
R11524 VPWR.n629 VPWR.n627 6.04494
R11525 VPWR.n633 VPWR.n631 6.04494
R11526 VPWR.n637 VPWR.n635 6.04494
R11527 VPWR.n639 VPWR.n578 6.04494
R11528 VPWR.n597 VPWR.n595 6.04494
R11529 VPWR.n2112 VPWR.n673 6.04494
R11530 VPWR.n2115 VPWR.n672 6.04494
R11531 VPWR.n2122 VPWR.n669 6.04494
R11532 VPWR.n2125 VPWR.n668 6.04494
R11533 VPWR.n2135 VPWR.n664 6.04494
R11534 VPWR.n2142 VPWR.n661 6.04494
R11535 VPWR.n2145 VPWR.n660 6.04494
R11536 VPWR.n2152 VPWR.n657 6.04494
R11537 VPWR.n2155 VPWR.n656 6.04494
R11538 VPWR.n2162 VPWR.n653 6.04494
R11539 VPWR.n2165 VPWR.n652 6.04494
R11540 VPWR.n2172 VPWR.n649 6.04494
R11541 VPWR.n2175 VPWR.n648 6.04494
R11542 VPWR.n2182 VPWR.n645 6.04494
R11543 VPWR.n2184 VPWR.n644 6.04494
R11544 VPWR.n2132 VPWR.n665 6.04494
R11545 VPWR.n735 VPWR.n674 6.04494
R11546 VPWR.n732 VPWR.n730 6.04494
R11547 VPWR.n728 VPWR.n726 6.04494
R11548 VPWR.n724 VPWR.n722 6.04494
R11549 VPWR.n716 VPWR.n714 6.04494
R11550 VPWR.n712 VPWR.n710 6.04494
R11551 VPWR.n708 VPWR.n706 6.04494
R11552 VPWR.n704 VPWR.n702 6.04494
R11553 VPWR.n700 VPWR.n698 6.04494
R11554 VPWR.n696 VPWR.n694 6.04494
R11555 VPWR.n692 VPWR.n690 6.04494
R11556 VPWR.n688 VPWR.n686 6.04494
R11557 VPWR.n684 VPWR.n682 6.04494
R11558 VPWR.n680 VPWR.n678 6.04494
R11559 VPWR.n677 VPWR.n675 6.04494
R11560 VPWR.n720 VPWR.n718 6.04494
R11561 VPWR.n2086 VPWR.n740 6.04494
R11562 VPWR.n2083 VPWR.n741 6.04494
R11563 VPWR.n2076 VPWR.n744 6.04494
R11564 VPWR.n2073 VPWR.n745 6.04494
R11565 VPWR.n2063 VPWR.n749 6.04494
R11566 VPWR.n2056 VPWR.n752 6.04494
R11567 VPWR.n2053 VPWR.n753 6.04494
R11568 VPWR.n2046 VPWR.n756 6.04494
R11569 VPWR.n2043 VPWR.n757 6.04494
R11570 VPWR.n2036 VPWR.n760 6.04494
R11571 VPWR.n2033 VPWR.n761 6.04494
R11572 VPWR.n2026 VPWR.n764 6.04494
R11573 VPWR.n2023 VPWR.n765 6.04494
R11574 VPWR.n2016 VPWR.n768 6.04494
R11575 VPWR.n2014 VPWR.n769 6.04494
R11576 VPWR.n2066 VPWR.n748 6.04494
R11577 VPWR.n773 VPWR.n771 6.04494
R11578 VPWR.n777 VPWR.n775 6.04494
R11579 VPWR.n781 VPWR.n779 6.04494
R11580 VPWR.n785 VPWR.n783 6.04494
R11581 VPWR.n793 VPWR.n791 6.04494
R11582 VPWR.n797 VPWR.n795 6.04494
R11583 VPWR.n801 VPWR.n799 6.04494
R11584 VPWR.n805 VPWR.n803 6.04494
R11585 VPWR.n809 VPWR.n807 6.04494
R11586 VPWR.n813 VPWR.n811 6.04494
R11587 VPWR.n817 VPWR.n815 6.04494
R11588 VPWR.n821 VPWR.n819 6.04494
R11589 VPWR.n825 VPWR.n823 6.04494
R11590 VPWR.n829 VPWR.n827 6.04494
R11591 VPWR.n831 VPWR.n770 6.04494
R11592 VPWR.n789 VPWR.n787 6.04494
R11593 VPWR.n1916 VPWR.n865 6.04494
R11594 VPWR.n1919 VPWR.n864 6.04494
R11595 VPWR.n1926 VPWR.n861 6.04494
R11596 VPWR.n1929 VPWR.n860 6.04494
R11597 VPWR.n1939 VPWR.n856 6.04494
R11598 VPWR.n1946 VPWR.n853 6.04494
R11599 VPWR.n1949 VPWR.n852 6.04494
R11600 VPWR.n1956 VPWR.n849 6.04494
R11601 VPWR.n1959 VPWR.n848 6.04494
R11602 VPWR.n1966 VPWR.n845 6.04494
R11603 VPWR.n1969 VPWR.n844 6.04494
R11604 VPWR.n1976 VPWR.n841 6.04494
R11605 VPWR.n1979 VPWR.n840 6.04494
R11606 VPWR.n1986 VPWR.n837 6.04494
R11607 VPWR.n1988 VPWR.n836 6.04494
R11608 VPWR.n1936 VPWR.n857 6.04494
R11609 VPWR.n927 VPWR.n866 6.04494
R11610 VPWR.n924 VPWR.n922 6.04494
R11611 VPWR.n920 VPWR.n918 6.04494
R11612 VPWR.n916 VPWR.n914 6.04494
R11613 VPWR.n908 VPWR.n906 6.04494
R11614 VPWR.n904 VPWR.n902 6.04494
R11615 VPWR.n900 VPWR.n898 6.04494
R11616 VPWR.n896 VPWR.n894 6.04494
R11617 VPWR.n892 VPWR.n890 6.04494
R11618 VPWR.n888 VPWR.n886 6.04494
R11619 VPWR.n884 VPWR.n882 6.04494
R11620 VPWR.n880 VPWR.n878 6.04494
R11621 VPWR.n876 VPWR.n874 6.04494
R11622 VPWR.n872 VPWR.n870 6.04494
R11623 VPWR.n869 VPWR.n867 6.04494
R11624 VPWR.n912 VPWR.n910 6.04494
R11625 VPWR.n1870 VPWR.n940 6.04494
R11626 VPWR.n981 VPWR.n979 6.04494
R11627 VPWR.n1494 VPWR.n1227 6.04494
R11628 VPWR.n1221 VPWR.n1179 6.04494
R11629 VPWR.n401 VPWR.n399 6.04494
R11630 VPWR.n2465 VPWR.n361 6.04494
R11631 VPWR.n340 VPWR.n338 6.04494
R11632 VPWR.n2520 VPWR.n92 6.04494
R11633 VPWR.n977 VPWR.n975 6.04494
R11634 VPWR.n1491 VPWR.n1485 6.04494
R11635 VPWR.n1184 VPWR.n1183 6.04494
R11636 VPWR.n1867 VPWR.n941 6.04494
R11637 VPWR.n985 VPWR.n983 6.04494
R11638 VPWR.n1505 VPWR.n1173 6.04494
R11639 VPWR.n1218 VPWR.n1217 6.04494
R11640 VPWR.n409 VPWR.n407 6.04494
R11641 VPWR.n417 VPWR.n415 6.04494
R11642 VPWR.n421 VPWR.n419 6.04494
R11643 VPWR.n425 VPWR.n423 6.04494
R11644 VPWR.n429 VPWR.n427 6.04494
R11645 VPWR.n433 VPWR.n431 6.04494
R11646 VPWR.n437 VPWR.n435 6.04494
R11647 VPWR.n441 VPWR.n439 6.04494
R11648 VPWR.n445 VPWR.n443 6.04494
R11649 VPWR.n447 VPWR.n386 6.04494
R11650 VPWR.n413 VPWR.n411 6.04494
R11651 VPWR.n2448 VPWR.n368 6.04494
R11652 VPWR.n328 VPWR.n326 6.04494
R11653 VPWR.n2541 VPWR.n81 6.04494
R11654 VPWR.n989 VPWR.n987 6.04494
R11655 VPWR.n1508 VPWR.n1169 6.04494
R11656 VPWR.n1215 VPWR.n1214 6.04494
R11657 VPWR.n1860 VPWR.n944 6.04494
R11658 VPWR.n1850 VPWR.n948 6.04494
R11659 VPWR.n1847 VPWR.n949 6.04494
R11660 VPWR.n1840 VPWR.n952 6.04494
R11661 VPWR.n1837 VPWR.n953 6.04494
R11662 VPWR.n1830 VPWR.n956 6.04494
R11663 VPWR.n1827 VPWR.n957 6.04494
R11664 VPWR.n1820 VPWR.n960 6.04494
R11665 VPWR.n1818 VPWR.n961 6.04494
R11666 VPWR.n1857 VPWR.n945 6.04494
R11667 VPWR.n993 VPWR.n991 6.04494
R11668 VPWR.n1519 VPWR.n1163 6.04494
R11669 VPWR.n1212 VPWR.n1206 6.04494
R11670 VPWR.n2468 VPWR.n360 6.04494
R11671 VPWR.n344 VPWR.n342 6.04494
R11672 VPWR.n2517 VPWR.n93 6.04494
R11673 VPWR.n1480 VPWR.n1479 6.04494
R11674 VPWR.n1181 VPWR.n1180 6.04494
R11675 VPWR.n997 VPWR.n995 6.04494
R11676 VPWR.n1522 VPWR.n1159 6.04494
R11677 VPWR.n1204 VPWR.n1203 6.04494
R11678 VPWR.n2438 VPWR.n372 6.04494
R11679 VPWR.n2428 VPWR.n376 6.04494
R11680 VPWR.n2425 VPWR.n377 6.04494
R11681 VPWR.n2418 VPWR.n380 6.04494
R11682 VPWR.n2415 VPWR.n381 6.04494
R11683 VPWR.n2408 VPWR.n384 6.04494
R11684 VPWR.n2406 VPWR.n385 6.04494
R11685 VPWR.n2435 VPWR.n373 6.04494
R11686 VPWR.n316 VPWR.n314 6.04494
R11687 VPWR.n2556 VPWR.n74 6.04494
R11688 VPWR.n1537 VPWR.n1149 6.04494
R11689 VPWR.n1201 VPWR.n1200 6.04494
R11690 VPWR.n1001 VPWR.n999 6.04494
R11691 VPWR.n1005 VPWR.n1003 6.04494
R11692 VPWR.n1009 VPWR.n1007 6.04494
R11693 VPWR.n1013 VPWR.n1011 6.04494
R11694 VPWR.n1017 VPWR.n1015 6.04494
R11695 VPWR.n1021 VPWR.n1019 6.04494
R11696 VPWR.n1023 VPWR.n962 6.04494
R11697 VPWR.n969 VPWR.n967 6.04494
R11698 VPWR.n1474 VPWR.n1472 6.04494
R11699 VPWR.n1592 VPWR.n1123 6.04494
R11700 VPWR.n312 VPWR.n310 6.04494
R11701 VPWR.n2565 VPWR.n69 6.04494
R11702 VPWR.n1198 VPWR.n1192 6.04494
R11703 VPWR.n1762 VPWR.n1049 6.04494
R11704 VPWR.n1190 VPWR.n1189 6.04494
R11705 VPWR.n308 VPWR.n306 6.04494
R11706 VPWR.n304 VPWR.n302 6.04494
R11707 VPWR.n296 VPWR.n294 6.04494
R11708 VPWR.n293 VPWR.n291 6.04494
R11709 VPWR.n300 VPWR.n298 6.04494
R11710 VPWR.n1741 VPWR.n1058 6.04494
R11711 VPWR.n1750 VPWR.n1748 6.04494
R11712 VPWR.n1790 VPWR.n1036 6.04494
R11713 VPWR.n1792 VPWR.n1032 6.04494
R11714 VPWR.n1759 VPWR.n1053 6.04494
R11715 VPWR.n1187 VPWR.n1186 6.04494
R11716 VPWR.n2577 VPWR.n63 6.04494
R11717 VPWR.n2580 VPWR.n62 6.04494
R11718 VPWR.n2589 VPWR.n57 6.04494
R11719 VPWR.n2591 VPWR.n56 6.04494
R11720 VPWR.n1738 VPWR.n1059 6.04494
R11721 VPWR.n1062 VPWR.n1061 6.04494
R11722 VPWR.n2785 VPWR.n2784 5.39628
R11723 VPWR.n2765 VPWR.n2764 5.39628
R11724 VPWR.n2746 VPWR.n2745 5.39628
R11725 VPWR.n54 VPWR 4.72593
R11726 VPWR.n52 VPWR 4.72593
R11727 VPWR.n50 VPWR 4.72593
R11728 VPWR.n48 VPWR 4.72593
R11729 VPWR.n46 VPWR 4.72593
R11730 VPWR.n44 VPWR 4.72593
R11731 VPWR.n42 VPWR 4.72593
R11732 VPWR.n40 VPWR 4.72593
R11733 VPWR.n38 VPWR 4.72593
R11734 VPWR.n36 VPWR 4.72593
R11735 VPWR.n34 VPWR 4.72593
R11736 VPWR.n32 VPWR 4.72593
R11737 VPWR.n30 VPWR 4.72593
R11738 VPWR.n28 VPWR 4.72593
R11739 VPWR.n26 VPWR 4.72593
R11740 VPWR.n1446 VPWR.n1445 4.55954
R11741 VPWR.n2571 VPWR.n2570 4.5005
R11742 VPWR.n2511 VPWR.n2510 4.5005
R11743 VPWR.n2551 VPWR.n2550 4.5005
R11744 VPWR.n319 VPWR.n77 4.5005
R11745 VPWR.n2547 VPWR.n2546 4.5005
R11746 VPWR.n323 VPWR.n78 4.5005
R11747 VPWR.n2535 VPWR.n2534 4.5005
R11748 VPWR.n331 VPWR.n84 4.5005
R11749 VPWR.n2454 VPWR.n2453 4.5005
R11750 VPWR.n2527 VPWR.n2526 4.5005
R11751 VPWR.n335 VPWR.n89 4.5005
R11752 VPWR.n2460 VPWR.n2459 4.5005
R11753 VPWR.n1498 VPWR.n1223 4.5005
R11754 VPWR.n1497 VPWR.n1495 4.5005
R11755 VPWR.n980 VPWR.n939 4.5005
R11756 VPWR.n1872 VPWR.n1871 4.5005
R11757 VPWR.n911 VPWR.n858 4.5005
R11758 VPWR.n1935 VPWR.n1934 4.5005
R11759 VPWR.n788 VPWR.n747 4.5005
R11760 VPWR.n2068 VPWR.n2067 4.5005
R11761 VPWR.n719 VPWR.n666 4.5005
R11762 VPWR.n2131 VPWR.n2130 4.5005
R11763 VPWR.n596 VPWR.n555 4.5005
R11764 VPWR.n2264 VPWR.n2263 4.5005
R11765 VPWR.n527 VPWR.n474 4.5005
R11766 VPWR.n2327 VPWR.n2326 4.5005
R11767 VPWR.n404 VPWR.n363 4.5005
R11768 VPWR.n2523 VPWR.n2522 4.5005
R11769 VPWR.n339 VPWR.n90 4.5005
R11770 VPWR.n2464 VPWR.n2463 4.5005
R11771 VPWR.n400 VPWR.n362 4.5005
R11772 VPWR.n2323 VPWR.n2322 4.5005
R11773 VPWR.n531 VPWR.n475 4.5005
R11774 VPWR.n2268 VPWR.n2267 4.5005
R11775 VPWR.n592 VPWR.n554 4.5005
R11776 VPWR.n2127 VPWR.n2126 4.5005
R11777 VPWR.n723 VPWR.n667 4.5005
R11778 VPWR.n2072 VPWR.n2071 4.5005
R11779 VPWR.n784 VPWR.n746 4.5005
R11780 VPWR.n1931 VPWR.n1930 4.5005
R11781 VPWR.n915 VPWR.n859 4.5005
R11782 VPWR.n1488 VPWR.n1486 4.5005
R11783 VPWR.n1490 VPWR.n1489 4.5005
R11784 VPWR.n976 VPWR.n938 4.5005
R11785 VPWR.n1876 VPWR.n1875 4.5005
R11786 VPWR.n1501 VPWR.n1174 4.5005
R11787 VPWR.n1504 VPWR.n1503 4.5005
R11788 VPWR.n984 VPWR.n942 4.5005
R11789 VPWR.n1866 VPWR.n1865 4.5005
R11790 VPWR.n907 VPWR.n855 4.5005
R11791 VPWR.n1941 VPWR.n1940 4.5005
R11792 VPWR.n792 VPWR.n750 4.5005
R11793 VPWR.n2062 VPWR.n2061 4.5005
R11794 VPWR.n715 VPWR.n663 4.5005
R11795 VPWR.n2137 VPWR.n2136 4.5005
R11796 VPWR.n600 VPWR.n558 4.5005
R11797 VPWR.n2258 VPWR.n2257 4.5005
R11798 VPWR.n523 VPWR.n471 4.5005
R11799 VPWR.n2333 VPWR.n2332 4.5005
R11800 VPWR.n408 VPWR.n366 4.5005
R11801 VPWR.n2539 VPWR.n2538 4.5005
R11802 VPWR.n327 VPWR.n83 4.5005
R11803 VPWR.n2450 VPWR.n2449 4.5005
R11804 VPWR.n412 VPWR.n367 4.5005
R11805 VPWR.n2337 VPWR.n2336 4.5005
R11806 VPWR.n519 VPWR.n470 4.5005
R11807 VPWR.n2254 VPWR.n2253 4.5005
R11808 VPWR.n604 VPWR.n559 4.5005
R11809 VPWR.n2141 VPWR.n2140 4.5005
R11810 VPWR.n711 VPWR.n662 4.5005
R11811 VPWR.n2058 VPWR.n2057 4.5005
R11812 VPWR.n796 VPWR.n751 4.5005
R11813 VPWR.n1945 VPWR.n1944 4.5005
R11814 VPWR.n903 VPWR.n854 4.5005
R11815 VPWR.n1512 VPWR.n1165 4.5005
R11816 VPWR.n1511 VPWR.n1509 4.5005
R11817 VPWR.n988 VPWR.n943 4.5005
R11818 VPWR.n1862 VPWR.n1861 4.5005
R11819 VPWR.n1515 VPWR.n1164 4.5005
R11820 VPWR.n1518 VPWR.n1517 4.5005
R11821 VPWR.n992 VPWR.n946 4.5005
R11822 VPWR.n1856 VPWR.n1855 4.5005
R11823 VPWR.n899 VPWR.n851 4.5005
R11824 VPWR.n1951 VPWR.n1950 4.5005
R11825 VPWR.n800 VPWR.n754 4.5005
R11826 VPWR.n2052 VPWR.n2051 4.5005
R11827 VPWR.n707 VPWR.n659 4.5005
R11828 VPWR.n2147 VPWR.n2146 4.5005
R11829 VPWR.n608 VPWR.n562 4.5005
R11830 VPWR.n2248 VPWR.n2247 4.5005
R11831 VPWR.n515 VPWR.n467 4.5005
R11832 VPWR.n2343 VPWR.n2342 4.5005
R11833 VPWR.n416 VPWR.n370 4.5005
R11834 VPWR.n2444 VPWR.n2443 4.5005
R11835 VPWR.n2515 VPWR.n2514 4.5005
R11836 VPWR.n343 VPWR.n95 4.5005
R11837 VPWR.n2470 VPWR.n2469 4.5005
R11838 VPWR.n396 VPWR.n359 4.5005
R11839 VPWR.n2317 VPWR.n2316 4.5005
R11840 VPWR.n535 VPWR.n478 4.5005
R11841 VPWR.n2274 VPWR.n2273 4.5005
R11842 VPWR.n588 VPWR.n551 4.5005
R11843 VPWR.n2121 VPWR.n2120 4.5005
R11844 VPWR.n727 VPWR.n670 4.5005
R11845 VPWR.n2078 VPWR.n2077 4.5005
R11846 VPWR.n780 VPWR.n743 4.5005
R11847 VPWR.n1925 VPWR.n1924 4.5005
R11848 VPWR.n919 VPWR.n862 4.5005
R11849 VPWR.n1882 VPWR.n1881 4.5005
R11850 VPWR.n1586 VPWR.n1129 4.5005
R11851 VPWR.n1585 VPWR.n1130 4.5005
R11852 VPWR.n972 VPWR.n935 4.5005
R11853 VPWR.n1526 VPWR.n1155 4.5005
R11854 VPWR.n1525 VPWR.n1523 4.5005
R11855 VPWR.n996 VPWR.n947 4.5005
R11856 VPWR.n1852 VPWR.n1851 4.5005
R11857 VPWR.n895 VPWR.n850 4.5005
R11858 VPWR.n1955 VPWR.n1954 4.5005
R11859 VPWR.n804 VPWR.n755 4.5005
R11860 VPWR.n2048 VPWR.n2047 4.5005
R11861 VPWR.n703 VPWR.n658 4.5005
R11862 VPWR.n2151 VPWR.n2150 4.5005
R11863 VPWR.n612 VPWR.n563 4.5005
R11864 VPWR.n2244 VPWR.n2243 4.5005
R11865 VPWR.n511 VPWR.n466 4.5005
R11866 VPWR.n2347 VPWR.n2346 4.5005
R11867 VPWR.n420 VPWR.n371 4.5005
R11868 VPWR.n2440 VPWR.n2439 4.5005
R11869 VPWR.n2559 VPWR.n2558 4.5005
R11870 VPWR.n315 VPWR.n72 4.5005
R11871 VPWR.n2434 VPWR.n2433 4.5005
R11872 VPWR.n424 VPWR.n374 4.5005
R11873 VPWR.n2353 VPWR.n2352 4.5005
R11874 VPWR.n507 VPWR.n463 4.5005
R11875 VPWR.n2238 VPWR.n2237 4.5005
R11876 VPWR.n616 VPWR.n566 4.5005
R11877 VPWR.n2157 VPWR.n2156 4.5005
R11878 VPWR.n699 VPWR.n655 4.5005
R11879 VPWR.n2042 VPWR.n2041 4.5005
R11880 VPWR.n808 VPWR.n758 4.5005
R11881 VPWR.n1961 VPWR.n1960 4.5005
R11882 VPWR.n891 VPWR.n847 4.5005
R11883 VPWR.n1846 VPWR.n1845 4.5005
R11884 VPWR.n1145 VPWR.n1144 4.5005
R11885 VPWR.n1539 VPWR.n1538 4.5005
R11886 VPWR.n1000 VPWR.n950 4.5005
R11887 VPWR.n1590 VPWR.n1589 4.5005
R11888 VPWR.n1473 VPWR.n1128 4.5005
R11889 VPWR.n968 VPWR.n934 4.5005
R11890 VPWR.n1886 VPWR.n1885 4.5005
R11891 VPWR.n923 VPWR.n863 4.5005
R11892 VPWR.n1921 VPWR.n1920 4.5005
R11893 VPWR.n776 VPWR.n742 4.5005
R11894 VPWR.n2082 VPWR.n2081 4.5005
R11895 VPWR.n731 VPWR.n671 4.5005
R11896 VPWR.n2117 VPWR.n2116 4.5005
R11897 VPWR.n584 VPWR.n550 4.5005
R11898 VPWR.n2278 VPWR.n2277 4.5005
R11899 VPWR.n539 VPWR.n479 4.5005
R11900 VPWR.n2313 VPWR.n2312 4.5005
R11901 VPWR.n392 VPWR.n358 4.5005
R11902 VPWR.n2474 VPWR.n2473 4.5005
R11903 VPWR.n347 VPWR.n96 4.5005
R11904 VPWR.n2563 VPWR.n2562 4.5005
R11905 VPWR.n311 VPWR.n71 4.5005
R11906 VPWR.n2430 VPWR.n2429 4.5005
R11907 VPWR.n428 VPWR.n375 4.5005
R11908 VPWR.n2357 VPWR.n2356 4.5005
R11909 VPWR.n503 VPWR.n462 4.5005
R11910 VPWR.n2234 VPWR.n2233 4.5005
R11911 VPWR.n620 VPWR.n567 4.5005
R11912 VPWR.n2161 VPWR.n2160 4.5005
R11913 VPWR.n695 VPWR.n654 4.5005
R11914 VPWR.n2038 VPWR.n2037 4.5005
R11915 VPWR.n812 VPWR.n759 4.5005
R11916 VPWR.n1965 VPWR.n1964 4.5005
R11917 VPWR.n887 VPWR.n846 4.5005
R11918 VPWR.n1842 VPWR.n1841 4.5005
R11919 VPWR.n1004 VPWR.n951 4.5005
R11920 VPWR.n1531 VPWR.n1154 4.5005
R11921 VPWR.n1533 VPWR.n1532 4.5005
R11922 VPWR.n1073 VPWR.n1045 4.5005
R11923 VPWR.n1764 VPWR.n1763 4.5005
R11924 VPWR.n1008 VPWR.n954 4.5005
R11925 VPWR.n1836 VPWR.n1835 4.5005
R11926 VPWR.n883 VPWR.n843 4.5005
R11927 VPWR.n1971 VPWR.n1970 4.5005
R11928 VPWR.n816 VPWR.n762 4.5005
R11929 VPWR.n2032 VPWR.n2031 4.5005
R11930 VPWR.n691 VPWR.n651 4.5005
R11931 VPWR.n2167 VPWR.n2166 4.5005
R11932 VPWR.n624 VPWR.n570 4.5005
R11933 VPWR.n2228 VPWR.n2227 4.5005
R11934 VPWR.n499 VPWR.n459 4.5005
R11935 VPWR.n2363 VPWR.n2362 4.5005
R11936 VPWR.n432 VPWR.n378 4.5005
R11937 VPWR.n2424 VPWR.n2423 4.5005
R11938 VPWR.n307 VPWR.n66 4.5005
R11939 VPWR.n299 VPWR.n60 4.5005
R11940 VPWR.n2414 VPWR.n2413 4.5005
R11941 VPWR.n440 VPWR.n382 4.5005
R11942 VPWR.n2373 VPWR.n2372 4.5005
R11943 VPWR.n491 VPWR.n455 4.5005
R11944 VPWR.n2218 VPWR.n2217 4.5005
R11945 VPWR.n632 VPWR.n574 4.5005
R11946 VPWR.n2177 VPWR.n2176 4.5005
R11947 VPWR.n683 VPWR.n647 4.5005
R11948 VPWR.n2022 VPWR.n2021 4.5005
R11949 VPWR.n824 VPWR.n766 4.5005
R11950 VPWR.n1981 VPWR.n1980 4.5005
R11951 VPWR.n875 VPWR.n839 4.5005
R11952 VPWR.n1826 VPWR.n1825 4.5005
R11953 VPWR.n1016 VPWR.n958 4.5005
R11954 VPWR.n1753 VPWR.n1743 4.5005
R11955 VPWR.n1752 VPWR.n1751 4.5005
R11956 VPWR.n1756 VPWR.n1054 4.5005
R11957 VPWR.n1758 VPWR.n1757 4.5005
R11958 VPWR.n1012 VPWR.n955 4.5005
R11959 VPWR.n1832 VPWR.n1831 4.5005
R11960 VPWR.n879 VPWR.n842 4.5005
R11961 VPWR.n1975 VPWR.n1974 4.5005
R11962 VPWR.n820 VPWR.n763 4.5005
R11963 VPWR.n2028 VPWR.n2027 4.5005
R11964 VPWR.n687 VPWR.n650 4.5005
R11965 VPWR.n2171 VPWR.n2170 4.5005
R11966 VPWR.n628 VPWR.n571 4.5005
R11967 VPWR.n2224 VPWR.n2223 4.5005
R11968 VPWR.n495 VPWR.n458 4.5005
R11969 VPWR.n2367 VPWR.n2366 4.5005
R11970 VPWR.n436 VPWR.n379 4.5005
R11971 VPWR.n2420 VPWR.n2419 4.5005
R11972 VPWR.n303 VPWR.n65 4.5005
R11973 VPWR.n2575 VPWR.n2574 4.5005
R11974 VPWR.n2583 VPWR.n2582 4.5005
R11975 VPWR.n2587 VPWR.n2586 4.5005
R11976 VPWR.n295 VPWR.n59 4.5005
R11977 VPWR.n2410 VPWR.n2409 4.5005
R11978 VPWR.n444 VPWR.n383 4.5005
R11979 VPWR.n2377 VPWR.n2376 4.5005
R11980 VPWR.n487 VPWR.n454 4.5005
R11981 VPWR.n2214 VPWR.n2213 4.5005
R11982 VPWR.n636 VPWR.n575 4.5005
R11983 VPWR.n2181 VPWR.n2180 4.5005
R11984 VPWR.n679 VPWR.n646 4.5005
R11985 VPWR.n2018 VPWR.n2017 4.5005
R11986 VPWR.n828 VPWR.n767 4.5005
R11987 VPWR.n1985 VPWR.n1984 4.5005
R11988 VPWR.n871 VPWR.n838 4.5005
R11989 VPWR.n1822 VPWR.n1821 4.5005
R11990 VPWR.n1020 VPWR.n959 4.5005
R11991 VPWR.n1789 VPWR.n1788 4.5005
R11992 VPWR.n1736 VPWR.n1037 4.5005
R11993 VPWR.n1232 VPWR.n1121 4.5005
R11994 VPWR.n1466 VPWR.n1465 4.5005
R11995 VPWR.n964 VPWR.n931 4.5005
R11996 VPWR.n1892 VPWR.n1891 4.5005
R11997 VPWR.n929 VPWR.n928 4.5005
R11998 VPWR.n1915 VPWR.n1914 4.5005
R11999 VPWR.n772 VPWR.n739 4.5005
R12000 VPWR.n2088 VPWR.n2087 4.5005
R12001 VPWR.n737 VPWR.n736 4.5005
R12002 VPWR.n2111 VPWR.n2110 4.5005
R12003 VPWR.n580 VPWR.n547 4.5005
R12004 VPWR.n2284 VPWR.n2283 4.5005
R12005 VPWR.n545 VPWR.n544 4.5005
R12006 VPWR.n2307 VPWR.n2306 4.5005
R12007 VPWR.n388 VPWR.n355 4.5005
R12008 VPWR.n2480 VPWR.n2479 4.5005
R12009 VPWR.n353 VPWR.n352 4.5005
R12010 VPWR.n2503 VPWR.n2502 4.5005
R12011 VPWR.n2594 VPWR.n2593 4.5005
R12012 VPWR.n292 VPWR.n22 4.5005
R12013 VPWR.n2405 VPWR.n2404 4.5005
R12014 VPWR.n449 VPWR.n448 4.5005
R12015 VPWR.n2382 VPWR.n2381 4.5005
R12016 VPWR.n484 VPWR.n451 4.5005
R12017 VPWR.n2209 VPWR.n2208 4.5005
R12018 VPWR.n641 VPWR.n640 4.5005
R12019 VPWR.n2186 VPWR.n2185 4.5005
R12020 VPWR.n676 VPWR.n643 4.5005
R12021 VPWR.n2013 VPWR.n2012 4.5005
R12022 VPWR.n833 VPWR.n832 4.5005
R12023 VPWR.n1990 VPWR.n1989 4.5005
R12024 VPWR.n868 VPWR.n835 4.5005
R12025 VPWR.n1817 VPWR.n1816 4.5005
R12026 VPWR.n1025 VPWR.n1024 4.5005
R12027 VPWR.n1794 VPWR.n1793 4.5005
R12028 VPWR.n1060 VPWR.n1028 4.5005
R12029 VPWR.n2628 VPWR 4.49965
R12030 VPWR.n19 VPWR.n18 4.20017
R12031 VPWR.n1255 VPWR.n1254 4.20017
R12032 VPWR.n1279 VPWR.n1278 4.20017
R12033 VPWR.n1302 VPWR.n1301 4.20017
R12034 VPWR.n1337 VPWR.n1336 4.20017
R12035 VPWR.n1376 VPWR.n1375 4.20017
R12036 VPWR.n1414 VPWR.n1413 4.20017
R12037 VPWR.n2813 VPWR 4.14027
R12038 VPWR.n2797 VPWR 4.14027
R12039 VPWR.n2778 VPWR 4.14027
R12040 VPWR.n2758 VPWR 4.14027
R12041 VPWR.n2739 VPWR 4.14027
R12042 VPWR.n2703 VPWR 4.14027
R12043 VPWR.n2665 VPWR 4.14027
R12044 VPWR.n55 VPWR.n54 4.0005
R12045 VPWR.n2716 VPWR.n2713 3.76521
R12046 VPWR.n2680 VPWR.n2676 3.76521
R12047 VPWR.n2643 VPWR.n2639 3.76521
R12048 VPWR.n2611 VPWR.n2610 3.76521
R12049 VPWR.n1906 VPWR.n858 3.4105
R12050 VPWR.n1934 VPWR.n1933 3.4105
R12051 VPWR.n1997 VPWR.n747 3.4105
R12052 VPWR.n2069 VPWR.n2068 3.4105
R12053 VPWR.n2102 VPWR.n666 3.4105
R12054 VPWR.n2130 VPWR.n2129 3.4105
R12055 VPWR.n2193 VPWR.n555 3.4105
R12056 VPWR.n2265 VPWR.n2264 3.4105
R12057 VPWR.n2298 VPWR.n474 3.4105
R12058 VPWR.n2326 VPWR.n2325 3.4105
R12059 VPWR.n2389 VPWR.n363 3.4105
R12060 VPWR.n2388 VPWR.n362 3.4105
R12061 VPWR.n2324 VPWR.n2323 3.4105
R12062 VPWR.n2299 VPWR.n475 3.4105
R12063 VPWR.n2267 VPWR.n2266 3.4105
R12064 VPWR.n2192 VPWR.n554 3.4105
R12065 VPWR.n2128 VPWR.n2127 3.4105
R12066 VPWR.n2103 VPWR.n667 3.4105
R12067 VPWR.n2071 VPWR.n2070 3.4105
R12068 VPWR.n1996 VPWR.n746 3.4105
R12069 VPWR.n1932 VPWR.n1931 3.4105
R12070 VPWR.n1907 VPWR.n859 3.4105
R12071 VPWR.n1875 VPWR.n1874 3.4105
R12072 VPWR.n1873 VPWR.n1872 3.4105
R12073 VPWR.n1865 VPWR.n1864 3.4105
R12074 VPWR.n1905 VPWR.n855 3.4105
R12075 VPWR.n1942 VPWR.n1941 3.4105
R12076 VPWR.n1998 VPWR.n750 3.4105
R12077 VPWR.n2061 VPWR.n2060 3.4105
R12078 VPWR.n2101 VPWR.n663 3.4105
R12079 VPWR.n2138 VPWR.n2137 3.4105
R12080 VPWR.n2194 VPWR.n558 3.4105
R12081 VPWR.n2257 VPWR.n2256 3.4105
R12082 VPWR.n2297 VPWR.n471 3.4105
R12083 VPWR.n2334 VPWR.n2333 3.4105
R12084 VPWR.n2390 VPWR.n366 3.4105
R12085 VPWR.n2391 VPWR.n367 3.4105
R12086 VPWR.n2336 VPWR.n2335 3.4105
R12087 VPWR.n2296 VPWR.n470 3.4105
R12088 VPWR.n2255 VPWR.n2254 3.4105
R12089 VPWR.n2195 VPWR.n559 3.4105
R12090 VPWR.n2140 VPWR.n2139 3.4105
R12091 VPWR.n2100 VPWR.n662 3.4105
R12092 VPWR.n2059 VPWR.n2058 3.4105
R12093 VPWR.n1999 VPWR.n751 3.4105
R12094 VPWR.n1944 VPWR.n1943 3.4105
R12095 VPWR.n1904 VPWR.n854 3.4105
R12096 VPWR.n1863 VPWR.n1862 3.4105
R12097 VPWR.n1855 VPWR.n1854 3.4105
R12098 VPWR.n1903 VPWR.n851 3.4105
R12099 VPWR.n1952 VPWR.n1951 3.4105
R12100 VPWR.n2000 VPWR.n754 3.4105
R12101 VPWR.n2051 VPWR.n2050 3.4105
R12102 VPWR.n2099 VPWR.n659 3.4105
R12103 VPWR.n2148 VPWR.n2147 3.4105
R12104 VPWR.n2196 VPWR.n562 3.4105
R12105 VPWR.n2247 VPWR.n2246 3.4105
R12106 VPWR.n2295 VPWR.n467 3.4105
R12107 VPWR.n2344 VPWR.n2343 3.4105
R12108 VPWR.n2392 VPWR.n370 3.4105
R12109 VPWR.n2443 VPWR.n2442 3.4105
R12110 VPWR.n2451 VPWR.n2450 3.4105
R12111 VPWR.n2453 VPWR.n2452 3.4105
R12112 VPWR.n2461 VPWR.n2460 3.4105
R12113 VPWR.n2463 VPWR.n2462 3.4105
R12114 VPWR.n2471 VPWR.n2470 3.4105
R12115 VPWR.n2387 VPWR.n359 3.4105
R12116 VPWR.n2316 VPWR.n2315 3.4105
R12117 VPWR.n2300 VPWR.n478 3.4105
R12118 VPWR.n2275 VPWR.n2274 3.4105
R12119 VPWR.n2191 VPWR.n551 3.4105
R12120 VPWR.n2120 VPWR.n2119 3.4105
R12121 VPWR.n2104 VPWR.n670 3.4105
R12122 VPWR.n2079 VPWR.n2078 3.4105
R12123 VPWR.n1995 VPWR.n743 3.4105
R12124 VPWR.n1924 VPWR.n1923 3.4105
R12125 VPWR.n1908 VPWR.n862 3.4105
R12126 VPWR.n1883 VPWR.n1882 3.4105
R12127 VPWR.n1799 VPWR.n935 3.4105
R12128 VPWR.n1800 VPWR.n938 3.4105
R12129 VPWR.n1801 VPWR.n939 3.4105
R12130 VPWR.n1802 VPWR.n942 3.4105
R12131 VPWR.n1803 VPWR.n943 3.4105
R12132 VPWR.n1804 VPWR.n946 3.4105
R12133 VPWR.n1805 VPWR.n947 3.4105
R12134 VPWR.n1853 VPWR.n1852 3.4105
R12135 VPWR.n1902 VPWR.n850 3.4105
R12136 VPWR.n1954 VPWR.n1953 3.4105
R12137 VPWR.n2001 VPWR.n755 3.4105
R12138 VPWR.n2049 VPWR.n2048 3.4105
R12139 VPWR.n2098 VPWR.n658 3.4105
R12140 VPWR.n2150 VPWR.n2149 3.4105
R12141 VPWR.n2197 VPWR.n563 3.4105
R12142 VPWR.n2245 VPWR.n2244 3.4105
R12143 VPWR.n2294 VPWR.n466 3.4105
R12144 VPWR.n2346 VPWR.n2345 3.4105
R12145 VPWR.n2393 VPWR.n371 3.4105
R12146 VPWR.n2441 VPWR.n2440 3.4105
R12147 VPWR.n2433 VPWR.n2432 3.4105
R12148 VPWR.n2394 VPWR.n374 3.4105
R12149 VPWR.n2354 VPWR.n2353 3.4105
R12150 VPWR.n2293 VPWR.n463 3.4105
R12151 VPWR.n2237 VPWR.n2236 3.4105
R12152 VPWR.n2198 VPWR.n566 3.4105
R12153 VPWR.n2158 VPWR.n2157 3.4105
R12154 VPWR.n2097 VPWR.n655 3.4105
R12155 VPWR.n2041 VPWR.n2040 3.4105
R12156 VPWR.n2002 VPWR.n758 3.4105
R12157 VPWR.n1962 VPWR.n1961 3.4105
R12158 VPWR.n1901 VPWR.n847 3.4105
R12159 VPWR.n1845 VPWR.n1844 3.4105
R12160 VPWR.n1806 VPWR.n950 3.4105
R12161 VPWR.n1798 VPWR.n934 3.4105
R12162 VPWR.n1885 VPWR.n1884 3.4105
R12163 VPWR.n1909 VPWR.n863 3.4105
R12164 VPWR.n1922 VPWR.n1921 3.4105
R12165 VPWR.n1994 VPWR.n742 3.4105
R12166 VPWR.n2081 VPWR.n2080 3.4105
R12167 VPWR.n2105 VPWR.n671 3.4105
R12168 VPWR.n2118 VPWR.n2117 3.4105
R12169 VPWR.n2190 VPWR.n550 3.4105
R12170 VPWR.n2277 VPWR.n2276 3.4105
R12171 VPWR.n2301 VPWR.n479 3.4105
R12172 VPWR.n2314 VPWR.n2313 3.4105
R12173 VPWR.n2386 VPWR.n358 3.4105
R12174 VPWR.n2473 VPWR.n2472 3.4105
R12175 VPWR.n2497 VPWR.n96 3.4105
R12176 VPWR.n2496 VPWR.n95 3.4105
R12177 VPWR.n2495 VPWR.n90 3.4105
R12178 VPWR.n2494 VPWR.n89 3.4105
R12179 VPWR.n2493 VPWR.n84 3.4105
R12180 VPWR.n2492 VPWR.n83 3.4105
R12181 VPWR.n2491 VPWR.n78 3.4105
R12182 VPWR.n2490 VPWR.n77 3.4105
R12183 VPWR.n2489 VPWR.n72 3.4105
R12184 VPWR.n2488 VPWR.n71 3.4105
R12185 VPWR.n2431 VPWR.n2430 3.4105
R12186 VPWR.n2395 VPWR.n375 3.4105
R12187 VPWR.n2356 VPWR.n2355 3.4105
R12188 VPWR.n2292 VPWR.n462 3.4105
R12189 VPWR.n2235 VPWR.n2234 3.4105
R12190 VPWR.n2199 VPWR.n567 3.4105
R12191 VPWR.n2160 VPWR.n2159 3.4105
R12192 VPWR.n2096 VPWR.n654 3.4105
R12193 VPWR.n2039 VPWR.n2038 3.4105
R12194 VPWR.n2003 VPWR.n759 3.4105
R12195 VPWR.n1964 VPWR.n1963 3.4105
R12196 VPWR.n1900 VPWR.n846 3.4105
R12197 VPWR.n1843 VPWR.n1842 3.4105
R12198 VPWR.n1807 VPWR.n951 3.4105
R12199 VPWR.n1532 VPWR.n1143 3.4105
R12200 VPWR.n1540 VPWR.n1539 3.4105
R12201 VPWR.n1525 VPWR.n1524 3.4105
R12202 VPWR.n1517 VPWR.n1516 3.4105
R12203 VPWR.n1511 VPWR.n1510 3.4105
R12204 VPWR.n1503 VPWR.n1502 3.4105
R12205 VPWR.n1497 VPWR.n1496 3.4105
R12206 VPWR.n1489 VPWR.n1132 3.4105
R12207 VPWR.n1585 VPWR.n1584 3.4105
R12208 VPWR.n1452 VPWR.n1128 3.4105
R12209 VPWR.n1765 VPWR.n1764 3.4105
R12210 VPWR.n1808 VPWR.n954 3.4105
R12211 VPWR.n1835 VPWR.n1834 3.4105
R12212 VPWR.n1899 VPWR.n843 3.4105
R12213 VPWR.n1972 VPWR.n1971 3.4105
R12214 VPWR.n2004 VPWR.n762 3.4105
R12215 VPWR.n2031 VPWR.n2030 3.4105
R12216 VPWR.n2095 VPWR.n651 3.4105
R12217 VPWR.n2168 VPWR.n2167 3.4105
R12218 VPWR.n2200 VPWR.n570 3.4105
R12219 VPWR.n2227 VPWR.n2226 3.4105
R12220 VPWR.n2291 VPWR.n459 3.4105
R12221 VPWR.n2364 VPWR.n2363 3.4105
R12222 VPWR.n2396 VPWR.n378 3.4105
R12223 VPWR.n2423 VPWR.n2422 3.4105
R12224 VPWR.n2487 VPWR.n66 3.4105
R12225 VPWR.n2485 VPWR.n60 3.4105
R12226 VPWR.n2413 VPWR.n2412 3.4105
R12227 VPWR.n2398 VPWR.n382 3.4105
R12228 VPWR.n2374 VPWR.n2373 3.4105
R12229 VPWR.n2289 VPWR.n455 3.4105
R12230 VPWR.n2217 VPWR.n2216 3.4105
R12231 VPWR.n2202 VPWR.n574 3.4105
R12232 VPWR.n2178 VPWR.n2177 3.4105
R12233 VPWR.n2093 VPWR.n647 3.4105
R12234 VPWR.n2021 VPWR.n2020 3.4105
R12235 VPWR.n2006 VPWR.n766 3.4105
R12236 VPWR.n1982 VPWR.n1981 3.4105
R12237 VPWR.n1897 VPWR.n839 3.4105
R12238 VPWR.n1825 VPWR.n1824 3.4105
R12239 VPWR.n1810 VPWR.n958 3.4105
R12240 VPWR.n1752 VPWR.n1744 3.4105
R12241 VPWR.n1757 VPWR.n1043 3.4105
R12242 VPWR.n1809 VPWR.n955 3.4105
R12243 VPWR.n1833 VPWR.n1832 3.4105
R12244 VPWR.n1898 VPWR.n842 3.4105
R12245 VPWR.n1974 VPWR.n1973 3.4105
R12246 VPWR.n2005 VPWR.n763 3.4105
R12247 VPWR.n2029 VPWR.n2028 3.4105
R12248 VPWR.n2094 VPWR.n650 3.4105
R12249 VPWR.n2170 VPWR.n2169 3.4105
R12250 VPWR.n2201 VPWR.n571 3.4105
R12251 VPWR.n2225 VPWR.n2224 3.4105
R12252 VPWR.n2290 VPWR.n458 3.4105
R12253 VPWR.n2366 VPWR.n2365 3.4105
R12254 VPWR.n2397 VPWR.n379 3.4105
R12255 VPWR.n2421 VPWR.n2420 3.4105
R12256 VPWR.n2486 VPWR.n65 3.4105
R12257 VPWR.n2484 VPWR.n59 3.4105
R12258 VPWR.n2411 VPWR.n2410 3.4105
R12259 VPWR.n2399 VPWR.n383 3.4105
R12260 VPWR.n2376 VPWR.n2375 3.4105
R12261 VPWR.n2288 VPWR.n454 3.4105
R12262 VPWR.n2215 VPWR.n2214 3.4105
R12263 VPWR.n2203 VPWR.n575 3.4105
R12264 VPWR.n2180 VPWR.n2179 3.4105
R12265 VPWR.n2092 VPWR.n646 3.4105
R12266 VPWR.n2019 VPWR.n2018 3.4105
R12267 VPWR.n2007 VPWR.n767 3.4105
R12268 VPWR.n1984 VPWR.n1983 3.4105
R12269 VPWR.n1896 VPWR.n838 3.4105
R12270 VPWR.n1823 VPWR.n1822 3.4105
R12271 VPWR.n1811 VPWR.n959 3.4105
R12272 VPWR.n1788 VPWR.n1787 3.4105
R12273 VPWR.n1465 VPWR.n1464 3.4105
R12274 VPWR.n1797 VPWR.n931 3.4105
R12275 VPWR.n1893 VPWR.n1892 3.4105
R12276 VPWR.n1910 VPWR.n929 3.4105
R12277 VPWR.n1914 VPWR.n1913 3.4105
R12278 VPWR.n1993 VPWR.n739 3.4105
R12279 VPWR.n2089 VPWR.n2088 3.4105
R12280 VPWR.n2106 VPWR.n737 3.4105
R12281 VPWR.n2110 VPWR.n2109 3.4105
R12282 VPWR.n2189 VPWR.n547 3.4105
R12283 VPWR.n2285 VPWR.n2284 3.4105
R12284 VPWR.n2302 VPWR.n545 3.4105
R12285 VPWR.n2306 VPWR.n2305 3.4105
R12286 VPWR.n2385 VPWR.n355 3.4105
R12287 VPWR.n2481 VPWR.n2480 3.4105
R12288 VPWR.n2498 VPWR.n353 3.4105
R12289 VPWR.n2502 VPWR.n2501 3.4105
R12290 VPWR.n2512 VPWR.n2511 3.4105
R12291 VPWR.n2514 VPWR.n2513 3.4105
R12292 VPWR.n2524 VPWR.n2523 3.4105
R12293 VPWR.n2526 VPWR.n2525 3.4105
R12294 VPWR.n2536 VPWR.n2535 3.4105
R12295 VPWR.n2538 VPWR.n2537 3.4105
R12296 VPWR.n2548 VPWR.n2547 3.4105
R12297 VPWR.n2550 VPWR.n2549 3.4105
R12298 VPWR.n2560 VPWR.n2559 3.4105
R12299 VPWR.n2562 VPWR.n2561 3.4105
R12300 VPWR.n2572 VPWR.n2571 3.4105
R12301 VPWR.n2574 VPWR.n2573 3.4105
R12302 VPWR.n2584 VPWR.n2583 3.4105
R12303 VPWR.n2586 VPWR.n2585 3.4105
R12304 VPWR.n2595 VPWR.n2594 3.4105
R12305 VPWR.n2483 VPWR.n22 3.4105
R12306 VPWR.n2404 VPWR.n2403 3.4105
R12307 VPWR.n2400 VPWR.n449 3.4105
R12308 VPWR.n2383 VPWR.n2382 3.4105
R12309 VPWR.n2287 VPWR.n451 3.4105
R12310 VPWR.n2208 VPWR.n2207 3.4105
R12311 VPWR.n2204 VPWR.n641 3.4105
R12312 VPWR.n2187 VPWR.n2186 3.4105
R12313 VPWR.n2091 VPWR.n643 3.4105
R12314 VPWR.n2012 VPWR.n2011 3.4105
R12315 VPWR.n2008 VPWR.n833 3.4105
R12316 VPWR.n1991 VPWR.n1990 3.4105
R12317 VPWR.n1895 VPWR.n835 3.4105
R12318 VPWR.n1816 VPWR.n1815 3.4105
R12319 VPWR.n1812 VPWR.n1025 3.4105
R12320 VPWR.n1795 VPWR.n1794 3.4105
R12321 VPWR.n1055 VPWR.n1028 3.4105
R12322 VPWR.n1056 VPWR.n1037 3.4105
R12323 VPWR.n1754 VPWR.n1753 3.4105
R12324 VPWR.n1756 VPWR.n1755 3.4105
R12325 VPWR.n1529 VPWR.n1045 3.4105
R12326 VPWR.n1531 VPWR.n1530 3.4105
R12327 VPWR.n1528 VPWR.n1145 3.4105
R12328 VPWR.n1527 VPWR.n1526 3.4105
R12329 VPWR.n1515 VPWR.n1514 3.4105
R12330 VPWR.n1513 VPWR.n1512 3.4105
R12331 VPWR.n1501 VPWR.n1500 3.4105
R12332 VPWR.n1499 VPWR.n1498 3.4105
R12333 VPWR.n1488 VPWR.n1487 3.4105
R12334 VPWR.n1587 VPWR.n1586 3.4105
R12335 VPWR.n1589 VPWR.n1588 3.4105
R12336 VPWR.n1448 VPWR.n1232 3.4105
R12337 VPWR.n1345 VPWR.n1341 3.38874
R12338 VPWR.n1384 VPWR.n1380 3.38874
R12339 VPWR.n1421 VPWR.n1417 3.38874
R12340 VPWR.n28 VPWR.n26 3.36211
R12341 VPWR.n30 VPWR.n28 3.36211
R12342 VPWR.n32 VPWR.n30 3.36211
R12343 VPWR.n34 VPWR.n32 3.36211
R12344 VPWR.n36 VPWR.n34 3.36211
R12345 VPWR.n38 VPWR.n36 3.36211
R12346 VPWR.n40 VPWR.n38 3.36211
R12347 VPWR.n42 VPWR.n40 3.36211
R12348 VPWR.n44 VPWR.n42 3.36211
R12349 VPWR.n46 VPWR.n44 3.36211
R12350 VPWR.n48 VPWR.n46 3.36211
R12351 VPWR.n50 VPWR.n48 3.36211
R12352 VPWR.n52 VPWR.n50 3.36211
R12353 VPWR.n54 VPWR.n52 3.36211
R12354 VPWR.t1744 VPWR.t950 3.35739
R12355 VPWR.t941 VPWR.t1266 3.35739
R12356 VPWR.n2571 VPWR.n66 3.28012
R12357 VPWR.n2511 VPWR.n96 3.28012
R12358 VPWR.n2550 VPWR.n77 3.28012
R12359 VPWR.n2440 VPWR.n77 3.28012
R12360 VPWR.n2547 VPWR.n78 3.28012
R12361 VPWR.n2443 VPWR.n78 3.28012
R12362 VPWR.n2535 VPWR.n84 3.28012
R12363 VPWR.n2453 VPWR.n84 3.28012
R12364 VPWR.n2453 VPWR.n366 3.28012
R12365 VPWR.n2526 VPWR.n89 3.28012
R12366 VPWR.n2460 VPWR.n89 3.28012
R12367 VPWR.n2460 VPWR.n363 3.28012
R12368 VPWR.n1498 VPWR.n1497 3.28012
R12369 VPWR.n1497 VPWR.n939 3.28012
R12370 VPWR.n1872 VPWR.n939 3.28012
R12371 VPWR.n1872 VPWR.n858 3.28012
R12372 VPWR.n1934 VPWR.n858 3.28012
R12373 VPWR.n1934 VPWR.n747 3.28012
R12374 VPWR.n2068 VPWR.n747 3.28012
R12375 VPWR.n2068 VPWR.n666 3.28012
R12376 VPWR.n2130 VPWR.n666 3.28012
R12377 VPWR.n2130 VPWR.n555 3.28012
R12378 VPWR.n2264 VPWR.n555 3.28012
R12379 VPWR.n2264 VPWR.n474 3.28012
R12380 VPWR.n2326 VPWR.n474 3.28012
R12381 VPWR.n2326 VPWR.n363 3.28012
R12382 VPWR.n2523 VPWR.n90 3.28012
R12383 VPWR.n2463 VPWR.n90 3.28012
R12384 VPWR.n2463 VPWR.n362 3.28012
R12385 VPWR.n2323 VPWR.n362 3.28012
R12386 VPWR.n2323 VPWR.n475 3.28012
R12387 VPWR.n2267 VPWR.n475 3.28012
R12388 VPWR.n2267 VPWR.n554 3.28012
R12389 VPWR.n2127 VPWR.n554 3.28012
R12390 VPWR.n2127 VPWR.n667 3.28012
R12391 VPWR.n2071 VPWR.n667 3.28012
R12392 VPWR.n2071 VPWR.n746 3.28012
R12393 VPWR.n1931 VPWR.n746 3.28012
R12394 VPWR.n1931 VPWR.n859 3.28012
R12395 VPWR.n1875 VPWR.n859 3.28012
R12396 VPWR.n1489 VPWR.n1488 3.28012
R12397 VPWR.n1489 VPWR.n938 3.28012
R12398 VPWR.n1875 VPWR.n938 3.28012
R12399 VPWR.n1503 VPWR.n1501 3.28012
R12400 VPWR.n1503 VPWR.n942 3.28012
R12401 VPWR.n1865 VPWR.n942 3.28012
R12402 VPWR.n1865 VPWR.n855 3.28012
R12403 VPWR.n1941 VPWR.n855 3.28012
R12404 VPWR.n1941 VPWR.n750 3.28012
R12405 VPWR.n2061 VPWR.n750 3.28012
R12406 VPWR.n2061 VPWR.n663 3.28012
R12407 VPWR.n2137 VPWR.n663 3.28012
R12408 VPWR.n2137 VPWR.n558 3.28012
R12409 VPWR.n2257 VPWR.n558 3.28012
R12410 VPWR.n2257 VPWR.n471 3.28012
R12411 VPWR.n2333 VPWR.n471 3.28012
R12412 VPWR.n2333 VPWR.n366 3.28012
R12413 VPWR.n2538 VPWR.n83 3.28012
R12414 VPWR.n2450 VPWR.n83 3.28012
R12415 VPWR.n2450 VPWR.n367 3.28012
R12416 VPWR.n2336 VPWR.n367 3.28012
R12417 VPWR.n2336 VPWR.n470 3.28012
R12418 VPWR.n2254 VPWR.n470 3.28012
R12419 VPWR.n2254 VPWR.n559 3.28012
R12420 VPWR.n2140 VPWR.n559 3.28012
R12421 VPWR.n2140 VPWR.n662 3.28012
R12422 VPWR.n2058 VPWR.n662 3.28012
R12423 VPWR.n2058 VPWR.n751 3.28012
R12424 VPWR.n1944 VPWR.n751 3.28012
R12425 VPWR.n1944 VPWR.n854 3.28012
R12426 VPWR.n1862 VPWR.n854 3.28012
R12427 VPWR.n1512 VPWR.n1511 3.28012
R12428 VPWR.n1511 VPWR.n943 3.28012
R12429 VPWR.n1862 VPWR.n943 3.28012
R12430 VPWR.n1517 VPWR.n1515 3.28012
R12431 VPWR.n1517 VPWR.n946 3.28012
R12432 VPWR.n1855 VPWR.n946 3.28012
R12433 VPWR.n1855 VPWR.n851 3.28012
R12434 VPWR.n1951 VPWR.n851 3.28012
R12435 VPWR.n1951 VPWR.n754 3.28012
R12436 VPWR.n2051 VPWR.n754 3.28012
R12437 VPWR.n2051 VPWR.n659 3.28012
R12438 VPWR.n2147 VPWR.n659 3.28012
R12439 VPWR.n2147 VPWR.n562 3.28012
R12440 VPWR.n2247 VPWR.n562 3.28012
R12441 VPWR.n2247 VPWR.n467 3.28012
R12442 VPWR.n2343 VPWR.n467 3.28012
R12443 VPWR.n2343 VPWR.n370 3.28012
R12444 VPWR.n2443 VPWR.n370 3.28012
R12445 VPWR.n2514 VPWR.n95 3.28012
R12446 VPWR.n2470 VPWR.n95 3.28012
R12447 VPWR.n2470 VPWR.n359 3.28012
R12448 VPWR.n2316 VPWR.n359 3.28012
R12449 VPWR.n2316 VPWR.n478 3.28012
R12450 VPWR.n2274 VPWR.n478 3.28012
R12451 VPWR.n2274 VPWR.n551 3.28012
R12452 VPWR.n2120 VPWR.n551 3.28012
R12453 VPWR.n2120 VPWR.n670 3.28012
R12454 VPWR.n2078 VPWR.n670 3.28012
R12455 VPWR.n2078 VPWR.n743 3.28012
R12456 VPWR.n1924 VPWR.n743 3.28012
R12457 VPWR.n1924 VPWR.n862 3.28012
R12458 VPWR.n1882 VPWR.n862 3.28012
R12459 VPWR.n1882 VPWR.n935 3.28012
R12460 VPWR.n1586 VPWR.n1585 3.28012
R12461 VPWR.n1585 VPWR.n935 3.28012
R12462 VPWR.n1526 VPWR.n1525 3.28012
R12463 VPWR.n1525 VPWR.n947 3.28012
R12464 VPWR.n1852 VPWR.n947 3.28012
R12465 VPWR.n1852 VPWR.n850 3.28012
R12466 VPWR.n1954 VPWR.n850 3.28012
R12467 VPWR.n1954 VPWR.n755 3.28012
R12468 VPWR.n2048 VPWR.n755 3.28012
R12469 VPWR.n2048 VPWR.n658 3.28012
R12470 VPWR.n2150 VPWR.n658 3.28012
R12471 VPWR.n2150 VPWR.n563 3.28012
R12472 VPWR.n2244 VPWR.n563 3.28012
R12473 VPWR.n2244 VPWR.n466 3.28012
R12474 VPWR.n2346 VPWR.n466 3.28012
R12475 VPWR.n2346 VPWR.n371 3.28012
R12476 VPWR.n2440 VPWR.n371 3.28012
R12477 VPWR.n2559 VPWR.n72 3.28012
R12478 VPWR.n2433 VPWR.n72 3.28012
R12479 VPWR.n2433 VPWR.n374 3.28012
R12480 VPWR.n2353 VPWR.n374 3.28012
R12481 VPWR.n2353 VPWR.n463 3.28012
R12482 VPWR.n2237 VPWR.n463 3.28012
R12483 VPWR.n2237 VPWR.n566 3.28012
R12484 VPWR.n2157 VPWR.n566 3.28012
R12485 VPWR.n2157 VPWR.n655 3.28012
R12486 VPWR.n2041 VPWR.n655 3.28012
R12487 VPWR.n2041 VPWR.n758 3.28012
R12488 VPWR.n1961 VPWR.n758 3.28012
R12489 VPWR.n1961 VPWR.n847 3.28012
R12490 VPWR.n1845 VPWR.n847 3.28012
R12491 VPWR.n1845 VPWR.n950 3.28012
R12492 VPWR.n1539 VPWR.n1145 3.28012
R12493 VPWR.n1539 VPWR.n950 3.28012
R12494 VPWR.n1589 VPWR.n1128 3.28012
R12495 VPWR.n1128 VPWR.n934 3.28012
R12496 VPWR.n1885 VPWR.n934 3.28012
R12497 VPWR.n1885 VPWR.n863 3.28012
R12498 VPWR.n1921 VPWR.n863 3.28012
R12499 VPWR.n1921 VPWR.n742 3.28012
R12500 VPWR.n2081 VPWR.n742 3.28012
R12501 VPWR.n2081 VPWR.n671 3.28012
R12502 VPWR.n2117 VPWR.n671 3.28012
R12503 VPWR.n2117 VPWR.n550 3.28012
R12504 VPWR.n2277 VPWR.n550 3.28012
R12505 VPWR.n2277 VPWR.n479 3.28012
R12506 VPWR.n2313 VPWR.n479 3.28012
R12507 VPWR.n2313 VPWR.n358 3.28012
R12508 VPWR.n2473 VPWR.n358 3.28012
R12509 VPWR.n2473 VPWR.n96 3.28012
R12510 VPWR.n2562 VPWR.n71 3.28012
R12511 VPWR.n2430 VPWR.n71 3.28012
R12512 VPWR.n2430 VPWR.n375 3.28012
R12513 VPWR.n2356 VPWR.n375 3.28012
R12514 VPWR.n2356 VPWR.n462 3.28012
R12515 VPWR.n2234 VPWR.n462 3.28012
R12516 VPWR.n2234 VPWR.n567 3.28012
R12517 VPWR.n2160 VPWR.n567 3.28012
R12518 VPWR.n2160 VPWR.n654 3.28012
R12519 VPWR.n2038 VPWR.n654 3.28012
R12520 VPWR.n2038 VPWR.n759 3.28012
R12521 VPWR.n1964 VPWR.n759 3.28012
R12522 VPWR.n1964 VPWR.n846 3.28012
R12523 VPWR.n1842 VPWR.n846 3.28012
R12524 VPWR.n1842 VPWR.n951 3.28012
R12525 VPWR.n1532 VPWR.n951 3.28012
R12526 VPWR.n1532 VPWR.n1531 3.28012
R12527 VPWR.n1764 VPWR.n1045 3.28012
R12528 VPWR.n1764 VPWR.n954 3.28012
R12529 VPWR.n1835 VPWR.n954 3.28012
R12530 VPWR.n1835 VPWR.n843 3.28012
R12531 VPWR.n1971 VPWR.n843 3.28012
R12532 VPWR.n1971 VPWR.n762 3.28012
R12533 VPWR.n2031 VPWR.n762 3.28012
R12534 VPWR.n2031 VPWR.n651 3.28012
R12535 VPWR.n2167 VPWR.n651 3.28012
R12536 VPWR.n2167 VPWR.n570 3.28012
R12537 VPWR.n2227 VPWR.n570 3.28012
R12538 VPWR.n2227 VPWR.n459 3.28012
R12539 VPWR.n2363 VPWR.n459 3.28012
R12540 VPWR.n2363 VPWR.n378 3.28012
R12541 VPWR.n2423 VPWR.n378 3.28012
R12542 VPWR.n2423 VPWR.n66 3.28012
R12543 VPWR.n2583 VPWR.n60 3.28012
R12544 VPWR.n2413 VPWR.n60 3.28012
R12545 VPWR.n2413 VPWR.n382 3.28012
R12546 VPWR.n2373 VPWR.n382 3.28012
R12547 VPWR.n2373 VPWR.n455 3.28012
R12548 VPWR.n2217 VPWR.n455 3.28012
R12549 VPWR.n2217 VPWR.n574 3.28012
R12550 VPWR.n2177 VPWR.n574 3.28012
R12551 VPWR.n2177 VPWR.n647 3.28012
R12552 VPWR.n2021 VPWR.n647 3.28012
R12553 VPWR.n2021 VPWR.n766 3.28012
R12554 VPWR.n1981 VPWR.n766 3.28012
R12555 VPWR.n1981 VPWR.n839 3.28012
R12556 VPWR.n1825 VPWR.n839 3.28012
R12557 VPWR.n1825 VPWR.n958 3.28012
R12558 VPWR.n1752 VPWR.n958 3.28012
R12559 VPWR.n1753 VPWR.n1752 3.28012
R12560 VPWR.n1757 VPWR.n1756 3.28012
R12561 VPWR.n1757 VPWR.n955 3.28012
R12562 VPWR.n1832 VPWR.n955 3.28012
R12563 VPWR.n1832 VPWR.n842 3.28012
R12564 VPWR.n1974 VPWR.n842 3.28012
R12565 VPWR.n1974 VPWR.n763 3.28012
R12566 VPWR.n2028 VPWR.n763 3.28012
R12567 VPWR.n2028 VPWR.n650 3.28012
R12568 VPWR.n2170 VPWR.n650 3.28012
R12569 VPWR.n2170 VPWR.n571 3.28012
R12570 VPWR.n2224 VPWR.n571 3.28012
R12571 VPWR.n2224 VPWR.n458 3.28012
R12572 VPWR.n2366 VPWR.n458 3.28012
R12573 VPWR.n2366 VPWR.n379 3.28012
R12574 VPWR.n2420 VPWR.n379 3.28012
R12575 VPWR.n2420 VPWR.n65 3.28012
R12576 VPWR.n2574 VPWR.n65 3.28012
R12577 VPWR.n2586 VPWR.n59 3.28012
R12578 VPWR.n2410 VPWR.n59 3.28012
R12579 VPWR.n2410 VPWR.n383 3.28012
R12580 VPWR.n2376 VPWR.n383 3.28012
R12581 VPWR.n2376 VPWR.n454 3.28012
R12582 VPWR.n2214 VPWR.n454 3.28012
R12583 VPWR.n2214 VPWR.n575 3.28012
R12584 VPWR.n2180 VPWR.n575 3.28012
R12585 VPWR.n2180 VPWR.n646 3.28012
R12586 VPWR.n2018 VPWR.n646 3.28012
R12587 VPWR.n2018 VPWR.n767 3.28012
R12588 VPWR.n1984 VPWR.n767 3.28012
R12589 VPWR.n1984 VPWR.n838 3.28012
R12590 VPWR.n1822 VPWR.n838 3.28012
R12591 VPWR.n1822 VPWR.n959 3.28012
R12592 VPWR.n1788 VPWR.n959 3.28012
R12593 VPWR.n1788 VPWR.n1037 3.28012
R12594 VPWR.n1465 VPWR.n1232 3.28012
R12595 VPWR.n1465 VPWR.n931 3.28012
R12596 VPWR.n1892 VPWR.n931 3.28012
R12597 VPWR.n1892 VPWR.n929 3.28012
R12598 VPWR.n1914 VPWR.n929 3.28012
R12599 VPWR.n1914 VPWR.n739 3.28012
R12600 VPWR.n2088 VPWR.n739 3.28012
R12601 VPWR.n2088 VPWR.n737 3.28012
R12602 VPWR.n2110 VPWR.n737 3.28012
R12603 VPWR.n2110 VPWR.n547 3.28012
R12604 VPWR.n2284 VPWR.n547 3.28012
R12605 VPWR.n2284 VPWR.n545 3.28012
R12606 VPWR.n2306 VPWR.n545 3.28012
R12607 VPWR.n2306 VPWR.n355 3.28012
R12608 VPWR.n2480 VPWR.n355 3.28012
R12609 VPWR.n2480 VPWR.n353 3.28012
R12610 VPWR.n2502 VPWR.n353 3.28012
R12611 VPWR.n2404 VPWR.n22 3.28012
R12612 VPWR.n2404 VPWR.n449 3.28012
R12613 VPWR.n2382 VPWR.n449 3.28012
R12614 VPWR.n2382 VPWR.n451 3.28012
R12615 VPWR.n2208 VPWR.n451 3.28012
R12616 VPWR.n2208 VPWR.n641 3.28012
R12617 VPWR.n2186 VPWR.n641 3.28012
R12618 VPWR.n2186 VPWR.n643 3.28012
R12619 VPWR.n2012 VPWR.n643 3.28012
R12620 VPWR.n2012 VPWR.n833 3.28012
R12621 VPWR.n1990 VPWR.n833 3.28012
R12622 VPWR.n1990 VPWR.n835 3.28012
R12623 VPWR.n1816 VPWR.n835 3.28012
R12624 VPWR.n1816 VPWR.n1025 3.28012
R12625 VPWR.n1794 VPWR.n1025 3.28012
R12626 VPWR.n1794 VPWR.n1028 3.28012
R12627 VPWR.n2594 VPWR.n22 3.26393
R12628 VPWR.n2832 VPWR.n2831 3.1005
R12629 VPWR.n2826 VPWR.n2825 3.1005
R12630 VPWR.n2846 VPWR.n2815 3.1005
R12631 VPWR.n1324 VPWR.n1322 3.01226
R12632 VPWR.n2863 VPWR 2.83761
R12633 VPWR.n1328 VPWR.n1304 2.63579
R12634 VPWR.n2731 VPWR.n2730 2.25932
R12635 VPWR.n1447 VPWR.n1446 2.01514
R12636 VPWR.n1447 VPWR.n1026 1.65255
R12637 VPWR.n2384 VPWR.n2383 1.32852
R12638 VPWR.n2287 VPWR.n450 1.32852
R12639 VPWR.n2207 VPWR.n2206 1.32852
R12640 VPWR.n2205 VPWR.n2204 1.32852
R12641 VPWR.n2188 VPWR.n2187 1.32852
R12642 VPWR.n2091 VPWR.n642 1.32852
R12643 VPWR.n2011 VPWR.n2010 1.32852
R12644 VPWR.n2009 VPWR.n2008 1.32852
R12645 VPWR.n1992 VPWR.n1991 1.32852
R12646 VPWR.n1895 VPWR.n834 1.32852
R12647 VPWR.n2401 VPWR.n2400 1.32852
R12648 VPWR.n1815 VPWR.n1814 1.32852
R12649 VPWR.n2403 VPWR.n2402 1.32852
R12650 VPWR.n1813 VPWR.n1812 1.32852
R12651 VPWR.n2483 VPWR.n21 1.32852
R12652 VPWR.n1796 VPWR.n1795 1.32852
R12653 VPWR.n2596 VPWR.n2595 1.32852
R12654 VPWR.n1055 VPWR.n1026 1.32852
R12655 VPWR.n2482 VPWR 1.25994
R12656 VPWR VPWR.n354 1.25994
R12657 VPWR VPWR.n2304 1.25994
R12658 VPWR.n2303 VPWR 1.25994
R12659 VPWR.n2286 VPWR 1.25994
R12660 VPWR VPWR.n546 1.25994
R12661 VPWR VPWR.n2108 1.25994
R12662 VPWR.n2107 VPWR 1.25994
R12663 VPWR.n2090 VPWR 1.25994
R12664 VPWR VPWR.n738 1.25994
R12665 VPWR VPWR.n1912 1.25994
R12666 VPWR.n1911 VPWR 1.25994
R12667 VPWR.n1894 VPWR 1.25994
R12668 VPWR VPWR.n930 1.25994
R12669 VPWR.n2499 VPWR 1.25994
R12670 VPWR VPWR.n1450 1.25994
R12671 VPWR VPWR.n2500 1.25994
R12672 VPWR.n1449 VPWR 1.25994
R12673 VPWR.n2597 VPWR.n2596 1.144
R12674 VPWR.n2861 VPWR.n2860 0.936724
R12675 VPWR.n2592 VPWR 0.925943
R12676 VPWR VPWR.n1063 0.925943
R12677 VPWR.n2860 VPWR.n2816 0.925245
R12678 VPWR.n2569 VPWR.n67 0.904391
R12679 VPWR.n2509 VPWR.n97 0.904391
R12680 VPWR.n2552 VPWR.n76 0.904391
R12681 VPWR.n2545 VPWR.n79 0.904391
R12682 VPWR.n2533 VPWR.n85 0.904391
R12683 VPWR.n2528 VPWR.n88 0.904391
R12684 VPWR.n1222 VPWR.n1178 0.904391
R12685 VPWR.n2521 VPWR.n91 0.904391
R12686 VPWR.n1624 VPWR.n1102 0.904391
R12687 VPWR.n1640 VPWR.n1094 0.904391
R12688 VPWR.n2540 VPWR.n82 0.904391
R12689 VPWR.n1651 VPWR.n1092 0.904391
R12690 VPWR.n1211 VPWR.n1210 0.904391
R12691 VPWR.n2516 VPWR.n94 0.904391
R12692 VPWR.n1613 VPWR.n1104 0.904391
R12693 VPWR.n1667 VPWR.n1084 0.904391
R12694 VPWR.n2557 VPWR.n73 0.904391
R12695 VPWR.n1678 VPWR.n1082 0.904391
R12696 VPWR.n1591 VPWR.n1127 0.904391
R12697 VPWR.n2564 VPWR.n70 0.904391
R12698 VPWR.n1197 VPWR.n1196 0.904391
R12699 VPWR.n1694 VPWR.n1074 0.904391
R12700 VPWR.n1742 VPWR.n1057 0.904391
R12701 VPWR.n1705 VPWR.n1071 0.904391
R12702 VPWR.n2581 VPWR.n61 0.904391
R12703 VPWR.n2588 VPWR.n58 0.904391
R12704 VPWR.n1737 VPWR.n1735 0.904391
R12705 VPWR.n1597 VPWR.n1596 0.904391
R12706 VPWR.n2504 VPWR.n289 0.904391
R12707 VPWR.n2576 VPWR.n64 0.904391
R12708 VPWR VPWR.n2863 0.812229
R12709 VPWR.n140 VPWR.n64 0.675548
R12710 VPWR.n152 VPWR.n67 0.675548
R12711 VPWR.n164 VPWR.n70 0.675548
R12712 VPWR.n176 VPWR.n73 0.675548
R12713 VPWR.n188 VPWR.n76 0.675548
R12714 VPWR.n200 VPWR.n79 0.675548
R12715 VPWR.n212 VPWR.n82 0.675548
R12716 VPWR.n224 VPWR.n85 0.675548
R12717 VPWR.n236 VPWR.n88 0.675548
R12718 VPWR.n248 VPWR.n91 0.675548
R12719 VPWR.n260 VPWR.n94 0.675548
R12720 VPWR.n272 VPWR.n97 0.675548
R12721 VPWR.n289 VPWR.n288 0.675548
R12722 VPWR.n128 VPWR.n61 0.675548
R12723 VPWR.n117 VPWR.n58 0.675548
R12724 VPWR.n1735 VPWR.n1734 0.675548
R12725 VPWR.n1719 VPWR.n1057 0.675548
R12726 VPWR.n1707 VPWR.n1705 0.675548
R12727 VPWR.n1696 VPWR.n1694 0.675548
R12728 VPWR.n1196 VPWR.n1195 0.675548
R12729 VPWR.n1680 VPWR.n1678 0.675548
R12730 VPWR.n1669 VPWR.n1667 0.675548
R12731 VPWR.n1210 VPWR.n1209 0.675548
R12732 VPWR.n1653 VPWR.n1651 0.675548
R12733 VPWR.n1642 VPWR.n1640 0.675548
R12734 VPWR.n1178 VPWR.n1177 0.675548
R12735 VPWR.n1626 VPWR.n1624 0.675548
R12736 VPWR.n1615 VPWR.n1613 0.675548
R12737 VPWR.n1127 VPWR.n1126 0.675548
R12738 VPWR.n1599 VPWR.n1597 0.675548
R12739 VPWR.n2806 VPWR.n2805 0.672385
R12740 VPWR.n2790 VPWR.n2785 0.672385
R12741 VPWR.n2770 VPWR.n2765 0.672385
R12742 VPWR.n2751 VPWR.n2746 0.672385
R12743 VPWR.n7 VPWR 0.63497
R12744 VPWR.n1242 VPWR 0.63497
R12745 VPWR.n1265 VPWR 0.63497
R12746 VPWR.n1289 VPWR 0.63497
R12747 VPWR.n24 VPWR 0.499542
R12748 VPWR.n2814 VPWR.n2813 0.442692
R12749 VPWR.n1120 VPWR.n1118 0.404056
R12750 VPWR.n144 VPWR.n138 0.404056
R12751 VPWR.n156 VPWR.n150 0.404056
R12752 VPWR.n168 VPWR.n162 0.404056
R12753 VPWR.n180 VPWR.n174 0.404056
R12754 VPWR.n192 VPWR.n186 0.404056
R12755 VPWR.n204 VPWR.n198 0.404056
R12756 VPWR.n216 VPWR.n210 0.404056
R12757 VPWR.n228 VPWR.n222 0.404056
R12758 VPWR.n240 VPWR.n234 0.404056
R12759 VPWR.n252 VPWR.n246 0.404056
R12760 VPWR.n264 VPWR.n258 0.404056
R12761 VPWR.n276 VPWR.n270 0.404056
R12762 VPWR.n283 VPWR.n101 0.404056
R12763 VPWR.n110 VPWR.n105 0.404056
R12764 VPWR.n132 VPWR.n126 0.404056
R12765 VPWR.n121 VPWR.n115 0.404056
R12766 VPWR.n1729 VPWR.n1065 0.404056
R12767 VPWR.n1723 VPWR.n1717 0.404056
R12768 VPWR.n1711 VPWR.n1070 0.404056
R12769 VPWR.n1704 VPWR.n1702 0.404056
R12770 VPWR.n1693 VPWR.n1691 0.404056
R12771 VPWR.n1684 VPWR.n1081 0.404056
R12772 VPWR.n1677 VPWR.n1675 0.404056
R12773 VPWR.n1666 VPWR.n1664 0.404056
R12774 VPWR.n1657 VPWR.n1091 0.404056
R12775 VPWR.n1650 VPWR.n1648 0.404056
R12776 VPWR.n1639 VPWR.n1637 0.404056
R12777 VPWR.n1630 VPWR.n1101 0.404056
R12778 VPWR.n1623 VPWR.n1621 0.404056
R12779 VPWR.n1612 VPWR.n1610 0.404056
R12780 VPWR.n1603 VPWR.n1111 0.404056
R12781 VPWR.n2860 VPWR.n2859 0.388
R12782 VPWR.n1608 VPWR.n1607 0.349144
R12783 VPWR.n1608 VPWR.n1099 0.349144
R12784 VPWR.n1634 VPWR.n1099 0.349144
R12785 VPWR.n1635 VPWR.n1634 0.349144
R12786 VPWR.n1635 VPWR.n1089 0.349144
R12787 VPWR.n1661 VPWR.n1089 0.349144
R12788 VPWR.n1662 VPWR.n1661 0.349144
R12789 VPWR.n1662 VPWR.n1079 0.349144
R12790 VPWR.n1688 VPWR.n1079 0.349144
R12791 VPWR.n1689 VPWR.n1688 0.349144
R12792 VPWR.n1689 VPWR.n1068 0.349144
R12793 VPWR.n1715 VPWR.n1068 0.349144
R12794 VPWR.n1727 VPWR.n1715 0.349144
R12795 VPWR.n281 VPWR.n280 0.349144
R12796 VPWR.n280 VPWR.n268 0.349144
R12797 VPWR.n268 VPWR.n256 0.349144
R12798 VPWR.n256 VPWR.n244 0.349144
R12799 VPWR.n244 VPWR.n232 0.349144
R12800 VPWR.n232 VPWR.n220 0.349144
R12801 VPWR.n220 VPWR.n208 0.349144
R12802 VPWR.n208 VPWR.n196 0.349144
R12803 VPWR.n196 VPWR.n184 0.349144
R12804 VPWR.n184 VPWR.n172 0.349144
R12805 VPWR.n172 VPWR.n160 0.349144
R12806 VPWR.n160 VPWR.n148 0.349144
R12807 VPWR.n148 VPWR.n136 0.349144
R12808 VPWR.n1462 VPWR.n1456 0.346131
R12809 VPWR.n1461 VPWR.n1457 0.346131
R12810 VPWR.n1582 VPWR.n1136 0.346131
R12811 VPWR.n1581 VPWR.n1577 0.346131
R12812 VPWR.n1576 VPWR.n1572 0.346131
R12813 VPWR.n1571 VPWR.n1567 0.346131
R12814 VPWR.n1566 VPWR.n1562 0.346131
R12815 VPWR.n1561 VPWR.n1557 0.346131
R12816 VPWR.n1556 VPWR.n1552 0.346131
R12817 VPWR.n1551 VPWR.n1547 0.346131
R12818 VPWR.n1546 VPWR.n1542 0.346131
R12819 VPWR.n1767 VPWR.n1042 0.346131
R12820 VPWR.n1784 VPWR.n1780 0.346131
R12821 VPWR.n1785 VPWR.n1776 0.346131
R12822 VPWR.n1772 VPWR.n1771 0.346131
R12823 VPWR.n2862 VPWR.n2861 0.304571
R12824 VPWR.n2594 VPWR.n55 0.300179
R12825 VPWR.n1118 VPWR.n1113 0.286958
R12826 VPWR.n145 VPWR.n144 0.286958
R12827 VPWR.n157 VPWR.n156 0.286958
R12828 VPWR.n169 VPWR.n168 0.286958
R12829 VPWR.n181 VPWR.n180 0.286958
R12830 VPWR.n193 VPWR.n192 0.286958
R12831 VPWR.n205 VPWR.n204 0.286958
R12832 VPWR.n217 VPWR.n216 0.286958
R12833 VPWR.n229 VPWR.n228 0.286958
R12834 VPWR.n241 VPWR.n240 0.286958
R12835 VPWR.n253 VPWR.n252 0.286958
R12836 VPWR.n265 VPWR.n264 0.286958
R12837 VPWR.n277 VPWR.n276 0.286958
R12838 VPWR.n283 VPWR.n102 0.286958
R12839 VPWR.n111 VPWR.n110 0.286958
R12840 VPWR.n133 VPWR.n132 0.286958
R12841 VPWR.n122 VPWR.n121 0.286958
R12842 VPWR.n1729 VPWR.n1066 0.286958
R12843 VPWR.n1724 VPWR.n1723 0.286958
R12844 VPWR.n1712 VPWR.n1711 0.286958
R12845 VPWR.n1702 VPWR.n1072 0.286958
R12846 VPWR.n1691 VPWR.n1075 0.286958
R12847 VPWR.n1685 VPWR.n1684 0.286958
R12848 VPWR.n1675 VPWR.n1083 0.286958
R12849 VPWR.n1664 VPWR.n1085 0.286958
R12850 VPWR.n1658 VPWR.n1657 0.286958
R12851 VPWR.n1648 VPWR.n1093 0.286958
R12852 VPWR.n1637 VPWR.n1095 0.286958
R12853 VPWR.n1631 VPWR.n1630 0.286958
R12854 VPWR.n1621 VPWR.n1103 0.286958
R12855 VPWR.n1610 VPWR.n1105 0.286958
R12856 VPWR.n1604 VPWR.n1603 0.286958
R12857 VPWR.n55 VPWR 0.2505
R12858 VPWR VPWR.n2481 0.249238
R12859 VPWR.n2472 VPWR 0.249238
R12860 VPWR VPWR.n2471 0.249238
R12861 VPWR.n2385 VPWR 0.249238
R12862 VPWR.n2386 VPWR 0.249238
R12863 VPWR.n2387 VPWR 0.249238
R12864 VPWR.n2388 VPWR 0.249238
R12865 VPWR.n2305 VPWR 0.249238
R12866 VPWR.n2314 VPWR 0.249238
R12867 VPWR.n2315 VPWR 0.249238
R12868 VPWR.n2324 VPWR 0.249238
R12869 VPWR.n2325 VPWR 0.249238
R12870 VPWR.n2383 VPWR 0.249238
R12871 VPWR.n2375 VPWR 0.249238
R12872 VPWR.n2374 VPWR 0.249238
R12873 VPWR.n2365 VPWR 0.249238
R12874 VPWR.n2364 VPWR 0.249238
R12875 VPWR.n2355 VPWR 0.249238
R12876 VPWR.n2354 VPWR 0.249238
R12877 VPWR.n2345 VPWR 0.249238
R12878 VPWR.n2344 VPWR 0.249238
R12879 VPWR.n2335 VPWR 0.249238
R12880 VPWR.n2334 VPWR 0.249238
R12881 VPWR VPWR.n2302 0.249238
R12882 VPWR VPWR.n2301 0.249238
R12883 VPWR VPWR.n2300 0.249238
R12884 VPWR VPWR.n2299 0.249238
R12885 VPWR VPWR.n2298 0.249238
R12886 VPWR VPWR.n2287 0.249238
R12887 VPWR VPWR.n2288 0.249238
R12888 VPWR VPWR.n2289 0.249238
R12889 VPWR VPWR.n2290 0.249238
R12890 VPWR VPWR.n2291 0.249238
R12891 VPWR VPWR.n2292 0.249238
R12892 VPWR VPWR.n2293 0.249238
R12893 VPWR VPWR.n2294 0.249238
R12894 VPWR VPWR.n2295 0.249238
R12895 VPWR VPWR.n2296 0.249238
R12896 VPWR VPWR.n2297 0.249238
R12897 VPWR VPWR.n2285 0.249238
R12898 VPWR.n2276 VPWR 0.249238
R12899 VPWR VPWR.n2275 0.249238
R12900 VPWR.n2266 VPWR 0.249238
R12901 VPWR VPWR.n2265 0.249238
R12902 VPWR.n2207 VPWR 0.249238
R12903 VPWR VPWR.n2215 0.249238
R12904 VPWR.n2216 VPWR 0.249238
R12905 VPWR VPWR.n2225 0.249238
R12906 VPWR.n2226 VPWR 0.249238
R12907 VPWR VPWR.n2235 0.249238
R12908 VPWR.n2236 VPWR 0.249238
R12909 VPWR VPWR.n2245 0.249238
R12910 VPWR.n2246 VPWR 0.249238
R12911 VPWR VPWR.n2255 0.249238
R12912 VPWR.n2256 VPWR 0.249238
R12913 VPWR.n2189 VPWR 0.249238
R12914 VPWR.n2190 VPWR 0.249238
R12915 VPWR.n2191 VPWR 0.249238
R12916 VPWR.n2192 VPWR 0.249238
R12917 VPWR.n2193 VPWR 0.249238
R12918 VPWR.n2204 VPWR 0.249238
R12919 VPWR.n2203 VPWR 0.249238
R12920 VPWR.n2202 VPWR 0.249238
R12921 VPWR.n2201 VPWR 0.249238
R12922 VPWR.n2200 VPWR 0.249238
R12923 VPWR.n2199 VPWR 0.249238
R12924 VPWR.n2198 VPWR 0.249238
R12925 VPWR.n2197 VPWR 0.249238
R12926 VPWR.n2196 VPWR 0.249238
R12927 VPWR.n2195 VPWR 0.249238
R12928 VPWR.n2194 VPWR 0.249238
R12929 VPWR.n2109 VPWR 0.249238
R12930 VPWR.n2118 VPWR 0.249238
R12931 VPWR.n2119 VPWR 0.249238
R12932 VPWR.n2128 VPWR 0.249238
R12933 VPWR.n2129 VPWR 0.249238
R12934 VPWR.n2187 VPWR 0.249238
R12935 VPWR.n2179 VPWR 0.249238
R12936 VPWR.n2178 VPWR 0.249238
R12937 VPWR.n2169 VPWR 0.249238
R12938 VPWR.n2168 VPWR 0.249238
R12939 VPWR.n2159 VPWR 0.249238
R12940 VPWR.n2158 VPWR 0.249238
R12941 VPWR.n2149 VPWR 0.249238
R12942 VPWR.n2148 VPWR 0.249238
R12943 VPWR.n2139 VPWR 0.249238
R12944 VPWR.n2138 VPWR 0.249238
R12945 VPWR VPWR.n2106 0.249238
R12946 VPWR VPWR.n2105 0.249238
R12947 VPWR VPWR.n2104 0.249238
R12948 VPWR VPWR.n2103 0.249238
R12949 VPWR VPWR.n2102 0.249238
R12950 VPWR VPWR.n2091 0.249238
R12951 VPWR VPWR.n2092 0.249238
R12952 VPWR VPWR.n2093 0.249238
R12953 VPWR VPWR.n2094 0.249238
R12954 VPWR VPWR.n2095 0.249238
R12955 VPWR VPWR.n2096 0.249238
R12956 VPWR VPWR.n2097 0.249238
R12957 VPWR VPWR.n2098 0.249238
R12958 VPWR VPWR.n2099 0.249238
R12959 VPWR VPWR.n2100 0.249238
R12960 VPWR VPWR.n2101 0.249238
R12961 VPWR VPWR.n2089 0.249238
R12962 VPWR.n2080 VPWR 0.249238
R12963 VPWR VPWR.n2079 0.249238
R12964 VPWR.n2070 VPWR 0.249238
R12965 VPWR VPWR.n2069 0.249238
R12966 VPWR.n2011 VPWR 0.249238
R12967 VPWR VPWR.n2019 0.249238
R12968 VPWR.n2020 VPWR 0.249238
R12969 VPWR VPWR.n2029 0.249238
R12970 VPWR.n2030 VPWR 0.249238
R12971 VPWR VPWR.n2039 0.249238
R12972 VPWR.n2040 VPWR 0.249238
R12973 VPWR VPWR.n2049 0.249238
R12974 VPWR.n2050 VPWR 0.249238
R12975 VPWR VPWR.n2059 0.249238
R12976 VPWR.n2060 VPWR 0.249238
R12977 VPWR.n1993 VPWR 0.249238
R12978 VPWR.n1994 VPWR 0.249238
R12979 VPWR.n1995 VPWR 0.249238
R12980 VPWR.n1996 VPWR 0.249238
R12981 VPWR.n1997 VPWR 0.249238
R12982 VPWR.n2008 VPWR 0.249238
R12983 VPWR.n2007 VPWR 0.249238
R12984 VPWR.n2006 VPWR 0.249238
R12985 VPWR.n2005 VPWR 0.249238
R12986 VPWR.n2004 VPWR 0.249238
R12987 VPWR.n2003 VPWR 0.249238
R12988 VPWR.n2002 VPWR 0.249238
R12989 VPWR.n2001 VPWR 0.249238
R12990 VPWR.n2000 VPWR 0.249238
R12991 VPWR.n1999 VPWR 0.249238
R12992 VPWR.n1998 VPWR 0.249238
R12993 VPWR.n1913 VPWR 0.249238
R12994 VPWR.n1922 VPWR 0.249238
R12995 VPWR.n1923 VPWR 0.249238
R12996 VPWR.n1932 VPWR 0.249238
R12997 VPWR.n1933 VPWR 0.249238
R12998 VPWR.n1991 VPWR 0.249238
R12999 VPWR.n1983 VPWR 0.249238
R13000 VPWR.n1982 VPWR 0.249238
R13001 VPWR.n1973 VPWR 0.249238
R13002 VPWR.n1972 VPWR 0.249238
R13003 VPWR.n1963 VPWR 0.249238
R13004 VPWR.n1962 VPWR 0.249238
R13005 VPWR.n1953 VPWR 0.249238
R13006 VPWR.n1952 VPWR 0.249238
R13007 VPWR.n1943 VPWR 0.249238
R13008 VPWR.n1942 VPWR 0.249238
R13009 VPWR VPWR.n1910 0.249238
R13010 VPWR VPWR.n1909 0.249238
R13011 VPWR VPWR.n1908 0.249238
R13012 VPWR VPWR.n1907 0.249238
R13013 VPWR VPWR.n1906 0.249238
R13014 VPWR VPWR.n1895 0.249238
R13015 VPWR VPWR.n1896 0.249238
R13016 VPWR VPWR.n1897 0.249238
R13017 VPWR VPWR.n1898 0.249238
R13018 VPWR VPWR.n1899 0.249238
R13019 VPWR VPWR.n1900 0.249238
R13020 VPWR VPWR.n1901 0.249238
R13021 VPWR VPWR.n1902 0.249238
R13022 VPWR VPWR.n1903 0.249238
R13023 VPWR VPWR.n1904 0.249238
R13024 VPWR VPWR.n1905 0.249238
R13025 VPWR.n2400 VPWR 0.249238
R13026 VPWR.n2399 VPWR 0.249238
R13027 VPWR.n2398 VPWR 0.249238
R13028 VPWR.n2397 VPWR 0.249238
R13029 VPWR.n2396 VPWR 0.249238
R13030 VPWR.n2395 VPWR 0.249238
R13031 VPWR.n2394 VPWR 0.249238
R13032 VPWR.n2393 VPWR 0.249238
R13033 VPWR.n2392 VPWR 0.249238
R13034 VPWR.n2391 VPWR 0.249238
R13035 VPWR.n2390 VPWR 0.249238
R13036 VPWR.n2389 VPWR 0.249238
R13037 VPWR VPWR.n1893 0.249238
R13038 VPWR.n1884 VPWR 0.249238
R13039 VPWR VPWR.n1883 0.249238
R13040 VPWR.n1874 VPWR 0.249238
R13041 VPWR VPWR.n1873 0.249238
R13042 VPWR.n1864 VPWR 0.249238
R13043 VPWR.n1815 VPWR 0.249238
R13044 VPWR VPWR.n1823 0.249238
R13045 VPWR.n1824 VPWR 0.249238
R13046 VPWR VPWR.n1833 0.249238
R13047 VPWR.n1834 VPWR 0.249238
R13048 VPWR VPWR.n1843 0.249238
R13049 VPWR.n1844 VPWR 0.249238
R13050 VPWR VPWR.n1853 0.249238
R13051 VPWR.n1854 VPWR 0.249238
R13052 VPWR VPWR.n1863 0.249238
R13053 VPWR.n2403 VPWR 0.249238
R13054 VPWR VPWR.n2411 0.249238
R13055 VPWR.n2412 VPWR 0.249238
R13056 VPWR VPWR.n2421 0.249238
R13057 VPWR.n2422 VPWR 0.249238
R13058 VPWR VPWR.n2431 0.249238
R13059 VPWR.n2432 VPWR 0.249238
R13060 VPWR VPWR.n2441 0.249238
R13061 VPWR.n2442 VPWR 0.249238
R13062 VPWR VPWR.n2451 0.249238
R13063 VPWR.n2452 VPWR 0.249238
R13064 VPWR VPWR.n2461 0.249238
R13065 VPWR.n2462 VPWR 0.249238
R13066 VPWR.n1797 VPWR 0.249238
R13067 VPWR.n1798 VPWR 0.249238
R13068 VPWR.n1799 VPWR 0.249238
R13069 VPWR.n1800 VPWR 0.249238
R13070 VPWR.n1801 VPWR 0.249238
R13071 VPWR.n1802 VPWR 0.249238
R13072 VPWR.n1803 VPWR 0.249238
R13073 VPWR.n1804 VPWR 0.249238
R13074 VPWR.n1805 VPWR 0.249238
R13075 VPWR.n1812 VPWR 0.249238
R13076 VPWR.n1811 VPWR 0.249238
R13077 VPWR.n1810 VPWR 0.249238
R13078 VPWR.n1809 VPWR 0.249238
R13079 VPWR.n1808 VPWR 0.249238
R13080 VPWR.n1807 VPWR 0.249238
R13081 VPWR.n1806 VPWR 0.249238
R13082 VPWR VPWR.n2498 0.249238
R13083 VPWR VPWR.n2497 0.249238
R13084 VPWR VPWR.n2496 0.249238
R13085 VPWR VPWR.n2495 0.249238
R13086 VPWR VPWR.n2494 0.249238
R13087 VPWR VPWR.n2493 0.249238
R13088 VPWR VPWR.n2492 0.249238
R13089 VPWR VPWR.n2491 0.249238
R13090 VPWR VPWR.n2490 0.249238
R13091 VPWR VPWR.n2489 0.249238
R13092 VPWR VPWR.n2488 0.249238
R13093 VPWR VPWR.n2483 0.249238
R13094 VPWR VPWR.n2484 0.249238
R13095 VPWR VPWR.n2485 0.249238
R13096 VPWR VPWR.n2486 0.249238
R13097 VPWR VPWR.n2487 0.249238
R13098 VPWR.n2501 VPWR 0.249238
R13099 VPWR.n2512 VPWR 0.249238
R13100 VPWR.n2513 VPWR 0.249238
R13101 VPWR.n2524 VPWR 0.249238
R13102 VPWR.n2525 VPWR 0.249238
R13103 VPWR.n2536 VPWR 0.249238
R13104 VPWR.n2537 VPWR 0.249238
R13105 VPWR.n2548 VPWR 0.249238
R13106 VPWR.n2549 VPWR 0.249238
R13107 VPWR.n2560 VPWR 0.249238
R13108 VPWR.n2561 VPWR 0.249238
R13109 VPWR.n2572 VPWR 0.249238
R13110 VPWR.n2573 VPWR 0.249238
R13111 VPWR.n2584 VPWR 0.249238
R13112 VPWR.n2585 VPWR 0.249238
R13113 VPWR.n2595 VPWR 0.249238
R13114 VPWR VPWR.n1055 0.249238
R13115 VPWR VPWR.n1056 0.249238
R13116 VPWR VPWR.n1754 0.249238
R13117 VPWR.n1755 VPWR 0.249238
R13118 VPWR VPWR.n1529 0.249238
R13119 VPWR.n1530 VPWR 0.249238
R13120 VPWR.n1528 VPWR 0.249238
R13121 VPWR.n1527 VPWR 0.249238
R13122 VPWR.n1514 VPWR 0.249238
R13123 VPWR.n1513 VPWR 0.249238
R13124 VPWR.n1500 VPWR 0.249238
R13125 VPWR.n1499 VPWR 0.249238
R13126 VPWR.n1487 VPWR 0.249238
R13127 VPWR VPWR.n1587 0.249238
R13128 VPWR.n1588 VPWR 0.249238
R13129 VPWR VPWR.n1448 0.249238
R13130 VPWR.n2861 VPWR.n2815 0.245065
R13131 VPWR.n2813 VPWR.n2797 0.213567
R13132 VPWR.n2797 VPWR.n2778 0.213567
R13133 VPWR.n2778 VPWR.n2758 0.213567
R13134 VPWR.n2758 VPWR.n2739 0.213567
R13135 VPWR.n2739 VPWR.n2703 0.213567
R13136 VPWR.n2703 VPWR.n2665 0.213567
R13137 VPWR.n2665 VPWR.n2628 0.213567
R13138 VPWR.n1446 VPWR.n1414 0.213567
R13139 VPWR.n1414 VPWR.n1376 0.213567
R13140 VPWR.n1376 VPWR.n1337 0.213567
R13141 VPWR.n1337 VPWR.n1302 0.213567
R13142 VPWR.n1302 VPWR.n1279 0.213567
R13143 VPWR.n1279 VPWR.n1255 0.213567
R13144 VPWR.n1255 VPWR.n19 0.213567
R13145 VPWR VPWR.n2862 0.204304
R13146 VPWR.n1449 VPWR.n1447 0.182233
R13147 VPWR.n1450 VPWR.n1449 0.154425
R13148 VPWR.n1450 VPWR.n930 0.154425
R13149 VPWR.n1894 VPWR.n930 0.154425
R13150 VPWR.n1911 VPWR.n1894 0.154425
R13151 VPWR.n1912 VPWR.n1911 0.154425
R13152 VPWR.n1912 VPWR.n738 0.154425
R13153 VPWR.n2090 VPWR.n738 0.154425
R13154 VPWR.n2107 VPWR.n2090 0.154425
R13155 VPWR.n2108 VPWR.n2107 0.154425
R13156 VPWR.n2108 VPWR.n546 0.154425
R13157 VPWR.n2286 VPWR.n546 0.154425
R13158 VPWR.n2303 VPWR.n2286 0.154425
R13159 VPWR.n2304 VPWR.n2303 0.154425
R13160 VPWR.n2304 VPWR.n354 0.154425
R13161 VPWR.n2482 VPWR.n354 0.154425
R13162 VPWR.n2499 VPWR.n2482 0.154425
R13163 VPWR.n2500 VPWR.n2499 0.154425
R13164 VPWR.n1796 VPWR.n1026 0.154425
R13165 VPWR.n1813 VPWR.n1796 0.154425
R13166 VPWR.n1814 VPWR.n1813 0.154425
R13167 VPWR.n1814 VPWR.n834 0.154425
R13168 VPWR.n1992 VPWR.n834 0.154425
R13169 VPWR.n2009 VPWR.n1992 0.154425
R13170 VPWR.n2010 VPWR.n2009 0.154425
R13171 VPWR.n2010 VPWR.n642 0.154425
R13172 VPWR.n2188 VPWR.n642 0.154425
R13173 VPWR.n2205 VPWR.n2188 0.154425
R13174 VPWR.n2206 VPWR.n2205 0.154425
R13175 VPWR.n2206 VPWR.n450 0.154425
R13176 VPWR.n2384 VPWR.n450 0.154425
R13177 VPWR.n2401 VPWR.n2384 0.154425
R13178 VPWR.n2402 VPWR.n2401 0.154425
R13179 VPWR.n2402 VPWR.n21 0.154425
R13180 VPWR.n2596 VPWR.n21 0.154425
R13181 VPWR.n8 VPWR.n7 0.147771
R13182 VPWR.n1243 VPWR.n1242 0.147771
R13183 VPWR.n1266 VPWR.n1265 0.147771
R13184 VPWR.n1290 VPWR.n1289 0.147771
R13185 VPWR.n1113 VPWR 0.135917
R13186 VPWR.n145 VPWR 0.135917
R13187 VPWR.n157 VPWR 0.135917
R13188 VPWR.n169 VPWR 0.135917
R13189 VPWR.n181 VPWR 0.135917
R13190 VPWR.n193 VPWR 0.135917
R13191 VPWR.n205 VPWR 0.135917
R13192 VPWR.n217 VPWR 0.135917
R13193 VPWR.n229 VPWR 0.135917
R13194 VPWR.n241 VPWR 0.135917
R13195 VPWR.n253 VPWR 0.135917
R13196 VPWR.n265 VPWR 0.135917
R13197 VPWR.n277 VPWR 0.135917
R13198 VPWR.n102 VPWR 0.135917
R13199 VPWR.n111 VPWR 0.135917
R13200 VPWR.n133 VPWR 0.135917
R13201 VPWR.n122 VPWR 0.135917
R13202 VPWR.n1066 VPWR 0.135917
R13203 VPWR.n1724 VPWR 0.135917
R13204 VPWR.n1712 VPWR 0.135917
R13205 VPWR.n1072 VPWR 0.135917
R13206 VPWR.n1075 VPWR 0.135917
R13207 VPWR.n1685 VPWR 0.135917
R13208 VPWR.n1083 VPWR 0.135917
R13209 VPWR.n1085 VPWR 0.135917
R13210 VPWR.n1658 VPWR 0.135917
R13211 VPWR.n1093 VPWR 0.135917
R13212 VPWR.n1095 VPWR 0.135917
R13213 VPWR.n1631 VPWR 0.135917
R13214 VPWR.n1103 VPWR 0.135917
R13215 VPWR.n1105 VPWR 0.135917
R13216 VPWR.n1604 VPWR 0.135917
R13217 VPWR.n2863 VPWR.n2814 0.127988
R13218 VPWR.n2825 VPWR.n2816 0.1255
R13219 VPWR.n2831 VPWR.n2816 0.1255
R13220 VPWR.n18 VPWR.n0 0.120292
R13221 VPWR.n14 VPWR.n0 0.120292
R13222 VPWR.n9 VPWR.n8 0.120292
R13223 VPWR.n1254 VPWR.n1233 0.120292
R13224 VPWR.n1250 VPWR.n1233 0.120292
R13225 VPWR.n1244 VPWR.n1243 0.120292
R13226 VPWR.n1278 VPWR.n1256 0.120292
R13227 VPWR.n1273 VPWR.n1256 0.120292
R13228 VPWR.n1267 VPWR.n1266 0.120292
R13229 VPWR.n1301 VPWR.n1280 0.120292
R13230 VPWR.n1297 VPWR.n1280 0.120292
R13231 VPWR.n1291 VPWR.n1290 0.120292
R13232 VPWR.n1333 VPWR.n1332 0.120292
R13233 VPWR.n1326 VPWR.n1305 0.120292
R13234 VPWR.n1319 VPWR.n1305 0.120292
R13235 VPWR.n1319 VPWR.n1318 0.120292
R13236 VPWR.n1317 VPWR.n1309 0.120292
R13237 VPWR.n1312 VPWR.n1309 0.120292
R13238 VPWR.n1312 VPWR.n1311 0.120292
R13239 VPWR.n1371 VPWR.n1370 0.120292
R13240 VPWR.n1364 VPWR.n1363 0.120292
R13241 VPWR.n1363 VPWR.n1340 0.120292
R13242 VPWR.n1356 VPWR.n1340 0.120292
R13243 VPWR.n1356 VPWR.n1355 0.120292
R13244 VPWR.n1355 VPWR.n1354 0.120292
R13245 VPWR.n1354 VPWR.n1342 0.120292
R13246 VPWR.n1348 VPWR.n1342 0.120292
R13247 VPWR.n1348 VPWR.n1347 0.120292
R13248 VPWR.n1410 VPWR.n1409 0.120292
R13249 VPWR.n1403 VPWR.n1402 0.120292
R13250 VPWR.n1402 VPWR.n1379 0.120292
R13251 VPWR.n1395 VPWR.n1379 0.120292
R13252 VPWR.n1395 VPWR.n1394 0.120292
R13253 VPWR.n1394 VPWR.n1393 0.120292
R13254 VPWR.n1393 VPWR.n1381 0.120292
R13255 VPWR.n1387 VPWR.n1381 0.120292
R13256 VPWR.n1387 VPWR.n1386 0.120292
R13257 VPWR.n1440 VPWR.n1439 0.120292
R13258 VPWR.n1439 VPWR.n1416 0.120292
R13259 VPWR.n1432 VPWR.n1416 0.120292
R13260 VPWR.n1432 VPWR.n1431 0.120292
R13261 VPWR.n1431 VPWR.n1430 0.120292
R13262 VPWR.n1430 VPWR.n1418 0.120292
R13263 VPWR.n1424 VPWR.n1418 0.120292
R13264 VPWR.n1424 VPWR.n1423 0.120292
R13265 VPWR.n2812 VPWR.n2798 0.120292
R13266 VPWR.n2796 VPWR.n2779 0.120292
R13267 VPWR.n2777 VPWR.n2759 0.120292
R13268 VPWR.n2757 VPWR.n2740 0.120292
R13269 VPWR.n2719 VPWR.n2718 0.120292
R13270 VPWR.n2720 VPWR.n2719 0.120292
R13271 VPWR.n2720 VPWR.n2711 0.120292
R13272 VPWR.n2725 VPWR.n2711 0.120292
R13273 VPWR.n2726 VPWR.n2725 0.120292
R13274 VPWR.n2726 VPWR.n2707 0.120292
R13275 VPWR.n2732 VPWR.n2707 0.120292
R13276 VPWR.n2734 VPWR.n2704 0.120292
R13277 VPWR.n2738 VPWR.n2704 0.120292
R13278 VPWR.n2683 VPWR.n2682 0.120292
R13279 VPWR.n2684 VPWR.n2683 0.120292
R13280 VPWR.n2684 VPWR.n2673 0.120292
R13281 VPWR.n2689 VPWR.n2673 0.120292
R13282 VPWR.n2690 VPWR.n2689 0.120292
R13283 VPWR.n2690 VPWR.n2669 0.120292
R13284 VPWR.n2695 VPWR.n2669 0.120292
R13285 VPWR.n2697 VPWR.n2666 0.120292
R13286 VPWR.n2702 VPWR.n2666 0.120292
R13287 VPWR.n2646 VPWR.n2645 0.120292
R13288 VPWR.n2647 VPWR.n2646 0.120292
R13289 VPWR.n2647 VPWR.n2636 0.120292
R13290 VPWR.n2652 VPWR.n2636 0.120292
R13291 VPWR.n2653 VPWR.n2652 0.120292
R13292 VPWR.n2653 VPWR.n2632 0.120292
R13293 VPWR.n2658 VPWR.n2632 0.120292
R13294 VPWR.n2660 VPWR.n2629 0.120292
R13295 VPWR.n2664 VPWR.n2629 0.120292
R13296 VPWR.n2608 VPWR.n2604 0.120292
R13297 VPWR.n2616 VPWR.n2604 0.120292
R13298 VPWR.n2617 VPWR.n2616 0.120292
R13299 VPWR.n2618 VPWR.n2617 0.120292
R13300 VPWR.n2618 VPWR.n2600 0.120292
R13301 VPWR.n2623 VPWR.n2600 0.120292
R13302 VPWR.n2624 VPWR.n2623 0.120292
R13303 VPWR.n1605 VPWR 0.118556
R13304 VPWR.n1108 VPWR 0.118556
R13305 VPWR.n1619 VPWR 0.118556
R13306 VPWR.n1632 VPWR 0.118556
R13307 VPWR.n1098 VPWR 0.118556
R13308 VPWR.n1646 VPWR 0.118556
R13309 VPWR.n1659 VPWR 0.118556
R13310 VPWR.n1088 VPWR 0.118556
R13311 VPWR.n1673 VPWR 0.118556
R13312 VPWR.n1686 VPWR 0.118556
R13313 VPWR.n1078 VPWR 0.118556
R13314 VPWR.n1700 VPWR 0.118556
R13315 VPWR.n1713 VPWR 0.118556
R13316 VPWR.n1725 VPWR 0.118556
R13317 VPWR VPWR.n1112 0.118556
R13318 VPWR.n1067 VPWR 0.118556
R13319 VPWR.n123 VPWR 0.118556
R13320 VPWR.n112 VPWR 0.118556
R13321 VPWR.n103 VPWR 0.118556
R13322 VPWR.n278 VPWR 0.118556
R13323 VPWR.n266 VPWR 0.118556
R13324 VPWR.n254 VPWR 0.118556
R13325 VPWR.n242 VPWR 0.118556
R13326 VPWR.n230 VPWR 0.118556
R13327 VPWR.n218 VPWR 0.118556
R13328 VPWR.n206 VPWR 0.118556
R13329 VPWR.n194 VPWR 0.118556
R13330 VPWR.n182 VPWR 0.118556
R13331 VPWR.n170 VPWR 0.118556
R13332 VPWR.n158 VPWR 0.118556
R13333 VPWR.n146 VPWR 0.118556
R13334 VPWR.n134 VPWR 0.118556
R13335 VPWR.n1765 VPWR.n1044 0.108238
R13336 VPWR.n1541 VPWR.n1143 0.108238
R13337 VPWR.n1540 VPWR.n1142 0.108238
R13338 VPWR.n1524 VPWR.n1141 0.108238
R13339 VPWR.n1516 VPWR.n1140 0.108238
R13340 VPWR.n1510 VPWR.n1139 0.108238
R13341 VPWR.n1502 VPWR.n1138 0.108238
R13342 VPWR.n1496 VPWR.n1137 0.108238
R13343 VPWR.n1583 VPWR.n1132 0.108238
R13344 VPWR.n1584 VPWR.n1131 0.108238
R13345 VPWR.n1463 VPWR.n1452 0.108238
R13346 VPWR.n1464 VPWR.n1451 0.108238
R13347 VPWR.n1795 VPWR.n1027 0.108238
R13348 VPWR.n1766 VPWR.n1043 0.108238
R13349 VPWR.n1744 VPWR.n1038 0.108238
R13350 VPWR.n1787 VPWR.n1786 0.108238
R13351 VPWR.n2481 VPWR 0.100405
R13352 VPWR.n2472 VPWR 0.100405
R13353 VPWR VPWR.n2385 0.100405
R13354 VPWR VPWR.n2386 0.100405
R13355 VPWR VPWR.n2387 0.100405
R13356 VPWR.n2305 VPWR 0.100405
R13357 VPWR VPWR.n2314 0.100405
R13358 VPWR.n2315 VPWR 0.100405
R13359 VPWR VPWR.n2324 0.100405
R13360 VPWR.n2375 VPWR 0.100405
R13361 VPWR VPWR.n2374 0.100405
R13362 VPWR.n2365 VPWR 0.100405
R13363 VPWR VPWR.n2364 0.100405
R13364 VPWR.n2355 VPWR 0.100405
R13365 VPWR VPWR.n2354 0.100405
R13366 VPWR.n2345 VPWR 0.100405
R13367 VPWR VPWR.n2344 0.100405
R13368 VPWR.n2335 VPWR 0.100405
R13369 VPWR VPWR.n2334 0.100405
R13370 VPWR.n2325 VPWR 0.100405
R13371 VPWR.n2302 VPWR 0.100405
R13372 VPWR.n2301 VPWR 0.100405
R13373 VPWR.n2300 VPWR 0.100405
R13374 VPWR.n2299 VPWR 0.100405
R13375 VPWR.n2288 VPWR 0.100405
R13376 VPWR.n2289 VPWR 0.100405
R13377 VPWR.n2290 VPWR 0.100405
R13378 VPWR.n2291 VPWR 0.100405
R13379 VPWR.n2292 VPWR 0.100405
R13380 VPWR.n2293 VPWR 0.100405
R13381 VPWR.n2294 VPWR 0.100405
R13382 VPWR.n2295 VPWR 0.100405
R13383 VPWR.n2296 VPWR 0.100405
R13384 VPWR.n2297 VPWR 0.100405
R13385 VPWR.n2298 VPWR 0.100405
R13386 VPWR.n2285 VPWR 0.100405
R13387 VPWR.n2276 VPWR 0.100405
R13388 VPWR.n2275 VPWR 0.100405
R13389 VPWR.n2266 VPWR 0.100405
R13390 VPWR.n2215 VPWR 0.100405
R13391 VPWR.n2216 VPWR 0.100405
R13392 VPWR.n2225 VPWR 0.100405
R13393 VPWR.n2226 VPWR 0.100405
R13394 VPWR.n2235 VPWR 0.100405
R13395 VPWR.n2236 VPWR 0.100405
R13396 VPWR.n2245 VPWR 0.100405
R13397 VPWR.n2246 VPWR 0.100405
R13398 VPWR.n2255 VPWR 0.100405
R13399 VPWR.n2256 VPWR 0.100405
R13400 VPWR.n2265 VPWR 0.100405
R13401 VPWR VPWR.n2189 0.100405
R13402 VPWR VPWR.n2190 0.100405
R13403 VPWR VPWR.n2191 0.100405
R13404 VPWR VPWR.n2192 0.100405
R13405 VPWR VPWR.n2203 0.100405
R13406 VPWR VPWR.n2202 0.100405
R13407 VPWR VPWR.n2201 0.100405
R13408 VPWR VPWR.n2200 0.100405
R13409 VPWR VPWR.n2199 0.100405
R13410 VPWR VPWR.n2198 0.100405
R13411 VPWR VPWR.n2197 0.100405
R13412 VPWR VPWR.n2196 0.100405
R13413 VPWR VPWR.n2195 0.100405
R13414 VPWR VPWR.n2194 0.100405
R13415 VPWR VPWR.n2193 0.100405
R13416 VPWR.n2109 VPWR 0.100405
R13417 VPWR VPWR.n2118 0.100405
R13418 VPWR.n2119 VPWR 0.100405
R13419 VPWR VPWR.n2128 0.100405
R13420 VPWR.n2179 VPWR 0.100405
R13421 VPWR VPWR.n2178 0.100405
R13422 VPWR.n2169 VPWR 0.100405
R13423 VPWR VPWR.n2168 0.100405
R13424 VPWR.n2159 VPWR 0.100405
R13425 VPWR VPWR.n2158 0.100405
R13426 VPWR.n2149 VPWR 0.100405
R13427 VPWR VPWR.n2148 0.100405
R13428 VPWR.n2139 VPWR 0.100405
R13429 VPWR VPWR.n2138 0.100405
R13430 VPWR.n2129 VPWR 0.100405
R13431 VPWR.n2106 VPWR 0.100405
R13432 VPWR.n2105 VPWR 0.100405
R13433 VPWR.n2104 VPWR 0.100405
R13434 VPWR.n2103 VPWR 0.100405
R13435 VPWR.n2092 VPWR 0.100405
R13436 VPWR.n2093 VPWR 0.100405
R13437 VPWR.n2094 VPWR 0.100405
R13438 VPWR.n2095 VPWR 0.100405
R13439 VPWR.n2096 VPWR 0.100405
R13440 VPWR.n2097 VPWR 0.100405
R13441 VPWR.n2098 VPWR 0.100405
R13442 VPWR.n2099 VPWR 0.100405
R13443 VPWR.n2100 VPWR 0.100405
R13444 VPWR.n2101 VPWR 0.100405
R13445 VPWR.n2102 VPWR 0.100405
R13446 VPWR.n2089 VPWR 0.100405
R13447 VPWR.n2080 VPWR 0.100405
R13448 VPWR.n2079 VPWR 0.100405
R13449 VPWR.n2070 VPWR 0.100405
R13450 VPWR.n2019 VPWR 0.100405
R13451 VPWR.n2020 VPWR 0.100405
R13452 VPWR.n2029 VPWR 0.100405
R13453 VPWR.n2030 VPWR 0.100405
R13454 VPWR.n2039 VPWR 0.100405
R13455 VPWR.n2040 VPWR 0.100405
R13456 VPWR.n2049 VPWR 0.100405
R13457 VPWR.n2050 VPWR 0.100405
R13458 VPWR.n2059 VPWR 0.100405
R13459 VPWR.n2060 VPWR 0.100405
R13460 VPWR.n2069 VPWR 0.100405
R13461 VPWR VPWR.n1993 0.100405
R13462 VPWR VPWR.n1994 0.100405
R13463 VPWR VPWR.n1995 0.100405
R13464 VPWR VPWR.n1996 0.100405
R13465 VPWR VPWR.n2007 0.100405
R13466 VPWR VPWR.n2006 0.100405
R13467 VPWR VPWR.n2005 0.100405
R13468 VPWR VPWR.n2004 0.100405
R13469 VPWR VPWR.n2003 0.100405
R13470 VPWR VPWR.n2002 0.100405
R13471 VPWR VPWR.n2001 0.100405
R13472 VPWR VPWR.n2000 0.100405
R13473 VPWR VPWR.n1999 0.100405
R13474 VPWR VPWR.n1998 0.100405
R13475 VPWR VPWR.n1997 0.100405
R13476 VPWR.n1913 VPWR 0.100405
R13477 VPWR VPWR.n1922 0.100405
R13478 VPWR.n1923 VPWR 0.100405
R13479 VPWR VPWR.n1932 0.100405
R13480 VPWR.n1983 VPWR 0.100405
R13481 VPWR VPWR.n1982 0.100405
R13482 VPWR.n1973 VPWR 0.100405
R13483 VPWR VPWR.n1972 0.100405
R13484 VPWR.n1963 VPWR 0.100405
R13485 VPWR VPWR.n1962 0.100405
R13486 VPWR.n1953 VPWR 0.100405
R13487 VPWR VPWR.n1952 0.100405
R13488 VPWR.n1943 VPWR 0.100405
R13489 VPWR VPWR.n1942 0.100405
R13490 VPWR.n1933 VPWR 0.100405
R13491 VPWR.n1910 VPWR 0.100405
R13492 VPWR.n1909 VPWR 0.100405
R13493 VPWR.n1908 VPWR 0.100405
R13494 VPWR.n1907 VPWR 0.100405
R13495 VPWR.n1896 VPWR 0.100405
R13496 VPWR.n1897 VPWR 0.100405
R13497 VPWR.n1898 VPWR 0.100405
R13498 VPWR.n1899 VPWR 0.100405
R13499 VPWR.n1900 VPWR 0.100405
R13500 VPWR.n1901 VPWR 0.100405
R13501 VPWR.n1902 VPWR 0.100405
R13502 VPWR.n1903 VPWR 0.100405
R13503 VPWR.n1904 VPWR 0.100405
R13504 VPWR.n1905 VPWR 0.100405
R13505 VPWR.n1906 VPWR 0.100405
R13506 VPWR VPWR.n2399 0.100405
R13507 VPWR VPWR.n2398 0.100405
R13508 VPWR VPWR.n2397 0.100405
R13509 VPWR VPWR.n2396 0.100405
R13510 VPWR VPWR.n2395 0.100405
R13511 VPWR VPWR.n2394 0.100405
R13512 VPWR VPWR.n2393 0.100405
R13513 VPWR VPWR.n2392 0.100405
R13514 VPWR VPWR.n2391 0.100405
R13515 VPWR VPWR.n2390 0.100405
R13516 VPWR VPWR.n2389 0.100405
R13517 VPWR VPWR.n2388 0.100405
R13518 VPWR.n1893 VPWR 0.100405
R13519 VPWR.n1884 VPWR 0.100405
R13520 VPWR.n1883 VPWR 0.100405
R13521 VPWR.n1874 VPWR 0.100405
R13522 VPWR.n1873 VPWR 0.100405
R13523 VPWR.n1823 VPWR 0.100405
R13524 VPWR.n1824 VPWR 0.100405
R13525 VPWR.n1833 VPWR 0.100405
R13526 VPWR.n1834 VPWR 0.100405
R13527 VPWR.n1843 VPWR 0.100405
R13528 VPWR.n1844 VPWR 0.100405
R13529 VPWR.n1853 VPWR 0.100405
R13530 VPWR.n1854 VPWR 0.100405
R13531 VPWR.n1863 VPWR 0.100405
R13532 VPWR.n1864 VPWR 0.100405
R13533 VPWR.n2411 VPWR 0.100405
R13534 VPWR.n2412 VPWR 0.100405
R13535 VPWR.n2421 VPWR 0.100405
R13536 VPWR.n2422 VPWR 0.100405
R13537 VPWR.n2431 VPWR 0.100405
R13538 VPWR.n2432 VPWR 0.100405
R13539 VPWR.n2441 VPWR 0.100405
R13540 VPWR.n2442 VPWR 0.100405
R13541 VPWR.n2451 VPWR 0.100405
R13542 VPWR.n2452 VPWR 0.100405
R13543 VPWR.n2461 VPWR 0.100405
R13544 VPWR.n2462 VPWR 0.100405
R13545 VPWR.n2471 VPWR 0.100405
R13546 VPWR VPWR.n1797 0.100405
R13547 VPWR VPWR.n1798 0.100405
R13548 VPWR VPWR.n1799 0.100405
R13549 VPWR VPWR.n1800 0.100405
R13550 VPWR VPWR.n1801 0.100405
R13551 VPWR VPWR.n1802 0.100405
R13552 VPWR VPWR.n1803 0.100405
R13553 VPWR VPWR.n1804 0.100405
R13554 VPWR VPWR.n1811 0.100405
R13555 VPWR VPWR.n1810 0.100405
R13556 VPWR VPWR.n1809 0.100405
R13557 VPWR VPWR.n1808 0.100405
R13558 VPWR VPWR.n1807 0.100405
R13559 VPWR VPWR.n1806 0.100405
R13560 VPWR VPWR.n1805 0.100405
R13561 VPWR.n2498 VPWR 0.100405
R13562 VPWR.n2497 VPWR 0.100405
R13563 VPWR.n2496 VPWR 0.100405
R13564 VPWR.n2495 VPWR 0.100405
R13565 VPWR.n2494 VPWR 0.100405
R13566 VPWR.n2493 VPWR 0.100405
R13567 VPWR.n2492 VPWR 0.100405
R13568 VPWR.n2491 VPWR 0.100405
R13569 VPWR.n2490 VPWR 0.100405
R13570 VPWR.n2489 VPWR 0.100405
R13571 VPWR.n2484 VPWR 0.100405
R13572 VPWR.n2485 VPWR 0.100405
R13573 VPWR.n2486 VPWR 0.100405
R13574 VPWR.n2487 VPWR 0.100405
R13575 VPWR.n2488 VPWR 0.100405
R13576 VPWR.n1143 VPWR 0.100405
R13577 VPWR VPWR.n1540 0.100405
R13578 VPWR.n1524 VPWR 0.100405
R13579 VPWR.n1516 VPWR 0.100405
R13580 VPWR.n1510 VPWR 0.100405
R13581 VPWR.n1502 VPWR 0.100405
R13582 VPWR.n1496 VPWR 0.100405
R13583 VPWR VPWR.n1132 0.100405
R13584 VPWR.n1584 VPWR 0.100405
R13585 VPWR.n1452 VPWR 0.100405
R13586 VPWR.n1464 VPWR 0.100405
R13587 VPWR.n1043 VPWR 0.100405
R13588 VPWR.n1744 VPWR 0.100405
R13589 VPWR.n1787 VPWR 0.100405
R13590 VPWR VPWR.n1765 0.100405
R13591 VPWR.n2501 VPWR 0.100405
R13592 VPWR VPWR.n2512 0.100405
R13593 VPWR.n2513 VPWR 0.100405
R13594 VPWR VPWR.n2524 0.100405
R13595 VPWR.n2525 VPWR 0.100405
R13596 VPWR VPWR.n2536 0.100405
R13597 VPWR.n2537 VPWR 0.100405
R13598 VPWR VPWR.n2548 0.100405
R13599 VPWR.n2549 VPWR 0.100405
R13600 VPWR VPWR.n2560 0.100405
R13601 VPWR.n2561 VPWR 0.100405
R13602 VPWR VPWR.n2572 0.100405
R13603 VPWR.n2573 VPWR 0.100405
R13604 VPWR VPWR.n2584 0.100405
R13605 VPWR.n2585 VPWR 0.100405
R13606 VPWR.n1056 VPWR 0.100405
R13607 VPWR.n1754 VPWR 0.100405
R13608 VPWR.n1755 VPWR 0.100405
R13609 VPWR.n1529 VPWR 0.100405
R13610 VPWR.n1530 VPWR 0.100405
R13611 VPWR VPWR.n1528 0.100405
R13612 VPWR VPWR.n1527 0.100405
R13613 VPWR.n1514 VPWR 0.100405
R13614 VPWR VPWR.n1513 0.100405
R13615 VPWR.n1500 VPWR 0.100405
R13616 VPWR VPWR.n1499 0.100405
R13617 VPWR.n1487 VPWR 0.100405
R13618 VPWR.n1587 VPWR 0.100405
R13619 VPWR.n1588 VPWR 0.100405
R13620 VPWR.n1448 VPWR 0.100405
R13621 VPWR VPWR.n2798 0.0994583
R13622 VPWR VPWR.n2779 0.0994583
R13623 VPWR VPWR.n1326 0.0981562
R13624 VPWR.n1371 VPWR 0.0981562
R13625 VPWR.n1410 VPWR 0.0981562
R13626 VPWR.n9 VPWR 0.0968542
R13627 VPWR.n1244 VPWR 0.0968542
R13628 VPWR.n1267 VPWR 0.0968542
R13629 VPWR.n1291 VPWR 0.0968542
R13630 VPWR.n1333 VPWR 0.0968542
R13631 VPWR VPWR.n2759 0.0968542
R13632 VPWR VPWR.n2740 0.0968542
R13633 VPWR.n2718 VPWR 0.0968542
R13634 VPWR.n2682 VPWR 0.0968542
R13635 VPWR.n2645 VPWR 0.0968542
R13636 VPWR.n2608 VPWR 0.0968542
R13637 VPWR VPWR.n1044 0.0945
R13638 VPWR.n1541 VPWR 0.0945
R13639 VPWR VPWR.n1142 0.0945
R13640 VPWR VPWR.n1141 0.0945
R13641 VPWR VPWR.n1140 0.0945
R13642 VPWR VPWR.n1139 0.0945
R13643 VPWR VPWR.n1138 0.0945
R13644 VPWR.n1137 VPWR 0.0945
R13645 VPWR VPWR.n1583 0.0945
R13646 VPWR VPWR.n1131 0.0945
R13647 VPWR VPWR.n1463 0.0945
R13648 VPWR.n1451 VPWR 0.0945
R13649 VPWR VPWR.n1038 0.0945
R13650 VPWR.n1786 VPWR 0.0945
R13651 VPWR VPWR.n1027 0.0945
R13652 VPWR.n1766 VPWR 0.0945
R13653 VPWR.n1117 VPWR 0.093504
R13654 VPWR.n109 VPWR 0.093504
R13655 VPWR.n143 VPWR 0.093504
R13656 VPWR.n155 VPWR 0.093504
R13657 VPWR.n167 VPWR 0.093504
R13658 VPWR.n179 VPWR 0.093504
R13659 VPWR.n191 VPWR 0.093504
R13660 VPWR.n203 VPWR 0.093504
R13661 VPWR.n215 VPWR 0.093504
R13662 VPWR.n227 VPWR 0.093504
R13663 VPWR.n239 VPWR 0.093504
R13664 VPWR.n251 VPWR 0.093504
R13665 VPWR.n263 VPWR 0.093504
R13666 VPWR.n275 VPWR 0.093504
R13667 VPWR VPWR.n285 0.093504
R13668 VPWR.n131 VPWR 0.093504
R13669 VPWR.n120 VPWR 0.093504
R13670 VPWR VPWR.n1731 0.093504
R13671 VPWR.n1722 VPWR 0.093504
R13672 VPWR.n1710 VPWR 0.093504
R13673 VPWR.n1699 VPWR 0.093504
R13674 VPWR VPWR.n1077 0.093504
R13675 VPWR.n1683 VPWR 0.093504
R13676 VPWR.n1672 VPWR 0.093504
R13677 VPWR VPWR.n1087 0.093504
R13678 VPWR.n1656 VPWR 0.093504
R13679 VPWR.n1645 VPWR 0.093504
R13680 VPWR VPWR.n1097 0.093504
R13681 VPWR.n1629 VPWR 0.093504
R13682 VPWR.n1618 VPWR 0.093504
R13683 VPWR VPWR.n1107 0.093504
R13684 VPWR.n1602 VPWR 0.093504
R13685 VPWR.n2598 VPWR 0.0849042
R13686 VPWR.n1112 VPWR.n1109 0.0845517
R13687 VPWR.n147 VPWR.n146 0.0845517
R13688 VPWR.n159 VPWR.n158 0.0845517
R13689 VPWR.n171 VPWR.n170 0.0845517
R13690 VPWR.n183 VPWR.n182 0.0845517
R13691 VPWR.n195 VPWR.n194 0.0845517
R13692 VPWR.n207 VPWR.n206 0.0845517
R13693 VPWR.n219 VPWR.n218 0.0845517
R13694 VPWR.n231 VPWR.n230 0.0845517
R13695 VPWR.n243 VPWR.n242 0.0845517
R13696 VPWR.n255 VPWR.n254 0.0845517
R13697 VPWR.n267 VPWR.n266 0.0845517
R13698 VPWR.n279 VPWR.n278 0.0845517
R13699 VPWR.n282 VPWR.n103 0.0845517
R13700 VPWR.n113 VPWR.n112 0.0845517
R13701 VPWR.n135 VPWR.n134 0.0845517
R13702 VPWR.n124 VPWR.n123 0.0845517
R13703 VPWR.n1728 VPWR.n1067 0.0845517
R13704 VPWR.n1726 VPWR.n1725 0.0845517
R13705 VPWR.n1714 VPWR.n1713 0.0845517
R13706 VPWR.n1701 VPWR.n1700 0.0845517
R13707 VPWR.n1690 VPWR.n1078 0.0845517
R13708 VPWR.n1687 VPWR.n1686 0.0845517
R13709 VPWR.n1674 VPWR.n1673 0.0845517
R13710 VPWR.n1663 VPWR.n1088 0.0845517
R13711 VPWR.n1660 VPWR.n1659 0.0845517
R13712 VPWR.n1647 VPWR.n1646 0.0845517
R13713 VPWR.n1636 VPWR.n1098 0.0845517
R13714 VPWR.n1633 VPWR.n1632 0.0845517
R13715 VPWR.n1620 VPWR.n1619 0.0845517
R13716 VPWR.n1609 VPWR.n1108 0.0845517
R13717 VPWR.n1606 VPWR.n1605 0.0845517
R13718 VPWR.n1456 VPWR.n1451 0.0740128
R13719 VPWR.n1542 VPWR.n1044 0.071
R13720 VPWR.n1547 VPWR.n1541 0.071
R13721 VPWR.n1552 VPWR.n1142 0.071
R13722 VPWR.n1557 VPWR.n1141 0.071
R13723 VPWR.n1562 VPWR.n1140 0.071
R13724 VPWR.n1567 VPWR.n1139 0.071
R13725 VPWR.n1572 VPWR.n1138 0.071
R13726 VPWR.n1577 VPWR.n1137 0.071
R13727 VPWR.n1583 VPWR.n1582 0.071
R13728 VPWR.n1457 VPWR.n1131 0.071
R13729 VPWR.n1463 VPWR.n1462 0.071
R13730 VPWR.n1772 VPWR.n1038 0.071
R13731 VPWR.n1786 VPWR.n1785 0.071
R13732 VPWR.n1780 VPWR.n1027 0.071
R13733 VPWR.n1767 VPWR.n1766 0.071
R13734 VPWR VPWR.n1115 0.0678077
R13735 VPWR VPWR.n107 0.0678077
R13736 VPWR VPWR.n141 0.0678077
R13737 VPWR VPWR.n153 0.0678077
R13738 VPWR VPWR.n165 0.0678077
R13739 VPWR VPWR.n177 0.0678077
R13740 VPWR VPWR.n189 0.0678077
R13741 VPWR VPWR.n201 0.0678077
R13742 VPWR VPWR.n213 0.0678077
R13743 VPWR VPWR.n225 0.0678077
R13744 VPWR VPWR.n237 0.0678077
R13745 VPWR VPWR.n249 0.0678077
R13746 VPWR VPWR.n261 0.0678077
R13747 VPWR VPWR.n273 0.0678077
R13748 VPWR.n286 VPWR 0.0678077
R13749 VPWR VPWR.n129 0.0678077
R13750 VPWR VPWR.n118 0.0678077
R13751 VPWR.n1732 VPWR 0.0678077
R13752 VPWR VPWR.n1720 0.0678077
R13753 VPWR VPWR.n1708 0.0678077
R13754 VPWR VPWR.n1697 0.0678077
R13755 VPWR.n1193 VPWR 0.0678077
R13756 VPWR VPWR.n1681 0.0678077
R13757 VPWR VPWR.n1670 0.0678077
R13758 VPWR.n1207 VPWR 0.0678077
R13759 VPWR VPWR.n1654 0.0678077
R13760 VPWR VPWR.n1643 0.0678077
R13761 VPWR.n1175 VPWR 0.0678077
R13762 VPWR VPWR.n1627 0.0678077
R13763 VPWR VPWR.n1616 0.0678077
R13764 VPWR.n1124 VPWR 0.0678077
R13765 VPWR VPWR.n1600 0.0678077
R13766 VPWR.n150 VPWR 0.063
R13767 VPWR.n162 VPWR 0.063
R13768 VPWR.n174 VPWR 0.063
R13769 VPWR.n186 VPWR 0.063
R13770 VPWR.n198 VPWR 0.063
R13771 VPWR.n210 VPWR 0.063
R13772 VPWR.n222 VPWR 0.063
R13773 VPWR.n234 VPWR 0.063
R13774 VPWR.n246 VPWR 0.063
R13775 VPWR.n258 VPWR 0.063
R13776 VPWR.n270 VPWR 0.063
R13777 VPWR.n101 VPWR 0.063
R13778 VPWR.n105 VPWR 0.063
R13779 VPWR.n138 VPWR 0.063
R13780 VPWR.n115 VPWR 0.063
R13781 VPWR.n126 VPWR 0.063
R13782 VPWR.n1065 VPWR 0.063
R13783 VPWR.n1717 VPWR 0.063
R13784 VPWR.n1070 VPWR 0.063
R13785 VPWR VPWR.n1704 0.063
R13786 VPWR VPWR.n1693 0.063
R13787 VPWR VPWR.n1081 0.063
R13788 VPWR VPWR.n1677 0.063
R13789 VPWR VPWR.n1666 0.063
R13790 VPWR VPWR.n1091 0.063
R13791 VPWR VPWR.n1650 0.063
R13792 VPWR VPWR.n1639 0.063
R13793 VPWR VPWR.n1101 0.063
R13794 VPWR VPWR.n1623 0.063
R13795 VPWR VPWR.n1612 0.063
R13796 VPWR VPWR.n1111 0.063
R13797 VPWR VPWR.n1120 0.063
R13798 VPWR.n1115 VPWR 0.0608448
R13799 VPWR.n107 VPWR 0.0608448
R13800 VPWR.n141 VPWR 0.0608448
R13801 VPWR.n153 VPWR 0.0608448
R13802 VPWR.n165 VPWR 0.0608448
R13803 VPWR.n177 VPWR 0.0608448
R13804 VPWR.n189 VPWR 0.0608448
R13805 VPWR.n201 VPWR 0.0608448
R13806 VPWR.n213 VPWR 0.0608448
R13807 VPWR.n225 VPWR 0.0608448
R13808 VPWR.n237 VPWR 0.0608448
R13809 VPWR.n249 VPWR 0.0608448
R13810 VPWR.n261 VPWR 0.0608448
R13811 VPWR.n273 VPWR 0.0608448
R13812 VPWR.n286 VPWR 0.0608448
R13813 VPWR.n129 VPWR 0.0608448
R13814 VPWR.n118 VPWR 0.0608448
R13815 VPWR.n1732 VPWR 0.0608448
R13816 VPWR.n1720 VPWR 0.0608448
R13817 VPWR.n1708 VPWR 0.0608448
R13818 VPWR.n1697 VPWR 0.0608448
R13819 VPWR.n1193 VPWR 0.0608448
R13820 VPWR.n1681 VPWR 0.0608448
R13821 VPWR.n1670 VPWR 0.0608448
R13822 VPWR.n1207 VPWR 0.0608448
R13823 VPWR.n1654 VPWR 0.0608448
R13824 VPWR.n1643 VPWR 0.0608448
R13825 VPWR.n1175 VPWR 0.0608448
R13826 VPWR.n1627 VPWR 0.0608448
R13827 VPWR.n1616 VPWR 0.0608448
R13828 VPWR.n1124 VPWR 0.0608448
R13829 VPWR.n1600 VPWR 0.0608448
R13830 VPWR VPWR.n13 0.0603958
R13831 VPWR VPWR.n12 0.0603958
R13832 VPWR VPWR.n1249 0.0603958
R13833 VPWR VPWR.n1248 0.0603958
R13834 VPWR VPWR.n1272 0.0603958
R13835 VPWR VPWR.n1271 0.0603958
R13836 VPWR VPWR.n1296 0.0603958
R13837 VPWR VPWR.n1295 0.0603958
R13838 VPWR.n1332 VPWR 0.0603958
R13839 VPWR VPWR.n1331 0.0603958
R13840 VPWR.n1327 VPWR 0.0603958
R13841 VPWR.n1318 VPWR 0.0603958
R13842 VPWR VPWR.n1317 0.0603958
R13843 VPWR.n1370 VPWR 0.0603958
R13844 VPWR VPWR.n1369 0.0603958
R13845 VPWR.n1364 VPWR 0.0603958
R13846 VPWR.n1409 VPWR 0.0603958
R13847 VPWR VPWR.n1408 0.0603958
R13848 VPWR.n1403 VPWR 0.0603958
R13849 VPWR.n1440 VPWR 0.0603958
R13850 VPWR VPWR.n2800 0.0603958
R13851 VPWR VPWR.n2799 0.0603958
R13852 VPWR VPWR.n2812 0.0603958
R13853 VPWR.n2791 VPWR 0.0603958
R13854 VPWR.n2792 VPWR 0.0603958
R13855 VPWR VPWR.n2796 0.0603958
R13856 VPWR.n2771 VPWR 0.0603958
R13857 VPWR.n2772 VPWR 0.0603958
R13858 VPWR VPWR.n2777 0.0603958
R13859 VPWR.n2752 VPWR 0.0603958
R13860 VPWR.n2753 VPWR 0.0603958
R13861 VPWR VPWR.n2757 0.0603958
R13862 VPWR.n2733 VPWR 0.0603958
R13863 VPWR.n2734 VPWR 0.0603958
R13864 VPWR VPWR.n2695 0.0603958
R13865 VPWR.n2696 VPWR 0.0603958
R13866 VPWR.n2697 VPWR 0.0603958
R13867 VPWR VPWR.n2658 0.0603958
R13868 VPWR.n2659 VPWR 0.0603958
R13869 VPWR.n2660 VPWR 0.0603958
R13870 VPWR.n2624 VPWR 0.0603958
R13871 VPWR.n2627 VPWR 0.0603958
R13872 VPWR.n1770 VPWR.n1769 0.0599512
R13873 VPWR.n1041 VPWR.n1040 0.0599512
R13874 VPWR.n1545 VPWR.n1544 0.0599512
R13875 VPWR.n1550 VPWR.n1549 0.0599512
R13876 VPWR.n1555 VPWR.n1554 0.0599512
R13877 VPWR.n1560 VPWR.n1559 0.0599512
R13878 VPWR.n1565 VPWR.n1564 0.0599512
R13879 VPWR.n1570 VPWR.n1569 0.0599512
R13880 VPWR.n1575 VPWR.n1574 0.0599512
R13881 VPWR.n1580 VPWR.n1579 0.0599512
R13882 VPWR.n1135 VPWR.n1134 0.0599512
R13883 VPWR.n1460 VPWR.n1459 0.0599512
R13884 VPWR.n1455 VPWR.n1454 0.0599512
R13885 VPWR.n1775 VPWR.n1774 0.0599512
R13886 VPWR.n1783 VPWR.n1782 0.0599512
R13887 VPWR.n1779 VPWR.n1778 0.0599512
R13888 VPWR.n1118 VPWR.n1117 0.0565345
R13889 VPWR.n1112 VPWR 0.0565345
R13890 VPWR.n144 VPWR.n143 0.0565345
R13891 VPWR.n146 VPWR 0.0565345
R13892 VPWR.n156 VPWR.n155 0.0565345
R13893 VPWR.n158 VPWR 0.0565345
R13894 VPWR.n168 VPWR.n167 0.0565345
R13895 VPWR.n170 VPWR 0.0565345
R13896 VPWR.n180 VPWR.n179 0.0565345
R13897 VPWR.n182 VPWR 0.0565345
R13898 VPWR.n192 VPWR.n191 0.0565345
R13899 VPWR.n194 VPWR 0.0565345
R13900 VPWR.n204 VPWR.n203 0.0565345
R13901 VPWR.n206 VPWR 0.0565345
R13902 VPWR.n216 VPWR.n215 0.0565345
R13903 VPWR.n218 VPWR 0.0565345
R13904 VPWR.n228 VPWR.n227 0.0565345
R13905 VPWR.n230 VPWR 0.0565345
R13906 VPWR.n240 VPWR.n239 0.0565345
R13907 VPWR.n242 VPWR 0.0565345
R13908 VPWR.n252 VPWR.n251 0.0565345
R13909 VPWR.n254 VPWR 0.0565345
R13910 VPWR.n264 VPWR.n263 0.0565345
R13911 VPWR.n266 VPWR 0.0565345
R13912 VPWR.n276 VPWR.n275 0.0565345
R13913 VPWR.n278 VPWR 0.0565345
R13914 VPWR.n285 VPWR.n283 0.0565345
R13915 VPWR.n103 VPWR 0.0565345
R13916 VPWR.n110 VPWR.n109 0.0565345
R13917 VPWR.n112 VPWR 0.0565345
R13918 VPWR.n132 VPWR.n131 0.0565345
R13919 VPWR.n134 VPWR 0.0565345
R13920 VPWR.n121 VPWR.n120 0.0565345
R13921 VPWR.n123 VPWR 0.0565345
R13922 VPWR.n1731 VPWR.n1729 0.0565345
R13923 VPWR.n1067 VPWR 0.0565345
R13924 VPWR.n1723 VPWR.n1722 0.0565345
R13925 VPWR.n1725 VPWR 0.0565345
R13926 VPWR.n1711 VPWR.n1710 0.0565345
R13927 VPWR.n1713 VPWR 0.0565345
R13928 VPWR.n1702 VPWR.n1699 0.0565345
R13929 VPWR.n1700 VPWR 0.0565345
R13930 VPWR.n1691 VPWR.n1077 0.0565345
R13931 VPWR.n1078 VPWR 0.0565345
R13932 VPWR.n1684 VPWR.n1683 0.0565345
R13933 VPWR.n1686 VPWR 0.0565345
R13934 VPWR.n1675 VPWR.n1672 0.0565345
R13935 VPWR.n1673 VPWR 0.0565345
R13936 VPWR.n1664 VPWR.n1087 0.0565345
R13937 VPWR.n1088 VPWR 0.0565345
R13938 VPWR.n1657 VPWR.n1656 0.0565345
R13939 VPWR.n1659 VPWR 0.0565345
R13940 VPWR.n1648 VPWR.n1645 0.0565345
R13941 VPWR.n1646 VPWR 0.0565345
R13942 VPWR.n1637 VPWR.n1097 0.0565345
R13943 VPWR.n1098 VPWR 0.0565345
R13944 VPWR.n1630 VPWR.n1629 0.0565345
R13945 VPWR.n1632 VPWR 0.0565345
R13946 VPWR.n1621 VPWR.n1618 0.0565345
R13947 VPWR.n1619 VPWR 0.0565345
R13948 VPWR.n1610 VPWR.n1107 0.0565345
R13949 VPWR.n1108 VPWR 0.0565345
R13950 VPWR.n1603 VPWR.n1602 0.0565345
R13951 VPWR.n1605 VPWR 0.0565345
R13952 VPWR.n1769 VPWR 0.0469286
R13953 VPWR.n1040 VPWR 0.0469286
R13954 VPWR.n1544 VPWR 0.0469286
R13955 VPWR.n1549 VPWR 0.0469286
R13956 VPWR.n1554 VPWR 0.0469286
R13957 VPWR.n1559 VPWR 0.0469286
R13958 VPWR.n1564 VPWR 0.0469286
R13959 VPWR.n1569 VPWR 0.0469286
R13960 VPWR.n1574 VPWR 0.0469286
R13961 VPWR.n1579 VPWR 0.0469286
R13962 VPWR.n1134 VPWR 0.0469286
R13963 VPWR.n1459 VPWR 0.0469286
R13964 VPWR.n1454 VPWR 0.0469286
R13965 VPWR.n1774 VPWR 0.0469286
R13966 VPWR.n1782 VPWR 0.0469286
R13967 VPWR.n1778 VPWR 0.0469286
R13968 VPWR.n1769 VPWR 0.0401341
R13969 VPWR.n1040 VPWR 0.0401341
R13970 VPWR.n1544 VPWR 0.0401341
R13971 VPWR.n1549 VPWR 0.0401341
R13972 VPWR.n1554 VPWR 0.0401341
R13973 VPWR.n1559 VPWR 0.0401341
R13974 VPWR.n1564 VPWR 0.0401341
R13975 VPWR.n1569 VPWR 0.0401341
R13976 VPWR.n1574 VPWR 0.0401341
R13977 VPWR.n1579 VPWR 0.0401341
R13978 VPWR.n1134 VPWR 0.0401341
R13979 VPWR.n1459 VPWR 0.0401341
R13980 VPWR.n1454 VPWR 0.0401341
R13981 VPWR.n1774 VPWR 0.0401341
R13982 VPWR.n1782 VPWR 0.0401341
R13983 VPWR.n1778 VPWR 0.0401341
R13984 VPWR.n13 VPWR 0.0382604
R13985 VPWR.n1249 VPWR 0.0382604
R13986 VPWR.n1272 VPWR 0.0382604
R13987 VPWR.n1296 VPWR 0.0382604
R13988 VPWR.n1331 VPWR 0.0382604
R13989 VPWR.n1369 VPWR 0.0382604
R13990 VPWR.n1408 VPWR 0.0382604
R13991 VPWR.n1445 VPWR 0.0382604
R13992 VPWR.n20 VPWR 0.0375125
R13993 VPWR.n20 VPWR 0.0373589
R13994 VPWR.n1118 VPWR.n1109 0.0349828
R13995 VPWR.n147 VPWR.n144 0.0349828
R13996 VPWR.n159 VPWR.n156 0.0349828
R13997 VPWR.n171 VPWR.n168 0.0349828
R13998 VPWR.n183 VPWR.n180 0.0349828
R13999 VPWR.n195 VPWR.n192 0.0349828
R14000 VPWR.n207 VPWR.n204 0.0349828
R14001 VPWR.n219 VPWR.n216 0.0349828
R14002 VPWR.n231 VPWR.n228 0.0349828
R14003 VPWR.n243 VPWR.n240 0.0349828
R14004 VPWR.n255 VPWR.n252 0.0349828
R14005 VPWR.n267 VPWR.n264 0.0349828
R14006 VPWR.n279 VPWR.n276 0.0349828
R14007 VPWR.n283 VPWR.n282 0.0349828
R14008 VPWR.n113 VPWR.n110 0.0349828
R14009 VPWR.n135 VPWR.n132 0.0349828
R14010 VPWR.n124 VPWR.n121 0.0349828
R14011 VPWR.n1729 VPWR.n1728 0.0349828
R14012 VPWR.n1726 VPWR.n1723 0.0349828
R14013 VPWR.n1714 VPWR.n1711 0.0349828
R14014 VPWR.n1702 VPWR.n1701 0.0349828
R14015 VPWR.n1691 VPWR.n1690 0.0349828
R14016 VPWR.n1687 VPWR.n1684 0.0349828
R14017 VPWR.n1675 VPWR.n1674 0.0349828
R14018 VPWR.n1664 VPWR.n1663 0.0349828
R14019 VPWR.n1660 VPWR.n1657 0.0349828
R14020 VPWR.n1648 VPWR.n1647 0.0349828
R14021 VPWR.n1637 VPWR.n1636 0.0349828
R14022 VPWR.n1633 VPWR.n1630 0.0349828
R14023 VPWR.n1621 VPWR.n1620 0.0349828
R14024 VPWR.n1610 VPWR.n1609 0.0349828
R14025 VPWR.n1606 VPWR.n1603 0.0349828
R14026 VPWR.n2504 VPWR.n2503 0.0340366
R14027 VPWR.n2570 VPWR.n2569 0.0340366
R14028 VPWR.n2510 VPWR.n2509 0.0340366
R14029 VPWR.n2552 VPWR.n2551 0.0340366
R14030 VPWR.n2546 VPWR.n2545 0.0340366
R14031 VPWR.n2534 VPWR.n2533 0.0340366
R14032 VPWR.n2528 VPWR.n2527 0.0340366
R14033 VPWR.n1223 VPWR.n1222 0.0340366
R14034 VPWR.n2522 VPWR.n2521 0.0340366
R14035 VPWR.n1486 VPWR.n1102 0.0340366
R14036 VPWR.n1174 VPWR.n1094 0.0340366
R14037 VPWR.n2540 VPWR.n2539 0.0340366
R14038 VPWR.n1165 VPWR.n1092 0.0340366
R14039 VPWR.n1211 VPWR.n1164 0.0340366
R14040 VPWR.n2516 VPWR.n2515 0.0340366
R14041 VPWR.n1129 VPWR.n1104 0.0340366
R14042 VPWR.n1155 VPWR.n1084 0.0340366
R14043 VPWR.n2558 VPWR.n2557 0.0340366
R14044 VPWR.n1144 VPWR.n1082 0.0340366
R14045 VPWR.n1591 VPWR.n1590 0.0340366
R14046 VPWR.n2564 VPWR.n2563 0.0340366
R14047 VPWR.n1197 VPWR.n1154 0.0340366
R14048 VPWR.n1074 VPWR.n1073 0.0340366
R14049 VPWR.n1743 VPWR.n1742 0.0340366
R14050 VPWR.n1071 VPWR.n1054 0.0340366
R14051 VPWR.n2576 VPWR.n2575 0.0340366
R14052 VPWR.n2582 VPWR.n2581 0.0340366
R14053 VPWR.n2593 VPWR.n2592 0.0340366
R14054 VPWR.n2588 VPWR.n2587 0.0340366
R14055 VPWR.n1737 VPWR.n1736 0.0340366
R14056 VPWR.n1063 VPWR.n1060 0.0340366
R14057 VPWR.n1596 VPWR.n1121 0.0340366
R14058 VPWR.n2628 VPWR.n2598 0.0320292
R14059 VPWR.n2800 VPWR 0.03175
R14060 VPWR VPWR.n2791 0.03175
R14061 VPWR VPWR.n2771 0.03175
R14062 VPWR VPWR.n2752 0.03175
R14063 VPWR VPWR.n2733 0.03175
R14064 VPWR VPWR.n2696 0.03175
R14065 VPWR VPWR.n2659 0.03175
R14066 VPWR VPWR.n2627 0.03175
R14067 VPWR.n2598 VPWR.n2597 0.0240975
R14068 VPWR.n2597 VPWR.n20 0.0240975
R14069 VPWR.n2814 VPWR 0.024
R14070 VPWR.n14 VPWR 0.0239375
R14071 VPWR.n12 VPWR 0.0239375
R14072 VPWR.n1250 VPWR 0.0239375
R14073 VPWR.n1248 VPWR 0.0239375
R14074 VPWR.n1271 VPWR 0.0239375
R14075 VPWR.n1295 VPWR 0.0239375
R14076 VPWR.n2753 VPWR 0.0239375
R14077 VPWR.n2503 VPWR 0.0233659
R14078 VPWR.n1466 VPWR 0.0233659
R14079 VPWR.n352 VPWR 0.0233659
R14080 VPWR.n2570 VPWR 0.0233659
R14081 VPWR.n1533 VPWR 0.0233659
R14082 VPWR.n347 VPWR 0.0233659
R14083 VPWR.n2510 VPWR 0.0233659
R14084 VPWR.n964 VPWR 0.0233659
R14085 VPWR.n2479 VPWR 0.0233659
R14086 VPWR.n2474 VPWR 0.0233659
R14087 VPWR.n319 VPWR 0.0233659
R14088 VPWR.n2551 VPWR 0.0233659
R14089 VPWR.n972 VPWR 0.0233659
R14090 VPWR.n2444 VPWR 0.0233659
R14091 VPWR.n323 VPWR 0.0233659
R14092 VPWR.n2546 VPWR 0.0233659
R14093 VPWR.n1891 VPWR 0.0233659
R14094 VPWR.n1886 VPWR 0.0233659
R14095 VPWR.n1881 VPWR 0.0233659
R14096 VPWR.n388 VPWR 0.0233659
R14097 VPWR.n392 VPWR 0.0233659
R14098 VPWR.n396 VPWR 0.0233659
R14099 VPWR.n2454 VPWR 0.0233659
R14100 VPWR.n331 VPWR 0.0233659
R14101 VPWR.n2534 VPWR 0.0233659
R14102 VPWR.n1876 VPWR 0.0233659
R14103 VPWR.n404 VPWR 0.0233659
R14104 VPWR.n2459 VPWR 0.0233659
R14105 VPWR.n335 VPWR 0.0233659
R14106 VPWR.n2527 VPWR 0.0233659
R14107 VPWR.n2307 VPWR 0.0233659
R14108 VPWR.n2312 VPWR 0.0233659
R14109 VPWR.n2317 VPWR 0.0233659
R14110 VPWR.n2322 VPWR 0.0233659
R14111 VPWR.n2332 VPWR 0.0233659
R14112 VPWR.n2337 VPWR 0.0233659
R14113 VPWR.n2342 VPWR 0.0233659
R14114 VPWR.n2347 VPWR 0.0233659
R14115 VPWR.n2352 VPWR 0.0233659
R14116 VPWR.n2357 VPWR 0.0233659
R14117 VPWR.n2362 VPWR 0.0233659
R14118 VPWR.n2367 VPWR 0.0233659
R14119 VPWR.n2372 VPWR 0.0233659
R14120 VPWR.n2377 VPWR 0.0233659
R14121 VPWR.n2381 VPWR 0.0233659
R14122 VPWR.n2327 VPWR 0.0233659
R14123 VPWR.n544 VPWR 0.0233659
R14124 VPWR.n539 VPWR 0.0233659
R14125 VPWR.n535 VPWR 0.0233659
R14126 VPWR.n531 VPWR 0.0233659
R14127 VPWR.n523 VPWR 0.0233659
R14128 VPWR.n519 VPWR 0.0233659
R14129 VPWR.n515 VPWR 0.0233659
R14130 VPWR.n511 VPWR 0.0233659
R14131 VPWR.n507 VPWR 0.0233659
R14132 VPWR.n503 VPWR 0.0233659
R14133 VPWR.n499 VPWR 0.0233659
R14134 VPWR.n495 VPWR 0.0233659
R14135 VPWR.n491 VPWR 0.0233659
R14136 VPWR.n487 VPWR 0.0233659
R14137 VPWR.n484 VPWR 0.0233659
R14138 VPWR.n527 VPWR 0.0233659
R14139 VPWR.n2283 VPWR 0.0233659
R14140 VPWR.n2278 VPWR 0.0233659
R14141 VPWR.n2273 VPWR 0.0233659
R14142 VPWR.n2268 VPWR 0.0233659
R14143 VPWR.n2258 VPWR 0.0233659
R14144 VPWR.n2253 VPWR 0.0233659
R14145 VPWR.n2248 VPWR 0.0233659
R14146 VPWR.n2243 VPWR 0.0233659
R14147 VPWR.n2238 VPWR 0.0233659
R14148 VPWR.n2233 VPWR 0.0233659
R14149 VPWR.n2228 VPWR 0.0233659
R14150 VPWR.n2223 VPWR 0.0233659
R14151 VPWR.n2218 VPWR 0.0233659
R14152 VPWR.n2213 VPWR 0.0233659
R14153 VPWR.n2209 VPWR 0.0233659
R14154 VPWR.n2263 VPWR 0.0233659
R14155 VPWR.n580 VPWR 0.0233659
R14156 VPWR.n584 VPWR 0.0233659
R14157 VPWR.n588 VPWR 0.0233659
R14158 VPWR.n592 VPWR 0.0233659
R14159 VPWR.n600 VPWR 0.0233659
R14160 VPWR.n604 VPWR 0.0233659
R14161 VPWR.n608 VPWR 0.0233659
R14162 VPWR.n612 VPWR 0.0233659
R14163 VPWR.n616 VPWR 0.0233659
R14164 VPWR.n620 VPWR 0.0233659
R14165 VPWR.n624 VPWR 0.0233659
R14166 VPWR.n628 VPWR 0.0233659
R14167 VPWR.n632 VPWR 0.0233659
R14168 VPWR.n636 VPWR 0.0233659
R14169 VPWR.n640 VPWR 0.0233659
R14170 VPWR.n596 VPWR 0.0233659
R14171 VPWR.n2111 VPWR 0.0233659
R14172 VPWR.n2116 VPWR 0.0233659
R14173 VPWR.n2121 VPWR 0.0233659
R14174 VPWR.n2126 VPWR 0.0233659
R14175 VPWR.n2136 VPWR 0.0233659
R14176 VPWR.n2141 VPWR 0.0233659
R14177 VPWR.n2146 VPWR 0.0233659
R14178 VPWR.n2151 VPWR 0.0233659
R14179 VPWR.n2156 VPWR 0.0233659
R14180 VPWR.n2161 VPWR 0.0233659
R14181 VPWR.n2166 VPWR 0.0233659
R14182 VPWR.n2171 VPWR 0.0233659
R14183 VPWR.n2176 VPWR 0.0233659
R14184 VPWR.n2181 VPWR 0.0233659
R14185 VPWR.n2185 VPWR 0.0233659
R14186 VPWR.n2131 VPWR 0.0233659
R14187 VPWR.n736 VPWR 0.0233659
R14188 VPWR.n731 VPWR 0.0233659
R14189 VPWR.n727 VPWR 0.0233659
R14190 VPWR.n723 VPWR 0.0233659
R14191 VPWR.n715 VPWR 0.0233659
R14192 VPWR.n711 VPWR 0.0233659
R14193 VPWR.n707 VPWR 0.0233659
R14194 VPWR.n703 VPWR 0.0233659
R14195 VPWR.n699 VPWR 0.0233659
R14196 VPWR.n695 VPWR 0.0233659
R14197 VPWR.n691 VPWR 0.0233659
R14198 VPWR.n687 VPWR 0.0233659
R14199 VPWR.n683 VPWR 0.0233659
R14200 VPWR.n679 VPWR 0.0233659
R14201 VPWR.n676 VPWR 0.0233659
R14202 VPWR.n719 VPWR 0.0233659
R14203 VPWR.n2087 VPWR 0.0233659
R14204 VPWR.n2082 VPWR 0.0233659
R14205 VPWR.n2077 VPWR 0.0233659
R14206 VPWR.n2072 VPWR 0.0233659
R14207 VPWR.n2062 VPWR 0.0233659
R14208 VPWR.n2057 VPWR 0.0233659
R14209 VPWR.n2052 VPWR 0.0233659
R14210 VPWR.n2047 VPWR 0.0233659
R14211 VPWR.n2042 VPWR 0.0233659
R14212 VPWR.n2037 VPWR 0.0233659
R14213 VPWR.n2032 VPWR 0.0233659
R14214 VPWR.n2027 VPWR 0.0233659
R14215 VPWR.n2022 VPWR 0.0233659
R14216 VPWR.n2017 VPWR 0.0233659
R14217 VPWR.n2013 VPWR 0.0233659
R14218 VPWR.n2067 VPWR 0.0233659
R14219 VPWR.n772 VPWR 0.0233659
R14220 VPWR.n776 VPWR 0.0233659
R14221 VPWR.n780 VPWR 0.0233659
R14222 VPWR.n784 VPWR 0.0233659
R14223 VPWR.n792 VPWR 0.0233659
R14224 VPWR.n796 VPWR 0.0233659
R14225 VPWR.n800 VPWR 0.0233659
R14226 VPWR.n804 VPWR 0.0233659
R14227 VPWR.n808 VPWR 0.0233659
R14228 VPWR.n812 VPWR 0.0233659
R14229 VPWR.n816 VPWR 0.0233659
R14230 VPWR.n820 VPWR 0.0233659
R14231 VPWR.n824 VPWR 0.0233659
R14232 VPWR.n828 VPWR 0.0233659
R14233 VPWR.n832 VPWR 0.0233659
R14234 VPWR.n788 VPWR 0.0233659
R14235 VPWR.n1915 VPWR 0.0233659
R14236 VPWR.n1920 VPWR 0.0233659
R14237 VPWR.n1925 VPWR 0.0233659
R14238 VPWR.n1930 VPWR 0.0233659
R14239 VPWR.n1940 VPWR 0.0233659
R14240 VPWR.n1945 VPWR 0.0233659
R14241 VPWR.n1950 VPWR 0.0233659
R14242 VPWR.n1955 VPWR 0.0233659
R14243 VPWR.n1960 VPWR 0.0233659
R14244 VPWR.n1965 VPWR 0.0233659
R14245 VPWR.n1970 VPWR 0.0233659
R14246 VPWR.n1975 VPWR 0.0233659
R14247 VPWR.n1980 VPWR 0.0233659
R14248 VPWR.n1985 VPWR 0.0233659
R14249 VPWR.n1989 VPWR 0.0233659
R14250 VPWR.n1935 VPWR 0.0233659
R14251 VPWR.n928 VPWR 0.0233659
R14252 VPWR.n923 VPWR 0.0233659
R14253 VPWR.n919 VPWR 0.0233659
R14254 VPWR.n915 VPWR 0.0233659
R14255 VPWR.n907 VPWR 0.0233659
R14256 VPWR.n903 VPWR 0.0233659
R14257 VPWR.n899 VPWR 0.0233659
R14258 VPWR.n895 VPWR 0.0233659
R14259 VPWR.n891 VPWR 0.0233659
R14260 VPWR.n887 VPWR 0.0233659
R14261 VPWR.n883 VPWR 0.0233659
R14262 VPWR.n879 VPWR 0.0233659
R14263 VPWR.n875 VPWR 0.0233659
R14264 VPWR.n871 VPWR 0.0233659
R14265 VPWR.n868 VPWR 0.0233659
R14266 VPWR.n911 VPWR 0.0233659
R14267 VPWR.n1871 VPWR 0.0233659
R14268 VPWR.n980 VPWR 0.0233659
R14269 VPWR.n1495 VPWR 0.0233659
R14270 VPWR.n1223 VPWR 0.0233659
R14271 VPWR.n400 VPWR 0.0233659
R14272 VPWR.n2464 VPWR 0.0233659
R14273 VPWR.n339 VPWR 0.0233659
R14274 VPWR.n2522 VPWR 0.0233659
R14275 VPWR.n976 VPWR 0.0233659
R14276 VPWR.n1490 VPWR 0.0233659
R14277 VPWR.n1486 VPWR 0.0233659
R14278 VPWR.n1866 VPWR 0.0233659
R14279 VPWR.n984 VPWR 0.0233659
R14280 VPWR.n1504 VPWR 0.0233659
R14281 VPWR.n1174 VPWR 0.0233659
R14282 VPWR.n408 VPWR 0.0233659
R14283 VPWR.n416 VPWR 0.0233659
R14284 VPWR.n420 VPWR 0.0233659
R14285 VPWR.n424 VPWR 0.0233659
R14286 VPWR.n428 VPWR 0.0233659
R14287 VPWR.n432 VPWR 0.0233659
R14288 VPWR.n436 VPWR 0.0233659
R14289 VPWR.n440 VPWR 0.0233659
R14290 VPWR.n444 VPWR 0.0233659
R14291 VPWR.n448 VPWR 0.0233659
R14292 VPWR.n412 VPWR 0.0233659
R14293 VPWR.n2449 VPWR 0.0233659
R14294 VPWR.n327 VPWR 0.0233659
R14295 VPWR.n2539 VPWR 0.0233659
R14296 VPWR.n988 VPWR 0.0233659
R14297 VPWR.n1509 VPWR 0.0233659
R14298 VPWR.n1165 VPWR 0.0233659
R14299 VPWR.n1861 VPWR 0.0233659
R14300 VPWR.n1851 VPWR 0.0233659
R14301 VPWR.n1846 VPWR 0.0233659
R14302 VPWR.n1841 VPWR 0.0233659
R14303 VPWR.n1836 VPWR 0.0233659
R14304 VPWR.n1831 VPWR 0.0233659
R14305 VPWR.n1826 VPWR 0.0233659
R14306 VPWR.n1821 VPWR 0.0233659
R14307 VPWR.n1817 VPWR 0.0233659
R14308 VPWR.n1856 VPWR 0.0233659
R14309 VPWR.n992 VPWR 0.0233659
R14310 VPWR.n1518 VPWR 0.0233659
R14311 VPWR.n1164 VPWR 0.0233659
R14312 VPWR.n2469 VPWR 0.0233659
R14313 VPWR.n343 VPWR 0.0233659
R14314 VPWR.n2515 VPWR 0.0233659
R14315 VPWR.n1130 VPWR 0.0233659
R14316 VPWR.n1129 VPWR 0.0233659
R14317 VPWR.n996 VPWR 0.0233659
R14318 VPWR.n1523 VPWR 0.0233659
R14319 VPWR.n1155 VPWR 0.0233659
R14320 VPWR.n2439 VPWR 0.0233659
R14321 VPWR.n2429 VPWR 0.0233659
R14322 VPWR.n2424 VPWR 0.0233659
R14323 VPWR.n2419 VPWR 0.0233659
R14324 VPWR.n2414 VPWR 0.0233659
R14325 VPWR.n2409 VPWR 0.0233659
R14326 VPWR.n2405 VPWR 0.0233659
R14327 VPWR.n2434 VPWR 0.0233659
R14328 VPWR.n315 VPWR 0.0233659
R14329 VPWR.n2558 VPWR 0.0233659
R14330 VPWR.n1538 VPWR 0.0233659
R14331 VPWR.n1144 VPWR 0.0233659
R14332 VPWR.n1000 VPWR 0.0233659
R14333 VPWR.n1004 VPWR 0.0233659
R14334 VPWR.n1008 VPWR 0.0233659
R14335 VPWR.n1012 VPWR 0.0233659
R14336 VPWR.n1016 VPWR 0.0233659
R14337 VPWR.n1020 VPWR 0.0233659
R14338 VPWR.n1024 VPWR 0.0233659
R14339 VPWR.n968 VPWR 0.0233659
R14340 VPWR.n1473 VPWR 0.0233659
R14341 VPWR.n1590 VPWR 0.0233659
R14342 VPWR.n311 VPWR 0.0233659
R14343 VPWR.n2563 VPWR 0.0233659
R14344 VPWR.n1154 VPWR 0.0233659
R14345 VPWR.n1763 VPWR 0.0233659
R14346 VPWR.n1073 VPWR 0.0233659
R14347 VPWR.n307 VPWR 0.0233659
R14348 VPWR.n303 VPWR 0.0233659
R14349 VPWR.n295 VPWR 0.0233659
R14350 VPWR.n292 VPWR 0.0233659
R14351 VPWR.n299 VPWR 0.0233659
R14352 VPWR.n1743 VPWR 0.0233659
R14353 VPWR.n1751 VPWR 0.0233659
R14354 VPWR.n1789 VPWR 0.0233659
R14355 VPWR.n1793 VPWR 0.0233659
R14356 VPWR.n1758 VPWR 0.0233659
R14357 VPWR.n1054 VPWR 0.0233659
R14358 VPWR.n2575 VPWR 0.0233659
R14359 VPWR.n2582 VPWR 0.0233659
R14360 VPWR.n2593 VPWR 0.0233659
R14361 VPWR.n2587 VPWR 0.0233659
R14362 VPWR.n1736 VPWR 0.0233659
R14363 VPWR.n1060 VPWR 0.0233659
R14364 VPWR.n1121 VPWR 0.0233659
R14365 VPWR.n1336 VPWR 0.0226354
R14366 VPWR.n1327 VPWR 0.0226354
R14367 VPWR.n1413 VPWR 0.0226354
R14368 VPWR.n2772 VPWR 0.0226354
R14369 VPWR VPWR.n2732 0.0226354
R14370 VPWR VPWR.n2702 0.0226354
R14371 VPWR VPWR.n2664 0.0226354
R14372 VPWR VPWR.n64 0.0220517
R14373 VPWR VPWR.n67 0.0220517
R14374 VPWR VPWR.n70 0.0220517
R14375 VPWR VPWR.n73 0.0220517
R14376 VPWR VPWR.n76 0.0220517
R14377 VPWR VPWR.n79 0.0220517
R14378 VPWR VPWR.n82 0.0220517
R14379 VPWR VPWR.n85 0.0220517
R14380 VPWR VPWR.n88 0.0220517
R14381 VPWR VPWR.n91 0.0220517
R14382 VPWR VPWR.n94 0.0220517
R14383 VPWR VPWR.n97 0.0220517
R14384 VPWR.n289 VPWR 0.0220517
R14385 VPWR VPWR.n61 0.0220517
R14386 VPWR VPWR.n58 0.0220517
R14387 VPWR.n1735 VPWR 0.0220517
R14388 VPWR VPWR.n1057 0.0220517
R14389 VPWR.n1705 VPWR 0.0220517
R14390 VPWR.n1694 VPWR 0.0220517
R14391 VPWR.n1196 VPWR 0.0220517
R14392 VPWR.n1678 VPWR 0.0220517
R14393 VPWR.n1667 VPWR 0.0220517
R14394 VPWR.n1210 VPWR 0.0220517
R14395 VPWR.n1651 VPWR 0.0220517
R14396 VPWR.n1640 VPWR 0.0220517
R14397 VPWR.n1178 VPWR 0.0220517
R14398 VPWR.n1624 VPWR 0.0220517
R14399 VPWR.n1613 VPWR 0.0220517
R14400 VPWR.n1127 VPWR 0.0220517
R14401 VPWR.n1597 VPWR 0.0220517
R14402 VPWR.n1273 VPWR 0.0213333
R14403 VPWR.n1297 VPWR 0.0213333
R14404 VPWR.n1311 VPWR 0.0213333
R14405 VPWR.n1375 VPWR 0.0213333
R14406 VPWR.n1347 VPWR 0.0213333
R14407 VPWR.n1386 VPWR 0.0213333
R14408 VPWR.n1423 VPWR 0.0213333
R14409 VPWR.n2806 VPWR 0.0213333
R14410 VPWR.n2799 VPWR 0.0213333
R14411 VPWR VPWR.n2790 0.0213333
R14412 VPWR.n2792 VPWR 0.0213333
R14413 VPWR VPWR.n2770 0.0213333
R14414 VPWR VPWR.n2751 0.0213333
R14415 VPWR VPWR.n2738 0.0213333
R14416 VPWR.n2500 VPWR 0.0196917
R14417 VPWR.n24 VPWR 0.0143889
R14418 VPWR VPWR.n19 0.0099
R14419 VPWR VPWR.n1604 0.00397222
R14420 VPWR VPWR.n1105 0.00397222
R14421 VPWR VPWR.n1103 0.00397222
R14422 VPWR VPWR.n1631 0.00397222
R14423 VPWR VPWR.n1095 0.00397222
R14424 VPWR VPWR.n1093 0.00397222
R14425 VPWR VPWR.n1658 0.00397222
R14426 VPWR VPWR.n1085 0.00397222
R14427 VPWR VPWR.n1083 0.00397222
R14428 VPWR VPWR.n1685 0.00397222
R14429 VPWR VPWR.n1075 0.00397222
R14430 VPWR VPWR.n1072 0.00397222
R14431 VPWR VPWR.n1712 0.00397222
R14432 VPWR VPWR.n1724 0.00397222
R14433 VPWR.n1113 VPWR 0.00397222
R14434 VPWR VPWR.n1066 0.00397222
R14435 VPWR VPWR.n122 0.00397222
R14436 VPWR VPWR.n111 0.00397222
R14437 VPWR VPWR.n102 0.00397222
R14438 VPWR VPWR.n277 0.00397222
R14439 VPWR VPWR.n265 0.00397222
R14440 VPWR VPWR.n253 0.00397222
R14441 VPWR VPWR.n241 0.00397222
R14442 VPWR VPWR.n229 0.00397222
R14443 VPWR VPWR.n217 0.00397222
R14444 VPWR VPWR.n205 0.00397222
R14445 VPWR VPWR.n193 0.00397222
R14446 VPWR VPWR.n181 0.00397222
R14447 VPWR VPWR.n169 0.00397222
R14448 VPWR VPWR.n157 0.00397222
R14449 VPWR VPWR.n145 0.00397222
R14450 VPWR VPWR.n133 0.00397222
R14451 VPWR.n1462 VPWR.n1461 0.00351282
R14452 VPWR.n1457 VPWR.n1136 0.00351282
R14453 VPWR.n1582 VPWR.n1581 0.00351282
R14454 VPWR.n1577 VPWR.n1576 0.00351282
R14455 VPWR.n1572 VPWR.n1571 0.00351282
R14456 VPWR.n1567 VPWR.n1566 0.00351282
R14457 VPWR.n1562 VPWR.n1561 0.00351282
R14458 VPWR.n1557 VPWR.n1556 0.00351282
R14459 VPWR.n1552 VPWR.n1551 0.00351282
R14460 VPWR.n1547 VPWR.n1546 0.00351282
R14461 VPWR.n1542 VPWR.n1042 0.00351282
R14462 VPWR.n1785 VPWR.n1784 0.00351282
R14463 VPWR.n1776 VPWR.n1772 0.00351282
R14464 VPWR.n1771 VPWR.n1767 0.00351282
R14465 VPWR.n141 VPWR.n140 0.00265517
R14466 VPWR.n153 VPWR.n152 0.00265517
R14467 VPWR.n165 VPWR.n164 0.00265517
R14468 VPWR.n177 VPWR.n176 0.00265517
R14469 VPWR.n189 VPWR.n188 0.00265517
R14470 VPWR.n201 VPWR.n200 0.00265517
R14471 VPWR.n213 VPWR.n212 0.00265517
R14472 VPWR.n225 VPWR.n224 0.00265517
R14473 VPWR.n237 VPWR.n236 0.00265517
R14474 VPWR.n249 VPWR.n248 0.00265517
R14475 VPWR.n261 VPWR.n260 0.00265517
R14476 VPWR.n273 VPWR.n272 0.00265517
R14477 VPWR.n288 VPWR.n286 0.00265517
R14478 VPWR.n129 VPWR.n128 0.00265517
R14479 VPWR.n118 VPWR.n117 0.00265517
R14480 VPWR.n1734 VPWR.n1732 0.00265517
R14481 VPWR.n1720 VPWR.n1719 0.00265517
R14482 VPWR.n1708 VPWR.n1707 0.00265517
R14483 VPWR.n1697 VPWR.n1696 0.00265517
R14484 VPWR.n1195 VPWR.n1193 0.00265517
R14485 VPWR.n1681 VPWR.n1680 0.00265517
R14486 VPWR.n1670 VPWR.n1669 0.00265517
R14487 VPWR.n1209 VPWR.n1207 0.00265517
R14488 VPWR.n1654 VPWR.n1653 0.00265517
R14489 VPWR.n1643 VPWR.n1642 0.00265517
R14490 VPWR.n1177 VPWR.n1175 0.00265517
R14491 VPWR.n1627 VPWR.n1626 0.00265517
R14492 VPWR.n1616 VPWR.n1615 0.00265517
R14493 VPWR.n1126 VPWR.n1124 0.00265517
R14494 VPWR.n1600 VPWR.n1599 0.00265517
R14495 Iout.n1020 Iout.t21 239.927
R14496 Iout.n509 Iout.t124 239.927
R14497 Iout.n513 Iout.t11 239.927
R14498 Iout.n507 Iout.t131 239.927
R14499 Iout.n504 Iout.t126 239.927
R14500 Iout.n500 Iout.t147 239.927
R14501 Iout.n192 Iout.t236 239.927
R14502 Iout.n195 Iout.t242 239.927
R14503 Iout.n199 Iout.t95 239.927
R14504 Iout.n202 Iout.t14 239.927
R14505 Iout.n206 Iout.t99 239.927
R14506 Iout.n210 Iout.t37 239.927
R14507 Iout.n214 Iout.t34 239.927
R14508 Iout.n218 Iout.t134 239.927
R14509 Iout.n222 Iout.t127 239.927
R14510 Iout.n226 Iout.t28 239.927
R14511 Iout.n232 Iout.t84 239.927
R14512 Iout.n235 Iout.t82 239.927
R14513 Iout.n238 Iout.t220 239.927
R14514 Iout.n241 Iout.t213 239.927
R14515 Iout.n244 Iout.t216 239.927
R14516 Iout.n247 Iout.t86 239.927
R14517 Iout.n250 Iout.t238 239.927
R14518 Iout.n255 Iout.t161 239.927
R14519 Iout.n252 Iout.t45 239.927
R14520 Iout.n489 Iout.t69 239.927
R14521 Iout.n494 Iout.t192 239.927
R14522 Iout.n491 Iout.t91 239.927
R14523 Iout.n519 Iout.t83 239.927
R14524 Iout.n149 Iout.t61 239.927
R14525 Iout.n146 Iout.t105 239.927
R14526 Iout.n1010 Iout.t139 239.927
R14527 Iout.n1007 Iout.t56 239.927
R14528 Iout.n140 Iout.t63 239.927
R14529 Iout.n143 Iout.t181 239.927
R14530 Iout.n525 Iout.t146 239.927
R14531 Iout.n480 Iout.t80 239.927
R14532 Iout.n483 Iout.t55 239.927
R14533 Iout.n478 Iout.t4 239.927
R14534 Iout.n259 Iout.t203 239.927
R14535 Iout.n186 Iout.t255 239.927
R14536 Iout.n271 Iout.t130 239.927
R14537 Iout.n180 Iout.t7 239.927
R14538 Iout.n283 Iout.t42 239.927
R14539 Iout.n174 Iout.t29 239.927
R14540 Iout.n168 Iout.t6 239.927
R14541 Iout.n301 Iout.t2 239.927
R14542 Iout.n289 Iout.t102 239.927
R14543 Iout.n177 Iout.t98 239.927
R14544 Iout.n277 Iout.t19 239.927
R14545 Iout.n183 Iout.t177 239.927
R14546 Iout.n265 Iout.t41 239.927
R14547 Iout.n189 Iout.t123 239.927
R14548 Iout.n472 Iout.t219 239.927
R14549 Iout.n469 Iout.t151 239.927
R14550 Iout.n156 Iout.t253 239.927
R14551 Iout.n531 Iout.t79 239.927
R14552 Iout.n534 Iout.t113 239.927
R14553 Iout.n536 Iout.t172 239.927
R14554 Iout.n133 Iout.t145 239.927
R14555 Iout.n136 Iout.t47 239.927
R14556 Iout.n542 Iout.t233 239.927
R14557 Iout.n460 Iout.t65 239.927
R14558 Iout.n463 Iout.t16 239.927
R14559 Iout.n458 Iout.t149 239.927
R14560 Iout.n305 Iout.t136 239.927
R14561 Iout.n308 Iout.t221 239.927
R14562 Iout.n311 Iout.t81 239.927
R14563 Iout.n314 Iout.t173 239.927
R14564 Iout.n317 Iout.t77 239.927
R14565 Iout.n320 Iout.t183 239.927
R14566 Iout.n392 Iout.t23 239.927
R14567 Iout.n378 Iout.t120 239.927
R14568 Iout.n376 Iout.t153 239.927
R14569 Iout.n394 Iout.t67 239.927
R14570 Iout.n408 Iout.t150 239.927
R14571 Iout.n410 Iout.t222 239.927
R14572 Iout.n424 Iout.t191 239.927
R14573 Iout.n426 Iout.t157 239.927
R14574 Iout.n447 Iout.t169 239.927
R14575 Iout.n452 Iout.t66 239.927
R14576 Iout.n449 Iout.t251 239.927
R14577 Iout.n548 Iout.t25 239.927
R14578 Iout.n130 Iout.t194 239.927
R14579 Iout.n559 Iout.t121 239.927
R14580 Iout.n557 Iout.t223 239.927
R14581 Iout.n554 Iout.t72 239.927
R14582 Iout.n434 Iout.t187 239.927
R14583 Iout.n438 Iout.t208 239.927
R14584 Iout.n441 Iout.t162 239.927
R14585 Iout.n432 Iout.t20 239.927
R14586 Iout.n418 Iout.t109 239.927
R14587 Iout.n416 Iout.t38 239.927
R14588 Iout.n402 Iout.t68 239.927
R14589 Iout.n357 Iout.t57 239.927
R14590 Iout.n360 Iout.t160 239.927
R14591 Iout.n363 Iout.t165 239.927
R14592 Iout.n366 Iout.t245 239.927
R14593 Iout.n354 Iout.t248 239.927
R14594 Iout.n351 Iout.t143 239.927
R14595 Iout.n348 Iout.t179 239.927
R14596 Iout.n345 Iout.t33 239.927
R14597 Iout.n342 Iout.t185 239.927
R14598 Iout.n339 Iout.t115 239.927
R14599 Iout.n336 Iout.t73 239.927
R14600 Iout.n333 Iout.t180 239.927
R14601 Iout.n117 Iout.t128 239.927
R14602 Iout.n582 Iout.t50 239.927
R14603 Iout.n111 Iout.t70 239.927
R14604 Iout.n594 Iout.t218 239.927
R14605 Iout.n105 Iout.t111 239.927
R14606 Iout.n606 Iout.t85 239.927
R14607 Iout.n99 Iout.t164 239.927
R14608 Iout.n618 Iout.t119 239.927
R14609 Iout.n624 Iout.t27 239.927
R14610 Iout.n90 Iout.t199 239.927
R14611 Iout.n636 Iout.t103 239.927
R14612 Iout.n81 Iout.t51 239.927
R14613 Iout.n648 Iout.t125 239.927
R14614 Iout.n96 Iout.t43 239.927
R14615 Iout.n612 Iout.t10 239.927
R14616 Iout.n102 Iout.t40 239.927
R14617 Iout.n600 Iout.t171 239.927
R14618 Iout.n108 Iout.t158 239.927
R14619 Iout.n588 Iout.t239 239.927
R14620 Iout.n687 Iout.t237 239.927
R14621 Iout.n684 Iout.t156 239.927
R14622 Iout.n681 Iout.t64 239.927
R14623 Iout.n678 Iout.t22 239.927
R14624 Iout.n675 Iout.t226 239.927
R14625 Iout.n672 Iout.t229 239.927
R14626 Iout.n747 Iout.t230 239.927
R14627 Iout.n50 Iout.t206 239.927
R14628 Iout.n759 Iout.t167 239.927
R14629 Iout.n44 Iout.t201 239.927
R14630 Iout.n771 Iout.t89 239.927
R14631 Iout.n42 Iout.t205 239.927
R14632 Iout.n56 Iout.t53 239.927
R14633 Iout.n735 Iout.t17 239.927
R14634 Iout.n62 Iout.t108 239.927
R14635 Iout.n723 Iout.t247 239.927
R14636 Iout.n717 Iout.t231 239.927
R14637 Iout.n65 Iout.t212 239.927
R14638 Iout.n729 Iout.t243 239.927
R14639 Iout.n59 Iout.t249 239.927
R14640 Iout.n805 Iout.t154 239.927
R14641 Iout.n808 Iout.t114 239.927
R14642 Iout.n811 Iout.t202 239.927
R14643 Iout.n814 Iout.t141 239.927
R14644 Iout.n817 Iout.t15 239.927
R14645 Iout.n820 Iout.t228 239.927
R14646 Iout.n823 Iout.t235 239.927
R14647 Iout.n802 Iout.t76 239.927
R14648 Iout.n799 Iout.t100 239.927
R14649 Iout.n890 Iout.t117 239.927
R14650 Iout.n888 Iout.t112 239.927
R14651 Iout.n881 Iout.t168 239.927
R14652 Iout.n869 Iout.t52 239.927
R14653 Iout.n867 Iout.t32 239.927
R14654 Iout.n855 Iout.t178 239.927
R14655 Iout.n853 Iout.t142 239.927
R14656 Iout.n841 Iout.t174 239.927
R14657 Iout.n839 Iout.t97 239.927
R14658 Iout.n827 Iout.t182 239.927
R14659 Iout.n883 Iout.t92 239.927
R14660 Iout.n895 Iout.t204 239.927
R14661 Iout.n897 Iout.t8 239.927
R14662 Iout.n909 Iout.t170 239.927
R14663 Iout.n911 Iout.t227 239.927
R14664 Iout.n923 Iout.t0 239.927
R14665 Iout.n926 Iout.t118 239.927
R14666 Iout.n22 Iout.t224 239.927
R14667 Iout.n876 Iout.t159 239.927
R14668 Iout.n874 Iout.t200 239.927
R14669 Iout.n862 Iout.t197 239.927
R14670 Iout.n860 Iout.t54 239.927
R14671 Iout.n848 Iout.t217 239.927
R14672 Iout.n846 Iout.t232 239.927
R14673 Iout.n834 Iout.t110 239.927
R14674 Iout.n832 Iout.t244 239.927
R14675 Iout.n902 Iout.t24 239.927
R14676 Iout.n904 Iout.t198 239.927
R14677 Iout.n916 Iout.t135 239.927
R14678 Iout.n918 Iout.t246 239.927
R14679 Iout.n931 Iout.t211 239.927
R14680 Iout.n934 Iout.t78 239.927
R14681 Iout.n796 Iout.t49 239.927
R14682 Iout.n793 Iout.t195 239.927
R14683 Iout.n790 Iout.t186 239.927
R14684 Iout.n787 Iout.t39 239.927
R14685 Iout.n784 Iout.t26 239.927
R14686 Iout.n781 Iout.t215 239.927
R14687 Iout.n938 Iout.t9 239.927
R14688 Iout.n741 Iout.t94 239.927
R14689 Iout.n53 Iout.t188 239.927
R14690 Iout.n753 Iout.t31 239.927
R14691 Iout.n47 Iout.t189 239.927
R14692 Iout.n765 Iout.t62 239.927
R14693 Iout.n38 Iout.t46 239.927
R14694 Iout.n777 Iout.t129 239.927
R14695 Iout.n71 Iout.t144 239.927
R14696 Iout.n705 Iout.t152 239.927
R14697 Iout.n77 Iout.t184 239.927
R14698 Iout.n944 Iout.t3 239.927
R14699 Iout.n19 Iout.t116 239.927
R14700 Iout.n68 Iout.t210 239.927
R14701 Iout.n711 Iout.t175 239.927
R14702 Iout.n74 Iout.t166 239.927
R14703 Iout.n699 Iout.t101 239.927
R14704 Iout.n950 Iout.t104 239.927
R14705 Iout.n953 Iout.t252 239.927
R14706 Iout.n669 Iout.t138 239.927
R14707 Iout.n666 Iout.t59 239.927
R14708 Iout.n663 Iout.t35 239.927
R14709 Iout.n660 Iout.t254 239.927
R14710 Iout.n657 Iout.t241 239.927
R14711 Iout.n654 Iout.t1 239.927
R14712 Iout.n690 Iout.t75 239.927
R14713 Iout.n695 Iout.t107 239.927
R14714 Iout.n692 Iout.t193 239.927
R14715 Iout.n957 Iout.t44 239.927
R14716 Iout.n114 Iout.t163 239.927
R14717 Iout.n576 Iout.t90 239.927
R14718 Iout.n573 Iout.t88 239.927
R14719 Iout.n963 Iout.t176 239.927
R14720 Iout.n14 Iout.t132 239.927
R14721 Iout.n93 Iout.t71 239.927
R14722 Iout.n630 Iout.t36 239.927
R14723 Iout.n87 Iout.t13 239.927
R14724 Iout.n642 Iout.t122 239.927
R14725 Iout.n85 Iout.t58 239.927
R14726 Iout.n563 Iout.t106 239.927
R14727 Iout.n969 Iout.t18 239.927
R14728 Iout.n972 Iout.t5 239.927
R14729 Iout.n569 Iout.t12 239.927
R14730 Iout.n123 Iout.t148 239.927
R14731 Iout.n120 Iout.t48 239.927
R14732 Iout.n976 Iout.t140 239.927
R14733 Iout.n400 Iout.t133 239.927
R14734 Iout.n386 Iout.t155 239.927
R14735 Iout.n384 Iout.t250 239.927
R14736 Iout.n370 Iout.t240 239.927
R14737 Iout.n982 Iout.t190 239.927
R14738 Iout.n9 Iout.t196 239.927
R14739 Iout.n127 Iout.t207 239.927
R14740 Iout.n988 Iout.t30 239.927
R14741 Iout.n991 Iout.t137 239.927
R14742 Iout.n323 Iout.t209 239.927
R14743 Iout.n326 Iout.t93 239.927
R14744 Iout.n329 Iout.t74 239.927
R14745 Iout.n995 Iout.t234 239.927
R14746 Iout.n1001 Iout.t60 239.927
R14747 Iout.n4 Iout.t96 239.927
R14748 Iout.n295 Iout.t214 239.927
R14749 Iout.n172 Iout.t225 239.927
R14750 Iout.n1014 Iout.t87 239.927
R14751 Iout.n1021 Iout.n1020 7.9105
R14752 Iout.n510 Iout.n509 7.9105
R14753 Iout.n514 Iout.n513 7.9105
R14754 Iout.n508 Iout.n507 7.9105
R14755 Iout.n505 Iout.n504 7.9105
R14756 Iout.n501 Iout.n500 7.9105
R14757 Iout.n193 Iout.n192 7.9105
R14758 Iout.n196 Iout.n195 7.9105
R14759 Iout.n200 Iout.n199 7.9105
R14760 Iout.n203 Iout.n202 7.9105
R14761 Iout.n207 Iout.n206 7.9105
R14762 Iout.n211 Iout.n210 7.9105
R14763 Iout.n215 Iout.n214 7.9105
R14764 Iout.n219 Iout.n218 7.9105
R14765 Iout.n223 Iout.n222 7.9105
R14766 Iout.n227 Iout.n226 7.9105
R14767 Iout.n233 Iout.n232 7.9105
R14768 Iout.n236 Iout.n235 7.9105
R14769 Iout.n239 Iout.n238 7.9105
R14770 Iout.n242 Iout.n241 7.9105
R14771 Iout.n245 Iout.n244 7.9105
R14772 Iout.n248 Iout.n247 7.9105
R14773 Iout.n251 Iout.n250 7.9105
R14774 Iout.n256 Iout.n255 7.9105
R14775 Iout.n253 Iout.n252 7.9105
R14776 Iout.n490 Iout.n489 7.9105
R14777 Iout.n495 Iout.n494 7.9105
R14778 Iout.n492 Iout.n491 7.9105
R14779 Iout.n520 Iout.n519 7.9105
R14780 Iout.n150 Iout.n149 7.9105
R14781 Iout.n147 Iout.n146 7.9105
R14782 Iout.n1011 Iout.n1010 7.9105
R14783 Iout.n1008 Iout.n1007 7.9105
R14784 Iout.n141 Iout.n140 7.9105
R14785 Iout.n144 Iout.n143 7.9105
R14786 Iout.n526 Iout.n525 7.9105
R14787 Iout.n481 Iout.n480 7.9105
R14788 Iout.n484 Iout.n483 7.9105
R14789 Iout.n479 Iout.n478 7.9105
R14790 Iout.n260 Iout.n259 7.9105
R14791 Iout.n187 Iout.n186 7.9105
R14792 Iout.n272 Iout.n271 7.9105
R14793 Iout.n181 Iout.n180 7.9105
R14794 Iout.n284 Iout.n283 7.9105
R14795 Iout.n175 Iout.n174 7.9105
R14796 Iout.n169 Iout.n168 7.9105
R14797 Iout.n302 Iout.n301 7.9105
R14798 Iout.n290 Iout.n289 7.9105
R14799 Iout.n178 Iout.n177 7.9105
R14800 Iout.n278 Iout.n277 7.9105
R14801 Iout.n184 Iout.n183 7.9105
R14802 Iout.n266 Iout.n265 7.9105
R14803 Iout.n190 Iout.n189 7.9105
R14804 Iout.n473 Iout.n472 7.9105
R14805 Iout.n470 Iout.n469 7.9105
R14806 Iout.n157 Iout.n156 7.9105
R14807 Iout.n532 Iout.n531 7.9105
R14808 Iout.n535 Iout.n534 7.9105
R14809 Iout.n537 Iout.n536 7.9105
R14810 Iout.n134 Iout.n133 7.9105
R14811 Iout.n137 Iout.n136 7.9105
R14812 Iout.n543 Iout.n542 7.9105
R14813 Iout.n461 Iout.n460 7.9105
R14814 Iout.n464 Iout.n463 7.9105
R14815 Iout.n459 Iout.n458 7.9105
R14816 Iout.n306 Iout.n305 7.9105
R14817 Iout.n309 Iout.n308 7.9105
R14818 Iout.n312 Iout.n311 7.9105
R14819 Iout.n315 Iout.n314 7.9105
R14820 Iout.n318 Iout.n317 7.9105
R14821 Iout.n321 Iout.n320 7.9105
R14822 Iout.n393 Iout.n392 7.9105
R14823 Iout.n379 Iout.n378 7.9105
R14824 Iout.n377 Iout.n376 7.9105
R14825 Iout.n395 Iout.n394 7.9105
R14826 Iout.n409 Iout.n408 7.9105
R14827 Iout.n411 Iout.n410 7.9105
R14828 Iout.n425 Iout.n424 7.9105
R14829 Iout.n427 Iout.n426 7.9105
R14830 Iout.n448 Iout.n447 7.9105
R14831 Iout.n453 Iout.n452 7.9105
R14832 Iout.n450 Iout.n449 7.9105
R14833 Iout.n549 Iout.n548 7.9105
R14834 Iout.n131 Iout.n130 7.9105
R14835 Iout.n560 Iout.n559 7.9105
R14836 Iout.n558 Iout.n557 7.9105
R14837 Iout.n555 Iout.n554 7.9105
R14838 Iout.n435 Iout.n434 7.9105
R14839 Iout.n439 Iout.n438 7.9105
R14840 Iout.n442 Iout.n441 7.9105
R14841 Iout.n433 Iout.n432 7.9105
R14842 Iout.n419 Iout.n418 7.9105
R14843 Iout.n417 Iout.n416 7.9105
R14844 Iout.n403 Iout.n402 7.9105
R14845 Iout.n358 Iout.n357 7.9105
R14846 Iout.n361 Iout.n360 7.9105
R14847 Iout.n364 Iout.n363 7.9105
R14848 Iout.n367 Iout.n366 7.9105
R14849 Iout.n355 Iout.n354 7.9105
R14850 Iout.n352 Iout.n351 7.9105
R14851 Iout.n349 Iout.n348 7.9105
R14852 Iout.n346 Iout.n345 7.9105
R14853 Iout.n343 Iout.n342 7.9105
R14854 Iout.n340 Iout.n339 7.9105
R14855 Iout.n337 Iout.n336 7.9105
R14856 Iout.n334 Iout.n333 7.9105
R14857 Iout.n118 Iout.n117 7.9105
R14858 Iout.n583 Iout.n582 7.9105
R14859 Iout.n112 Iout.n111 7.9105
R14860 Iout.n595 Iout.n594 7.9105
R14861 Iout.n106 Iout.n105 7.9105
R14862 Iout.n607 Iout.n606 7.9105
R14863 Iout.n100 Iout.n99 7.9105
R14864 Iout.n619 Iout.n618 7.9105
R14865 Iout.n625 Iout.n624 7.9105
R14866 Iout.n91 Iout.n90 7.9105
R14867 Iout.n637 Iout.n636 7.9105
R14868 Iout.n82 Iout.n81 7.9105
R14869 Iout.n649 Iout.n648 7.9105
R14870 Iout.n97 Iout.n96 7.9105
R14871 Iout.n613 Iout.n612 7.9105
R14872 Iout.n103 Iout.n102 7.9105
R14873 Iout.n601 Iout.n600 7.9105
R14874 Iout.n109 Iout.n108 7.9105
R14875 Iout.n589 Iout.n588 7.9105
R14876 Iout.n688 Iout.n687 7.9105
R14877 Iout.n685 Iout.n684 7.9105
R14878 Iout.n682 Iout.n681 7.9105
R14879 Iout.n679 Iout.n678 7.9105
R14880 Iout.n676 Iout.n675 7.9105
R14881 Iout.n673 Iout.n672 7.9105
R14882 Iout.n748 Iout.n747 7.9105
R14883 Iout.n51 Iout.n50 7.9105
R14884 Iout.n760 Iout.n759 7.9105
R14885 Iout.n45 Iout.n44 7.9105
R14886 Iout.n772 Iout.n771 7.9105
R14887 Iout.n43 Iout.n42 7.9105
R14888 Iout.n57 Iout.n56 7.9105
R14889 Iout.n736 Iout.n735 7.9105
R14890 Iout.n63 Iout.n62 7.9105
R14891 Iout.n724 Iout.n723 7.9105
R14892 Iout.n718 Iout.n717 7.9105
R14893 Iout.n66 Iout.n65 7.9105
R14894 Iout.n730 Iout.n729 7.9105
R14895 Iout.n60 Iout.n59 7.9105
R14896 Iout.n806 Iout.n805 7.9105
R14897 Iout.n809 Iout.n808 7.9105
R14898 Iout.n812 Iout.n811 7.9105
R14899 Iout.n815 Iout.n814 7.9105
R14900 Iout.n818 Iout.n817 7.9105
R14901 Iout.n821 Iout.n820 7.9105
R14902 Iout.n824 Iout.n823 7.9105
R14903 Iout.n803 Iout.n802 7.9105
R14904 Iout.n800 Iout.n799 7.9105
R14905 Iout.n891 Iout.n890 7.9105
R14906 Iout.n889 Iout.n888 7.9105
R14907 Iout.n882 Iout.n881 7.9105
R14908 Iout.n870 Iout.n869 7.9105
R14909 Iout.n868 Iout.n867 7.9105
R14910 Iout.n856 Iout.n855 7.9105
R14911 Iout.n854 Iout.n853 7.9105
R14912 Iout.n842 Iout.n841 7.9105
R14913 Iout.n840 Iout.n839 7.9105
R14914 Iout.n828 Iout.n827 7.9105
R14915 Iout.n884 Iout.n883 7.9105
R14916 Iout.n896 Iout.n895 7.9105
R14917 Iout.n898 Iout.n897 7.9105
R14918 Iout.n910 Iout.n909 7.9105
R14919 Iout.n912 Iout.n911 7.9105
R14920 Iout.n924 Iout.n923 7.9105
R14921 Iout.n927 Iout.n926 7.9105
R14922 Iout.n23 Iout.n22 7.9105
R14923 Iout.n877 Iout.n876 7.9105
R14924 Iout.n875 Iout.n874 7.9105
R14925 Iout.n863 Iout.n862 7.9105
R14926 Iout.n861 Iout.n860 7.9105
R14927 Iout.n849 Iout.n848 7.9105
R14928 Iout.n847 Iout.n846 7.9105
R14929 Iout.n835 Iout.n834 7.9105
R14930 Iout.n833 Iout.n832 7.9105
R14931 Iout.n903 Iout.n902 7.9105
R14932 Iout.n905 Iout.n904 7.9105
R14933 Iout.n917 Iout.n916 7.9105
R14934 Iout.n919 Iout.n918 7.9105
R14935 Iout.n932 Iout.n931 7.9105
R14936 Iout.n935 Iout.n934 7.9105
R14937 Iout.n797 Iout.n796 7.9105
R14938 Iout.n794 Iout.n793 7.9105
R14939 Iout.n791 Iout.n790 7.9105
R14940 Iout.n788 Iout.n787 7.9105
R14941 Iout.n785 Iout.n784 7.9105
R14942 Iout.n782 Iout.n781 7.9105
R14943 Iout.n939 Iout.n938 7.9105
R14944 Iout.n742 Iout.n741 7.9105
R14945 Iout.n54 Iout.n53 7.9105
R14946 Iout.n754 Iout.n753 7.9105
R14947 Iout.n48 Iout.n47 7.9105
R14948 Iout.n766 Iout.n765 7.9105
R14949 Iout.n39 Iout.n38 7.9105
R14950 Iout.n778 Iout.n777 7.9105
R14951 Iout.n72 Iout.n71 7.9105
R14952 Iout.n706 Iout.n705 7.9105
R14953 Iout.n78 Iout.n77 7.9105
R14954 Iout.n945 Iout.n944 7.9105
R14955 Iout.n20 Iout.n19 7.9105
R14956 Iout.n69 Iout.n68 7.9105
R14957 Iout.n712 Iout.n711 7.9105
R14958 Iout.n75 Iout.n74 7.9105
R14959 Iout.n700 Iout.n699 7.9105
R14960 Iout.n951 Iout.n950 7.9105
R14961 Iout.n954 Iout.n953 7.9105
R14962 Iout.n670 Iout.n669 7.9105
R14963 Iout.n667 Iout.n666 7.9105
R14964 Iout.n664 Iout.n663 7.9105
R14965 Iout.n661 Iout.n660 7.9105
R14966 Iout.n658 Iout.n657 7.9105
R14967 Iout.n655 Iout.n654 7.9105
R14968 Iout.n691 Iout.n690 7.9105
R14969 Iout.n696 Iout.n695 7.9105
R14970 Iout.n693 Iout.n692 7.9105
R14971 Iout.n958 Iout.n957 7.9105
R14972 Iout.n115 Iout.n114 7.9105
R14973 Iout.n577 Iout.n576 7.9105
R14974 Iout.n574 Iout.n573 7.9105
R14975 Iout.n964 Iout.n963 7.9105
R14976 Iout.n15 Iout.n14 7.9105
R14977 Iout.n94 Iout.n93 7.9105
R14978 Iout.n631 Iout.n630 7.9105
R14979 Iout.n88 Iout.n87 7.9105
R14980 Iout.n643 Iout.n642 7.9105
R14981 Iout.n86 Iout.n85 7.9105
R14982 Iout.n564 Iout.n563 7.9105
R14983 Iout.n970 Iout.n969 7.9105
R14984 Iout.n973 Iout.n972 7.9105
R14985 Iout.n570 Iout.n569 7.9105
R14986 Iout.n124 Iout.n123 7.9105
R14987 Iout.n121 Iout.n120 7.9105
R14988 Iout.n977 Iout.n976 7.9105
R14989 Iout.n401 Iout.n400 7.9105
R14990 Iout.n387 Iout.n386 7.9105
R14991 Iout.n385 Iout.n384 7.9105
R14992 Iout.n371 Iout.n370 7.9105
R14993 Iout.n983 Iout.n982 7.9105
R14994 Iout.n10 Iout.n9 7.9105
R14995 Iout.n128 Iout.n127 7.9105
R14996 Iout.n989 Iout.n988 7.9105
R14997 Iout.n992 Iout.n991 7.9105
R14998 Iout.n324 Iout.n323 7.9105
R14999 Iout.n327 Iout.n326 7.9105
R15000 Iout.n330 Iout.n329 7.9105
R15001 Iout.n996 Iout.n995 7.9105
R15002 Iout.n1002 Iout.n1001 7.9105
R15003 Iout.n5 Iout.n4 7.9105
R15004 Iout.n296 Iout.n295 7.9105
R15005 Iout.n173 Iout.n172 7.9105
R15006 Iout.n1015 Iout.n1014 7.9105
R15007 Iout.n886 Iout.n885 3.86101
R15008 Iout.n880 Iout.n879 3.86101
R15009 Iout.n894 Iout.n893 3.86101
R15010 Iout.n872 Iout.n871 3.86101
R15011 Iout.n900 Iout.n899 3.86101
R15012 Iout.n866 Iout.n865 3.86101
R15013 Iout.n908 Iout.n907 3.86101
R15014 Iout.n858 Iout.n857 3.86101
R15015 Iout.n914 Iout.n913 3.86101
R15016 Iout.n852 Iout.n851 3.86101
R15017 Iout.n922 Iout.n921 3.86101
R15018 Iout.n844 Iout.n843 3.86101
R15019 Iout.n929 Iout.n928 3.86101
R15020 Iout.n838 Iout.n837 3.86101
R15021 Iout.n925 Iout.n21 3.86101
R15022 Iout.n830 Iout.n829 3.86101
R15023 Iout.n879 Iout.n878 3.4105
R15024 Iout.n887 Iout.n886 3.4105
R15025 Iout.n893 Iout.n892 3.4105
R15026 Iout.n798 Iout.n28 3.4105
R15027 Iout.n801 Iout.n29 3.4105
R15028 Iout.n804 Iout.n30 3.4105
R15029 Iout.n807 Iout.n31 3.4105
R15030 Iout.n873 Iout.n872 3.4105
R15031 Iout.n744 Iout.n743 3.4105
R15032 Iout.n740 Iout.n739 3.4105
R15033 Iout.n732 Iout.n731 3.4105
R15034 Iout.n728 Iout.n727 3.4105
R15035 Iout.n720 Iout.n719 3.4105
R15036 Iout.n795 Iout.n27 3.4105
R15037 Iout.n901 Iout.n900 3.4105
R15038 Iout.n722 Iout.n721 3.4105
R15039 Iout.n726 Iout.n725 3.4105
R15040 Iout.n734 Iout.n733 3.4105
R15041 Iout.n738 Iout.n737 3.4105
R15042 Iout.n746 Iout.n745 3.4105
R15043 Iout.n750 Iout.n749 3.4105
R15044 Iout.n752 Iout.n751 3.4105
R15045 Iout.n810 Iout.n32 3.4105
R15046 Iout.n865 Iout.n864 3.4105
R15047 Iout.n668 Iout.n55 3.4105
R15048 Iout.n671 Iout.n58 3.4105
R15049 Iout.n674 Iout.n61 3.4105
R15050 Iout.n677 Iout.n64 3.4105
R15051 Iout.n680 Iout.n67 3.4105
R15052 Iout.n683 Iout.n70 3.4105
R15053 Iout.n686 Iout.n73 3.4105
R15054 Iout.n714 Iout.n713 3.4105
R15055 Iout.n716 Iout.n715 3.4105
R15056 Iout.n792 Iout.n26 3.4105
R15057 Iout.n907 Iout.n906 3.4105
R15058 Iout.n587 Iout.n586 3.4105
R15059 Iout.n591 Iout.n590 3.4105
R15060 Iout.n599 Iout.n598 3.4105
R15061 Iout.n603 Iout.n602 3.4105
R15062 Iout.n611 Iout.n610 3.4105
R15063 Iout.n615 Iout.n614 3.4105
R15064 Iout.n623 Iout.n622 3.4105
R15065 Iout.n627 Iout.n626 3.4105
R15066 Iout.n665 Iout.n52 3.4105
R15067 Iout.n758 Iout.n757 3.4105
R15068 Iout.n756 Iout.n755 3.4105
R15069 Iout.n813 Iout.n33 3.4105
R15070 Iout.n859 Iout.n858 3.4105
R15071 Iout.n629 Iout.n628 3.4105
R15072 Iout.n621 Iout.n620 3.4105
R15073 Iout.n617 Iout.n616 3.4105
R15074 Iout.n609 Iout.n608 3.4105
R15075 Iout.n605 Iout.n604 3.4105
R15076 Iout.n597 Iout.n596 3.4105
R15077 Iout.n593 Iout.n592 3.4105
R15078 Iout.n585 Iout.n584 3.4105
R15079 Iout.n581 Iout.n580 3.4105
R15080 Iout.n579 Iout.n578 3.4105
R15081 Iout.n689 Iout.n76 3.4105
R15082 Iout.n710 Iout.n709 3.4105
R15083 Iout.n708 Iout.n707 3.4105
R15084 Iout.n789 Iout.n25 3.4105
R15085 Iout.n915 Iout.n914 3.4105
R15086 Iout.n572 Iout.n571 3.4105
R15087 Iout.n335 Iout.n116 3.4105
R15088 Iout.n338 Iout.n113 3.4105
R15089 Iout.n341 Iout.n110 3.4105
R15090 Iout.n344 Iout.n107 3.4105
R15091 Iout.n347 Iout.n104 3.4105
R15092 Iout.n350 Iout.n101 3.4105
R15093 Iout.n353 Iout.n98 3.4105
R15094 Iout.n356 Iout.n95 3.4105
R15095 Iout.n359 Iout.n92 3.4105
R15096 Iout.n633 Iout.n632 3.4105
R15097 Iout.n635 Iout.n634 3.4105
R15098 Iout.n662 Iout.n49 3.4105
R15099 Iout.n762 Iout.n761 3.4105
R15100 Iout.n764 Iout.n763 3.4105
R15101 Iout.n816 Iout.n34 3.4105
R15102 Iout.n851 Iout.n850 3.4105
R15103 Iout.n399 Iout.n398 3.4105
R15104 Iout.n405 Iout.n404 3.4105
R15105 Iout.n415 Iout.n414 3.4105
R15106 Iout.n421 Iout.n420 3.4105
R15107 Iout.n431 Iout.n430 3.4105
R15108 Iout.n444 Iout.n443 3.4105
R15109 Iout.n440 Iout.n159 3.4105
R15110 Iout.n437 Iout.n436 3.4105
R15111 Iout.n553 Iout.n552 3.4105
R15112 Iout.n556 Iout.n119 3.4105
R15113 Iout.n562 Iout.n561 3.4105
R15114 Iout.n568 Iout.n567 3.4105
R15115 Iout.n566 Iout.n565 3.4105
R15116 Iout.n575 Iout.n79 3.4105
R15117 Iout.n698 Iout.n697 3.4105
R15118 Iout.n702 Iout.n701 3.4105
R15119 Iout.n704 Iout.n703 3.4105
R15120 Iout.n786 Iout.n24 3.4105
R15121 Iout.n921 Iout.n920 3.4105
R15122 Iout.n129 Iout.n125 3.4105
R15123 Iout.n547 Iout.n546 3.4105
R15124 Iout.n551 Iout.n550 3.4105
R15125 Iout.n451 Iout.n158 3.4105
R15126 Iout.n455 Iout.n454 3.4105
R15127 Iout.n446 Iout.n445 3.4105
R15128 Iout.n429 Iout.n428 3.4105
R15129 Iout.n423 Iout.n422 3.4105
R15130 Iout.n413 Iout.n412 3.4105
R15131 Iout.n407 Iout.n406 3.4105
R15132 Iout.n397 Iout.n396 3.4105
R15133 Iout.n391 Iout.n390 3.4105
R15134 Iout.n389 Iout.n388 3.4105
R15135 Iout.n362 Iout.n89 3.4105
R15136 Iout.n641 Iout.n640 3.4105
R15137 Iout.n639 Iout.n638 3.4105
R15138 Iout.n659 Iout.n46 3.4105
R15139 Iout.n770 Iout.n769 3.4105
R15140 Iout.n768 Iout.n767 3.4105
R15141 Iout.n819 Iout.n35 3.4105
R15142 Iout.n845 Iout.n844 3.4105
R15143 Iout.n325 Iout.n165 3.4105
R15144 Iout.n322 Iout.n164 3.4105
R15145 Iout.n319 Iout.n163 3.4105
R15146 Iout.n316 Iout.n162 3.4105
R15147 Iout.n313 Iout.n161 3.4105
R15148 Iout.n310 Iout.n160 3.4105
R15149 Iout.n307 Iout.n155 3.4105
R15150 Iout.n457 Iout.n456 3.4105
R15151 Iout.n466 Iout.n465 3.4105
R15152 Iout.n462 Iout.n126 3.4105
R15153 Iout.n545 Iout.n544 3.4105
R15154 Iout.n541 Iout.n540 3.4105
R15155 Iout.n135 Iout.n3 3.4105
R15156 Iout.n987 Iout.n986 3.4105
R15157 Iout.n985 Iout.n984 3.4105
R15158 Iout.n122 Iout.n8 3.4105
R15159 Iout.n968 Iout.n967 3.4105
R15160 Iout.n966 Iout.n965 3.4105
R15161 Iout.n694 Iout.n13 3.4105
R15162 Iout.n949 Iout.n948 3.4105
R15163 Iout.n947 Iout.n946 3.4105
R15164 Iout.n783 Iout.n18 3.4105
R15165 Iout.n930 Iout.n929 3.4105
R15166 Iout.n1004 Iout.n1003 3.4105
R15167 Iout.n539 Iout.n538 3.4105
R15168 Iout.n533 Iout.n132 3.4105
R15169 Iout.n530 Iout.n529 3.4105
R15170 Iout.n468 Iout.n467 3.4105
R15171 Iout.n471 Iout.n153 3.4105
R15172 Iout.n475 Iout.n474 3.4105
R15173 Iout.n264 Iout.n263 3.4105
R15174 Iout.n268 Iout.n267 3.4105
R15175 Iout.n276 Iout.n275 3.4105
R15176 Iout.n280 Iout.n279 3.4105
R15177 Iout.n288 Iout.n287 3.4105
R15178 Iout.n292 Iout.n291 3.4105
R15179 Iout.n300 Iout.n299 3.4105
R15180 Iout.n328 Iout.n166 3.4105
R15181 Iout.n381 Iout.n380 3.4105
R15182 Iout.n383 Iout.n382 3.4105
R15183 Iout.n365 Iout.n83 3.4105
R15184 Iout.n645 Iout.n644 3.4105
R15185 Iout.n647 Iout.n646 3.4105
R15186 Iout.n656 Iout.n40 3.4105
R15187 Iout.n774 Iout.n773 3.4105
R15188 Iout.n776 Iout.n775 3.4105
R15189 Iout.n822 Iout.n36 3.4105
R15190 Iout.n837 Iout.n836 3.4105
R15191 Iout.n298 Iout.n297 3.4105
R15192 Iout.n294 Iout.n293 3.4105
R15193 Iout.n286 Iout.n285 3.4105
R15194 Iout.n282 Iout.n281 3.4105
R15195 Iout.n274 Iout.n273 3.4105
R15196 Iout.n270 Iout.n269 3.4105
R15197 Iout.n262 Iout.n261 3.4105
R15198 Iout.n477 Iout.n476 3.4105
R15199 Iout.n486 Iout.n485 3.4105
R15200 Iout.n482 Iout.n151 3.4105
R15201 Iout.n528 Iout.n527 3.4105
R15202 Iout.n524 Iout.n523 3.4105
R15203 Iout.n142 Iout.n138 3.4105
R15204 Iout.n1006 Iout.n1005 3.4105
R15205 Iout.n1009 Iout.n0 3.4105
R15206 Iout.n1000 Iout.n999 3.4105
R15207 Iout.n998 Iout.n997 3.4105
R15208 Iout.n990 Iout.n6 3.4105
R15209 Iout.n981 Iout.n980 3.4105
R15210 Iout.n979 Iout.n978 3.4105
R15211 Iout.n971 Iout.n11 3.4105
R15212 Iout.n962 Iout.n961 3.4105
R15213 Iout.n960 Iout.n959 3.4105
R15214 Iout.n952 Iout.n16 3.4105
R15215 Iout.n943 Iout.n942 3.4105
R15216 Iout.n941 Iout.n940 3.4105
R15217 Iout.n933 Iout.n21 3.4105
R15218 Iout.n1017 Iout.n1016 3.4105
R15219 Iout.n148 Iout.n2 3.4105
R15220 Iout.n518 Iout.n517 3.4105
R15221 Iout.n522 Iout.n521 3.4105
R15222 Iout.n493 Iout.n139 3.4105
R15223 Iout.n497 Iout.n496 3.4105
R15224 Iout.n488 Iout.n487 3.4105
R15225 Iout.n254 Iout.n154 3.4105
R15226 Iout.n258 Iout.n257 3.4105
R15227 Iout.n249 Iout.n188 3.4105
R15228 Iout.n246 Iout.n185 3.4105
R15229 Iout.n243 Iout.n182 3.4105
R15230 Iout.n240 Iout.n179 3.4105
R15231 Iout.n237 Iout.n176 3.4105
R15232 Iout.n234 Iout.n170 3.4105
R15233 Iout.n231 Iout.n230 3.4105
R15234 Iout.n171 Iout.n167 3.4105
R15235 Iout.n304 Iout.n303 3.4105
R15236 Iout.n332 Iout.n331 3.4105
R15237 Iout.n375 Iout.n374 3.4105
R15238 Iout.n373 Iout.n372 3.4105
R15239 Iout.n369 Iout.n368 3.4105
R15240 Iout.n84 Iout.n80 3.4105
R15241 Iout.n651 Iout.n650 3.4105
R15242 Iout.n653 Iout.n652 3.4105
R15243 Iout.n41 Iout.n37 3.4105
R15244 Iout.n780 Iout.n779 3.4105
R15245 Iout.n826 Iout.n825 3.4105
R15246 Iout.n831 Iout.n830 3.4105
R15247 Iout.n229 Iout.n228 3.4105
R15248 Iout.n225 Iout.n224 3.4105
R15249 Iout.n221 Iout.n220 3.4105
R15250 Iout.n217 Iout.n216 3.4105
R15251 Iout.n213 Iout.n212 3.4105
R15252 Iout.n209 Iout.n208 3.4105
R15253 Iout.n205 Iout.n204 3.4105
R15254 Iout.n201 Iout.n191 3.4105
R15255 Iout.n198 Iout.n197 3.4105
R15256 Iout.n194 Iout.n152 3.4105
R15257 Iout.n499 Iout.n498 3.4105
R15258 Iout.n503 Iout.n502 3.4105
R15259 Iout.n506 Iout.n145 3.4105
R15260 Iout.n516 Iout.n515 3.4105
R15261 Iout.n512 Iout.n511 3.4105
R15262 Iout.n1019 Iout.n1018 3.4105
R15263 Iout.n936 Iout.n23 1.43848
R15264 Iout.n936 Iout.n935 1.34612
R15265 Iout.n939 Iout.n937 1.34612
R15266 Iout.n20 Iout.n17 1.34612
R15267 Iout.n955 Iout.n954 1.34612
R15268 Iout.n958 Iout.n956 1.34612
R15269 Iout.n15 Iout.n12 1.34612
R15270 Iout.n974 Iout.n973 1.34612
R15271 Iout.n977 Iout.n975 1.34612
R15272 Iout.n10 Iout.n7 1.34612
R15273 Iout.n993 Iout.n992 1.34612
R15274 Iout.n996 Iout.n994 1.34612
R15275 Iout.n5 Iout.n1 1.34612
R15276 Iout.n1012 Iout.n1011 1.34612
R15277 Iout.n1015 Iout.n1013 1.34612
R15278 Iout.n1022 Iout.n1021 1.34612
R15279 Iout.n197 Iout.n154 0.451012
R15280 Iout.n476 Iout.n154 0.451012
R15281 Iout.n476 Iout.n475 0.451012
R15282 Iout.n475 Iout.n155 0.451012
R15283 Iout.n445 Iout.n155 0.451012
R15284 Iout.n445 Iout.n444 0.451012
R15285 Iout.n444 Iout.n107 0.451012
R15286 Iout.n604 Iout.n107 0.451012
R15287 Iout.n604 Iout.n603 0.451012
R15288 Iout.n603 Iout.n64 0.451012
R15289 Iout.n733 Iout.n64 0.451012
R15290 Iout.n733 Iout.n732 0.451012
R15291 Iout.n732 Iout.n29 0.451012
R15292 Iout.n886 Iout.n29 0.451012
R15293 Iout.n258 Iout.n191 0.451012
R15294 Iout.n262 Iout.n258 0.451012
R15295 Iout.n263 Iout.n262 0.451012
R15296 Iout.n263 Iout.n160 0.451012
R15297 Iout.n429 Iout.n160 0.451012
R15298 Iout.n430 Iout.n429 0.451012
R15299 Iout.n430 Iout.n104 0.451012
R15300 Iout.n609 Iout.n104 0.451012
R15301 Iout.n610 Iout.n609 0.451012
R15302 Iout.n610 Iout.n61 0.451012
R15303 Iout.n738 Iout.n61 0.451012
R15304 Iout.n739 Iout.n738 0.451012
R15305 Iout.n739 Iout.n30 0.451012
R15306 Iout.n879 Iout.n30 0.451012
R15307 Iout.n487 Iout.n152 0.451012
R15308 Iout.n487 Iout.n486 0.451012
R15309 Iout.n486 Iout.n153 0.451012
R15310 Iout.n456 Iout.n153 0.451012
R15311 Iout.n456 Iout.n455 0.451012
R15312 Iout.n455 Iout.n159 0.451012
R15313 Iout.n159 Iout.n110 0.451012
R15314 Iout.n597 Iout.n110 0.451012
R15315 Iout.n598 Iout.n597 0.451012
R15316 Iout.n598 Iout.n67 0.451012
R15317 Iout.n726 Iout.n67 0.451012
R15318 Iout.n727 Iout.n726 0.451012
R15319 Iout.n727 Iout.n28 0.451012
R15320 Iout.n893 Iout.n28 0.451012
R15321 Iout.n204 Iout.n188 0.451012
R15322 Iout.n269 Iout.n188 0.451012
R15323 Iout.n269 Iout.n268 0.451012
R15324 Iout.n268 Iout.n161 0.451012
R15325 Iout.n422 Iout.n161 0.451012
R15326 Iout.n422 Iout.n421 0.451012
R15327 Iout.n421 Iout.n101 0.451012
R15328 Iout.n616 Iout.n101 0.451012
R15329 Iout.n616 Iout.n615 0.451012
R15330 Iout.n615 Iout.n58 0.451012
R15331 Iout.n745 Iout.n58 0.451012
R15332 Iout.n745 Iout.n744 0.451012
R15333 Iout.n744 Iout.n31 0.451012
R15334 Iout.n872 Iout.n31 0.451012
R15335 Iout.n498 Iout.n497 0.451012
R15336 Iout.n497 Iout.n151 0.451012
R15337 Iout.n467 Iout.n151 0.451012
R15338 Iout.n467 Iout.n466 0.451012
R15339 Iout.n466 Iout.n158 0.451012
R15340 Iout.n436 Iout.n158 0.451012
R15341 Iout.n436 Iout.n113 0.451012
R15342 Iout.n592 Iout.n113 0.451012
R15343 Iout.n592 Iout.n591 0.451012
R15344 Iout.n591 Iout.n70 0.451012
R15345 Iout.n721 Iout.n70 0.451012
R15346 Iout.n721 Iout.n720 0.451012
R15347 Iout.n720 Iout.n27 0.451012
R15348 Iout.n900 Iout.n27 0.451012
R15349 Iout.n208 Iout.n185 0.451012
R15350 Iout.n274 Iout.n185 0.451012
R15351 Iout.n275 Iout.n274 0.451012
R15352 Iout.n275 Iout.n162 0.451012
R15353 Iout.n413 Iout.n162 0.451012
R15354 Iout.n414 Iout.n413 0.451012
R15355 Iout.n414 Iout.n98 0.451012
R15356 Iout.n621 Iout.n98 0.451012
R15357 Iout.n622 Iout.n621 0.451012
R15358 Iout.n622 Iout.n55 0.451012
R15359 Iout.n750 Iout.n55 0.451012
R15360 Iout.n751 Iout.n750 0.451012
R15361 Iout.n751 Iout.n32 0.451012
R15362 Iout.n865 Iout.n32 0.451012
R15363 Iout.n502 Iout.n139 0.451012
R15364 Iout.n528 Iout.n139 0.451012
R15365 Iout.n529 Iout.n528 0.451012
R15366 Iout.n529 Iout.n126 0.451012
R15367 Iout.n551 Iout.n126 0.451012
R15368 Iout.n552 Iout.n551 0.451012
R15369 Iout.n552 Iout.n116 0.451012
R15370 Iout.n585 Iout.n116 0.451012
R15371 Iout.n586 Iout.n585 0.451012
R15372 Iout.n586 Iout.n73 0.451012
R15373 Iout.n714 Iout.n73 0.451012
R15374 Iout.n715 Iout.n714 0.451012
R15375 Iout.n715 Iout.n26 0.451012
R15376 Iout.n907 Iout.n26 0.451012
R15377 Iout.n212 Iout.n182 0.451012
R15378 Iout.n281 Iout.n182 0.451012
R15379 Iout.n281 Iout.n280 0.451012
R15380 Iout.n280 Iout.n163 0.451012
R15381 Iout.n406 Iout.n163 0.451012
R15382 Iout.n406 Iout.n405 0.451012
R15383 Iout.n405 Iout.n95 0.451012
R15384 Iout.n628 Iout.n95 0.451012
R15385 Iout.n628 Iout.n627 0.451012
R15386 Iout.n627 Iout.n52 0.451012
R15387 Iout.n757 Iout.n52 0.451012
R15388 Iout.n757 Iout.n756 0.451012
R15389 Iout.n756 Iout.n33 0.451012
R15390 Iout.n858 Iout.n33 0.451012
R15391 Iout.n522 Iout.n145 0.451012
R15392 Iout.n523 Iout.n522 0.451012
R15393 Iout.n523 Iout.n132 0.451012
R15394 Iout.n545 Iout.n132 0.451012
R15395 Iout.n546 Iout.n545 0.451012
R15396 Iout.n546 Iout.n119 0.451012
R15397 Iout.n572 Iout.n119 0.451012
R15398 Iout.n580 Iout.n572 0.451012
R15399 Iout.n580 Iout.n579 0.451012
R15400 Iout.n579 Iout.n76 0.451012
R15401 Iout.n709 Iout.n76 0.451012
R15402 Iout.n709 Iout.n708 0.451012
R15403 Iout.n708 Iout.n25 0.451012
R15404 Iout.n914 Iout.n25 0.451012
R15405 Iout.n216 Iout.n179 0.451012
R15406 Iout.n286 Iout.n179 0.451012
R15407 Iout.n287 Iout.n286 0.451012
R15408 Iout.n287 Iout.n164 0.451012
R15409 Iout.n397 Iout.n164 0.451012
R15410 Iout.n398 Iout.n397 0.451012
R15411 Iout.n398 Iout.n92 0.451012
R15412 Iout.n633 Iout.n92 0.451012
R15413 Iout.n634 Iout.n633 0.451012
R15414 Iout.n634 Iout.n49 0.451012
R15415 Iout.n762 Iout.n49 0.451012
R15416 Iout.n763 Iout.n762 0.451012
R15417 Iout.n763 Iout.n34 0.451012
R15418 Iout.n851 Iout.n34 0.451012
R15419 Iout.n517 Iout.n516 0.451012
R15420 Iout.n517 Iout.n138 0.451012
R15421 Iout.n539 Iout.n138 0.451012
R15422 Iout.n540 Iout.n539 0.451012
R15423 Iout.n540 Iout.n125 0.451012
R15424 Iout.n562 Iout.n125 0.451012
R15425 Iout.n567 Iout.n562 0.451012
R15426 Iout.n567 Iout.n566 0.451012
R15427 Iout.n566 Iout.n79 0.451012
R15428 Iout.n698 Iout.n79 0.451012
R15429 Iout.n702 Iout.n698 0.451012
R15430 Iout.n703 Iout.n702 0.451012
R15431 Iout.n703 Iout.n24 0.451012
R15432 Iout.n921 Iout.n24 0.451012
R15433 Iout.n220 Iout.n176 0.451012
R15434 Iout.n293 Iout.n176 0.451012
R15435 Iout.n293 Iout.n292 0.451012
R15436 Iout.n292 Iout.n165 0.451012
R15437 Iout.n390 Iout.n165 0.451012
R15438 Iout.n390 Iout.n389 0.451012
R15439 Iout.n389 Iout.n89 0.451012
R15440 Iout.n640 Iout.n89 0.451012
R15441 Iout.n640 Iout.n639 0.451012
R15442 Iout.n639 Iout.n46 0.451012
R15443 Iout.n769 Iout.n46 0.451012
R15444 Iout.n769 Iout.n768 0.451012
R15445 Iout.n768 Iout.n35 0.451012
R15446 Iout.n844 Iout.n35 0.451012
R15447 Iout.n511 Iout.n2 0.451012
R15448 Iout.n1005 Iout.n2 0.451012
R15449 Iout.n1005 Iout.n1004 0.451012
R15450 Iout.n1004 Iout.n3 0.451012
R15451 Iout.n986 Iout.n3 0.451012
R15452 Iout.n986 Iout.n985 0.451012
R15453 Iout.n985 Iout.n8 0.451012
R15454 Iout.n967 Iout.n8 0.451012
R15455 Iout.n967 Iout.n966 0.451012
R15456 Iout.n966 Iout.n13 0.451012
R15457 Iout.n948 Iout.n13 0.451012
R15458 Iout.n948 Iout.n947 0.451012
R15459 Iout.n947 Iout.n18 0.451012
R15460 Iout.n929 Iout.n18 0.451012
R15461 Iout.n224 Iout.n170 0.451012
R15462 Iout.n298 Iout.n170 0.451012
R15463 Iout.n299 Iout.n298 0.451012
R15464 Iout.n299 Iout.n166 0.451012
R15465 Iout.n381 Iout.n166 0.451012
R15466 Iout.n382 Iout.n381 0.451012
R15467 Iout.n382 Iout.n83 0.451012
R15468 Iout.n645 Iout.n83 0.451012
R15469 Iout.n646 Iout.n645 0.451012
R15470 Iout.n646 Iout.n40 0.451012
R15471 Iout.n774 Iout.n40 0.451012
R15472 Iout.n775 Iout.n774 0.451012
R15473 Iout.n775 Iout.n36 0.451012
R15474 Iout.n837 Iout.n36 0.451012
R15475 Iout.n1018 Iout.n1017 0.451012
R15476 Iout.n1017 Iout.n0 0.451012
R15477 Iout.n999 Iout.n0 0.451012
R15478 Iout.n999 Iout.n998 0.451012
R15479 Iout.n998 Iout.n6 0.451012
R15480 Iout.n980 Iout.n6 0.451012
R15481 Iout.n980 Iout.n979 0.451012
R15482 Iout.n979 Iout.n11 0.451012
R15483 Iout.n961 Iout.n11 0.451012
R15484 Iout.n961 Iout.n960 0.451012
R15485 Iout.n960 Iout.n16 0.451012
R15486 Iout.n942 Iout.n16 0.451012
R15487 Iout.n942 Iout.n941 0.451012
R15488 Iout.n941 Iout.n21 0.451012
R15489 Iout.n230 Iout.n229 0.451012
R15490 Iout.n230 Iout.n167 0.451012
R15491 Iout.n304 Iout.n167 0.451012
R15492 Iout.n332 Iout.n304 0.451012
R15493 Iout.n374 Iout.n332 0.451012
R15494 Iout.n374 Iout.n373 0.451012
R15495 Iout.n373 Iout.n369 0.451012
R15496 Iout.n369 Iout.n80 0.451012
R15497 Iout.n651 Iout.n80 0.451012
R15498 Iout.n652 Iout.n651 0.451012
R15499 Iout.n652 Iout.n37 0.451012
R15500 Iout.n780 Iout.n37 0.451012
R15501 Iout.n826 Iout.n780 0.451012
R15502 Iout.n830 Iout.n826 0.451012
R15503 Iout.n231 Iout 0.2919
R15504 Iout.n303 Iout 0.2919
R15505 Iout Iout.n300 0.2919
R15506 Iout.n375 Iout 0.2919
R15507 Iout.n380 Iout 0.2919
R15508 Iout.n391 Iout 0.2919
R15509 Iout.n368 Iout 0.2919
R15510 Iout Iout.n365 0.2919
R15511 Iout Iout.n362 0.2919
R15512 Iout Iout.n359 0.2919
R15513 Iout.n650 Iout 0.2919
R15514 Iout Iout.n647 0.2919
R15515 Iout.n638 Iout 0.2919
R15516 Iout Iout.n635 0.2919
R15517 Iout.n626 Iout 0.2919
R15518 Iout.n41 Iout 0.2919
R15519 Iout.n773 Iout 0.2919
R15520 Iout Iout.n770 0.2919
R15521 Iout.n761 Iout 0.2919
R15522 Iout Iout.n758 0.2919
R15523 Iout.n749 Iout 0.2919
R15524 Iout.n825 Iout 0.2919
R15525 Iout Iout.n822 0.2919
R15526 Iout Iout.n819 0.2919
R15527 Iout Iout.n816 0.2919
R15528 Iout Iout.n813 0.2919
R15529 Iout Iout.n810 0.2919
R15530 Iout Iout.n807 0.2919
R15531 Iout.n829 Iout 0.2919
R15532 Iout.n838 Iout 0.2919
R15533 Iout.n843 Iout 0.2919
R15534 Iout.n852 Iout 0.2919
R15535 Iout.n857 Iout 0.2919
R15536 Iout.n866 Iout 0.2919
R15537 Iout.n871 Iout 0.2919
R15538 Iout.n880 Iout 0.2919
R15539 Iout Iout.n925 0.2919
R15540 Iout.n928 Iout 0.2919
R15541 Iout.n922 Iout 0.2919
R15542 Iout.n913 Iout 0.2919
R15543 Iout.n908 Iout 0.2919
R15544 Iout.n899 Iout 0.2919
R15545 Iout.n894 Iout 0.2919
R15546 Iout.n885 Iout 0.2919
R15547 Iout.n831 Iout 0.2919
R15548 Iout.n836 Iout 0.2919
R15549 Iout.n845 Iout 0.2919
R15550 Iout.n850 Iout 0.2919
R15551 Iout.n859 Iout 0.2919
R15552 Iout.n864 Iout 0.2919
R15553 Iout.n873 Iout 0.2919
R15554 Iout.n878 Iout 0.2919
R15555 Iout.n887 Iout 0.2919
R15556 Iout.n892 Iout 0.2919
R15557 Iout.n933 Iout 0.2919
R15558 Iout.n930 Iout 0.2919
R15559 Iout.n920 Iout 0.2919
R15560 Iout.n915 Iout 0.2919
R15561 Iout.n906 Iout 0.2919
R15562 Iout.n901 Iout 0.2919
R15563 Iout.n940 Iout 0.2919
R15564 Iout Iout.n783 0.2919
R15565 Iout Iout.n786 0.2919
R15566 Iout Iout.n789 0.2919
R15567 Iout Iout.n792 0.2919
R15568 Iout Iout.n795 0.2919
R15569 Iout Iout.n798 0.2919
R15570 Iout Iout.n801 0.2919
R15571 Iout Iout.n804 0.2919
R15572 Iout.n779 Iout 0.2919
R15573 Iout Iout.n776 0.2919
R15574 Iout.n767 Iout 0.2919
R15575 Iout Iout.n764 0.2919
R15576 Iout.n755 Iout 0.2919
R15577 Iout Iout.n752 0.2919
R15578 Iout.n743 Iout 0.2919
R15579 Iout Iout.n740 0.2919
R15580 Iout.n731 Iout 0.2919
R15581 Iout Iout.n728 0.2919
R15582 Iout.n719 Iout 0.2919
R15583 Iout Iout.n943 0.2919
R15584 Iout.n946 Iout 0.2919
R15585 Iout Iout.n704 0.2919
R15586 Iout.n707 Iout 0.2919
R15587 Iout Iout.n716 0.2919
R15588 Iout.n952 Iout 0.2919
R15589 Iout.n949 Iout 0.2919
R15590 Iout.n701 Iout 0.2919
R15591 Iout Iout.n710 0.2919
R15592 Iout.n713 Iout 0.2919
R15593 Iout Iout.n722 0.2919
R15594 Iout.n725 Iout 0.2919
R15595 Iout Iout.n734 0.2919
R15596 Iout.n737 Iout 0.2919
R15597 Iout Iout.n746 0.2919
R15598 Iout.n653 Iout 0.2919
R15599 Iout.n656 Iout 0.2919
R15600 Iout.n659 Iout 0.2919
R15601 Iout.n662 Iout 0.2919
R15602 Iout.n665 Iout 0.2919
R15603 Iout.n668 Iout 0.2919
R15604 Iout.n671 Iout 0.2919
R15605 Iout.n674 Iout 0.2919
R15606 Iout.n677 Iout 0.2919
R15607 Iout.n680 Iout 0.2919
R15608 Iout.n683 Iout 0.2919
R15609 Iout.n686 Iout 0.2919
R15610 Iout.n959 Iout 0.2919
R15611 Iout Iout.n694 0.2919
R15612 Iout.n697 Iout 0.2919
R15613 Iout.n689 Iout 0.2919
R15614 Iout Iout.n962 0.2919
R15615 Iout.n965 Iout 0.2919
R15616 Iout Iout.n575 0.2919
R15617 Iout.n578 Iout 0.2919
R15618 Iout Iout.n587 0.2919
R15619 Iout.n590 Iout 0.2919
R15620 Iout Iout.n599 0.2919
R15621 Iout.n602 Iout 0.2919
R15622 Iout Iout.n611 0.2919
R15623 Iout.n614 Iout 0.2919
R15624 Iout Iout.n623 0.2919
R15625 Iout.n84 Iout 0.2919
R15626 Iout.n644 Iout 0.2919
R15627 Iout Iout.n641 0.2919
R15628 Iout.n632 Iout 0.2919
R15629 Iout Iout.n629 0.2919
R15630 Iout.n620 Iout 0.2919
R15631 Iout Iout.n617 0.2919
R15632 Iout.n608 Iout 0.2919
R15633 Iout Iout.n605 0.2919
R15634 Iout.n596 Iout 0.2919
R15635 Iout Iout.n593 0.2919
R15636 Iout.n584 Iout 0.2919
R15637 Iout Iout.n581 0.2919
R15638 Iout.n971 Iout 0.2919
R15639 Iout.n968 Iout 0.2919
R15640 Iout.n565 Iout 0.2919
R15641 Iout.n978 Iout 0.2919
R15642 Iout Iout.n122 0.2919
R15643 Iout Iout.n568 0.2919
R15644 Iout.n571 Iout 0.2919
R15645 Iout Iout.n335 0.2919
R15646 Iout Iout.n338 0.2919
R15647 Iout Iout.n341 0.2919
R15648 Iout Iout.n344 0.2919
R15649 Iout Iout.n347 0.2919
R15650 Iout Iout.n350 0.2919
R15651 Iout Iout.n353 0.2919
R15652 Iout Iout.n356 0.2919
R15653 Iout.n372 Iout 0.2919
R15654 Iout.n383 Iout 0.2919
R15655 Iout.n388 Iout 0.2919
R15656 Iout.n399 Iout 0.2919
R15657 Iout.n404 Iout 0.2919
R15658 Iout.n415 Iout 0.2919
R15659 Iout.n420 Iout 0.2919
R15660 Iout.n431 Iout 0.2919
R15661 Iout.n443 Iout 0.2919
R15662 Iout Iout.n440 0.2919
R15663 Iout Iout.n437 0.2919
R15664 Iout.n553 Iout 0.2919
R15665 Iout.n556 Iout 0.2919
R15666 Iout.n561 Iout 0.2919
R15667 Iout Iout.n981 0.2919
R15668 Iout.n984 Iout 0.2919
R15669 Iout.n990 Iout 0.2919
R15670 Iout.n987 Iout 0.2919
R15671 Iout Iout.n129 0.2919
R15672 Iout Iout.n547 0.2919
R15673 Iout.n550 Iout 0.2919
R15674 Iout Iout.n451 0.2919
R15675 Iout.n454 Iout 0.2919
R15676 Iout.n446 Iout 0.2919
R15677 Iout.n428 Iout 0.2919
R15678 Iout.n423 Iout 0.2919
R15679 Iout.n412 Iout 0.2919
R15680 Iout.n407 Iout 0.2919
R15681 Iout.n396 Iout 0.2919
R15682 Iout.n331 Iout 0.2919
R15683 Iout Iout.n328 0.2919
R15684 Iout Iout.n325 0.2919
R15685 Iout Iout.n322 0.2919
R15686 Iout Iout.n319 0.2919
R15687 Iout Iout.n316 0.2919
R15688 Iout Iout.n313 0.2919
R15689 Iout Iout.n310 0.2919
R15690 Iout Iout.n307 0.2919
R15691 Iout.n457 Iout 0.2919
R15692 Iout.n465 Iout 0.2919
R15693 Iout Iout.n462 0.2919
R15694 Iout.n544 Iout 0.2919
R15695 Iout Iout.n541 0.2919
R15696 Iout Iout.n135 0.2919
R15697 Iout.n997 Iout 0.2919
R15698 Iout Iout.n1000 0.2919
R15699 Iout.n1003 Iout 0.2919
R15700 Iout.n538 Iout 0.2919
R15701 Iout.n533 Iout 0.2919
R15702 Iout.n530 Iout 0.2919
R15703 Iout Iout.n468 0.2919
R15704 Iout Iout.n471 0.2919
R15705 Iout.n474 Iout 0.2919
R15706 Iout Iout.n264 0.2919
R15707 Iout.n267 Iout 0.2919
R15708 Iout Iout.n276 0.2919
R15709 Iout.n279 Iout 0.2919
R15710 Iout Iout.n288 0.2919
R15711 Iout.n291 Iout 0.2919
R15712 Iout.n171 Iout 0.2919
R15713 Iout.n297 Iout 0.2919
R15714 Iout Iout.n294 0.2919
R15715 Iout.n285 Iout 0.2919
R15716 Iout Iout.n282 0.2919
R15717 Iout.n273 Iout 0.2919
R15718 Iout Iout.n270 0.2919
R15719 Iout.n261 Iout 0.2919
R15720 Iout.n477 Iout 0.2919
R15721 Iout.n485 Iout 0.2919
R15722 Iout Iout.n482 0.2919
R15723 Iout.n527 Iout 0.2919
R15724 Iout Iout.n524 0.2919
R15725 Iout Iout.n142 0.2919
R15726 Iout.n1006 Iout 0.2919
R15727 Iout.n1009 Iout 0.2919
R15728 Iout.n1016 Iout 0.2919
R15729 Iout Iout.n148 0.2919
R15730 Iout Iout.n518 0.2919
R15731 Iout.n521 Iout 0.2919
R15732 Iout Iout.n493 0.2919
R15733 Iout.n496 Iout 0.2919
R15734 Iout.n488 Iout 0.2919
R15735 Iout Iout.n254 0.2919
R15736 Iout.n257 Iout 0.2919
R15737 Iout.n249 Iout 0.2919
R15738 Iout.n246 Iout 0.2919
R15739 Iout.n243 Iout 0.2919
R15740 Iout.n240 Iout 0.2919
R15741 Iout.n237 Iout 0.2919
R15742 Iout.n234 Iout 0.2919
R15743 Iout.n228 Iout 0.2919
R15744 Iout Iout.n225 0.2919
R15745 Iout Iout.n221 0.2919
R15746 Iout Iout.n217 0.2919
R15747 Iout Iout.n213 0.2919
R15748 Iout Iout.n209 0.2919
R15749 Iout Iout.n205 0.2919
R15750 Iout Iout.n201 0.2919
R15751 Iout Iout.n198 0.2919
R15752 Iout Iout.n194 0.2919
R15753 Iout.n499 Iout 0.2919
R15754 Iout.n503 Iout 0.2919
R15755 Iout.n506 Iout 0.2919
R15756 Iout.n515 Iout 0.2919
R15757 Iout Iout.n512 0.2919
R15758 Iout.n1019 Iout 0.2919
R15759 Iout.n1013 Iout.n1012 0.092855
R15760 Iout.n1012 Iout.n1 0.092855
R15761 Iout.n994 Iout.n1 0.092855
R15762 Iout.n994 Iout.n993 0.092855
R15763 Iout.n993 Iout.n7 0.092855
R15764 Iout.n975 Iout.n7 0.092855
R15765 Iout.n975 Iout.n974 0.092855
R15766 Iout.n974 Iout.n12 0.092855
R15767 Iout.n956 Iout.n12 0.092855
R15768 Iout.n956 Iout.n955 0.092855
R15769 Iout.n955 Iout.n17 0.092855
R15770 Iout.n937 Iout.n17 0.092855
R15771 Iout.n937 Iout.n936 0.092855
R15772 Iout.n197 Iout 0.0818902
R15773 Iout.n191 Iout 0.0818902
R15774 Iout.n152 Iout 0.0818902
R15775 Iout.n204 Iout 0.0818902
R15776 Iout.n498 Iout 0.0818902
R15777 Iout.n208 Iout 0.0818902
R15778 Iout.n502 Iout 0.0818902
R15779 Iout.n212 Iout 0.0818902
R15780 Iout.n145 Iout 0.0818902
R15781 Iout.n216 Iout 0.0818902
R15782 Iout.n516 Iout 0.0818902
R15783 Iout.n220 Iout 0.0818902
R15784 Iout.n511 Iout 0.0818902
R15785 Iout.n224 Iout 0.0818902
R15786 Iout.n1018 Iout 0.0818902
R15787 Iout.n229 Iout 0.0818902
R15788 Iout.n1013 Iout 0.072645
R15789 Iout.n302 Iout 0.0532071
R15790 Iout Iout.n377 0.0532071
R15791 Iout.n379 Iout 0.0532071
R15792 Iout.n367 Iout 0.0532071
R15793 Iout.n364 Iout 0.0532071
R15794 Iout.n361 Iout 0.0532071
R15795 Iout.n649 Iout 0.0532071
R15796 Iout Iout.n82 0.0532071
R15797 Iout.n637 Iout 0.0532071
R15798 Iout Iout.n91 0.0532071
R15799 Iout Iout.n43 0.0532071
R15800 Iout.n772 Iout 0.0532071
R15801 Iout Iout.n45 0.0532071
R15802 Iout.n760 Iout 0.0532071
R15803 Iout Iout.n51 0.0532071
R15804 Iout.n824 Iout 0.0532071
R15805 Iout.n821 Iout 0.0532071
R15806 Iout.n818 Iout 0.0532071
R15807 Iout.n815 Iout 0.0532071
R15808 Iout.n812 Iout 0.0532071
R15809 Iout.n809 Iout 0.0532071
R15810 Iout.n828 Iout 0.0532071
R15811 Iout Iout.n840 0.0532071
R15812 Iout.n842 Iout 0.0532071
R15813 Iout Iout.n854 0.0532071
R15814 Iout.n856 Iout 0.0532071
R15815 Iout Iout.n868 0.0532071
R15816 Iout.n870 Iout 0.0532071
R15817 Iout.n927 Iout 0.0532071
R15818 Iout Iout.n924 0.0532071
R15819 Iout.n912 Iout 0.0532071
R15820 Iout Iout.n910 0.0532071
R15821 Iout.n898 Iout 0.0532071
R15822 Iout Iout.n896 0.0532071
R15823 Iout.n884 Iout 0.0532071
R15824 Iout Iout.n882 0.0532071
R15825 Iout Iout.n833 0.0532071
R15826 Iout.n835 Iout 0.0532071
R15827 Iout Iout.n847 0.0532071
R15828 Iout.n849 Iout 0.0532071
R15829 Iout Iout.n861 0.0532071
R15830 Iout.n863 Iout 0.0532071
R15831 Iout Iout.n875 0.0532071
R15832 Iout.n877 Iout 0.0532071
R15833 Iout Iout.n889 0.0532071
R15834 Iout Iout.n932 0.0532071
R15835 Iout.n919 Iout 0.0532071
R15836 Iout Iout.n917 0.0532071
R15837 Iout.n905 Iout 0.0532071
R15838 Iout Iout.n903 0.0532071
R15839 Iout.n891 Iout 0.0532071
R15840 Iout.n782 Iout 0.0532071
R15841 Iout.n785 Iout 0.0532071
R15842 Iout.n788 Iout 0.0532071
R15843 Iout.n791 Iout 0.0532071
R15844 Iout.n794 Iout 0.0532071
R15845 Iout.n797 Iout 0.0532071
R15846 Iout.n800 Iout 0.0532071
R15847 Iout.n803 Iout 0.0532071
R15848 Iout.n806 Iout 0.0532071
R15849 Iout.n778 Iout 0.0532071
R15850 Iout Iout.n39 0.0532071
R15851 Iout.n766 Iout 0.0532071
R15852 Iout Iout.n48 0.0532071
R15853 Iout.n754 Iout 0.0532071
R15854 Iout Iout.n54 0.0532071
R15855 Iout.n742 Iout 0.0532071
R15856 Iout Iout.n60 0.0532071
R15857 Iout.n730 Iout 0.0532071
R15858 Iout Iout.n66 0.0532071
R15859 Iout.n945 Iout 0.0532071
R15860 Iout.n78 Iout 0.0532071
R15861 Iout.n706 Iout 0.0532071
R15862 Iout Iout.n72 0.0532071
R15863 Iout.n718 Iout 0.0532071
R15864 Iout Iout.n951 0.0532071
R15865 Iout.n700 Iout 0.0532071
R15866 Iout Iout.n75 0.0532071
R15867 Iout.n712 Iout 0.0532071
R15868 Iout Iout.n69 0.0532071
R15869 Iout.n724 Iout 0.0532071
R15870 Iout Iout.n63 0.0532071
R15871 Iout.n736 Iout 0.0532071
R15872 Iout Iout.n57 0.0532071
R15873 Iout.n748 Iout 0.0532071
R15874 Iout Iout.n655 0.0532071
R15875 Iout Iout.n658 0.0532071
R15876 Iout Iout.n661 0.0532071
R15877 Iout Iout.n664 0.0532071
R15878 Iout Iout.n667 0.0532071
R15879 Iout Iout.n670 0.0532071
R15880 Iout Iout.n673 0.0532071
R15881 Iout Iout.n676 0.0532071
R15882 Iout Iout.n679 0.0532071
R15883 Iout Iout.n682 0.0532071
R15884 Iout Iout.n685 0.0532071
R15885 Iout.n693 Iout 0.0532071
R15886 Iout.n696 Iout 0.0532071
R15887 Iout Iout.n691 0.0532071
R15888 Iout Iout.n688 0.0532071
R15889 Iout.n964 Iout 0.0532071
R15890 Iout.n574 Iout 0.0532071
R15891 Iout.n577 Iout 0.0532071
R15892 Iout Iout.n115 0.0532071
R15893 Iout.n589 Iout 0.0532071
R15894 Iout Iout.n109 0.0532071
R15895 Iout.n601 Iout 0.0532071
R15896 Iout Iout.n103 0.0532071
R15897 Iout.n613 Iout 0.0532071
R15898 Iout Iout.n97 0.0532071
R15899 Iout.n625 Iout 0.0532071
R15900 Iout Iout.n86 0.0532071
R15901 Iout.n643 Iout 0.0532071
R15902 Iout Iout.n88 0.0532071
R15903 Iout.n631 Iout 0.0532071
R15904 Iout Iout.n94 0.0532071
R15905 Iout.n619 Iout 0.0532071
R15906 Iout Iout.n100 0.0532071
R15907 Iout.n607 Iout 0.0532071
R15908 Iout Iout.n106 0.0532071
R15909 Iout.n595 Iout 0.0532071
R15910 Iout Iout.n112 0.0532071
R15911 Iout.n583 Iout 0.0532071
R15912 Iout Iout.n970 0.0532071
R15913 Iout.n564 Iout 0.0532071
R15914 Iout Iout.n118 0.0532071
R15915 Iout.n121 Iout 0.0532071
R15916 Iout.n124 Iout 0.0532071
R15917 Iout.n570 Iout 0.0532071
R15918 Iout.n334 Iout 0.0532071
R15919 Iout.n337 Iout 0.0532071
R15920 Iout.n340 Iout 0.0532071
R15921 Iout.n343 Iout 0.0532071
R15922 Iout.n346 Iout 0.0532071
R15923 Iout.n349 Iout 0.0532071
R15924 Iout.n352 Iout 0.0532071
R15925 Iout.n355 Iout 0.0532071
R15926 Iout.n358 Iout 0.0532071
R15927 Iout.n371 Iout 0.0532071
R15928 Iout Iout.n385 0.0532071
R15929 Iout.n387 Iout 0.0532071
R15930 Iout Iout.n401 0.0532071
R15931 Iout.n403 Iout 0.0532071
R15932 Iout Iout.n417 0.0532071
R15933 Iout.n419 Iout 0.0532071
R15934 Iout Iout.n433 0.0532071
R15935 Iout.n442 Iout 0.0532071
R15936 Iout.n439 Iout 0.0532071
R15937 Iout.n435 Iout 0.0532071
R15938 Iout Iout.n555 0.0532071
R15939 Iout Iout.n558 0.0532071
R15940 Iout.n983 Iout 0.0532071
R15941 Iout.n560 Iout 0.0532071
R15942 Iout Iout.n989 0.0532071
R15943 Iout.n128 Iout 0.0532071
R15944 Iout.n131 Iout 0.0532071
R15945 Iout.n549 Iout 0.0532071
R15946 Iout.n450 Iout 0.0532071
R15947 Iout.n453 Iout 0.0532071
R15948 Iout Iout.n448 0.0532071
R15949 Iout.n427 Iout 0.0532071
R15950 Iout Iout.n425 0.0532071
R15951 Iout.n411 Iout 0.0532071
R15952 Iout Iout.n409 0.0532071
R15953 Iout.n395 Iout 0.0532071
R15954 Iout Iout.n393 0.0532071
R15955 Iout.n330 Iout 0.0532071
R15956 Iout.n327 Iout 0.0532071
R15957 Iout.n324 Iout 0.0532071
R15958 Iout.n321 Iout 0.0532071
R15959 Iout.n318 Iout 0.0532071
R15960 Iout.n315 Iout 0.0532071
R15961 Iout.n312 Iout 0.0532071
R15962 Iout.n309 Iout 0.0532071
R15963 Iout.n306 Iout 0.0532071
R15964 Iout Iout.n459 0.0532071
R15965 Iout.n464 Iout 0.0532071
R15966 Iout.n461 Iout 0.0532071
R15967 Iout.n543 Iout 0.0532071
R15968 Iout.n137 Iout 0.0532071
R15969 Iout.n134 Iout 0.0532071
R15970 Iout.n1002 Iout 0.0532071
R15971 Iout.n537 Iout 0.0532071
R15972 Iout Iout.n535 0.0532071
R15973 Iout Iout.n532 0.0532071
R15974 Iout.n157 Iout 0.0532071
R15975 Iout.n470 Iout 0.0532071
R15976 Iout.n473 Iout 0.0532071
R15977 Iout.n190 Iout 0.0532071
R15978 Iout.n266 Iout 0.0532071
R15979 Iout Iout.n184 0.0532071
R15980 Iout.n278 Iout 0.0532071
R15981 Iout Iout.n178 0.0532071
R15982 Iout.n290 Iout 0.0532071
R15983 Iout Iout.n169 0.0532071
R15984 Iout Iout.n173 0.0532071
R15985 Iout.n296 Iout 0.0532071
R15986 Iout Iout.n175 0.0532071
R15987 Iout.n284 Iout 0.0532071
R15988 Iout Iout.n181 0.0532071
R15989 Iout.n272 Iout 0.0532071
R15990 Iout Iout.n187 0.0532071
R15991 Iout.n260 Iout 0.0532071
R15992 Iout Iout.n479 0.0532071
R15993 Iout.n484 Iout 0.0532071
R15994 Iout.n481 Iout 0.0532071
R15995 Iout.n526 Iout 0.0532071
R15996 Iout.n144 Iout 0.0532071
R15997 Iout.n141 Iout 0.0532071
R15998 Iout Iout.n1008 0.0532071
R15999 Iout.n147 Iout 0.0532071
R16000 Iout.n150 Iout 0.0532071
R16001 Iout.n520 Iout 0.0532071
R16002 Iout.n492 Iout 0.0532071
R16003 Iout.n495 Iout 0.0532071
R16004 Iout Iout.n490 0.0532071
R16005 Iout.n253 Iout 0.0532071
R16006 Iout.n256 Iout 0.0532071
R16007 Iout Iout.n251 0.0532071
R16008 Iout Iout.n248 0.0532071
R16009 Iout Iout.n245 0.0532071
R16010 Iout Iout.n242 0.0532071
R16011 Iout Iout.n239 0.0532071
R16012 Iout Iout.n236 0.0532071
R16013 Iout Iout.n233 0.0532071
R16014 Iout.n227 Iout 0.0532071
R16015 Iout.n223 Iout 0.0532071
R16016 Iout.n219 Iout 0.0532071
R16017 Iout.n215 Iout 0.0532071
R16018 Iout.n211 Iout 0.0532071
R16019 Iout.n207 Iout 0.0532071
R16020 Iout.n203 Iout 0.0532071
R16021 Iout.n200 Iout 0.0532071
R16022 Iout.n196 Iout 0.0532071
R16023 Iout.n193 Iout 0.0532071
R16024 Iout Iout.n501 0.0532071
R16025 Iout Iout.n505 0.0532071
R16026 Iout Iout.n508 0.0532071
R16027 Iout.n514 Iout 0.0532071
R16028 Iout.n510 Iout 0.0532071
R16029 Iout.n1020 Iout 0.03925
R16030 Iout.n509 Iout 0.03925
R16031 Iout.n513 Iout 0.03925
R16032 Iout.n507 Iout 0.03925
R16033 Iout.n504 Iout 0.03925
R16034 Iout.n500 Iout 0.03925
R16035 Iout.n192 Iout 0.03925
R16036 Iout.n195 Iout 0.03925
R16037 Iout.n199 Iout 0.03925
R16038 Iout.n202 Iout 0.03925
R16039 Iout.n206 Iout 0.03925
R16040 Iout.n210 Iout 0.03925
R16041 Iout.n214 Iout 0.03925
R16042 Iout.n218 Iout 0.03925
R16043 Iout.n222 Iout 0.03925
R16044 Iout.n226 Iout 0.03925
R16045 Iout.n232 Iout 0.03925
R16046 Iout.n235 Iout 0.03925
R16047 Iout.n238 Iout 0.03925
R16048 Iout.n241 Iout 0.03925
R16049 Iout.n244 Iout 0.03925
R16050 Iout.n247 Iout 0.03925
R16051 Iout.n250 Iout 0.03925
R16052 Iout.n255 Iout 0.03925
R16053 Iout.n252 Iout 0.03925
R16054 Iout.n489 Iout 0.03925
R16055 Iout.n494 Iout 0.03925
R16056 Iout.n491 Iout 0.03925
R16057 Iout.n519 Iout 0.03925
R16058 Iout.n149 Iout 0.03925
R16059 Iout.n146 Iout 0.03925
R16060 Iout.n1010 Iout 0.03925
R16061 Iout.n1007 Iout 0.03925
R16062 Iout.n140 Iout 0.03925
R16063 Iout.n143 Iout 0.03925
R16064 Iout.n525 Iout 0.03925
R16065 Iout.n480 Iout 0.03925
R16066 Iout.n483 Iout 0.03925
R16067 Iout.n478 Iout 0.03925
R16068 Iout.n259 Iout 0.03925
R16069 Iout.n186 Iout 0.03925
R16070 Iout.n271 Iout 0.03925
R16071 Iout.n180 Iout 0.03925
R16072 Iout.n283 Iout 0.03925
R16073 Iout.n174 Iout 0.03925
R16074 Iout.n168 Iout 0.03925
R16075 Iout.n301 Iout 0.03925
R16076 Iout.n289 Iout 0.03925
R16077 Iout.n177 Iout 0.03925
R16078 Iout.n277 Iout 0.03925
R16079 Iout.n183 Iout 0.03925
R16080 Iout.n265 Iout 0.03925
R16081 Iout.n189 Iout 0.03925
R16082 Iout.n472 Iout 0.03925
R16083 Iout.n469 Iout 0.03925
R16084 Iout.n156 Iout 0.03925
R16085 Iout.n531 Iout 0.03925
R16086 Iout.n534 Iout 0.03925
R16087 Iout.n536 Iout 0.03925
R16088 Iout.n133 Iout 0.03925
R16089 Iout.n136 Iout 0.03925
R16090 Iout.n542 Iout 0.03925
R16091 Iout.n460 Iout 0.03925
R16092 Iout.n463 Iout 0.03925
R16093 Iout.n458 Iout 0.03925
R16094 Iout.n305 Iout 0.03925
R16095 Iout.n308 Iout 0.03925
R16096 Iout.n311 Iout 0.03925
R16097 Iout.n314 Iout 0.03925
R16098 Iout.n317 Iout 0.03925
R16099 Iout.n320 Iout 0.03925
R16100 Iout.n392 Iout 0.03925
R16101 Iout.n378 Iout 0.03925
R16102 Iout.n376 Iout 0.03925
R16103 Iout.n394 Iout 0.03925
R16104 Iout.n408 Iout 0.03925
R16105 Iout.n410 Iout 0.03925
R16106 Iout.n424 Iout 0.03925
R16107 Iout.n426 Iout 0.03925
R16108 Iout.n447 Iout 0.03925
R16109 Iout.n452 Iout 0.03925
R16110 Iout.n449 Iout 0.03925
R16111 Iout.n548 Iout 0.03925
R16112 Iout.n130 Iout 0.03925
R16113 Iout.n559 Iout 0.03925
R16114 Iout.n557 Iout 0.03925
R16115 Iout.n554 Iout 0.03925
R16116 Iout.n434 Iout 0.03925
R16117 Iout.n438 Iout 0.03925
R16118 Iout.n441 Iout 0.03925
R16119 Iout.n432 Iout 0.03925
R16120 Iout.n418 Iout 0.03925
R16121 Iout.n416 Iout 0.03925
R16122 Iout.n402 Iout 0.03925
R16123 Iout.n357 Iout 0.03925
R16124 Iout.n360 Iout 0.03925
R16125 Iout.n363 Iout 0.03925
R16126 Iout.n366 Iout 0.03925
R16127 Iout.n354 Iout 0.03925
R16128 Iout.n351 Iout 0.03925
R16129 Iout.n348 Iout 0.03925
R16130 Iout.n345 Iout 0.03925
R16131 Iout.n342 Iout 0.03925
R16132 Iout.n339 Iout 0.03925
R16133 Iout.n336 Iout 0.03925
R16134 Iout.n333 Iout 0.03925
R16135 Iout.n117 Iout 0.03925
R16136 Iout.n582 Iout 0.03925
R16137 Iout.n111 Iout 0.03925
R16138 Iout.n594 Iout 0.03925
R16139 Iout.n105 Iout 0.03925
R16140 Iout.n606 Iout 0.03925
R16141 Iout.n99 Iout 0.03925
R16142 Iout.n618 Iout 0.03925
R16143 Iout.n624 Iout 0.03925
R16144 Iout.n90 Iout 0.03925
R16145 Iout.n636 Iout 0.03925
R16146 Iout.n81 Iout 0.03925
R16147 Iout.n648 Iout 0.03925
R16148 Iout.n96 Iout 0.03925
R16149 Iout.n612 Iout 0.03925
R16150 Iout.n102 Iout 0.03925
R16151 Iout.n600 Iout 0.03925
R16152 Iout.n108 Iout 0.03925
R16153 Iout.n588 Iout 0.03925
R16154 Iout.n687 Iout 0.03925
R16155 Iout.n684 Iout 0.03925
R16156 Iout.n681 Iout 0.03925
R16157 Iout.n678 Iout 0.03925
R16158 Iout.n675 Iout 0.03925
R16159 Iout.n672 Iout 0.03925
R16160 Iout.n747 Iout 0.03925
R16161 Iout.n50 Iout 0.03925
R16162 Iout.n759 Iout 0.03925
R16163 Iout.n44 Iout 0.03925
R16164 Iout.n771 Iout 0.03925
R16165 Iout.n42 Iout 0.03925
R16166 Iout.n56 Iout 0.03925
R16167 Iout.n735 Iout 0.03925
R16168 Iout.n62 Iout 0.03925
R16169 Iout.n723 Iout 0.03925
R16170 Iout.n717 Iout 0.03925
R16171 Iout.n65 Iout 0.03925
R16172 Iout.n729 Iout 0.03925
R16173 Iout.n59 Iout 0.03925
R16174 Iout.n805 Iout 0.03925
R16175 Iout.n808 Iout 0.03925
R16176 Iout.n811 Iout 0.03925
R16177 Iout.n814 Iout 0.03925
R16178 Iout.n817 Iout 0.03925
R16179 Iout.n820 Iout 0.03925
R16180 Iout.n823 Iout 0.03925
R16181 Iout.n802 Iout 0.03925
R16182 Iout.n799 Iout 0.03925
R16183 Iout.n890 Iout 0.03925
R16184 Iout.n888 Iout 0.03925
R16185 Iout.n881 Iout 0.03925
R16186 Iout.n869 Iout 0.03925
R16187 Iout.n867 Iout 0.03925
R16188 Iout.n855 Iout 0.03925
R16189 Iout.n853 Iout 0.03925
R16190 Iout.n841 Iout 0.03925
R16191 Iout.n839 Iout 0.03925
R16192 Iout.n827 Iout 0.03925
R16193 Iout.n883 Iout 0.03925
R16194 Iout.n895 Iout 0.03925
R16195 Iout.n897 Iout 0.03925
R16196 Iout.n909 Iout 0.03925
R16197 Iout.n911 Iout 0.03925
R16198 Iout.n923 Iout 0.03925
R16199 Iout.n926 Iout 0.03925
R16200 Iout.n22 Iout 0.03925
R16201 Iout.n876 Iout 0.03925
R16202 Iout.n874 Iout 0.03925
R16203 Iout.n862 Iout 0.03925
R16204 Iout.n860 Iout 0.03925
R16205 Iout.n848 Iout 0.03925
R16206 Iout.n846 Iout 0.03925
R16207 Iout.n834 Iout 0.03925
R16208 Iout.n832 Iout 0.03925
R16209 Iout.n902 Iout 0.03925
R16210 Iout.n904 Iout 0.03925
R16211 Iout.n916 Iout 0.03925
R16212 Iout.n918 Iout 0.03925
R16213 Iout.n931 Iout 0.03925
R16214 Iout.n934 Iout 0.03925
R16215 Iout.n796 Iout 0.03925
R16216 Iout.n793 Iout 0.03925
R16217 Iout.n790 Iout 0.03925
R16218 Iout.n787 Iout 0.03925
R16219 Iout.n784 Iout 0.03925
R16220 Iout.n781 Iout 0.03925
R16221 Iout.n938 Iout 0.03925
R16222 Iout.n741 Iout 0.03925
R16223 Iout.n53 Iout 0.03925
R16224 Iout.n753 Iout 0.03925
R16225 Iout.n47 Iout 0.03925
R16226 Iout.n765 Iout 0.03925
R16227 Iout.n38 Iout 0.03925
R16228 Iout.n777 Iout 0.03925
R16229 Iout.n71 Iout 0.03925
R16230 Iout.n705 Iout 0.03925
R16231 Iout.n77 Iout 0.03925
R16232 Iout.n944 Iout 0.03925
R16233 Iout.n19 Iout 0.03925
R16234 Iout.n68 Iout 0.03925
R16235 Iout.n711 Iout 0.03925
R16236 Iout.n74 Iout 0.03925
R16237 Iout.n699 Iout 0.03925
R16238 Iout.n950 Iout 0.03925
R16239 Iout.n953 Iout 0.03925
R16240 Iout.n669 Iout 0.03925
R16241 Iout.n666 Iout 0.03925
R16242 Iout.n663 Iout 0.03925
R16243 Iout.n660 Iout 0.03925
R16244 Iout.n657 Iout 0.03925
R16245 Iout.n654 Iout 0.03925
R16246 Iout.n690 Iout 0.03925
R16247 Iout.n695 Iout 0.03925
R16248 Iout.n692 Iout 0.03925
R16249 Iout.n957 Iout 0.03925
R16250 Iout.n114 Iout 0.03925
R16251 Iout.n576 Iout 0.03925
R16252 Iout.n573 Iout 0.03925
R16253 Iout.n963 Iout 0.03925
R16254 Iout.n14 Iout 0.03925
R16255 Iout.n93 Iout 0.03925
R16256 Iout.n630 Iout 0.03925
R16257 Iout.n87 Iout 0.03925
R16258 Iout.n642 Iout 0.03925
R16259 Iout.n85 Iout 0.03925
R16260 Iout.n563 Iout 0.03925
R16261 Iout.n969 Iout 0.03925
R16262 Iout.n972 Iout 0.03925
R16263 Iout.n569 Iout 0.03925
R16264 Iout.n123 Iout 0.03925
R16265 Iout.n120 Iout 0.03925
R16266 Iout.n976 Iout 0.03925
R16267 Iout.n400 Iout 0.03925
R16268 Iout.n386 Iout 0.03925
R16269 Iout.n384 Iout 0.03925
R16270 Iout.n370 Iout 0.03925
R16271 Iout.n982 Iout 0.03925
R16272 Iout.n9 Iout 0.03925
R16273 Iout.n127 Iout 0.03925
R16274 Iout.n988 Iout 0.03925
R16275 Iout.n991 Iout 0.03925
R16276 Iout.n323 Iout 0.03925
R16277 Iout.n326 Iout 0.03925
R16278 Iout.n329 Iout 0.03925
R16279 Iout.n995 Iout 0.03925
R16280 Iout.n1001 Iout 0.03925
R16281 Iout.n4 Iout 0.03925
R16282 Iout.n295 Iout 0.03925
R16283 Iout.n172 Iout 0.03925
R16284 Iout.n1014 Iout 0.03925
R16285 Iout.n1022 Iout 0.02071
R16286 Iout Iout.n1022 0.00379
R16287 Iout.n303 Iout.n302 0.00105952
R16288 Iout.n377 Iout.n375 0.00105952
R16289 Iout.n380 Iout.n379 0.00105952
R16290 Iout.n368 Iout.n367 0.00105952
R16291 Iout.n365 Iout.n364 0.00105952
R16292 Iout.n362 Iout.n361 0.00105952
R16293 Iout.n650 Iout.n649 0.00105952
R16294 Iout.n647 Iout.n82 0.00105952
R16295 Iout.n638 Iout.n637 0.00105952
R16296 Iout.n635 Iout.n91 0.00105952
R16297 Iout.n43 Iout.n41 0.00105952
R16298 Iout.n773 Iout.n772 0.00105952
R16299 Iout.n770 Iout.n45 0.00105952
R16300 Iout.n761 Iout.n760 0.00105952
R16301 Iout.n758 Iout.n51 0.00105952
R16302 Iout.n825 Iout.n824 0.00105952
R16303 Iout.n822 Iout.n821 0.00105952
R16304 Iout.n819 Iout.n818 0.00105952
R16305 Iout.n816 Iout.n815 0.00105952
R16306 Iout.n813 Iout.n812 0.00105952
R16307 Iout.n810 Iout.n809 0.00105952
R16308 Iout.n829 Iout.n828 0.00105952
R16309 Iout.n840 Iout.n838 0.00105952
R16310 Iout.n843 Iout.n842 0.00105952
R16311 Iout.n854 Iout.n852 0.00105952
R16312 Iout.n857 Iout.n856 0.00105952
R16313 Iout.n868 Iout.n866 0.00105952
R16314 Iout.n871 Iout.n870 0.00105952
R16315 Iout.n925 Iout.n23 0.00105952
R16316 Iout.n928 Iout.n927 0.00105952
R16317 Iout.n924 Iout.n922 0.00105952
R16318 Iout.n913 Iout.n912 0.00105952
R16319 Iout.n910 Iout.n908 0.00105952
R16320 Iout.n899 Iout.n898 0.00105952
R16321 Iout.n896 Iout.n894 0.00105952
R16322 Iout.n885 Iout.n884 0.00105952
R16323 Iout.n882 Iout.n880 0.00105952
R16324 Iout.n833 Iout.n831 0.00105952
R16325 Iout.n836 Iout.n835 0.00105952
R16326 Iout.n847 Iout.n845 0.00105952
R16327 Iout.n850 Iout.n849 0.00105952
R16328 Iout.n861 Iout.n859 0.00105952
R16329 Iout.n864 Iout.n863 0.00105952
R16330 Iout.n875 Iout.n873 0.00105952
R16331 Iout.n878 Iout.n877 0.00105952
R16332 Iout.n889 Iout.n887 0.00105952
R16333 Iout.n935 Iout.n933 0.00105952
R16334 Iout.n932 Iout.n930 0.00105952
R16335 Iout.n920 Iout.n919 0.00105952
R16336 Iout.n917 Iout.n915 0.00105952
R16337 Iout.n906 Iout.n905 0.00105952
R16338 Iout.n903 Iout.n901 0.00105952
R16339 Iout.n892 Iout.n891 0.00105952
R16340 Iout.n940 Iout.n939 0.00105952
R16341 Iout.n783 Iout.n782 0.00105952
R16342 Iout.n786 Iout.n785 0.00105952
R16343 Iout.n789 Iout.n788 0.00105952
R16344 Iout.n792 Iout.n791 0.00105952
R16345 Iout.n795 Iout.n794 0.00105952
R16346 Iout.n798 Iout.n797 0.00105952
R16347 Iout.n801 Iout.n800 0.00105952
R16348 Iout.n804 Iout.n803 0.00105952
R16349 Iout.n807 Iout.n806 0.00105952
R16350 Iout.n779 Iout.n778 0.00105952
R16351 Iout.n776 Iout.n39 0.00105952
R16352 Iout.n767 Iout.n766 0.00105952
R16353 Iout.n764 Iout.n48 0.00105952
R16354 Iout.n755 Iout.n754 0.00105952
R16355 Iout.n752 Iout.n54 0.00105952
R16356 Iout.n743 Iout.n742 0.00105952
R16357 Iout.n740 Iout.n60 0.00105952
R16358 Iout.n731 Iout.n730 0.00105952
R16359 Iout.n728 Iout.n66 0.00105952
R16360 Iout.n943 Iout.n20 0.00105952
R16361 Iout.n946 Iout.n945 0.00105952
R16362 Iout.n704 Iout.n78 0.00105952
R16363 Iout.n707 Iout.n706 0.00105952
R16364 Iout.n716 Iout.n72 0.00105952
R16365 Iout.n719 Iout.n718 0.00105952
R16366 Iout.n954 Iout.n952 0.00105952
R16367 Iout.n951 Iout.n949 0.00105952
R16368 Iout.n701 Iout.n700 0.00105952
R16369 Iout.n710 Iout.n75 0.00105952
R16370 Iout.n713 Iout.n712 0.00105952
R16371 Iout.n722 Iout.n69 0.00105952
R16372 Iout.n725 Iout.n724 0.00105952
R16373 Iout.n734 Iout.n63 0.00105952
R16374 Iout.n737 Iout.n736 0.00105952
R16375 Iout.n746 Iout.n57 0.00105952
R16376 Iout.n749 Iout.n748 0.00105952
R16377 Iout.n655 Iout.n653 0.00105952
R16378 Iout.n658 Iout.n656 0.00105952
R16379 Iout.n661 Iout.n659 0.00105952
R16380 Iout.n664 Iout.n662 0.00105952
R16381 Iout.n667 Iout.n665 0.00105952
R16382 Iout.n670 Iout.n668 0.00105952
R16383 Iout.n673 Iout.n671 0.00105952
R16384 Iout.n676 Iout.n674 0.00105952
R16385 Iout.n679 Iout.n677 0.00105952
R16386 Iout.n682 Iout.n680 0.00105952
R16387 Iout.n685 Iout.n683 0.00105952
R16388 Iout.n959 Iout.n958 0.00105952
R16389 Iout.n694 Iout.n693 0.00105952
R16390 Iout.n697 Iout.n696 0.00105952
R16391 Iout.n691 Iout.n689 0.00105952
R16392 Iout.n688 Iout.n686 0.00105952
R16393 Iout.n962 Iout.n15 0.00105952
R16394 Iout.n965 Iout.n964 0.00105952
R16395 Iout.n575 Iout.n574 0.00105952
R16396 Iout.n578 Iout.n577 0.00105952
R16397 Iout.n587 Iout.n115 0.00105952
R16398 Iout.n590 Iout.n589 0.00105952
R16399 Iout.n599 Iout.n109 0.00105952
R16400 Iout.n602 Iout.n601 0.00105952
R16401 Iout.n611 Iout.n103 0.00105952
R16402 Iout.n614 Iout.n613 0.00105952
R16403 Iout.n623 Iout.n97 0.00105952
R16404 Iout.n626 Iout.n625 0.00105952
R16405 Iout.n86 Iout.n84 0.00105952
R16406 Iout.n644 Iout.n643 0.00105952
R16407 Iout.n641 Iout.n88 0.00105952
R16408 Iout.n632 Iout.n631 0.00105952
R16409 Iout.n629 Iout.n94 0.00105952
R16410 Iout.n620 Iout.n619 0.00105952
R16411 Iout.n617 Iout.n100 0.00105952
R16412 Iout.n608 Iout.n607 0.00105952
R16413 Iout.n605 Iout.n106 0.00105952
R16414 Iout.n596 Iout.n595 0.00105952
R16415 Iout.n593 Iout.n112 0.00105952
R16416 Iout.n584 Iout.n583 0.00105952
R16417 Iout.n973 Iout.n971 0.00105952
R16418 Iout.n970 Iout.n968 0.00105952
R16419 Iout.n565 Iout.n564 0.00105952
R16420 Iout.n581 Iout.n118 0.00105952
R16421 Iout.n978 Iout.n977 0.00105952
R16422 Iout.n122 Iout.n121 0.00105952
R16423 Iout.n568 Iout.n124 0.00105952
R16424 Iout.n571 Iout.n570 0.00105952
R16425 Iout.n335 Iout.n334 0.00105952
R16426 Iout.n338 Iout.n337 0.00105952
R16427 Iout.n341 Iout.n340 0.00105952
R16428 Iout.n344 Iout.n343 0.00105952
R16429 Iout.n347 Iout.n346 0.00105952
R16430 Iout.n350 Iout.n349 0.00105952
R16431 Iout.n353 Iout.n352 0.00105952
R16432 Iout.n356 Iout.n355 0.00105952
R16433 Iout.n359 Iout.n358 0.00105952
R16434 Iout.n372 Iout.n371 0.00105952
R16435 Iout.n385 Iout.n383 0.00105952
R16436 Iout.n388 Iout.n387 0.00105952
R16437 Iout.n401 Iout.n399 0.00105952
R16438 Iout.n404 Iout.n403 0.00105952
R16439 Iout.n417 Iout.n415 0.00105952
R16440 Iout.n420 Iout.n419 0.00105952
R16441 Iout.n433 Iout.n431 0.00105952
R16442 Iout.n443 Iout.n442 0.00105952
R16443 Iout.n440 Iout.n439 0.00105952
R16444 Iout.n437 Iout.n435 0.00105952
R16445 Iout.n555 Iout.n553 0.00105952
R16446 Iout.n558 Iout.n556 0.00105952
R16447 Iout.n981 Iout.n10 0.00105952
R16448 Iout.n984 Iout.n983 0.00105952
R16449 Iout.n561 Iout.n560 0.00105952
R16450 Iout.n992 Iout.n990 0.00105952
R16451 Iout.n989 Iout.n987 0.00105952
R16452 Iout.n129 Iout.n128 0.00105952
R16453 Iout.n547 Iout.n131 0.00105952
R16454 Iout.n550 Iout.n549 0.00105952
R16455 Iout.n451 Iout.n450 0.00105952
R16456 Iout.n454 Iout.n453 0.00105952
R16457 Iout.n448 Iout.n446 0.00105952
R16458 Iout.n428 Iout.n427 0.00105952
R16459 Iout.n425 Iout.n423 0.00105952
R16460 Iout.n412 Iout.n411 0.00105952
R16461 Iout.n409 Iout.n407 0.00105952
R16462 Iout.n396 Iout.n395 0.00105952
R16463 Iout.n393 Iout.n391 0.00105952
R16464 Iout.n331 Iout.n330 0.00105952
R16465 Iout.n328 Iout.n327 0.00105952
R16466 Iout.n325 Iout.n324 0.00105952
R16467 Iout.n322 Iout.n321 0.00105952
R16468 Iout.n319 Iout.n318 0.00105952
R16469 Iout.n316 Iout.n315 0.00105952
R16470 Iout.n313 Iout.n312 0.00105952
R16471 Iout.n310 Iout.n309 0.00105952
R16472 Iout.n307 Iout.n306 0.00105952
R16473 Iout.n459 Iout.n457 0.00105952
R16474 Iout.n465 Iout.n464 0.00105952
R16475 Iout.n462 Iout.n461 0.00105952
R16476 Iout.n544 Iout.n543 0.00105952
R16477 Iout.n541 Iout.n137 0.00105952
R16478 Iout.n997 Iout.n996 0.00105952
R16479 Iout.n135 Iout.n134 0.00105952
R16480 Iout.n1000 Iout.n5 0.00105952
R16481 Iout.n1003 Iout.n1002 0.00105952
R16482 Iout.n538 Iout.n537 0.00105952
R16483 Iout.n535 Iout.n533 0.00105952
R16484 Iout.n532 Iout.n530 0.00105952
R16485 Iout.n468 Iout.n157 0.00105952
R16486 Iout.n471 Iout.n470 0.00105952
R16487 Iout.n474 Iout.n473 0.00105952
R16488 Iout.n264 Iout.n190 0.00105952
R16489 Iout.n267 Iout.n266 0.00105952
R16490 Iout.n276 Iout.n184 0.00105952
R16491 Iout.n279 Iout.n278 0.00105952
R16492 Iout.n288 Iout.n178 0.00105952
R16493 Iout.n291 Iout.n290 0.00105952
R16494 Iout.n300 Iout.n169 0.00105952
R16495 Iout.n173 Iout.n171 0.00105952
R16496 Iout.n297 Iout.n296 0.00105952
R16497 Iout.n294 Iout.n175 0.00105952
R16498 Iout.n285 Iout.n284 0.00105952
R16499 Iout.n282 Iout.n181 0.00105952
R16500 Iout.n273 Iout.n272 0.00105952
R16501 Iout.n270 Iout.n187 0.00105952
R16502 Iout.n261 Iout.n260 0.00105952
R16503 Iout.n479 Iout.n477 0.00105952
R16504 Iout.n485 Iout.n484 0.00105952
R16505 Iout.n482 Iout.n481 0.00105952
R16506 Iout.n527 Iout.n526 0.00105952
R16507 Iout.n524 Iout.n144 0.00105952
R16508 Iout.n142 Iout.n141 0.00105952
R16509 Iout.n1008 Iout.n1006 0.00105952
R16510 Iout.n1011 Iout.n1009 0.00105952
R16511 Iout.n1016 Iout.n1015 0.00105952
R16512 Iout.n148 Iout.n147 0.00105952
R16513 Iout.n518 Iout.n150 0.00105952
R16514 Iout.n521 Iout.n520 0.00105952
R16515 Iout.n493 Iout.n492 0.00105952
R16516 Iout.n496 Iout.n495 0.00105952
R16517 Iout.n490 Iout.n488 0.00105952
R16518 Iout.n254 Iout.n253 0.00105952
R16519 Iout.n257 Iout.n256 0.00105952
R16520 Iout.n251 Iout.n249 0.00105952
R16521 Iout.n248 Iout.n246 0.00105952
R16522 Iout.n245 Iout.n243 0.00105952
R16523 Iout.n242 Iout.n240 0.00105952
R16524 Iout.n239 Iout.n237 0.00105952
R16525 Iout.n236 Iout.n234 0.00105952
R16526 Iout.n233 Iout.n231 0.00105952
R16527 Iout.n228 Iout.n227 0.00105952
R16528 Iout.n225 Iout.n223 0.00105952
R16529 Iout.n221 Iout.n219 0.00105952
R16530 Iout.n217 Iout.n215 0.00105952
R16531 Iout.n213 Iout.n211 0.00105952
R16532 Iout.n209 Iout.n207 0.00105952
R16533 Iout.n205 Iout.n203 0.00105952
R16534 Iout.n201 Iout.n200 0.00105952
R16535 Iout.n198 Iout.n196 0.00105952
R16536 Iout.n194 Iout.n193 0.00105952
R16537 Iout.n501 Iout.n499 0.00105952
R16538 Iout.n505 Iout.n503 0.00105952
R16539 Iout.n508 Iout.n506 0.00105952
R16540 Iout.n515 Iout.n514 0.00105952
R16541 Iout.n512 Iout.n510 0.00105952
R16542 Iout.n1021 Iout.n1019 0.00105952
R16543 XThC.Tn[10].n71 XThC.Tn[10].n70 256.104
R16544 XThC.Tn[10].n75 XThC.Tn[10].n74 243.679
R16545 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16546 XThC.Tn[10].n75 XThC.Tn[10].n73 205.28
R16547 XThC.Tn[10].n71 XThC.Tn[10].n69 202.095
R16548 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16549 XThC.Tn[10].n65 XThC.Tn[10].n63 161.365
R16550 XThC.Tn[10].n61 XThC.Tn[10].n59 161.365
R16551 XThC.Tn[10].n57 XThC.Tn[10].n55 161.365
R16552 XThC.Tn[10].n53 XThC.Tn[10].n51 161.365
R16553 XThC.Tn[10].n49 XThC.Tn[10].n47 161.365
R16554 XThC.Tn[10].n45 XThC.Tn[10].n43 161.365
R16555 XThC.Tn[10].n41 XThC.Tn[10].n39 161.365
R16556 XThC.Tn[10].n37 XThC.Tn[10].n35 161.365
R16557 XThC.Tn[10].n33 XThC.Tn[10].n31 161.365
R16558 XThC.Tn[10].n29 XThC.Tn[10].n27 161.365
R16559 XThC.Tn[10].n25 XThC.Tn[10].n23 161.365
R16560 XThC.Tn[10].n21 XThC.Tn[10].n19 161.365
R16561 XThC.Tn[10].n17 XThC.Tn[10].n15 161.365
R16562 XThC.Tn[10].n13 XThC.Tn[10].n11 161.365
R16563 XThC.Tn[10].n9 XThC.Tn[10].n7 161.365
R16564 XThC.Tn[10].n6 XThC.Tn[10].n4 161.365
R16565 XThC.Tn[10].n63 XThC.Tn[10].t42 161.202
R16566 XThC.Tn[10].n59 XThC.Tn[10].t32 161.202
R16567 XThC.Tn[10].n55 XThC.Tn[10].t19 161.202
R16568 XThC.Tn[10].n51 XThC.Tn[10].t16 161.202
R16569 XThC.Tn[10].n47 XThC.Tn[10].t40 161.202
R16570 XThC.Tn[10].n43 XThC.Tn[10].t27 161.202
R16571 XThC.Tn[10].n39 XThC.Tn[10].t26 161.202
R16572 XThC.Tn[10].n35 XThC.Tn[10].t39 161.202
R16573 XThC.Tn[10].n31 XThC.Tn[10].t37 161.202
R16574 XThC.Tn[10].n27 XThC.Tn[10].t28 161.202
R16575 XThC.Tn[10].n23 XThC.Tn[10].t15 161.202
R16576 XThC.Tn[10].n19 XThC.Tn[10].t14 161.202
R16577 XThC.Tn[10].n15 XThC.Tn[10].t25 161.202
R16578 XThC.Tn[10].n11 XThC.Tn[10].t23 161.202
R16579 XThC.Tn[10].n7 XThC.Tn[10].t21 161.202
R16580 XThC.Tn[10].n4 XThC.Tn[10].t36 161.202
R16581 XThC.Tn[10].n63 XThC.Tn[10].t13 145.137
R16582 XThC.Tn[10].n59 XThC.Tn[10].t35 145.137
R16583 XThC.Tn[10].n55 XThC.Tn[10].t22 145.137
R16584 XThC.Tn[10].n51 XThC.Tn[10].t20 145.137
R16585 XThC.Tn[10].n47 XThC.Tn[10].t12 145.137
R16586 XThC.Tn[10].n43 XThC.Tn[10].t33 145.137
R16587 XThC.Tn[10].n39 XThC.Tn[10].t31 145.137
R16588 XThC.Tn[10].n35 XThC.Tn[10].t43 145.137
R16589 XThC.Tn[10].n31 XThC.Tn[10].t41 145.137
R16590 XThC.Tn[10].n27 XThC.Tn[10].t34 145.137
R16591 XThC.Tn[10].n23 XThC.Tn[10].t18 145.137
R16592 XThC.Tn[10].n19 XThC.Tn[10].t17 145.137
R16593 XThC.Tn[10].n15 XThC.Tn[10].t30 145.137
R16594 XThC.Tn[10].n11 XThC.Tn[10].t29 145.137
R16595 XThC.Tn[10].n7 XThC.Tn[10].t24 145.137
R16596 XThC.Tn[10].n4 XThC.Tn[10].t38 145.137
R16597 XThC.Tn[10].n69 XThC.Tn[10].t7 26.5955
R16598 XThC.Tn[10].n69 XThC.Tn[10].t6 26.5955
R16599 XThC.Tn[10].n70 XThC.Tn[10].t2 26.5955
R16600 XThC.Tn[10].n70 XThC.Tn[10].t10 26.5955
R16601 XThC.Tn[10].n73 XThC.Tn[10].t8 26.5955
R16602 XThC.Tn[10].n73 XThC.Tn[10].t9 26.5955
R16603 XThC.Tn[10].n74 XThC.Tn[10].t0 26.5955
R16604 XThC.Tn[10].n74 XThC.Tn[10].t11 26.5955
R16605 XThC.Tn[10].n1 XThC.Tn[10].t3 24.9236
R16606 XThC.Tn[10].n1 XThC.Tn[10].t5 24.9236
R16607 XThC.Tn[10].n0 XThC.Tn[10].t4 24.9236
R16608 XThC.Tn[10].n0 XThC.Tn[10].t1 24.9236
R16609 XThC.Tn[10] XThC.Tn[10].n75 22.9652
R16610 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16611 XThC.Tn[10].n72 XThC.Tn[10].n71 13.9299
R16612 XThC.Tn[10] XThC.Tn[10].n72 13.9299
R16613 XThC.Tn[10] XThC.Tn[10].n6 8.0245
R16614 XThC.Tn[10].n66 XThC.Tn[10].n65 7.9105
R16615 XThC.Tn[10].n62 XThC.Tn[10].n61 7.9105
R16616 XThC.Tn[10].n58 XThC.Tn[10].n57 7.9105
R16617 XThC.Tn[10].n54 XThC.Tn[10].n53 7.9105
R16618 XThC.Tn[10].n50 XThC.Tn[10].n49 7.9105
R16619 XThC.Tn[10].n46 XThC.Tn[10].n45 7.9105
R16620 XThC.Tn[10].n42 XThC.Tn[10].n41 7.9105
R16621 XThC.Tn[10].n38 XThC.Tn[10].n37 7.9105
R16622 XThC.Tn[10].n34 XThC.Tn[10].n33 7.9105
R16623 XThC.Tn[10].n30 XThC.Tn[10].n29 7.9105
R16624 XThC.Tn[10].n26 XThC.Tn[10].n25 7.9105
R16625 XThC.Tn[10].n22 XThC.Tn[10].n21 7.9105
R16626 XThC.Tn[10].n18 XThC.Tn[10].n17 7.9105
R16627 XThC.Tn[10].n14 XThC.Tn[10].n13 7.9105
R16628 XThC.Tn[10].n10 XThC.Tn[10].n9 7.9105
R16629 XThC.Tn[10].n68 XThC.Tn[10].n67 7.40985
R16630 XThC.Tn[10].n67 XThC.Tn[10] 4.38575
R16631 XThC.Tn[10].n72 XThC.Tn[10].n68 2.99115
R16632 XThC.Tn[10].n72 XThC.Tn[10] 2.87153
R16633 XThC.Tn[10].n3 XThC.Tn[10] 2.688
R16634 XThC.Tn[10].n68 XThC.Tn[10] 2.2734
R16635 XThC.Tn[10].n67 XThC.Tn[10].n3 0.244922
R16636 XThC.Tn[10].n10 XThC.Tn[10] 0.235138
R16637 XThC.Tn[10].n14 XThC.Tn[10] 0.235138
R16638 XThC.Tn[10].n18 XThC.Tn[10] 0.235138
R16639 XThC.Tn[10].n22 XThC.Tn[10] 0.235138
R16640 XThC.Tn[10].n26 XThC.Tn[10] 0.235138
R16641 XThC.Tn[10].n30 XThC.Tn[10] 0.235138
R16642 XThC.Tn[10].n34 XThC.Tn[10] 0.235138
R16643 XThC.Tn[10].n38 XThC.Tn[10] 0.235138
R16644 XThC.Tn[10].n42 XThC.Tn[10] 0.235138
R16645 XThC.Tn[10].n46 XThC.Tn[10] 0.235138
R16646 XThC.Tn[10].n50 XThC.Tn[10] 0.235138
R16647 XThC.Tn[10].n54 XThC.Tn[10] 0.235138
R16648 XThC.Tn[10].n58 XThC.Tn[10] 0.235138
R16649 XThC.Tn[10].n62 XThC.Tn[10] 0.235138
R16650 XThC.Tn[10].n66 XThC.Tn[10] 0.235138
R16651 XThC.Tn[10].n3 XThC.Tn[10] 0.141947
R16652 XThC.Tn[10] XThC.Tn[10].n10 0.114505
R16653 XThC.Tn[10] XThC.Tn[10].n14 0.114505
R16654 XThC.Tn[10] XThC.Tn[10].n18 0.114505
R16655 XThC.Tn[10] XThC.Tn[10].n22 0.114505
R16656 XThC.Tn[10] XThC.Tn[10].n26 0.114505
R16657 XThC.Tn[10] XThC.Tn[10].n30 0.114505
R16658 XThC.Tn[10] XThC.Tn[10].n34 0.114505
R16659 XThC.Tn[10] XThC.Tn[10].n38 0.114505
R16660 XThC.Tn[10] XThC.Tn[10].n42 0.114505
R16661 XThC.Tn[10] XThC.Tn[10].n46 0.114505
R16662 XThC.Tn[10] XThC.Tn[10].n50 0.114505
R16663 XThC.Tn[10] XThC.Tn[10].n54 0.114505
R16664 XThC.Tn[10] XThC.Tn[10].n58 0.114505
R16665 XThC.Tn[10] XThC.Tn[10].n62 0.114505
R16666 XThC.Tn[10] XThC.Tn[10].n66 0.114505
R16667 XThC.Tn[10].n65 XThC.Tn[10].n64 0.0599512
R16668 XThC.Tn[10].n61 XThC.Tn[10].n60 0.0599512
R16669 XThC.Tn[10].n57 XThC.Tn[10].n56 0.0599512
R16670 XThC.Tn[10].n53 XThC.Tn[10].n52 0.0599512
R16671 XThC.Tn[10].n49 XThC.Tn[10].n48 0.0599512
R16672 XThC.Tn[10].n45 XThC.Tn[10].n44 0.0599512
R16673 XThC.Tn[10].n41 XThC.Tn[10].n40 0.0599512
R16674 XThC.Tn[10].n37 XThC.Tn[10].n36 0.0599512
R16675 XThC.Tn[10].n33 XThC.Tn[10].n32 0.0599512
R16676 XThC.Tn[10].n29 XThC.Tn[10].n28 0.0599512
R16677 XThC.Tn[10].n25 XThC.Tn[10].n24 0.0599512
R16678 XThC.Tn[10].n21 XThC.Tn[10].n20 0.0599512
R16679 XThC.Tn[10].n17 XThC.Tn[10].n16 0.0599512
R16680 XThC.Tn[10].n13 XThC.Tn[10].n12 0.0599512
R16681 XThC.Tn[10].n9 XThC.Tn[10].n8 0.0599512
R16682 XThC.Tn[10].n6 XThC.Tn[10].n5 0.0599512
R16683 XThC.Tn[10].n64 XThC.Tn[10] 0.0469286
R16684 XThC.Tn[10].n60 XThC.Tn[10] 0.0469286
R16685 XThC.Tn[10].n56 XThC.Tn[10] 0.0469286
R16686 XThC.Tn[10].n52 XThC.Tn[10] 0.0469286
R16687 XThC.Tn[10].n48 XThC.Tn[10] 0.0469286
R16688 XThC.Tn[10].n44 XThC.Tn[10] 0.0469286
R16689 XThC.Tn[10].n40 XThC.Tn[10] 0.0469286
R16690 XThC.Tn[10].n36 XThC.Tn[10] 0.0469286
R16691 XThC.Tn[10].n32 XThC.Tn[10] 0.0469286
R16692 XThC.Tn[10].n28 XThC.Tn[10] 0.0469286
R16693 XThC.Tn[10].n24 XThC.Tn[10] 0.0469286
R16694 XThC.Tn[10].n20 XThC.Tn[10] 0.0469286
R16695 XThC.Tn[10].n16 XThC.Tn[10] 0.0469286
R16696 XThC.Tn[10].n12 XThC.Tn[10] 0.0469286
R16697 XThC.Tn[10].n8 XThC.Tn[10] 0.0469286
R16698 XThC.Tn[10].n5 XThC.Tn[10] 0.0469286
R16699 XThC.Tn[10].n64 XThC.Tn[10] 0.0401341
R16700 XThC.Tn[10].n60 XThC.Tn[10] 0.0401341
R16701 XThC.Tn[10].n56 XThC.Tn[10] 0.0401341
R16702 XThC.Tn[10].n52 XThC.Tn[10] 0.0401341
R16703 XThC.Tn[10].n48 XThC.Tn[10] 0.0401341
R16704 XThC.Tn[10].n44 XThC.Tn[10] 0.0401341
R16705 XThC.Tn[10].n40 XThC.Tn[10] 0.0401341
R16706 XThC.Tn[10].n36 XThC.Tn[10] 0.0401341
R16707 XThC.Tn[10].n32 XThC.Tn[10] 0.0401341
R16708 XThC.Tn[10].n28 XThC.Tn[10] 0.0401341
R16709 XThC.Tn[10].n24 XThC.Tn[10] 0.0401341
R16710 XThC.Tn[10].n20 XThC.Tn[10] 0.0401341
R16711 XThC.Tn[10].n16 XThC.Tn[10] 0.0401341
R16712 XThC.Tn[10].n12 XThC.Tn[10] 0.0401341
R16713 XThC.Tn[10].n8 XThC.Tn[10] 0.0401341
R16714 XThC.Tn[10].n5 XThC.Tn[10] 0.0401341
R16715 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R16716 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R16717 XThR.Tn[6] XThR.Tn[6].n82 161.363
R16718 XThR.Tn[6] XThR.Tn[6].n77 161.363
R16719 XThR.Tn[6] XThR.Tn[6].n72 161.363
R16720 XThR.Tn[6] XThR.Tn[6].n67 161.363
R16721 XThR.Tn[6] XThR.Tn[6].n62 161.363
R16722 XThR.Tn[6] XThR.Tn[6].n57 161.363
R16723 XThR.Tn[6] XThR.Tn[6].n52 161.363
R16724 XThR.Tn[6] XThR.Tn[6].n47 161.363
R16725 XThR.Tn[6] XThR.Tn[6].n42 161.363
R16726 XThR.Tn[6] XThR.Tn[6].n37 161.363
R16727 XThR.Tn[6] XThR.Tn[6].n32 161.363
R16728 XThR.Tn[6] XThR.Tn[6].n27 161.363
R16729 XThR.Tn[6] XThR.Tn[6].n22 161.363
R16730 XThR.Tn[6] XThR.Tn[6].n17 161.363
R16731 XThR.Tn[6] XThR.Tn[6].n12 161.363
R16732 XThR.Tn[6] XThR.Tn[6].n10 161.363
R16733 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R16734 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R16735 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R16736 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R16737 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R16738 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R16739 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R16740 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R16741 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R16742 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R16743 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R16744 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R16745 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R16746 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R16747 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R16748 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R16749 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R16750 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R16751 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R16752 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R16753 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R16754 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R16755 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R16756 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R16757 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R16758 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R16759 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R16760 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R16761 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R16762 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R16763 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R16764 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R16765 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R16766 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R16767 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R16768 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R16769 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R16770 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R16771 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R16772 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R16773 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R16774 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R16775 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R16776 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R16777 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R16778 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R16779 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R16780 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R16781 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R16782 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R16783 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R16784 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R16785 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R16786 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R16787 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R16788 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R16789 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R16790 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R16791 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R16792 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R16793 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R16794 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R16795 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R16796 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R16797 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R16798 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R16799 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R16800 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R16801 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R16802 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R16803 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R16804 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R16805 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R16806 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R16807 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R16808 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R16809 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R16810 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R16811 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R16812 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R16813 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R16814 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R16815 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R16816 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R16817 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R16818 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R16819 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R16820 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R16821 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R16822 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R16823 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R16824 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R16825 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R16826 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R16827 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R16828 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R16829 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R16830 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R16831 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R16832 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R16833 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R16834 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R16835 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R16836 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R16837 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R16838 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R16839 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R16840 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R16841 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R16842 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R16843 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R16844 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R16845 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R16846 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R16847 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R16848 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R16849 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R16850 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R16851 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R16852 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R16853 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R16854 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R16855 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R16856 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R16857 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R16858 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R16859 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R16860 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R16861 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R16862 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R16863 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R16864 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R16865 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R16866 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R16867 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R16868 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R16869 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R16870 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R16871 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R16872 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R16873 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R16874 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R16875 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R16876 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R16877 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R16878 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R16879 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R16880 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R16881 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R16882 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R16883 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R16884 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R16885 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R16886 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R16887 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R16888 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R16889 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R16890 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R16891 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R16892 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R16893 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R16894 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R16895 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R16896 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R16897 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R16898 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R16899 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R16900 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R16901 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R16902 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R16903 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R16904 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R16905 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R16906 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R16907 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R16908 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R16909 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R16910 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R16911 XThR.Tn[6] XThR.Tn[6].n87 0.038
R16912 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R16913 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R16914 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R16915 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R16916 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R16917 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R16918 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R16919 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R16920 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R16921 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R16922 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R16923 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R16924 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R16925 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R16926 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R16927 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R16928 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R16929 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R16930 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R16931 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R16932 XThR.Tn[14].n87 XThR.Tn[14].n85 202.094
R16933 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R16934 XThR.Tn[14] XThR.Tn[14].n78 161.363
R16935 XThR.Tn[14] XThR.Tn[14].n73 161.363
R16936 XThR.Tn[14] XThR.Tn[14].n68 161.363
R16937 XThR.Tn[14] XThR.Tn[14].n63 161.363
R16938 XThR.Tn[14] XThR.Tn[14].n58 161.363
R16939 XThR.Tn[14] XThR.Tn[14].n53 161.363
R16940 XThR.Tn[14] XThR.Tn[14].n48 161.363
R16941 XThR.Tn[14] XThR.Tn[14].n43 161.363
R16942 XThR.Tn[14] XThR.Tn[14].n38 161.363
R16943 XThR.Tn[14] XThR.Tn[14].n33 161.363
R16944 XThR.Tn[14] XThR.Tn[14].n28 161.363
R16945 XThR.Tn[14] XThR.Tn[14].n23 161.363
R16946 XThR.Tn[14] XThR.Tn[14].n18 161.363
R16947 XThR.Tn[14] XThR.Tn[14].n13 161.363
R16948 XThR.Tn[14] XThR.Tn[14].n8 161.363
R16949 XThR.Tn[14] XThR.Tn[14].n6 161.363
R16950 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R16951 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R16952 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R16953 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R16954 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R16955 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R16956 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R16957 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R16958 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R16959 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R16960 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R16961 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R16962 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R16963 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R16964 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R16965 XThR.Tn[14].n78 XThR.Tn[14].t51 161.106
R16966 XThR.Tn[14].n73 XThR.Tn[14].t58 161.106
R16967 XThR.Tn[14].n68 XThR.Tn[14].t39 161.106
R16968 XThR.Tn[14].n63 XThR.Tn[14].t22 161.106
R16969 XThR.Tn[14].n58 XThR.Tn[14].t49 161.106
R16970 XThR.Tn[14].n53 XThR.Tn[14].t12 161.106
R16971 XThR.Tn[14].n48 XThR.Tn[14].t56 161.106
R16972 XThR.Tn[14].n43 XThR.Tn[14].t36 161.106
R16973 XThR.Tn[14].n38 XThR.Tn[14].t19 161.106
R16974 XThR.Tn[14].n33 XThR.Tn[14].t25 161.106
R16975 XThR.Tn[14].n28 XThR.Tn[14].t73 161.106
R16976 XThR.Tn[14].n23 XThR.Tn[14].t38 161.106
R16977 XThR.Tn[14].n18 XThR.Tn[14].t72 161.106
R16978 XThR.Tn[14].n13 XThR.Tn[14].t54 161.106
R16979 XThR.Tn[14].n8 XThR.Tn[14].t13 161.106
R16980 XThR.Tn[14].n6 XThR.Tn[14].t62 161.106
R16981 XThR.Tn[14].n79 XThR.Tn[14].t32 159.978
R16982 XThR.Tn[14].n74 XThR.Tn[14].t37 159.978
R16983 XThR.Tn[14].n69 XThR.Tn[14].t20 159.978
R16984 XThR.Tn[14].n64 XThR.Tn[14].t68 159.978
R16985 XThR.Tn[14].n59 XThR.Tn[14].t30 159.978
R16986 XThR.Tn[14].n54 XThR.Tn[14].t55 159.978
R16987 XThR.Tn[14].n49 XThR.Tn[14].t35 159.978
R16988 XThR.Tn[14].n44 XThR.Tn[14].t16 159.978
R16989 XThR.Tn[14].n39 XThR.Tn[14].t66 159.978
R16990 XThR.Tn[14].n34 XThR.Tn[14].t71 159.978
R16991 XThR.Tn[14].n29 XThR.Tn[14].t53 159.978
R16992 XThR.Tn[14].n24 XThR.Tn[14].t18 159.978
R16993 XThR.Tn[14].n19 XThR.Tn[14].t52 159.978
R16994 XThR.Tn[14].n14 XThR.Tn[14].t34 159.978
R16995 XThR.Tn[14].n9 XThR.Tn[14].t60 159.978
R16996 XThR.Tn[14].n78 XThR.Tn[14].t41 145.038
R16997 XThR.Tn[14].n73 XThR.Tn[14].t65 145.038
R16998 XThR.Tn[14].n68 XThR.Tn[14].t45 145.038
R16999 XThR.Tn[14].n63 XThR.Tn[14].t26 145.038
R17000 XThR.Tn[14].n58 XThR.Tn[14].t59 145.038
R17001 XThR.Tn[14].n53 XThR.Tn[14].t40 145.038
R17002 XThR.Tn[14].n48 XThR.Tn[14].t46 145.038
R17003 XThR.Tn[14].n43 XThR.Tn[14].t27 145.038
R17004 XThR.Tn[14].n38 XThR.Tn[14].t23 145.038
R17005 XThR.Tn[14].n33 XThR.Tn[14].t57 145.038
R17006 XThR.Tn[14].n28 XThR.Tn[14].t15 145.038
R17007 XThR.Tn[14].n23 XThR.Tn[14].t44 145.038
R17008 XThR.Tn[14].n18 XThR.Tn[14].t14 145.038
R17009 XThR.Tn[14].n13 XThR.Tn[14].t64 145.038
R17010 XThR.Tn[14].n8 XThR.Tn[14].t24 145.038
R17011 XThR.Tn[14].n6 XThR.Tn[14].t69 145.038
R17012 XThR.Tn[14].n79 XThR.Tn[14].t43 143.911
R17013 XThR.Tn[14].n74 XThR.Tn[14].t70 143.911
R17014 XThR.Tn[14].n69 XThR.Tn[14].t48 143.911
R17015 XThR.Tn[14].n64 XThR.Tn[14].t31 143.911
R17016 XThR.Tn[14].n59 XThR.Tn[14].t63 143.911
R17017 XThR.Tn[14].n54 XThR.Tn[14].t42 143.911
R17018 XThR.Tn[14].n49 XThR.Tn[14].t50 143.911
R17019 XThR.Tn[14].n44 XThR.Tn[14].t33 143.911
R17020 XThR.Tn[14].n39 XThR.Tn[14].t29 143.911
R17021 XThR.Tn[14].n34 XThR.Tn[14].t61 143.911
R17022 XThR.Tn[14].n29 XThR.Tn[14].t21 143.911
R17023 XThR.Tn[14].n24 XThR.Tn[14].t47 143.911
R17024 XThR.Tn[14].n19 XThR.Tn[14].t17 143.911
R17025 XThR.Tn[14].n14 XThR.Tn[14].t67 143.911
R17026 XThR.Tn[14].n9 XThR.Tn[14].t28 143.911
R17027 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17028 XThR.Tn[14].n86 XThR.Tn[14].t0 26.5955
R17029 XThR.Tn[14].n86 XThR.Tn[14].t1 26.5955
R17030 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R17031 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R17032 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R17033 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R17034 XThR.Tn[14].n85 XThR.Tn[14].t2 26.5955
R17035 XThR.Tn[14].n85 XThR.Tn[14].t3 26.5955
R17036 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R17037 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R17038 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R17039 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R17040 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R17041 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R17042 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R17043 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R17044 XThR.Tn[14] XThR.Tn[14].n7 5.34038
R17045 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R17046 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R17047 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R17048 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R17049 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R17050 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R17051 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R17052 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R17053 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R17054 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R17055 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R17056 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R17057 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R17058 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R17059 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R17060 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R17061 XThR.Tn[14].n12 XThR.Tn[14] 2.52282
R17062 XThR.Tn[14].n17 XThR.Tn[14] 2.52282
R17063 XThR.Tn[14].n22 XThR.Tn[14] 2.52282
R17064 XThR.Tn[14].n27 XThR.Tn[14] 2.52282
R17065 XThR.Tn[14].n32 XThR.Tn[14] 2.52282
R17066 XThR.Tn[14].n37 XThR.Tn[14] 2.52282
R17067 XThR.Tn[14].n42 XThR.Tn[14] 2.52282
R17068 XThR.Tn[14].n47 XThR.Tn[14] 2.52282
R17069 XThR.Tn[14].n52 XThR.Tn[14] 2.52282
R17070 XThR.Tn[14].n57 XThR.Tn[14] 2.52282
R17071 XThR.Tn[14].n62 XThR.Tn[14] 2.52282
R17072 XThR.Tn[14].n67 XThR.Tn[14] 2.52282
R17073 XThR.Tn[14].n72 XThR.Tn[14] 2.52282
R17074 XThR.Tn[14].n77 XThR.Tn[14] 2.52282
R17075 XThR.Tn[14].n82 XThR.Tn[14] 2.52282
R17076 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R17077 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R17078 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R17079 XThR.Tn[14].n80 XThR.Tn[14] 1.08677
R17080 XThR.Tn[14].n75 XThR.Tn[14] 1.08677
R17081 XThR.Tn[14].n70 XThR.Tn[14] 1.08677
R17082 XThR.Tn[14].n65 XThR.Tn[14] 1.08677
R17083 XThR.Tn[14].n60 XThR.Tn[14] 1.08677
R17084 XThR.Tn[14].n55 XThR.Tn[14] 1.08677
R17085 XThR.Tn[14].n50 XThR.Tn[14] 1.08677
R17086 XThR.Tn[14].n45 XThR.Tn[14] 1.08677
R17087 XThR.Tn[14].n40 XThR.Tn[14] 1.08677
R17088 XThR.Tn[14].n35 XThR.Tn[14] 1.08677
R17089 XThR.Tn[14].n30 XThR.Tn[14] 1.08677
R17090 XThR.Tn[14].n25 XThR.Tn[14] 1.08677
R17091 XThR.Tn[14].n20 XThR.Tn[14] 1.08677
R17092 XThR.Tn[14].n15 XThR.Tn[14] 1.08677
R17093 XThR.Tn[14].n10 XThR.Tn[14] 1.08677
R17094 XThR.Tn[14] XThR.Tn[14].n12 0.839786
R17095 XThR.Tn[14] XThR.Tn[14].n17 0.839786
R17096 XThR.Tn[14] XThR.Tn[14].n22 0.839786
R17097 XThR.Tn[14] XThR.Tn[14].n27 0.839786
R17098 XThR.Tn[14] XThR.Tn[14].n32 0.839786
R17099 XThR.Tn[14] XThR.Tn[14].n37 0.839786
R17100 XThR.Tn[14] XThR.Tn[14].n42 0.839786
R17101 XThR.Tn[14] XThR.Tn[14].n47 0.839786
R17102 XThR.Tn[14] XThR.Tn[14].n52 0.839786
R17103 XThR.Tn[14] XThR.Tn[14].n57 0.839786
R17104 XThR.Tn[14] XThR.Tn[14].n62 0.839786
R17105 XThR.Tn[14] XThR.Tn[14].n67 0.839786
R17106 XThR.Tn[14] XThR.Tn[14].n72 0.839786
R17107 XThR.Tn[14] XThR.Tn[14].n77 0.839786
R17108 XThR.Tn[14] XThR.Tn[14].n82 0.839786
R17109 XThR.Tn[14].n7 XThR.Tn[14] 0.499542
R17110 XThR.Tn[14].n81 XThR.Tn[14] 0.063
R17111 XThR.Tn[14].n76 XThR.Tn[14] 0.063
R17112 XThR.Tn[14].n71 XThR.Tn[14] 0.063
R17113 XThR.Tn[14].n66 XThR.Tn[14] 0.063
R17114 XThR.Tn[14].n61 XThR.Tn[14] 0.063
R17115 XThR.Tn[14].n56 XThR.Tn[14] 0.063
R17116 XThR.Tn[14].n51 XThR.Tn[14] 0.063
R17117 XThR.Tn[14].n46 XThR.Tn[14] 0.063
R17118 XThR.Tn[14].n41 XThR.Tn[14] 0.063
R17119 XThR.Tn[14].n36 XThR.Tn[14] 0.063
R17120 XThR.Tn[14].n31 XThR.Tn[14] 0.063
R17121 XThR.Tn[14].n26 XThR.Tn[14] 0.063
R17122 XThR.Tn[14].n21 XThR.Tn[14] 0.063
R17123 XThR.Tn[14].n16 XThR.Tn[14] 0.063
R17124 XThR.Tn[14].n11 XThR.Tn[14] 0.063
R17125 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R17126 XThR.Tn[14] XThR.Tn[14].n83 0.038
R17127 XThR.Tn[14].n7 XThR.Tn[14] 0.0143889
R17128 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00771154
R17129 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00771154
R17130 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00771154
R17131 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00771154
R17132 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00771154
R17133 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00771154
R17134 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00771154
R17135 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00771154
R17136 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00771154
R17137 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00771154
R17138 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00771154
R17139 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00771154
R17140 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00771154
R17141 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00771154
R17142 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00771154
R17143 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R17144 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R17145 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R17146 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R17147 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R17148 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R17149 XThR.Tn[12] XThR.Tn[12].n78 161.363
R17150 XThR.Tn[12] XThR.Tn[12].n73 161.363
R17151 XThR.Tn[12] XThR.Tn[12].n68 161.363
R17152 XThR.Tn[12] XThR.Tn[12].n63 161.363
R17153 XThR.Tn[12] XThR.Tn[12].n58 161.363
R17154 XThR.Tn[12] XThR.Tn[12].n53 161.363
R17155 XThR.Tn[12] XThR.Tn[12].n48 161.363
R17156 XThR.Tn[12] XThR.Tn[12].n43 161.363
R17157 XThR.Tn[12] XThR.Tn[12].n38 161.363
R17158 XThR.Tn[12] XThR.Tn[12].n33 161.363
R17159 XThR.Tn[12] XThR.Tn[12].n28 161.363
R17160 XThR.Tn[12] XThR.Tn[12].n23 161.363
R17161 XThR.Tn[12] XThR.Tn[12].n18 161.363
R17162 XThR.Tn[12] XThR.Tn[12].n13 161.363
R17163 XThR.Tn[12] XThR.Tn[12].n8 161.363
R17164 XThR.Tn[12] XThR.Tn[12].n6 161.363
R17165 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R17166 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R17167 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R17168 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R17169 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R17170 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R17171 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R17172 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R17173 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R17174 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R17175 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R17176 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R17177 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R17178 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R17179 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R17180 XThR.Tn[12].n78 XThR.Tn[12].t18 161.106
R17181 XThR.Tn[12].n73 XThR.Tn[12].t24 161.106
R17182 XThR.Tn[12].n68 XThR.Tn[12].t67 161.106
R17183 XThR.Tn[12].n63 XThR.Tn[12].t52 161.106
R17184 XThR.Tn[12].n58 XThR.Tn[12].t16 161.106
R17185 XThR.Tn[12].n53 XThR.Tn[12].t40 161.106
R17186 XThR.Tn[12].n48 XThR.Tn[12].t22 161.106
R17187 XThR.Tn[12].n43 XThR.Tn[12].t65 161.106
R17188 XThR.Tn[12].n38 XThR.Tn[12].t51 161.106
R17189 XThR.Tn[12].n33 XThR.Tn[12].t56 161.106
R17190 XThR.Tn[12].n28 XThR.Tn[12].t39 161.106
R17191 XThR.Tn[12].n23 XThR.Tn[12].t66 161.106
R17192 XThR.Tn[12].n18 XThR.Tn[12].t38 161.106
R17193 XThR.Tn[12].n13 XThR.Tn[12].t20 161.106
R17194 XThR.Tn[12].n8 XThR.Tn[12].t43 161.106
R17195 XThR.Tn[12].n6 XThR.Tn[12].t28 161.106
R17196 XThR.Tn[12].n79 XThR.Tn[12].t58 159.978
R17197 XThR.Tn[12].n74 XThR.Tn[12].t62 159.978
R17198 XThR.Tn[12].n69 XThR.Tn[12].t47 159.978
R17199 XThR.Tn[12].n64 XThR.Tn[12].t31 159.978
R17200 XThR.Tn[12].n59 XThR.Tn[12].t55 159.978
R17201 XThR.Tn[12].n54 XThR.Tn[12].t19 159.978
R17202 XThR.Tn[12].n49 XThR.Tn[12].t61 159.978
R17203 XThR.Tn[12].n44 XThR.Tn[12].t44 159.978
R17204 XThR.Tn[12].n39 XThR.Tn[12].t29 159.978
R17205 XThR.Tn[12].n34 XThR.Tn[12].t37 159.978
R17206 XThR.Tn[12].n29 XThR.Tn[12].t17 159.978
R17207 XThR.Tn[12].n24 XThR.Tn[12].t46 159.978
R17208 XThR.Tn[12].n19 XThR.Tn[12].t15 159.978
R17209 XThR.Tn[12].n14 XThR.Tn[12].t60 159.978
R17210 XThR.Tn[12].n9 XThR.Tn[12].t21 159.978
R17211 XThR.Tn[12].n78 XThR.Tn[12].t69 145.038
R17212 XThR.Tn[12].n73 XThR.Tn[12].t32 145.038
R17213 XThR.Tn[12].n68 XThR.Tn[12].t73 145.038
R17214 XThR.Tn[12].n63 XThR.Tn[12].t57 145.038
R17215 XThR.Tn[12].n58 XThR.Tn[12].t25 145.038
R17216 XThR.Tn[12].n53 XThR.Tn[12].t68 145.038
R17217 XThR.Tn[12].n48 XThR.Tn[12].t12 145.038
R17218 XThR.Tn[12].n43 XThR.Tn[12].t59 145.038
R17219 XThR.Tn[12].n38 XThR.Tn[12].t54 145.038
R17220 XThR.Tn[12].n33 XThR.Tn[12].t23 145.038
R17221 XThR.Tn[12].n28 XThR.Tn[12].t48 145.038
R17222 XThR.Tn[12].n23 XThR.Tn[12].t70 145.038
R17223 XThR.Tn[12].n18 XThR.Tn[12].t45 145.038
R17224 XThR.Tn[12].n13 XThR.Tn[12].t30 145.038
R17225 XThR.Tn[12].n8 XThR.Tn[12].t53 145.038
R17226 XThR.Tn[12].n6 XThR.Tn[12].t36 145.038
R17227 XThR.Tn[12].n79 XThR.Tn[12].t27 143.911
R17228 XThR.Tn[12].n74 XThR.Tn[12].t50 143.911
R17229 XThR.Tn[12].n69 XThR.Tn[12].t34 143.911
R17230 XThR.Tn[12].n64 XThR.Tn[12].t13 143.911
R17231 XThR.Tn[12].n59 XThR.Tn[12].t42 143.911
R17232 XThR.Tn[12].n54 XThR.Tn[12].t26 143.911
R17233 XThR.Tn[12].n49 XThR.Tn[12].t35 143.911
R17234 XThR.Tn[12].n44 XThR.Tn[12].t14 143.911
R17235 XThR.Tn[12].n39 XThR.Tn[12].t72 143.911
R17236 XThR.Tn[12].n34 XThR.Tn[12].t41 143.911
R17237 XThR.Tn[12].n29 XThR.Tn[12].t64 143.911
R17238 XThR.Tn[12].n24 XThR.Tn[12].t33 143.911
R17239 XThR.Tn[12].n19 XThR.Tn[12].t63 143.911
R17240 XThR.Tn[12].n14 XThR.Tn[12].t49 143.911
R17241 XThR.Tn[12].n9 XThR.Tn[12].t71 143.911
R17242 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17243 XThR.Tn[12].n85 XThR.Tn[12].t2 26.5955
R17244 XThR.Tn[12].n85 XThR.Tn[12].t0 26.5955
R17245 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R17246 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R17247 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R17248 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R17249 XThR.Tn[12].n86 XThR.Tn[12].t3 26.5955
R17250 XThR.Tn[12].n86 XThR.Tn[12].t1 26.5955
R17251 XThR.Tn[12].n4 XThR.Tn[12].t6 24.9236
R17252 XThR.Tn[12].n4 XThR.Tn[12].t4 24.9236
R17253 XThR.Tn[12].n3 XThR.Tn[12].t7 24.9236
R17254 XThR.Tn[12].n3 XThR.Tn[12].t5 24.9236
R17255 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R17256 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R17257 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R17258 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R17259 XThR.Tn[12] XThR.Tn[12].n7 5.34038
R17260 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R17261 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R17262 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R17263 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R17264 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R17265 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R17266 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R17267 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R17268 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R17269 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R17270 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R17271 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R17272 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R17273 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R17274 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R17275 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R17276 XThR.Tn[12].n12 XThR.Tn[12] 2.52282
R17277 XThR.Tn[12].n17 XThR.Tn[12] 2.52282
R17278 XThR.Tn[12].n22 XThR.Tn[12] 2.52282
R17279 XThR.Tn[12].n27 XThR.Tn[12] 2.52282
R17280 XThR.Tn[12].n32 XThR.Tn[12] 2.52282
R17281 XThR.Tn[12].n37 XThR.Tn[12] 2.52282
R17282 XThR.Tn[12].n42 XThR.Tn[12] 2.52282
R17283 XThR.Tn[12].n47 XThR.Tn[12] 2.52282
R17284 XThR.Tn[12].n52 XThR.Tn[12] 2.52282
R17285 XThR.Tn[12].n57 XThR.Tn[12] 2.52282
R17286 XThR.Tn[12].n62 XThR.Tn[12] 2.52282
R17287 XThR.Tn[12].n67 XThR.Tn[12] 2.52282
R17288 XThR.Tn[12].n72 XThR.Tn[12] 2.52282
R17289 XThR.Tn[12].n77 XThR.Tn[12] 2.52282
R17290 XThR.Tn[12].n82 XThR.Tn[12] 2.52282
R17291 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R17292 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R17293 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R17294 XThR.Tn[12].n80 XThR.Tn[12] 1.08677
R17295 XThR.Tn[12].n75 XThR.Tn[12] 1.08677
R17296 XThR.Tn[12].n70 XThR.Tn[12] 1.08677
R17297 XThR.Tn[12].n65 XThR.Tn[12] 1.08677
R17298 XThR.Tn[12].n60 XThR.Tn[12] 1.08677
R17299 XThR.Tn[12].n55 XThR.Tn[12] 1.08677
R17300 XThR.Tn[12].n50 XThR.Tn[12] 1.08677
R17301 XThR.Tn[12].n45 XThR.Tn[12] 1.08677
R17302 XThR.Tn[12].n40 XThR.Tn[12] 1.08677
R17303 XThR.Tn[12].n35 XThR.Tn[12] 1.08677
R17304 XThR.Tn[12].n30 XThR.Tn[12] 1.08677
R17305 XThR.Tn[12].n25 XThR.Tn[12] 1.08677
R17306 XThR.Tn[12].n20 XThR.Tn[12] 1.08677
R17307 XThR.Tn[12].n15 XThR.Tn[12] 1.08677
R17308 XThR.Tn[12].n10 XThR.Tn[12] 1.08677
R17309 XThR.Tn[12] XThR.Tn[12].n12 0.839786
R17310 XThR.Tn[12] XThR.Tn[12].n17 0.839786
R17311 XThR.Tn[12] XThR.Tn[12].n22 0.839786
R17312 XThR.Tn[12] XThR.Tn[12].n27 0.839786
R17313 XThR.Tn[12] XThR.Tn[12].n32 0.839786
R17314 XThR.Tn[12] XThR.Tn[12].n37 0.839786
R17315 XThR.Tn[12] XThR.Tn[12].n42 0.839786
R17316 XThR.Tn[12] XThR.Tn[12].n47 0.839786
R17317 XThR.Tn[12] XThR.Tn[12].n52 0.839786
R17318 XThR.Tn[12] XThR.Tn[12].n57 0.839786
R17319 XThR.Tn[12] XThR.Tn[12].n62 0.839786
R17320 XThR.Tn[12] XThR.Tn[12].n67 0.839786
R17321 XThR.Tn[12] XThR.Tn[12].n72 0.839786
R17322 XThR.Tn[12] XThR.Tn[12].n77 0.839786
R17323 XThR.Tn[12] XThR.Tn[12].n82 0.839786
R17324 XThR.Tn[12].n7 XThR.Tn[12] 0.499542
R17325 XThR.Tn[12].n81 XThR.Tn[12] 0.063
R17326 XThR.Tn[12].n76 XThR.Tn[12] 0.063
R17327 XThR.Tn[12].n71 XThR.Tn[12] 0.063
R17328 XThR.Tn[12].n66 XThR.Tn[12] 0.063
R17329 XThR.Tn[12].n61 XThR.Tn[12] 0.063
R17330 XThR.Tn[12].n56 XThR.Tn[12] 0.063
R17331 XThR.Tn[12].n51 XThR.Tn[12] 0.063
R17332 XThR.Tn[12].n46 XThR.Tn[12] 0.063
R17333 XThR.Tn[12].n41 XThR.Tn[12] 0.063
R17334 XThR.Tn[12].n36 XThR.Tn[12] 0.063
R17335 XThR.Tn[12].n31 XThR.Tn[12] 0.063
R17336 XThR.Tn[12].n26 XThR.Tn[12] 0.063
R17337 XThR.Tn[12].n21 XThR.Tn[12] 0.063
R17338 XThR.Tn[12].n16 XThR.Tn[12] 0.063
R17339 XThR.Tn[12].n11 XThR.Tn[12] 0.063
R17340 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R17341 XThR.Tn[12] XThR.Tn[12].n83 0.038
R17342 XThR.Tn[12].n7 XThR.Tn[12] 0.0143889
R17343 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00771154
R17344 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00771154
R17345 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00771154
R17346 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00771154
R17347 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00771154
R17348 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00771154
R17349 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00771154
R17350 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00771154
R17351 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00771154
R17352 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00771154
R17353 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00771154
R17354 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00771154
R17355 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00771154
R17356 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00771154
R17357 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00771154
R17358 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R17359 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R17360 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R17361 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R17362 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R17363 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R17364 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R17365 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R17366 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R17367 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R17368 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R17369 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R17370 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R17371 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R17372 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R17373 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R17374 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R17375 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R17376 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R17377 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R17378 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R17379 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R17380 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R17381 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R17382 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R17383 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R17384 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R17385 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R17386 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R17387 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R17388 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R17389 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R17390 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R17391 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R17392 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R17393 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R17394 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R17395 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R17396 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R17397 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R17398 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R17399 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R17400 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R17401 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R17402 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R17403 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R17404 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R17405 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R17406 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R17407 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R17408 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R17409 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R17410 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R17411 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R17412 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R17413 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R17414 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R17415 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R17416 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R17417 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R17418 XThC.XTBN.Y.n192 XThC.XTBN.Y.n191 208.964
R17419 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R17420 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R17421 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R17422 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R17423 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R17424 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R17425 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R17426 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R17427 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R17428 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R17429 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R17430 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R17431 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R17432 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R17433 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R17434 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R17435 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R17436 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R17437 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R17438 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R17439 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R17440 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R17441 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R17442 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R17443 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R17444 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R17445 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R17446 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R17447 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R17448 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R17449 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R17450 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R17451 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R17452 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R17453 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R17454 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R17455 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R17456 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R17457 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R17458 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R17459 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R17460 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R17461 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R17462 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R17463 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R17464 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R17465 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R17466 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R17467 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R17468 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R17469 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R17470 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R17471 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R17472 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R17473 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R17474 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R17475 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R17476 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R17477 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R17478 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R17479 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R17480 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R17481 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R17482 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R17483 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R17484 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R17485 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R17486 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R17487 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R17488 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R17489 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R17490 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R17491 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R17492 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R17493 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R17494 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R17495 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R17496 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R17497 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R17498 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R17499 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R17500 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R17501 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R17502 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R17503 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R17504 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R17505 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R17506 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R17507 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R17508 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R17509 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R17510 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R17511 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R17512 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R17513 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R17514 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R17515 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R17516 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R17517 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R17518 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R17519 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R17520 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R17521 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R17522 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R17523 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R17524 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R17525 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R17526 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R17527 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R17528 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R17529 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R17530 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R17531 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R17532 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R17533 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R17534 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R17535 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R17536 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R17537 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R17538 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R17539 XThC.XTBN.Y XThC.XTBN.Y.n188 96.8352
R17540 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R17541 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R17542 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R17543 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R17544 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R17545 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R17546 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R17547 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R17548 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R17549 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R17550 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R17551 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R17552 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R17553 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R17554 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R17555 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R17556 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R17557 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R17558 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R17559 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R17560 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R17561 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R17562 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R17563 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R17564 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R17565 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R17566 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R17567 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R17568 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R17569 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R17570 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R17571 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R17572 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R17573 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R17574 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R17575 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R17576 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R17577 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R17578 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R17579 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R17580 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R17581 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R17582 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R17583 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R17584 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R17585 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R17586 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R17587 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R17588 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R17589 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R17590 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R17591 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R17592 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R17593 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R17594 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R17595 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R17596 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R17597 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R17598 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R17599 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R17600 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R17601 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R17602 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R17603 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R17604 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R17605 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R17606 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R17607 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R17608 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R17609 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R17610 XThC.XTBN.Y.n191 XThC.XTBN.Y.t0 26.5955
R17611 XThC.XTBN.Y.n191 XThC.XTBN.Y.t1 26.5955
R17612 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 24.9236
R17613 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 24.9236
R17614 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R17615 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R17616 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R17617 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R17618 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R17619 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R17620 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R17621 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R17622 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R17623 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R17624 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R17625 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R17626 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R17627 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R17628 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R17629 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R17630 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R17631 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R17632 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R17633 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R17634 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R17635 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R17636 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R17637 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R17638 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R17639 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R17640 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R17641 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R17642 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R17643 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R17644 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R17645 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R17646 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R17647 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R17648 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R17649 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R17650 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R17651 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R17652 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R17653 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R17654 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R17655 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R17656 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R17657 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R17658 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R17659 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R17660 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R17661 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R17662 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R17663 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R17664 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R17665 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R17666 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R17667 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R17668 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R17669 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R17670 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R17671 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R17672 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R17673 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R17674 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R17675 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R17676 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R17677 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R17678 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R17679 XThC.XTBN.Y XThC.XTBN.Y.n190 12.5445
R17680 XThC.XTBN.Y XThC.XTBN.Y.n189 11.2645
R17681 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R17682 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R17683 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R17684 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R17685 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R17686 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R17687 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R17688 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R17689 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R17690 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R17691 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R17692 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R17693 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R17694 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R17695 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R17696 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R17697 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R17698 XThC.XTBN.Y.n189 XThC.XTBN.Y 6.1445
R17699 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R17700 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R17701 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R17702 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R17703 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R17704 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R17705 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R17706 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R17707 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R17708 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R17709 XThC.XTBN.Y.n190 XThC.XTBN.Y 4.8645
R17710 XThC.XTBN.Y.n189 XThC.XTBN.Y 4.65505
R17711 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R17712 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R17713 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R17714 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R17715 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R17716 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R17717 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R17718 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R17719 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R17720 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R17721 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R17722 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R17723 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R17724 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R17725 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R17726 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R17727 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R17728 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R17729 XThC.XTBN.Y.n192 XThC.XTBN.Y 2.0485
R17730 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R17731 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R17732 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R17733 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R17734 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R17735 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R17736 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R17737 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R17738 XThC.XTBN.Y XThC.XTBN.Y.n192 1.55202
R17739 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R17740 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R17741 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R17742 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R17743 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R17744 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R17745 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R17746 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R17747 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R17748 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R17749 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R17750 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R17751 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R17752 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R17753 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R17754 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R17755 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R17756 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R17757 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R17758 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R17759 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R17760 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R17761 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R17762 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R17763 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R17764 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R17765 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R17766 XThC.Tn[6].n71 XThC.Tn[6].n69 161.365
R17767 XThC.Tn[6].n67 XThC.Tn[6].n65 161.365
R17768 XThC.Tn[6].n63 XThC.Tn[6].n61 161.365
R17769 XThC.Tn[6].n59 XThC.Tn[6].n57 161.365
R17770 XThC.Tn[6].n55 XThC.Tn[6].n53 161.365
R17771 XThC.Tn[6].n51 XThC.Tn[6].n49 161.365
R17772 XThC.Tn[6].n47 XThC.Tn[6].n45 161.365
R17773 XThC.Tn[6].n43 XThC.Tn[6].n41 161.365
R17774 XThC.Tn[6].n39 XThC.Tn[6].n37 161.365
R17775 XThC.Tn[6].n35 XThC.Tn[6].n33 161.365
R17776 XThC.Tn[6].n31 XThC.Tn[6].n29 161.365
R17777 XThC.Tn[6].n27 XThC.Tn[6].n25 161.365
R17778 XThC.Tn[6].n23 XThC.Tn[6].n21 161.365
R17779 XThC.Tn[6].n19 XThC.Tn[6].n17 161.365
R17780 XThC.Tn[6].n15 XThC.Tn[6].n13 161.365
R17781 XThC.Tn[6].n12 XThC.Tn[6].n10 161.365
R17782 XThC.Tn[6].n69 XThC.Tn[6].t34 161.202
R17783 XThC.Tn[6].n65 XThC.Tn[6].t24 161.202
R17784 XThC.Tn[6].n61 XThC.Tn[6].t43 161.202
R17785 XThC.Tn[6].n57 XThC.Tn[6].t41 161.202
R17786 XThC.Tn[6].n53 XThC.Tn[6].t32 161.202
R17787 XThC.Tn[6].n49 XThC.Tn[6].t21 161.202
R17788 XThC.Tn[6].n45 XThC.Tn[6].t19 161.202
R17789 XThC.Tn[6].n41 XThC.Tn[6].t31 161.202
R17790 XThC.Tn[6].n37 XThC.Tn[6].t29 161.202
R17791 XThC.Tn[6].n33 XThC.Tn[6].t22 161.202
R17792 XThC.Tn[6].n29 XThC.Tn[6].t38 161.202
R17793 XThC.Tn[6].n25 XThC.Tn[6].t37 161.202
R17794 XThC.Tn[6].n21 XThC.Tn[6].t18 161.202
R17795 XThC.Tn[6].n17 XThC.Tn[6].t17 161.202
R17796 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R17797 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R17798 XThC.Tn[6].n69 XThC.Tn[6].t30 145.137
R17799 XThC.Tn[6].n65 XThC.Tn[6].t20 145.137
R17800 XThC.Tn[6].n61 XThC.Tn[6].t39 145.137
R17801 XThC.Tn[6].n57 XThC.Tn[6].t36 145.137
R17802 XThC.Tn[6].n53 XThC.Tn[6].t28 145.137
R17803 XThC.Tn[6].n49 XThC.Tn[6].t15 145.137
R17804 XThC.Tn[6].n45 XThC.Tn[6].t14 145.137
R17805 XThC.Tn[6].n41 XThC.Tn[6].t27 145.137
R17806 XThC.Tn[6].n37 XThC.Tn[6].t25 145.137
R17807 XThC.Tn[6].n33 XThC.Tn[6].t16 145.137
R17808 XThC.Tn[6].n29 XThC.Tn[6].t35 145.137
R17809 XThC.Tn[6].n25 XThC.Tn[6].t33 145.137
R17810 XThC.Tn[6].n21 XThC.Tn[6].t12 145.137
R17811 XThC.Tn[6].n17 XThC.Tn[6].t42 145.137
R17812 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R17813 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R17814 XThC.Tn[6].n7 XThC.Tn[6].n6 135.248
R17815 XThC.Tn[6].n9 XThC.Tn[6].n3 98.982
R17816 XThC.Tn[6].n8 XThC.Tn[6].n4 98.982
R17817 XThC.Tn[6].n7 XThC.Tn[6].n5 98.982
R17818 XThC.Tn[6].n9 XThC.Tn[6].n8 36.2672
R17819 XThC.Tn[6].n8 XThC.Tn[6].n7 36.2672
R17820 XThC.Tn[6].n73 XThC.Tn[6].n9 32.6405
R17821 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R17822 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R17823 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R17824 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R17825 XThC.Tn[6].n3 XThC.Tn[6].t8 24.9236
R17826 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R17827 XThC.Tn[6].n4 XThC.Tn[6].t10 24.9236
R17828 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R17829 XThC.Tn[6].n5 XThC.Tn[6].t1 24.9236
R17830 XThC.Tn[6].n5 XThC.Tn[6].t0 24.9236
R17831 XThC.Tn[6].n6 XThC.Tn[6].t3 24.9236
R17832 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R17833 XThC.Tn[6].n74 XThC.Tn[6].n2 18.5605
R17834 XThC.Tn[6].n74 XThC.Tn[6].n73 11.5205
R17835 XThC.Tn[6] XThC.Tn[6].n12 8.0245
R17836 XThC.Tn[6].n72 XThC.Tn[6].n71 7.9105
R17837 XThC.Tn[6].n68 XThC.Tn[6].n67 7.9105
R17838 XThC.Tn[6].n64 XThC.Tn[6].n63 7.9105
R17839 XThC.Tn[6].n60 XThC.Tn[6].n59 7.9105
R17840 XThC.Tn[6].n56 XThC.Tn[6].n55 7.9105
R17841 XThC.Tn[6].n52 XThC.Tn[6].n51 7.9105
R17842 XThC.Tn[6].n48 XThC.Tn[6].n47 7.9105
R17843 XThC.Tn[6].n44 XThC.Tn[6].n43 7.9105
R17844 XThC.Tn[6].n40 XThC.Tn[6].n39 7.9105
R17845 XThC.Tn[6].n36 XThC.Tn[6].n35 7.9105
R17846 XThC.Tn[6].n32 XThC.Tn[6].n31 7.9105
R17847 XThC.Tn[6].n28 XThC.Tn[6].n27 7.9105
R17848 XThC.Tn[6].n24 XThC.Tn[6].n23 7.9105
R17849 XThC.Tn[6].n20 XThC.Tn[6].n19 7.9105
R17850 XThC.Tn[6].n16 XThC.Tn[6].n15 7.9105
R17851 XThC.Tn[6].n73 XThC.Tn[6] 5.42203
R17852 XThC.Tn[6] XThC.Tn[6].n74 0.6405
R17853 XThC.Tn[6].n16 XThC.Tn[6] 0.235138
R17854 XThC.Tn[6].n20 XThC.Tn[6] 0.235138
R17855 XThC.Tn[6].n24 XThC.Tn[6] 0.235138
R17856 XThC.Tn[6].n28 XThC.Tn[6] 0.235138
R17857 XThC.Tn[6].n32 XThC.Tn[6] 0.235138
R17858 XThC.Tn[6].n36 XThC.Tn[6] 0.235138
R17859 XThC.Tn[6].n40 XThC.Tn[6] 0.235138
R17860 XThC.Tn[6].n44 XThC.Tn[6] 0.235138
R17861 XThC.Tn[6].n48 XThC.Tn[6] 0.235138
R17862 XThC.Tn[6].n52 XThC.Tn[6] 0.235138
R17863 XThC.Tn[6].n56 XThC.Tn[6] 0.235138
R17864 XThC.Tn[6].n60 XThC.Tn[6] 0.235138
R17865 XThC.Tn[6].n64 XThC.Tn[6] 0.235138
R17866 XThC.Tn[6].n68 XThC.Tn[6] 0.235138
R17867 XThC.Tn[6].n72 XThC.Tn[6] 0.235138
R17868 XThC.Tn[6] XThC.Tn[6].n16 0.114505
R17869 XThC.Tn[6] XThC.Tn[6].n20 0.114505
R17870 XThC.Tn[6] XThC.Tn[6].n24 0.114505
R17871 XThC.Tn[6] XThC.Tn[6].n28 0.114505
R17872 XThC.Tn[6] XThC.Tn[6].n32 0.114505
R17873 XThC.Tn[6] XThC.Tn[6].n36 0.114505
R17874 XThC.Tn[6] XThC.Tn[6].n40 0.114505
R17875 XThC.Tn[6] XThC.Tn[6].n44 0.114505
R17876 XThC.Tn[6] XThC.Tn[6].n48 0.114505
R17877 XThC.Tn[6] XThC.Tn[6].n52 0.114505
R17878 XThC.Tn[6] XThC.Tn[6].n56 0.114505
R17879 XThC.Tn[6] XThC.Tn[6].n60 0.114505
R17880 XThC.Tn[6] XThC.Tn[6].n64 0.114505
R17881 XThC.Tn[6] XThC.Tn[6].n68 0.114505
R17882 XThC.Tn[6] XThC.Tn[6].n72 0.114505
R17883 XThC.Tn[6].n71 XThC.Tn[6].n70 0.0599512
R17884 XThC.Tn[6].n67 XThC.Tn[6].n66 0.0599512
R17885 XThC.Tn[6].n63 XThC.Tn[6].n62 0.0599512
R17886 XThC.Tn[6].n59 XThC.Tn[6].n58 0.0599512
R17887 XThC.Tn[6].n55 XThC.Tn[6].n54 0.0599512
R17888 XThC.Tn[6].n51 XThC.Tn[6].n50 0.0599512
R17889 XThC.Tn[6].n47 XThC.Tn[6].n46 0.0599512
R17890 XThC.Tn[6].n43 XThC.Tn[6].n42 0.0599512
R17891 XThC.Tn[6].n39 XThC.Tn[6].n38 0.0599512
R17892 XThC.Tn[6].n35 XThC.Tn[6].n34 0.0599512
R17893 XThC.Tn[6].n31 XThC.Tn[6].n30 0.0599512
R17894 XThC.Tn[6].n27 XThC.Tn[6].n26 0.0599512
R17895 XThC.Tn[6].n23 XThC.Tn[6].n22 0.0599512
R17896 XThC.Tn[6].n19 XThC.Tn[6].n18 0.0599512
R17897 XThC.Tn[6].n15 XThC.Tn[6].n14 0.0599512
R17898 XThC.Tn[6].n12 XThC.Tn[6].n11 0.0599512
R17899 XThC.Tn[6].n70 XThC.Tn[6] 0.0469286
R17900 XThC.Tn[6].n66 XThC.Tn[6] 0.0469286
R17901 XThC.Tn[6].n62 XThC.Tn[6] 0.0469286
R17902 XThC.Tn[6].n58 XThC.Tn[6] 0.0469286
R17903 XThC.Tn[6].n54 XThC.Tn[6] 0.0469286
R17904 XThC.Tn[6].n50 XThC.Tn[6] 0.0469286
R17905 XThC.Tn[6].n46 XThC.Tn[6] 0.0469286
R17906 XThC.Tn[6].n42 XThC.Tn[6] 0.0469286
R17907 XThC.Tn[6].n38 XThC.Tn[6] 0.0469286
R17908 XThC.Tn[6].n34 XThC.Tn[6] 0.0469286
R17909 XThC.Tn[6].n30 XThC.Tn[6] 0.0469286
R17910 XThC.Tn[6].n26 XThC.Tn[6] 0.0469286
R17911 XThC.Tn[6].n22 XThC.Tn[6] 0.0469286
R17912 XThC.Tn[6].n18 XThC.Tn[6] 0.0469286
R17913 XThC.Tn[6].n14 XThC.Tn[6] 0.0469286
R17914 XThC.Tn[6].n11 XThC.Tn[6] 0.0469286
R17915 XThC.Tn[6].n70 XThC.Tn[6] 0.0401341
R17916 XThC.Tn[6].n66 XThC.Tn[6] 0.0401341
R17917 XThC.Tn[6].n62 XThC.Tn[6] 0.0401341
R17918 XThC.Tn[6].n58 XThC.Tn[6] 0.0401341
R17919 XThC.Tn[6].n54 XThC.Tn[6] 0.0401341
R17920 XThC.Tn[6].n50 XThC.Tn[6] 0.0401341
R17921 XThC.Tn[6].n46 XThC.Tn[6] 0.0401341
R17922 XThC.Tn[6].n42 XThC.Tn[6] 0.0401341
R17923 XThC.Tn[6].n38 XThC.Tn[6] 0.0401341
R17924 XThC.Tn[6].n34 XThC.Tn[6] 0.0401341
R17925 XThC.Tn[6].n30 XThC.Tn[6] 0.0401341
R17926 XThC.Tn[6].n26 XThC.Tn[6] 0.0401341
R17927 XThC.Tn[6].n22 XThC.Tn[6] 0.0401341
R17928 XThC.Tn[6].n18 XThC.Tn[6] 0.0401341
R17929 XThC.Tn[6].n14 XThC.Tn[6] 0.0401341
R17930 XThC.Tn[6].n11 XThC.Tn[6] 0.0401341
R17931 XThR.Tn[9].n87 XThR.Tn[9].n86 256.103
R17932 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R17933 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R17934 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R17935 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R17936 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R17937 XThR.Tn[9] XThR.Tn[9].n78 161.363
R17938 XThR.Tn[9] XThR.Tn[9].n73 161.363
R17939 XThR.Tn[9] XThR.Tn[9].n68 161.363
R17940 XThR.Tn[9] XThR.Tn[9].n63 161.363
R17941 XThR.Tn[9] XThR.Tn[9].n58 161.363
R17942 XThR.Tn[9] XThR.Tn[9].n53 161.363
R17943 XThR.Tn[9] XThR.Tn[9].n48 161.363
R17944 XThR.Tn[9] XThR.Tn[9].n43 161.363
R17945 XThR.Tn[9] XThR.Tn[9].n38 161.363
R17946 XThR.Tn[9] XThR.Tn[9].n33 161.363
R17947 XThR.Tn[9] XThR.Tn[9].n28 161.363
R17948 XThR.Tn[9] XThR.Tn[9].n23 161.363
R17949 XThR.Tn[9] XThR.Tn[9].n18 161.363
R17950 XThR.Tn[9] XThR.Tn[9].n13 161.363
R17951 XThR.Tn[9] XThR.Tn[9].n8 161.363
R17952 XThR.Tn[9] XThR.Tn[9].n6 161.363
R17953 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R17954 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R17955 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R17956 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R17957 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R17958 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R17959 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R17960 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R17961 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R17962 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R17963 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R17964 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R17965 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R17966 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R17967 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R17968 XThR.Tn[9].n78 XThR.Tn[9].t63 161.106
R17969 XThR.Tn[9].n73 XThR.Tn[9].t69 161.106
R17970 XThR.Tn[9].n68 XThR.Tn[9].t47 161.106
R17971 XThR.Tn[9].n63 XThR.Tn[9].t34 161.106
R17972 XThR.Tn[9].n58 XThR.Tn[9].t62 161.106
R17973 XThR.Tn[9].n53 XThR.Tn[9].t24 161.106
R17974 XThR.Tn[9].n48 XThR.Tn[9].t66 161.106
R17975 XThR.Tn[9].n43 XThR.Tn[9].t45 161.106
R17976 XThR.Tn[9].n38 XThR.Tn[9].t32 161.106
R17977 XThR.Tn[9].n33 XThR.Tn[9].t37 161.106
R17978 XThR.Tn[9].n28 XThR.Tn[9].t23 161.106
R17979 XThR.Tn[9].n23 XThR.Tn[9].t46 161.106
R17980 XThR.Tn[9].n18 XThR.Tn[9].t21 161.106
R17981 XThR.Tn[9].n13 XThR.Tn[9].t64 161.106
R17982 XThR.Tn[9].n8 XThR.Tn[9].t28 161.106
R17983 XThR.Tn[9].n6 XThR.Tn[9].t71 161.106
R17984 XThR.Tn[9].n79 XThR.Tn[9].t54 159.978
R17985 XThR.Tn[9].n74 XThR.Tn[9].t61 159.978
R17986 XThR.Tn[9].n69 XThR.Tn[9].t43 159.978
R17987 XThR.Tn[9].n64 XThR.Tn[9].t27 159.978
R17988 XThR.Tn[9].n59 XThR.Tn[9].t52 159.978
R17989 XThR.Tn[9].n54 XThR.Tn[9].t18 159.978
R17990 XThR.Tn[9].n49 XThR.Tn[9].t60 159.978
R17991 XThR.Tn[9].n44 XThR.Tn[9].t40 159.978
R17992 XThR.Tn[9].n39 XThR.Tn[9].t25 159.978
R17993 XThR.Tn[9].n34 XThR.Tn[9].t33 159.978
R17994 XThR.Tn[9].n29 XThR.Tn[9].t16 159.978
R17995 XThR.Tn[9].n24 XThR.Tn[9].t42 159.978
R17996 XThR.Tn[9].n19 XThR.Tn[9].t15 159.978
R17997 XThR.Tn[9].n14 XThR.Tn[9].t59 159.978
R17998 XThR.Tn[9].n9 XThR.Tn[9].t19 159.978
R17999 XThR.Tn[9].n78 XThR.Tn[9].t49 145.038
R18000 XThR.Tn[9].n73 XThR.Tn[9].t14 145.038
R18001 XThR.Tn[9].n68 XThR.Tn[9].t57 145.038
R18002 XThR.Tn[9].n63 XThR.Tn[9].t38 145.038
R18003 XThR.Tn[9].n58 XThR.Tn[9].t70 145.038
R18004 XThR.Tn[9].n53 XThR.Tn[9].t48 145.038
R18005 XThR.Tn[9].n48 XThR.Tn[9].t58 145.038
R18006 XThR.Tn[9].n43 XThR.Tn[9].t39 145.038
R18007 XThR.Tn[9].n38 XThR.Tn[9].t36 145.038
R18008 XThR.Tn[9].n33 XThR.Tn[9].t67 145.038
R18009 XThR.Tn[9].n28 XThR.Tn[9].t31 145.038
R18010 XThR.Tn[9].n23 XThR.Tn[9].t56 145.038
R18011 XThR.Tn[9].n18 XThR.Tn[9].t29 145.038
R18012 XThR.Tn[9].n13 XThR.Tn[9].t72 145.038
R18013 XThR.Tn[9].n8 XThR.Tn[9].t35 145.038
R18014 XThR.Tn[9].n6 XThR.Tn[9].t17 145.038
R18015 XThR.Tn[9].n79 XThR.Tn[9].t68 143.911
R18016 XThR.Tn[9].n74 XThR.Tn[9].t30 143.911
R18017 XThR.Tn[9].n69 XThR.Tn[9].t12 143.911
R18018 XThR.Tn[9].n64 XThR.Tn[9].t53 143.911
R18019 XThR.Tn[9].n59 XThR.Tn[9].t22 143.911
R18020 XThR.Tn[9].n54 XThR.Tn[9].t65 143.911
R18021 XThR.Tn[9].n49 XThR.Tn[9].t13 143.911
R18022 XThR.Tn[9].n44 XThR.Tn[9].t55 143.911
R18023 XThR.Tn[9].n39 XThR.Tn[9].t51 143.911
R18024 XThR.Tn[9].n34 XThR.Tn[9].t20 143.911
R18025 XThR.Tn[9].n29 XThR.Tn[9].t44 143.911
R18026 XThR.Tn[9].n24 XThR.Tn[9].t73 143.911
R18027 XThR.Tn[9].n19 XThR.Tn[9].t41 143.911
R18028 XThR.Tn[9].n14 XThR.Tn[9].t26 143.911
R18029 XThR.Tn[9].n9 XThR.Tn[9].t50 143.911
R18030 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R18031 XThR.Tn[9].n85 XThR.Tn[9].t2 26.5955
R18032 XThR.Tn[9].n85 XThR.Tn[9].t0 26.5955
R18033 XThR.Tn[9].n0 XThR.Tn[9].t10 26.5955
R18034 XThR.Tn[9].n0 XThR.Tn[9].t8 26.5955
R18035 XThR.Tn[9].n1 XThR.Tn[9].t11 26.5955
R18036 XThR.Tn[9].n1 XThR.Tn[9].t9 26.5955
R18037 XThR.Tn[9].n86 XThR.Tn[9].t3 26.5955
R18038 XThR.Tn[9].n86 XThR.Tn[9].t1 26.5955
R18039 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R18040 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R18041 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R18042 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R18043 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R18044 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R18045 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R18046 XThR.Tn[9] XThR.Tn[9].n7 5.34038
R18047 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R18048 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R18049 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R18050 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R18051 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R18052 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R18053 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R18054 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R18055 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R18056 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R18057 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R18058 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R18059 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R18060 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R18061 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R18062 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R18063 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R18064 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R18065 XThR.Tn[9].n12 XThR.Tn[9] 2.52282
R18066 XThR.Tn[9].n17 XThR.Tn[9] 2.52282
R18067 XThR.Tn[9].n22 XThR.Tn[9] 2.52282
R18068 XThR.Tn[9].n27 XThR.Tn[9] 2.52282
R18069 XThR.Tn[9].n32 XThR.Tn[9] 2.52282
R18070 XThR.Tn[9].n37 XThR.Tn[9] 2.52282
R18071 XThR.Tn[9].n42 XThR.Tn[9] 2.52282
R18072 XThR.Tn[9].n47 XThR.Tn[9] 2.52282
R18073 XThR.Tn[9].n52 XThR.Tn[9] 2.52282
R18074 XThR.Tn[9].n57 XThR.Tn[9] 2.52282
R18075 XThR.Tn[9].n62 XThR.Tn[9] 2.52282
R18076 XThR.Tn[9].n67 XThR.Tn[9] 2.52282
R18077 XThR.Tn[9].n72 XThR.Tn[9] 2.52282
R18078 XThR.Tn[9].n77 XThR.Tn[9] 2.52282
R18079 XThR.Tn[9].n82 XThR.Tn[9] 2.52282
R18080 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R18081 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R18082 XThR.Tn[9].n80 XThR.Tn[9] 1.08677
R18083 XThR.Tn[9].n75 XThR.Tn[9] 1.08677
R18084 XThR.Tn[9].n70 XThR.Tn[9] 1.08677
R18085 XThR.Tn[9].n65 XThR.Tn[9] 1.08677
R18086 XThR.Tn[9].n60 XThR.Tn[9] 1.08677
R18087 XThR.Tn[9].n55 XThR.Tn[9] 1.08677
R18088 XThR.Tn[9].n50 XThR.Tn[9] 1.08677
R18089 XThR.Tn[9].n45 XThR.Tn[9] 1.08677
R18090 XThR.Tn[9].n40 XThR.Tn[9] 1.08677
R18091 XThR.Tn[9].n35 XThR.Tn[9] 1.08677
R18092 XThR.Tn[9].n30 XThR.Tn[9] 1.08677
R18093 XThR.Tn[9].n25 XThR.Tn[9] 1.08677
R18094 XThR.Tn[9].n20 XThR.Tn[9] 1.08677
R18095 XThR.Tn[9].n15 XThR.Tn[9] 1.08677
R18096 XThR.Tn[9].n10 XThR.Tn[9] 1.08677
R18097 XThR.Tn[9] XThR.Tn[9].n12 0.839786
R18098 XThR.Tn[9] XThR.Tn[9].n17 0.839786
R18099 XThR.Tn[9] XThR.Tn[9].n22 0.839786
R18100 XThR.Tn[9] XThR.Tn[9].n27 0.839786
R18101 XThR.Tn[9] XThR.Tn[9].n32 0.839786
R18102 XThR.Tn[9] XThR.Tn[9].n37 0.839786
R18103 XThR.Tn[9] XThR.Tn[9].n42 0.839786
R18104 XThR.Tn[9] XThR.Tn[9].n47 0.839786
R18105 XThR.Tn[9] XThR.Tn[9].n52 0.839786
R18106 XThR.Tn[9] XThR.Tn[9].n57 0.839786
R18107 XThR.Tn[9] XThR.Tn[9].n62 0.839786
R18108 XThR.Tn[9] XThR.Tn[9].n67 0.839786
R18109 XThR.Tn[9] XThR.Tn[9].n72 0.839786
R18110 XThR.Tn[9] XThR.Tn[9].n77 0.839786
R18111 XThR.Tn[9] XThR.Tn[9].n82 0.839786
R18112 XThR.Tn[9].n7 XThR.Tn[9] 0.499542
R18113 XThR.Tn[9].n81 XThR.Tn[9] 0.063
R18114 XThR.Tn[9].n76 XThR.Tn[9] 0.063
R18115 XThR.Tn[9].n71 XThR.Tn[9] 0.063
R18116 XThR.Tn[9].n66 XThR.Tn[9] 0.063
R18117 XThR.Tn[9].n61 XThR.Tn[9] 0.063
R18118 XThR.Tn[9].n56 XThR.Tn[9] 0.063
R18119 XThR.Tn[9].n51 XThR.Tn[9] 0.063
R18120 XThR.Tn[9].n46 XThR.Tn[9] 0.063
R18121 XThR.Tn[9].n41 XThR.Tn[9] 0.063
R18122 XThR.Tn[9].n36 XThR.Tn[9] 0.063
R18123 XThR.Tn[9].n31 XThR.Tn[9] 0.063
R18124 XThR.Tn[9].n26 XThR.Tn[9] 0.063
R18125 XThR.Tn[9].n21 XThR.Tn[9] 0.063
R18126 XThR.Tn[9].n16 XThR.Tn[9] 0.063
R18127 XThR.Tn[9].n11 XThR.Tn[9] 0.063
R18128 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R18129 XThR.Tn[9] XThR.Tn[9].n83 0.038
R18130 XThR.Tn[9].n7 XThR.Tn[9] 0.0143889
R18131 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00771154
R18132 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00771154
R18133 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00771154
R18134 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00771154
R18135 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00771154
R18136 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00771154
R18137 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00771154
R18138 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00771154
R18139 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00771154
R18140 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00771154
R18141 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00771154
R18142 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00771154
R18143 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00771154
R18144 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00771154
R18145 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00771154
R18146 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18147 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18148 XThC.Tn[5].n71 XThC.Tn[5].n69 161.365
R18149 XThC.Tn[5].n67 XThC.Tn[5].n65 161.365
R18150 XThC.Tn[5].n63 XThC.Tn[5].n61 161.365
R18151 XThC.Tn[5].n59 XThC.Tn[5].n57 161.365
R18152 XThC.Tn[5].n55 XThC.Tn[5].n53 161.365
R18153 XThC.Tn[5].n51 XThC.Tn[5].n49 161.365
R18154 XThC.Tn[5].n47 XThC.Tn[5].n45 161.365
R18155 XThC.Tn[5].n43 XThC.Tn[5].n41 161.365
R18156 XThC.Tn[5].n39 XThC.Tn[5].n37 161.365
R18157 XThC.Tn[5].n35 XThC.Tn[5].n33 161.365
R18158 XThC.Tn[5].n31 XThC.Tn[5].n29 161.365
R18159 XThC.Tn[5].n27 XThC.Tn[5].n25 161.365
R18160 XThC.Tn[5].n23 XThC.Tn[5].n21 161.365
R18161 XThC.Tn[5].n19 XThC.Tn[5].n17 161.365
R18162 XThC.Tn[5].n15 XThC.Tn[5].n13 161.365
R18163 XThC.Tn[5].n12 XThC.Tn[5].n10 161.365
R18164 XThC.Tn[5].n69 XThC.Tn[5].t41 161.202
R18165 XThC.Tn[5].n65 XThC.Tn[5].t30 161.202
R18166 XThC.Tn[5].n61 XThC.Tn[5].t18 161.202
R18167 XThC.Tn[5].n57 XThC.Tn[5].t16 161.202
R18168 XThC.Tn[5].n53 XThC.Tn[5].t39 161.202
R18169 XThC.Tn[5].n49 XThC.Tn[5].t26 161.202
R18170 XThC.Tn[5].n45 XThC.Tn[5].t25 161.202
R18171 XThC.Tn[5].n41 XThC.Tn[5].t37 161.202
R18172 XThC.Tn[5].n37 XThC.Tn[5].t35 161.202
R18173 XThC.Tn[5].n33 XThC.Tn[5].t27 161.202
R18174 XThC.Tn[5].n29 XThC.Tn[5].t14 161.202
R18175 XThC.Tn[5].n25 XThC.Tn[5].t13 161.202
R18176 XThC.Tn[5].n21 XThC.Tn[5].t24 161.202
R18177 XThC.Tn[5].n17 XThC.Tn[5].t23 161.202
R18178 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18179 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18180 XThC.Tn[5].n69 XThC.Tn[5].t22 145.137
R18181 XThC.Tn[5].n65 XThC.Tn[5].t12 145.137
R18182 XThC.Tn[5].n61 XThC.Tn[5].t32 145.137
R18183 XThC.Tn[5].n57 XThC.Tn[5].t31 145.137
R18184 XThC.Tn[5].n53 XThC.Tn[5].t21 145.137
R18185 XThC.Tn[5].n49 XThC.Tn[5].t42 145.137
R18186 XThC.Tn[5].n45 XThC.Tn[5].t40 145.137
R18187 XThC.Tn[5].n41 XThC.Tn[5].t20 145.137
R18188 XThC.Tn[5].n37 XThC.Tn[5].t17 145.137
R18189 XThC.Tn[5].n33 XThC.Tn[5].t43 145.137
R18190 XThC.Tn[5].n29 XThC.Tn[5].t29 145.137
R18191 XThC.Tn[5].n25 XThC.Tn[5].t28 145.137
R18192 XThC.Tn[5].n21 XThC.Tn[5].t38 145.137
R18193 XThC.Tn[5].n17 XThC.Tn[5].t36 145.137
R18194 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18195 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18196 XThC.Tn[5].n7 XThC.Tn[5].n6 135.249
R18197 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18198 XThC.Tn[5].n8 XThC.Tn[5].n4 98.981
R18199 XThC.Tn[5].n7 XThC.Tn[5].n5 98.981
R18200 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18201 XThC.Tn[5].n8 XThC.Tn[5].n7 36.2672
R18202 XThC.Tn[5].n73 XThC.Tn[5].n9 32.6405
R18203 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R18204 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R18205 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R18206 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R18207 XThC.Tn[5].n3 XThC.Tn[5].t9 24.9236
R18208 XThC.Tn[5].n3 XThC.Tn[5].t8 24.9236
R18209 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R18210 XThC.Tn[5].n4 XThC.Tn[5].t10 24.9236
R18211 XThC.Tn[5].n5 XThC.Tn[5].t2 24.9236
R18212 XThC.Tn[5].n5 XThC.Tn[5].t1 24.9236
R18213 XThC.Tn[5].n6 XThC.Tn[5].t0 24.9236
R18214 XThC.Tn[5].n6 XThC.Tn[5].t3 24.9236
R18215 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18216 XThC.Tn[5] XThC.Tn[5].n12 8.0245
R18217 XThC.Tn[5].n72 XThC.Tn[5].n71 7.9105
R18218 XThC.Tn[5].n68 XThC.Tn[5].n67 7.9105
R18219 XThC.Tn[5].n64 XThC.Tn[5].n63 7.9105
R18220 XThC.Tn[5].n60 XThC.Tn[5].n59 7.9105
R18221 XThC.Tn[5].n56 XThC.Tn[5].n55 7.9105
R18222 XThC.Tn[5].n52 XThC.Tn[5].n51 7.9105
R18223 XThC.Tn[5].n48 XThC.Tn[5].n47 7.9105
R18224 XThC.Tn[5].n44 XThC.Tn[5].n43 7.9105
R18225 XThC.Tn[5].n40 XThC.Tn[5].n39 7.9105
R18226 XThC.Tn[5].n36 XThC.Tn[5].n35 7.9105
R18227 XThC.Tn[5].n32 XThC.Tn[5].n31 7.9105
R18228 XThC.Tn[5].n28 XThC.Tn[5].n27 7.9105
R18229 XThC.Tn[5].n24 XThC.Tn[5].n23 7.9105
R18230 XThC.Tn[5].n20 XThC.Tn[5].n19 7.9105
R18231 XThC.Tn[5].n16 XThC.Tn[5].n15 7.9105
R18232 XThC.Tn[5] XThC.Tn[5].n73 6.7205
R18233 XThC.Tn[5].n73 XThC.Tn[5] 5.69842
R18234 XThC.Tn[5].n16 XThC.Tn[5] 0.235138
R18235 XThC.Tn[5].n20 XThC.Tn[5] 0.235138
R18236 XThC.Tn[5].n24 XThC.Tn[5] 0.235138
R18237 XThC.Tn[5].n28 XThC.Tn[5] 0.235138
R18238 XThC.Tn[5].n32 XThC.Tn[5] 0.235138
R18239 XThC.Tn[5].n36 XThC.Tn[5] 0.235138
R18240 XThC.Tn[5].n40 XThC.Tn[5] 0.235138
R18241 XThC.Tn[5].n44 XThC.Tn[5] 0.235138
R18242 XThC.Tn[5].n48 XThC.Tn[5] 0.235138
R18243 XThC.Tn[5].n52 XThC.Tn[5] 0.235138
R18244 XThC.Tn[5].n56 XThC.Tn[5] 0.235138
R18245 XThC.Tn[5].n60 XThC.Tn[5] 0.235138
R18246 XThC.Tn[5].n64 XThC.Tn[5] 0.235138
R18247 XThC.Tn[5].n68 XThC.Tn[5] 0.235138
R18248 XThC.Tn[5].n72 XThC.Tn[5] 0.235138
R18249 XThC.Tn[5] XThC.Tn[5].n16 0.114505
R18250 XThC.Tn[5] XThC.Tn[5].n20 0.114505
R18251 XThC.Tn[5] XThC.Tn[5].n24 0.114505
R18252 XThC.Tn[5] XThC.Tn[5].n28 0.114505
R18253 XThC.Tn[5] XThC.Tn[5].n32 0.114505
R18254 XThC.Tn[5] XThC.Tn[5].n36 0.114505
R18255 XThC.Tn[5] XThC.Tn[5].n40 0.114505
R18256 XThC.Tn[5] XThC.Tn[5].n44 0.114505
R18257 XThC.Tn[5] XThC.Tn[5].n48 0.114505
R18258 XThC.Tn[5] XThC.Tn[5].n52 0.114505
R18259 XThC.Tn[5] XThC.Tn[5].n56 0.114505
R18260 XThC.Tn[5] XThC.Tn[5].n60 0.114505
R18261 XThC.Tn[5] XThC.Tn[5].n64 0.114505
R18262 XThC.Tn[5] XThC.Tn[5].n68 0.114505
R18263 XThC.Tn[5] XThC.Tn[5].n72 0.114505
R18264 XThC.Tn[5].n71 XThC.Tn[5].n70 0.0599512
R18265 XThC.Tn[5].n67 XThC.Tn[5].n66 0.0599512
R18266 XThC.Tn[5].n63 XThC.Tn[5].n62 0.0599512
R18267 XThC.Tn[5].n59 XThC.Tn[5].n58 0.0599512
R18268 XThC.Tn[5].n55 XThC.Tn[5].n54 0.0599512
R18269 XThC.Tn[5].n51 XThC.Tn[5].n50 0.0599512
R18270 XThC.Tn[5].n47 XThC.Tn[5].n46 0.0599512
R18271 XThC.Tn[5].n43 XThC.Tn[5].n42 0.0599512
R18272 XThC.Tn[5].n39 XThC.Tn[5].n38 0.0599512
R18273 XThC.Tn[5].n35 XThC.Tn[5].n34 0.0599512
R18274 XThC.Tn[5].n31 XThC.Tn[5].n30 0.0599512
R18275 XThC.Tn[5].n27 XThC.Tn[5].n26 0.0599512
R18276 XThC.Tn[5].n23 XThC.Tn[5].n22 0.0599512
R18277 XThC.Tn[5].n19 XThC.Tn[5].n18 0.0599512
R18278 XThC.Tn[5].n15 XThC.Tn[5].n14 0.0599512
R18279 XThC.Tn[5].n12 XThC.Tn[5].n11 0.0599512
R18280 XThC.Tn[5].n70 XThC.Tn[5] 0.0469286
R18281 XThC.Tn[5].n66 XThC.Tn[5] 0.0469286
R18282 XThC.Tn[5].n62 XThC.Tn[5] 0.0469286
R18283 XThC.Tn[5].n58 XThC.Tn[5] 0.0469286
R18284 XThC.Tn[5].n54 XThC.Tn[5] 0.0469286
R18285 XThC.Tn[5].n50 XThC.Tn[5] 0.0469286
R18286 XThC.Tn[5].n46 XThC.Tn[5] 0.0469286
R18287 XThC.Tn[5].n42 XThC.Tn[5] 0.0469286
R18288 XThC.Tn[5].n38 XThC.Tn[5] 0.0469286
R18289 XThC.Tn[5].n34 XThC.Tn[5] 0.0469286
R18290 XThC.Tn[5].n30 XThC.Tn[5] 0.0469286
R18291 XThC.Tn[5].n26 XThC.Tn[5] 0.0469286
R18292 XThC.Tn[5].n22 XThC.Tn[5] 0.0469286
R18293 XThC.Tn[5].n18 XThC.Tn[5] 0.0469286
R18294 XThC.Tn[5].n14 XThC.Tn[5] 0.0469286
R18295 XThC.Tn[5].n11 XThC.Tn[5] 0.0469286
R18296 XThC.Tn[5].n70 XThC.Tn[5] 0.0401341
R18297 XThC.Tn[5].n66 XThC.Tn[5] 0.0401341
R18298 XThC.Tn[5].n62 XThC.Tn[5] 0.0401341
R18299 XThC.Tn[5].n58 XThC.Tn[5] 0.0401341
R18300 XThC.Tn[5].n54 XThC.Tn[5] 0.0401341
R18301 XThC.Tn[5].n50 XThC.Tn[5] 0.0401341
R18302 XThC.Tn[5].n46 XThC.Tn[5] 0.0401341
R18303 XThC.Tn[5].n42 XThC.Tn[5] 0.0401341
R18304 XThC.Tn[5].n38 XThC.Tn[5] 0.0401341
R18305 XThC.Tn[5].n34 XThC.Tn[5] 0.0401341
R18306 XThC.Tn[5].n30 XThC.Tn[5] 0.0401341
R18307 XThC.Tn[5].n26 XThC.Tn[5] 0.0401341
R18308 XThC.Tn[5].n22 XThC.Tn[5] 0.0401341
R18309 XThC.Tn[5].n18 XThC.Tn[5] 0.0401341
R18310 XThC.Tn[5].n14 XThC.Tn[5] 0.0401341
R18311 XThC.Tn[5].n11 XThC.Tn[5] 0.0401341
R18312 XThC.Tn[9].n70 XThC.Tn[9].n69 265.341
R18313 XThC.Tn[9].n74 XThC.Tn[9].n72 243.68
R18314 XThC.Tn[9].n2 XThC.Tn[9].n0 241.847
R18315 XThC.Tn[9].n74 XThC.Tn[9].n73 205.28
R18316 XThC.Tn[9].n70 XThC.Tn[9].n68 202.094
R18317 XThC.Tn[9].n2 XThC.Tn[9].n1 185
R18318 XThC.Tn[9].n64 XThC.Tn[9].n62 161.365
R18319 XThC.Tn[9].n60 XThC.Tn[9].n58 161.365
R18320 XThC.Tn[9].n56 XThC.Tn[9].n54 161.365
R18321 XThC.Tn[9].n52 XThC.Tn[9].n50 161.365
R18322 XThC.Tn[9].n48 XThC.Tn[9].n46 161.365
R18323 XThC.Tn[9].n44 XThC.Tn[9].n42 161.365
R18324 XThC.Tn[9].n40 XThC.Tn[9].n38 161.365
R18325 XThC.Tn[9].n36 XThC.Tn[9].n34 161.365
R18326 XThC.Tn[9].n32 XThC.Tn[9].n30 161.365
R18327 XThC.Tn[9].n28 XThC.Tn[9].n26 161.365
R18328 XThC.Tn[9].n24 XThC.Tn[9].n22 161.365
R18329 XThC.Tn[9].n20 XThC.Tn[9].n18 161.365
R18330 XThC.Tn[9].n16 XThC.Tn[9].n14 161.365
R18331 XThC.Tn[9].n12 XThC.Tn[9].n10 161.365
R18332 XThC.Tn[9].n8 XThC.Tn[9].n6 161.365
R18333 XThC.Tn[9].n5 XThC.Tn[9].n3 161.365
R18334 XThC.Tn[9].n62 XThC.Tn[9].t20 161.202
R18335 XThC.Tn[9].n58 XThC.Tn[9].t41 161.202
R18336 XThC.Tn[9].n54 XThC.Tn[9].t29 161.202
R18337 XThC.Tn[9].n50 XThC.Tn[9].t27 161.202
R18338 XThC.Tn[9].n46 XThC.Tn[9].t18 161.202
R18339 XThC.Tn[9].n42 XThC.Tn[9].t37 161.202
R18340 XThC.Tn[9].n38 XThC.Tn[9].t36 161.202
R18341 XThC.Tn[9].n34 XThC.Tn[9].t16 161.202
R18342 XThC.Tn[9].n30 XThC.Tn[9].t14 161.202
R18343 XThC.Tn[9].n26 XThC.Tn[9].t38 161.202
R18344 XThC.Tn[9].n22 XThC.Tn[9].t25 161.202
R18345 XThC.Tn[9].n18 XThC.Tn[9].t24 161.202
R18346 XThC.Tn[9].n14 XThC.Tn[9].t35 161.202
R18347 XThC.Tn[9].n10 XThC.Tn[9].t34 161.202
R18348 XThC.Tn[9].n6 XThC.Tn[9].t30 161.202
R18349 XThC.Tn[9].n3 XThC.Tn[9].t12 161.202
R18350 XThC.Tn[9].n62 XThC.Tn[9].t33 145.137
R18351 XThC.Tn[9].n58 XThC.Tn[9].t23 145.137
R18352 XThC.Tn[9].n54 XThC.Tn[9].t43 145.137
R18353 XThC.Tn[9].n50 XThC.Tn[9].t42 145.137
R18354 XThC.Tn[9].n46 XThC.Tn[9].t32 145.137
R18355 XThC.Tn[9].n42 XThC.Tn[9].t21 145.137
R18356 XThC.Tn[9].n38 XThC.Tn[9].t19 145.137
R18357 XThC.Tn[9].n34 XThC.Tn[9].t31 145.137
R18358 XThC.Tn[9].n30 XThC.Tn[9].t28 145.137
R18359 XThC.Tn[9].n26 XThC.Tn[9].t22 145.137
R18360 XThC.Tn[9].n22 XThC.Tn[9].t40 145.137
R18361 XThC.Tn[9].n18 XThC.Tn[9].t39 145.137
R18362 XThC.Tn[9].n14 XThC.Tn[9].t17 145.137
R18363 XThC.Tn[9].n10 XThC.Tn[9].t15 145.137
R18364 XThC.Tn[9].n6 XThC.Tn[9].t13 145.137
R18365 XThC.Tn[9].n3 XThC.Tn[9].t26 145.137
R18366 XThC.Tn[9].n72 XThC.Tn[9].t1 26.5955
R18367 XThC.Tn[9].n72 XThC.Tn[9].t0 26.5955
R18368 XThC.Tn[9].n69 XThC.Tn[9].t6 26.5955
R18369 XThC.Tn[9].n69 XThC.Tn[9].t5 26.5955
R18370 XThC.Tn[9].n68 XThC.Tn[9].t4 26.5955
R18371 XThC.Tn[9].n68 XThC.Tn[9].t7 26.5955
R18372 XThC.Tn[9].n73 XThC.Tn[9].t3 26.5955
R18373 XThC.Tn[9].n73 XThC.Tn[9].t2 26.5955
R18374 XThC.Tn[9].n1 XThC.Tn[9].t10 24.9236
R18375 XThC.Tn[9].n1 XThC.Tn[9].t11 24.9236
R18376 XThC.Tn[9].n0 XThC.Tn[9].t9 24.9236
R18377 XThC.Tn[9].n0 XThC.Tn[9].t8 24.9236
R18378 XThC.Tn[9] XThC.Tn[9].n74 22.9652
R18379 XThC.Tn[9] XThC.Tn[9].n2 18.8943
R18380 XThC.Tn[9].n71 XThC.Tn[9].n70 13.9299
R18381 XThC.Tn[9] XThC.Tn[9].n71 13.9299
R18382 XThC.Tn[9] XThC.Tn[9].n5 8.0245
R18383 XThC.Tn[9].n65 XThC.Tn[9].n64 7.9105
R18384 XThC.Tn[9].n61 XThC.Tn[9].n60 7.9105
R18385 XThC.Tn[9].n57 XThC.Tn[9].n56 7.9105
R18386 XThC.Tn[9].n53 XThC.Tn[9].n52 7.9105
R18387 XThC.Tn[9].n49 XThC.Tn[9].n48 7.9105
R18388 XThC.Tn[9].n45 XThC.Tn[9].n44 7.9105
R18389 XThC.Tn[9].n41 XThC.Tn[9].n40 7.9105
R18390 XThC.Tn[9].n37 XThC.Tn[9].n36 7.9105
R18391 XThC.Tn[9].n33 XThC.Tn[9].n32 7.9105
R18392 XThC.Tn[9].n29 XThC.Tn[9].n28 7.9105
R18393 XThC.Tn[9].n25 XThC.Tn[9].n24 7.9105
R18394 XThC.Tn[9].n21 XThC.Tn[9].n20 7.9105
R18395 XThC.Tn[9].n17 XThC.Tn[9].n16 7.9105
R18396 XThC.Tn[9].n13 XThC.Tn[9].n12 7.9105
R18397 XThC.Tn[9].n9 XThC.Tn[9].n8 7.9105
R18398 XThC.Tn[9].n67 XThC.Tn[9].n66 7.44831
R18399 XThC.Tn[9].n67 XThC.Tn[9] 6.34069
R18400 XThC.Tn[9].n66 XThC.Tn[9] 4.25199
R18401 XThC.Tn[9] XThC.Tn[9].n67 1.79489
R18402 XThC.Tn[9].n71 XThC.Tn[9] 1.19676
R18403 XThC.Tn[9].n66 XThC.Tn[9] 0.657022
R18404 XThC.Tn[9].n9 XThC.Tn[9] 0.235138
R18405 XThC.Tn[9].n13 XThC.Tn[9] 0.235138
R18406 XThC.Tn[9].n17 XThC.Tn[9] 0.235138
R18407 XThC.Tn[9].n21 XThC.Tn[9] 0.235138
R18408 XThC.Tn[9].n25 XThC.Tn[9] 0.235138
R18409 XThC.Tn[9].n29 XThC.Tn[9] 0.235138
R18410 XThC.Tn[9].n33 XThC.Tn[9] 0.235138
R18411 XThC.Tn[9].n37 XThC.Tn[9] 0.235138
R18412 XThC.Tn[9].n41 XThC.Tn[9] 0.235138
R18413 XThC.Tn[9].n45 XThC.Tn[9] 0.235138
R18414 XThC.Tn[9].n49 XThC.Tn[9] 0.235138
R18415 XThC.Tn[9].n53 XThC.Tn[9] 0.235138
R18416 XThC.Tn[9].n57 XThC.Tn[9] 0.235138
R18417 XThC.Tn[9].n61 XThC.Tn[9] 0.235138
R18418 XThC.Tn[9].n65 XThC.Tn[9] 0.235138
R18419 XThC.Tn[9] XThC.Tn[9].n9 0.114505
R18420 XThC.Tn[9] XThC.Tn[9].n13 0.114505
R18421 XThC.Tn[9] XThC.Tn[9].n17 0.114505
R18422 XThC.Tn[9] XThC.Tn[9].n21 0.114505
R18423 XThC.Tn[9] XThC.Tn[9].n25 0.114505
R18424 XThC.Tn[9] XThC.Tn[9].n29 0.114505
R18425 XThC.Tn[9] XThC.Tn[9].n33 0.114505
R18426 XThC.Tn[9] XThC.Tn[9].n37 0.114505
R18427 XThC.Tn[9] XThC.Tn[9].n41 0.114505
R18428 XThC.Tn[9] XThC.Tn[9].n45 0.114505
R18429 XThC.Tn[9] XThC.Tn[9].n49 0.114505
R18430 XThC.Tn[9] XThC.Tn[9].n53 0.114505
R18431 XThC.Tn[9] XThC.Tn[9].n57 0.114505
R18432 XThC.Tn[9] XThC.Tn[9].n61 0.114505
R18433 XThC.Tn[9] XThC.Tn[9].n65 0.114505
R18434 XThC.Tn[9].n64 XThC.Tn[9].n63 0.0599512
R18435 XThC.Tn[9].n60 XThC.Tn[9].n59 0.0599512
R18436 XThC.Tn[9].n56 XThC.Tn[9].n55 0.0599512
R18437 XThC.Tn[9].n52 XThC.Tn[9].n51 0.0599512
R18438 XThC.Tn[9].n48 XThC.Tn[9].n47 0.0599512
R18439 XThC.Tn[9].n44 XThC.Tn[9].n43 0.0599512
R18440 XThC.Tn[9].n40 XThC.Tn[9].n39 0.0599512
R18441 XThC.Tn[9].n36 XThC.Tn[9].n35 0.0599512
R18442 XThC.Tn[9].n32 XThC.Tn[9].n31 0.0599512
R18443 XThC.Tn[9].n28 XThC.Tn[9].n27 0.0599512
R18444 XThC.Tn[9].n24 XThC.Tn[9].n23 0.0599512
R18445 XThC.Tn[9].n20 XThC.Tn[9].n19 0.0599512
R18446 XThC.Tn[9].n16 XThC.Tn[9].n15 0.0599512
R18447 XThC.Tn[9].n12 XThC.Tn[9].n11 0.0599512
R18448 XThC.Tn[9].n8 XThC.Tn[9].n7 0.0599512
R18449 XThC.Tn[9].n5 XThC.Tn[9].n4 0.0599512
R18450 XThC.Tn[9].n63 XThC.Tn[9] 0.0469286
R18451 XThC.Tn[9].n59 XThC.Tn[9] 0.0469286
R18452 XThC.Tn[9].n55 XThC.Tn[9] 0.0469286
R18453 XThC.Tn[9].n51 XThC.Tn[9] 0.0469286
R18454 XThC.Tn[9].n47 XThC.Tn[9] 0.0469286
R18455 XThC.Tn[9].n43 XThC.Tn[9] 0.0469286
R18456 XThC.Tn[9].n39 XThC.Tn[9] 0.0469286
R18457 XThC.Tn[9].n35 XThC.Tn[9] 0.0469286
R18458 XThC.Tn[9].n31 XThC.Tn[9] 0.0469286
R18459 XThC.Tn[9].n27 XThC.Tn[9] 0.0469286
R18460 XThC.Tn[9].n23 XThC.Tn[9] 0.0469286
R18461 XThC.Tn[9].n19 XThC.Tn[9] 0.0469286
R18462 XThC.Tn[9].n15 XThC.Tn[9] 0.0469286
R18463 XThC.Tn[9].n11 XThC.Tn[9] 0.0469286
R18464 XThC.Tn[9].n7 XThC.Tn[9] 0.0469286
R18465 XThC.Tn[9].n4 XThC.Tn[9] 0.0469286
R18466 XThC.Tn[9].n63 XThC.Tn[9] 0.0401341
R18467 XThC.Tn[9].n59 XThC.Tn[9] 0.0401341
R18468 XThC.Tn[9].n55 XThC.Tn[9] 0.0401341
R18469 XThC.Tn[9].n51 XThC.Tn[9] 0.0401341
R18470 XThC.Tn[9].n47 XThC.Tn[9] 0.0401341
R18471 XThC.Tn[9].n43 XThC.Tn[9] 0.0401341
R18472 XThC.Tn[9].n39 XThC.Tn[9] 0.0401341
R18473 XThC.Tn[9].n35 XThC.Tn[9] 0.0401341
R18474 XThC.Tn[9].n31 XThC.Tn[9] 0.0401341
R18475 XThC.Tn[9].n27 XThC.Tn[9] 0.0401341
R18476 XThC.Tn[9].n23 XThC.Tn[9] 0.0401341
R18477 XThC.Tn[9].n19 XThC.Tn[9] 0.0401341
R18478 XThC.Tn[9].n15 XThC.Tn[9] 0.0401341
R18479 XThC.Tn[9].n11 XThC.Tn[9] 0.0401341
R18480 XThC.Tn[9].n7 XThC.Tn[9] 0.0401341
R18481 XThC.Tn[9].n4 XThC.Tn[9] 0.0401341
R18482 XThC.Tn[11].n70 XThC.Tn[11].n69 265.341
R18483 XThC.Tn[11].n74 XThC.Tn[11].n73 243.68
R18484 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R18485 XThC.Tn[11].n74 XThC.Tn[11].n72 205.28
R18486 XThC.Tn[11].n70 XThC.Tn[11].n68 202.094
R18487 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R18488 XThC.Tn[11].n64 XThC.Tn[11].n62 161.365
R18489 XThC.Tn[11].n60 XThC.Tn[11].n58 161.365
R18490 XThC.Tn[11].n56 XThC.Tn[11].n54 161.365
R18491 XThC.Tn[11].n52 XThC.Tn[11].n50 161.365
R18492 XThC.Tn[11].n48 XThC.Tn[11].n46 161.365
R18493 XThC.Tn[11].n44 XThC.Tn[11].n42 161.365
R18494 XThC.Tn[11].n40 XThC.Tn[11].n38 161.365
R18495 XThC.Tn[11].n36 XThC.Tn[11].n34 161.365
R18496 XThC.Tn[11].n32 XThC.Tn[11].n30 161.365
R18497 XThC.Tn[11].n28 XThC.Tn[11].n26 161.365
R18498 XThC.Tn[11].n24 XThC.Tn[11].n22 161.365
R18499 XThC.Tn[11].n20 XThC.Tn[11].n18 161.365
R18500 XThC.Tn[11].n16 XThC.Tn[11].n14 161.365
R18501 XThC.Tn[11].n12 XThC.Tn[11].n10 161.365
R18502 XThC.Tn[11].n8 XThC.Tn[11].n6 161.365
R18503 XThC.Tn[11].n5 XThC.Tn[11].n3 161.365
R18504 XThC.Tn[11].n62 XThC.Tn[11].t24 161.202
R18505 XThC.Tn[11].n58 XThC.Tn[11].t14 161.202
R18506 XThC.Tn[11].n54 XThC.Tn[11].t33 161.202
R18507 XThC.Tn[11].n50 XThC.Tn[11].t30 161.202
R18508 XThC.Tn[11].n46 XThC.Tn[11].t22 161.202
R18509 XThC.Tn[11].n42 XThC.Tn[11].t41 161.202
R18510 XThC.Tn[11].n38 XThC.Tn[11].t40 161.202
R18511 XThC.Tn[11].n34 XThC.Tn[11].t21 161.202
R18512 XThC.Tn[11].n30 XThC.Tn[11].t19 161.202
R18513 XThC.Tn[11].n26 XThC.Tn[11].t42 161.202
R18514 XThC.Tn[11].n22 XThC.Tn[11].t29 161.202
R18515 XThC.Tn[11].n18 XThC.Tn[11].t28 161.202
R18516 XThC.Tn[11].n14 XThC.Tn[11].t39 161.202
R18517 XThC.Tn[11].n10 XThC.Tn[11].t37 161.202
R18518 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R18519 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R18520 XThC.Tn[11].n62 XThC.Tn[11].t27 145.137
R18521 XThC.Tn[11].n58 XThC.Tn[11].t17 145.137
R18522 XThC.Tn[11].n54 XThC.Tn[11].t36 145.137
R18523 XThC.Tn[11].n50 XThC.Tn[11].t34 145.137
R18524 XThC.Tn[11].n46 XThC.Tn[11].t26 145.137
R18525 XThC.Tn[11].n42 XThC.Tn[11].t15 145.137
R18526 XThC.Tn[11].n38 XThC.Tn[11].t13 145.137
R18527 XThC.Tn[11].n34 XThC.Tn[11].t25 145.137
R18528 XThC.Tn[11].n30 XThC.Tn[11].t23 145.137
R18529 XThC.Tn[11].n26 XThC.Tn[11].t16 145.137
R18530 XThC.Tn[11].n22 XThC.Tn[11].t32 145.137
R18531 XThC.Tn[11].n18 XThC.Tn[11].t31 145.137
R18532 XThC.Tn[11].n14 XThC.Tn[11].t12 145.137
R18533 XThC.Tn[11].n10 XThC.Tn[11].t43 145.137
R18534 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R18535 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R18536 XThC.Tn[11].n69 XThC.Tn[11].t6 26.5955
R18537 XThC.Tn[11].n69 XThC.Tn[11].t8 26.5955
R18538 XThC.Tn[11].n68 XThC.Tn[11].t4 26.5955
R18539 XThC.Tn[11].n68 XThC.Tn[11].t9 26.5955
R18540 XThC.Tn[11].n72 XThC.Tn[11].t2 26.5955
R18541 XThC.Tn[11].n72 XThC.Tn[11].t1 26.5955
R18542 XThC.Tn[11].n73 XThC.Tn[11].t0 26.5955
R18543 XThC.Tn[11].n73 XThC.Tn[11].t3 26.5955
R18544 XThC.Tn[11].n1 XThC.Tn[11].t5 24.9236
R18545 XThC.Tn[11].n1 XThC.Tn[11].t11 24.9236
R18546 XThC.Tn[11].n0 XThC.Tn[11].t7 24.9236
R18547 XThC.Tn[11].n0 XThC.Tn[11].t10 24.9236
R18548 XThC.Tn[11] XThC.Tn[11].n74 22.9652
R18549 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R18550 XThC.Tn[11].n71 XThC.Tn[11].n70 13.9299
R18551 XThC.Tn[11] XThC.Tn[11].n71 13.9299
R18552 XThC.Tn[11] XThC.Tn[11].n5 8.0245
R18553 XThC.Tn[11].n65 XThC.Tn[11].n64 7.9105
R18554 XThC.Tn[11].n61 XThC.Tn[11].n60 7.9105
R18555 XThC.Tn[11].n57 XThC.Tn[11].n56 7.9105
R18556 XThC.Tn[11].n53 XThC.Tn[11].n52 7.9105
R18557 XThC.Tn[11].n49 XThC.Tn[11].n48 7.9105
R18558 XThC.Tn[11].n45 XThC.Tn[11].n44 7.9105
R18559 XThC.Tn[11].n41 XThC.Tn[11].n40 7.9105
R18560 XThC.Tn[11].n37 XThC.Tn[11].n36 7.9105
R18561 XThC.Tn[11].n33 XThC.Tn[11].n32 7.9105
R18562 XThC.Tn[11].n29 XThC.Tn[11].n28 7.9105
R18563 XThC.Tn[11].n25 XThC.Tn[11].n24 7.9105
R18564 XThC.Tn[11].n21 XThC.Tn[11].n20 7.9105
R18565 XThC.Tn[11].n17 XThC.Tn[11].n16 7.9105
R18566 XThC.Tn[11].n13 XThC.Tn[11].n12 7.9105
R18567 XThC.Tn[11].n9 XThC.Tn[11].n8 7.9105
R18568 XThC.Tn[11].n67 XThC.Tn[11].n66 7.44831
R18569 XThC.Tn[11].n67 XThC.Tn[11] 6.34069
R18570 XThC.Tn[11].n66 XThC.Tn[11] 4.37928
R18571 XThC.Tn[11] XThC.Tn[11].n67 1.79489
R18572 XThC.Tn[11].n71 XThC.Tn[11] 1.19676
R18573 XThC.Tn[11].n66 XThC.Tn[11] 1.0918
R18574 XThC.Tn[11].n9 XThC.Tn[11] 0.235138
R18575 XThC.Tn[11].n13 XThC.Tn[11] 0.235138
R18576 XThC.Tn[11].n17 XThC.Tn[11] 0.235138
R18577 XThC.Tn[11].n21 XThC.Tn[11] 0.235138
R18578 XThC.Tn[11].n25 XThC.Tn[11] 0.235138
R18579 XThC.Tn[11].n29 XThC.Tn[11] 0.235138
R18580 XThC.Tn[11].n33 XThC.Tn[11] 0.235138
R18581 XThC.Tn[11].n37 XThC.Tn[11] 0.235138
R18582 XThC.Tn[11].n41 XThC.Tn[11] 0.235138
R18583 XThC.Tn[11].n45 XThC.Tn[11] 0.235138
R18584 XThC.Tn[11].n49 XThC.Tn[11] 0.235138
R18585 XThC.Tn[11].n53 XThC.Tn[11] 0.235138
R18586 XThC.Tn[11].n57 XThC.Tn[11] 0.235138
R18587 XThC.Tn[11].n61 XThC.Tn[11] 0.235138
R18588 XThC.Tn[11].n65 XThC.Tn[11] 0.235138
R18589 XThC.Tn[11] XThC.Tn[11].n9 0.114505
R18590 XThC.Tn[11] XThC.Tn[11].n13 0.114505
R18591 XThC.Tn[11] XThC.Tn[11].n17 0.114505
R18592 XThC.Tn[11] XThC.Tn[11].n21 0.114505
R18593 XThC.Tn[11] XThC.Tn[11].n25 0.114505
R18594 XThC.Tn[11] XThC.Tn[11].n29 0.114505
R18595 XThC.Tn[11] XThC.Tn[11].n33 0.114505
R18596 XThC.Tn[11] XThC.Tn[11].n37 0.114505
R18597 XThC.Tn[11] XThC.Tn[11].n41 0.114505
R18598 XThC.Tn[11] XThC.Tn[11].n45 0.114505
R18599 XThC.Tn[11] XThC.Tn[11].n49 0.114505
R18600 XThC.Tn[11] XThC.Tn[11].n53 0.114505
R18601 XThC.Tn[11] XThC.Tn[11].n57 0.114505
R18602 XThC.Tn[11] XThC.Tn[11].n61 0.114505
R18603 XThC.Tn[11] XThC.Tn[11].n65 0.114505
R18604 XThC.Tn[11].n64 XThC.Tn[11].n63 0.0599512
R18605 XThC.Tn[11].n60 XThC.Tn[11].n59 0.0599512
R18606 XThC.Tn[11].n56 XThC.Tn[11].n55 0.0599512
R18607 XThC.Tn[11].n52 XThC.Tn[11].n51 0.0599512
R18608 XThC.Tn[11].n48 XThC.Tn[11].n47 0.0599512
R18609 XThC.Tn[11].n44 XThC.Tn[11].n43 0.0599512
R18610 XThC.Tn[11].n40 XThC.Tn[11].n39 0.0599512
R18611 XThC.Tn[11].n36 XThC.Tn[11].n35 0.0599512
R18612 XThC.Tn[11].n32 XThC.Tn[11].n31 0.0599512
R18613 XThC.Tn[11].n28 XThC.Tn[11].n27 0.0599512
R18614 XThC.Tn[11].n24 XThC.Tn[11].n23 0.0599512
R18615 XThC.Tn[11].n20 XThC.Tn[11].n19 0.0599512
R18616 XThC.Tn[11].n16 XThC.Tn[11].n15 0.0599512
R18617 XThC.Tn[11].n12 XThC.Tn[11].n11 0.0599512
R18618 XThC.Tn[11].n8 XThC.Tn[11].n7 0.0599512
R18619 XThC.Tn[11].n5 XThC.Tn[11].n4 0.0599512
R18620 XThC.Tn[11].n63 XThC.Tn[11] 0.0469286
R18621 XThC.Tn[11].n59 XThC.Tn[11] 0.0469286
R18622 XThC.Tn[11].n55 XThC.Tn[11] 0.0469286
R18623 XThC.Tn[11].n51 XThC.Tn[11] 0.0469286
R18624 XThC.Tn[11].n47 XThC.Tn[11] 0.0469286
R18625 XThC.Tn[11].n43 XThC.Tn[11] 0.0469286
R18626 XThC.Tn[11].n39 XThC.Tn[11] 0.0469286
R18627 XThC.Tn[11].n35 XThC.Tn[11] 0.0469286
R18628 XThC.Tn[11].n31 XThC.Tn[11] 0.0469286
R18629 XThC.Tn[11].n27 XThC.Tn[11] 0.0469286
R18630 XThC.Tn[11].n23 XThC.Tn[11] 0.0469286
R18631 XThC.Tn[11].n19 XThC.Tn[11] 0.0469286
R18632 XThC.Tn[11].n15 XThC.Tn[11] 0.0469286
R18633 XThC.Tn[11].n11 XThC.Tn[11] 0.0469286
R18634 XThC.Tn[11].n7 XThC.Tn[11] 0.0469286
R18635 XThC.Tn[11].n4 XThC.Tn[11] 0.0469286
R18636 XThC.Tn[11].n63 XThC.Tn[11] 0.0401341
R18637 XThC.Tn[11].n59 XThC.Tn[11] 0.0401341
R18638 XThC.Tn[11].n55 XThC.Tn[11] 0.0401341
R18639 XThC.Tn[11].n51 XThC.Tn[11] 0.0401341
R18640 XThC.Tn[11].n47 XThC.Tn[11] 0.0401341
R18641 XThC.Tn[11].n43 XThC.Tn[11] 0.0401341
R18642 XThC.Tn[11].n39 XThC.Tn[11] 0.0401341
R18643 XThC.Tn[11].n35 XThC.Tn[11] 0.0401341
R18644 XThC.Tn[11].n31 XThC.Tn[11] 0.0401341
R18645 XThC.Tn[11].n27 XThC.Tn[11] 0.0401341
R18646 XThC.Tn[11].n23 XThC.Tn[11] 0.0401341
R18647 XThC.Tn[11].n19 XThC.Tn[11] 0.0401341
R18648 XThC.Tn[11].n15 XThC.Tn[11] 0.0401341
R18649 XThC.Tn[11].n11 XThC.Tn[11] 0.0401341
R18650 XThC.Tn[11].n7 XThC.Tn[11] 0.0401341
R18651 XThC.Tn[11].n4 XThC.Tn[11] 0.0401341
R18652 XThC.Tn[12].n70 XThC.Tn[12].n69 256.103
R18653 XThC.Tn[12].n74 XThC.Tn[12].n72 243.68
R18654 XThC.Tn[12].n2 XThC.Tn[12].n0 241.847
R18655 XThC.Tn[12].n74 XThC.Tn[12].n73 205.28
R18656 XThC.Tn[12].n70 XThC.Tn[12].n68 202.095
R18657 XThC.Tn[12].n2 XThC.Tn[12].n1 185
R18658 XThC.Tn[12].n64 XThC.Tn[12].n62 161.365
R18659 XThC.Tn[12].n60 XThC.Tn[12].n58 161.365
R18660 XThC.Tn[12].n56 XThC.Tn[12].n54 161.365
R18661 XThC.Tn[12].n52 XThC.Tn[12].n50 161.365
R18662 XThC.Tn[12].n48 XThC.Tn[12].n46 161.365
R18663 XThC.Tn[12].n44 XThC.Tn[12].n42 161.365
R18664 XThC.Tn[12].n40 XThC.Tn[12].n38 161.365
R18665 XThC.Tn[12].n36 XThC.Tn[12].n34 161.365
R18666 XThC.Tn[12].n32 XThC.Tn[12].n30 161.365
R18667 XThC.Tn[12].n28 XThC.Tn[12].n26 161.365
R18668 XThC.Tn[12].n24 XThC.Tn[12].n22 161.365
R18669 XThC.Tn[12].n20 XThC.Tn[12].n18 161.365
R18670 XThC.Tn[12].n16 XThC.Tn[12].n14 161.365
R18671 XThC.Tn[12].n12 XThC.Tn[12].n10 161.365
R18672 XThC.Tn[12].n8 XThC.Tn[12].n6 161.365
R18673 XThC.Tn[12].n5 XThC.Tn[12].n3 161.365
R18674 XThC.Tn[12].n62 XThC.Tn[12].t41 161.202
R18675 XThC.Tn[12].n58 XThC.Tn[12].t31 161.202
R18676 XThC.Tn[12].n54 XThC.Tn[12].t18 161.202
R18677 XThC.Tn[12].n50 XThC.Tn[12].t15 161.202
R18678 XThC.Tn[12].n46 XThC.Tn[12].t39 161.202
R18679 XThC.Tn[12].n42 XThC.Tn[12].t26 161.202
R18680 XThC.Tn[12].n38 XThC.Tn[12].t25 161.202
R18681 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R18682 XThC.Tn[12].n30 XThC.Tn[12].t36 161.202
R18683 XThC.Tn[12].n26 XThC.Tn[12].t27 161.202
R18684 XThC.Tn[12].n22 XThC.Tn[12].t14 161.202
R18685 XThC.Tn[12].n18 XThC.Tn[12].t13 161.202
R18686 XThC.Tn[12].n14 XThC.Tn[12].t24 161.202
R18687 XThC.Tn[12].n10 XThC.Tn[12].t22 161.202
R18688 XThC.Tn[12].n6 XThC.Tn[12].t20 161.202
R18689 XThC.Tn[12].n3 XThC.Tn[12].t35 161.202
R18690 XThC.Tn[12].n62 XThC.Tn[12].t12 145.137
R18691 XThC.Tn[12].n58 XThC.Tn[12].t34 145.137
R18692 XThC.Tn[12].n54 XThC.Tn[12].t21 145.137
R18693 XThC.Tn[12].n50 XThC.Tn[12].t19 145.137
R18694 XThC.Tn[12].n46 XThC.Tn[12].t43 145.137
R18695 XThC.Tn[12].n42 XThC.Tn[12].t32 145.137
R18696 XThC.Tn[12].n38 XThC.Tn[12].t30 145.137
R18697 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R18698 XThC.Tn[12].n30 XThC.Tn[12].t40 145.137
R18699 XThC.Tn[12].n26 XThC.Tn[12].t33 145.137
R18700 XThC.Tn[12].n22 XThC.Tn[12].t17 145.137
R18701 XThC.Tn[12].n18 XThC.Tn[12].t16 145.137
R18702 XThC.Tn[12].n14 XThC.Tn[12].t29 145.137
R18703 XThC.Tn[12].n10 XThC.Tn[12].t28 145.137
R18704 XThC.Tn[12].n6 XThC.Tn[12].t23 145.137
R18705 XThC.Tn[12].n3 XThC.Tn[12].t37 145.137
R18706 XThC.Tn[12].n68 XThC.Tn[12].t1 26.5955
R18707 XThC.Tn[12].n68 XThC.Tn[12].t2 26.5955
R18708 XThC.Tn[12].n72 XThC.Tn[12].t9 26.5955
R18709 XThC.Tn[12].n72 XThC.Tn[12].t8 26.5955
R18710 XThC.Tn[12].n73 XThC.Tn[12].t11 26.5955
R18711 XThC.Tn[12].n73 XThC.Tn[12].t10 26.5955
R18712 XThC.Tn[12].n69 XThC.Tn[12].t0 26.5955
R18713 XThC.Tn[12].n69 XThC.Tn[12].t3 26.5955
R18714 XThC.Tn[12].n1 XThC.Tn[12].t5 24.9236
R18715 XThC.Tn[12].n1 XThC.Tn[12].t4 24.9236
R18716 XThC.Tn[12].n0 XThC.Tn[12].t7 24.9236
R18717 XThC.Tn[12].n0 XThC.Tn[12].t6 24.9236
R18718 XThC.Tn[12] XThC.Tn[12].n74 22.9652
R18719 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R18720 XThC.Tn[12].n71 XThC.Tn[12].n70 13.9299
R18721 XThC.Tn[12] XThC.Tn[12].n71 13.9299
R18722 XThC.Tn[12] XThC.Tn[12].n5 8.0245
R18723 XThC.Tn[12].n65 XThC.Tn[12].n64 7.9105
R18724 XThC.Tn[12].n61 XThC.Tn[12].n60 7.9105
R18725 XThC.Tn[12].n57 XThC.Tn[12].n56 7.9105
R18726 XThC.Tn[12].n53 XThC.Tn[12].n52 7.9105
R18727 XThC.Tn[12].n49 XThC.Tn[12].n48 7.9105
R18728 XThC.Tn[12].n45 XThC.Tn[12].n44 7.9105
R18729 XThC.Tn[12].n41 XThC.Tn[12].n40 7.9105
R18730 XThC.Tn[12].n37 XThC.Tn[12].n36 7.9105
R18731 XThC.Tn[12].n33 XThC.Tn[12].n32 7.9105
R18732 XThC.Tn[12].n29 XThC.Tn[12].n28 7.9105
R18733 XThC.Tn[12].n25 XThC.Tn[12].n24 7.9105
R18734 XThC.Tn[12].n21 XThC.Tn[12].n20 7.9105
R18735 XThC.Tn[12].n17 XThC.Tn[12].n16 7.9105
R18736 XThC.Tn[12].n13 XThC.Tn[12].n12 7.9105
R18737 XThC.Tn[12].n9 XThC.Tn[12].n8 7.9105
R18738 XThC.Tn[12].n67 XThC.Tn[12].n66 7.4309
R18739 XThC.Tn[12].n66 XThC.Tn[12] 4.71945
R18740 XThC.Tn[12].n71 XThC.Tn[12].n67 2.99115
R18741 XThC.Tn[12].n71 XThC.Tn[12] 2.87153
R18742 XThC.Tn[12].n67 XThC.Tn[12] 2.2734
R18743 XThC.Tn[12].n66 XThC.Tn[12] 0.88175
R18744 XThC.Tn[12].n9 XThC.Tn[12] 0.235138
R18745 XThC.Tn[12].n13 XThC.Tn[12] 0.235138
R18746 XThC.Tn[12].n17 XThC.Tn[12] 0.235138
R18747 XThC.Tn[12].n21 XThC.Tn[12] 0.235138
R18748 XThC.Tn[12].n25 XThC.Tn[12] 0.235138
R18749 XThC.Tn[12].n29 XThC.Tn[12] 0.235138
R18750 XThC.Tn[12].n33 XThC.Tn[12] 0.235138
R18751 XThC.Tn[12].n37 XThC.Tn[12] 0.235138
R18752 XThC.Tn[12].n41 XThC.Tn[12] 0.235138
R18753 XThC.Tn[12].n45 XThC.Tn[12] 0.235138
R18754 XThC.Tn[12].n49 XThC.Tn[12] 0.235138
R18755 XThC.Tn[12].n53 XThC.Tn[12] 0.235138
R18756 XThC.Tn[12].n57 XThC.Tn[12] 0.235138
R18757 XThC.Tn[12].n61 XThC.Tn[12] 0.235138
R18758 XThC.Tn[12].n65 XThC.Tn[12] 0.235138
R18759 XThC.Tn[12] XThC.Tn[12].n9 0.114505
R18760 XThC.Tn[12] XThC.Tn[12].n13 0.114505
R18761 XThC.Tn[12] XThC.Tn[12].n17 0.114505
R18762 XThC.Tn[12] XThC.Tn[12].n21 0.114505
R18763 XThC.Tn[12] XThC.Tn[12].n25 0.114505
R18764 XThC.Tn[12] XThC.Tn[12].n29 0.114505
R18765 XThC.Tn[12] XThC.Tn[12].n33 0.114505
R18766 XThC.Tn[12] XThC.Tn[12].n37 0.114505
R18767 XThC.Tn[12] XThC.Tn[12].n41 0.114505
R18768 XThC.Tn[12] XThC.Tn[12].n45 0.114505
R18769 XThC.Tn[12] XThC.Tn[12].n49 0.114505
R18770 XThC.Tn[12] XThC.Tn[12].n53 0.114505
R18771 XThC.Tn[12] XThC.Tn[12].n57 0.114505
R18772 XThC.Tn[12] XThC.Tn[12].n61 0.114505
R18773 XThC.Tn[12] XThC.Tn[12].n65 0.114505
R18774 XThC.Tn[12].n64 XThC.Tn[12].n63 0.0599512
R18775 XThC.Tn[12].n60 XThC.Tn[12].n59 0.0599512
R18776 XThC.Tn[12].n56 XThC.Tn[12].n55 0.0599512
R18777 XThC.Tn[12].n52 XThC.Tn[12].n51 0.0599512
R18778 XThC.Tn[12].n48 XThC.Tn[12].n47 0.0599512
R18779 XThC.Tn[12].n44 XThC.Tn[12].n43 0.0599512
R18780 XThC.Tn[12].n40 XThC.Tn[12].n39 0.0599512
R18781 XThC.Tn[12].n36 XThC.Tn[12].n35 0.0599512
R18782 XThC.Tn[12].n32 XThC.Tn[12].n31 0.0599512
R18783 XThC.Tn[12].n28 XThC.Tn[12].n27 0.0599512
R18784 XThC.Tn[12].n24 XThC.Tn[12].n23 0.0599512
R18785 XThC.Tn[12].n20 XThC.Tn[12].n19 0.0599512
R18786 XThC.Tn[12].n16 XThC.Tn[12].n15 0.0599512
R18787 XThC.Tn[12].n12 XThC.Tn[12].n11 0.0599512
R18788 XThC.Tn[12].n8 XThC.Tn[12].n7 0.0599512
R18789 XThC.Tn[12].n5 XThC.Tn[12].n4 0.0599512
R18790 XThC.Tn[12].n63 XThC.Tn[12] 0.0469286
R18791 XThC.Tn[12].n59 XThC.Tn[12] 0.0469286
R18792 XThC.Tn[12].n55 XThC.Tn[12] 0.0469286
R18793 XThC.Tn[12].n51 XThC.Tn[12] 0.0469286
R18794 XThC.Tn[12].n47 XThC.Tn[12] 0.0469286
R18795 XThC.Tn[12].n43 XThC.Tn[12] 0.0469286
R18796 XThC.Tn[12].n39 XThC.Tn[12] 0.0469286
R18797 XThC.Tn[12].n35 XThC.Tn[12] 0.0469286
R18798 XThC.Tn[12].n31 XThC.Tn[12] 0.0469286
R18799 XThC.Tn[12].n27 XThC.Tn[12] 0.0469286
R18800 XThC.Tn[12].n23 XThC.Tn[12] 0.0469286
R18801 XThC.Tn[12].n19 XThC.Tn[12] 0.0469286
R18802 XThC.Tn[12].n15 XThC.Tn[12] 0.0469286
R18803 XThC.Tn[12].n11 XThC.Tn[12] 0.0469286
R18804 XThC.Tn[12].n7 XThC.Tn[12] 0.0469286
R18805 XThC.Tn[12].n4 XThC.Tn[12] 0.0469286
R18806 XThC.Tn[12].n63 XThC.Tn[12] 0.0401341
R18807 XThC.Tn[12].n59 XThC.Tn[12] 0.0401341
R18808 XThC.Tn[12].n55 XThC.Tn[12] 0.0401341
R18809 XThC.Tn[12].n51 XThC.Tn[12] 0.0401341
R18810 XThC.Tn[12].n47 XThC.Tn[12] 0.0401341
R18811 XThC.Tn[12].n43 XThC.Tn[12] 0.0401341
R18812 XThC.Tn[12].n39 XThC.Tn[12] 0.0401341
R18813 XThC.Tn[12].n35 XThC.Tn[12] 0.0401341
R18814 XThC.Tn[12].n31 XThC.Tn[12] 0.0401341
R18815 XThC.Tn[12].n27 XThC.Tn[12] 0.0401341
R18816 XThC.Tn[12].n23 XThC.Tn[12] 0.0401341
R18817 XThC.Tn[12].n19 XThC.Tn[12] 0.0401341
R18818 XThC.Tn[12].n15 XThC.Tn[12] 0.0401341
R18819 XThC.Tn[12].n11 XThC.Tn[12] 0.0401341
R18820 XThC.Tn[12].n7 XThC.Tn[12] 0.0401341
R18821 XThC.Tn[12].n4 XThC.Tn[12] 0.0401341
R18822 XThC.Tn[13].n70 XThC.Tn[13].n69 265.341
R18823 XThC.Tn[13].n74 XThC.Tn[13].n72 243.68
R18824 XThC.Tn[13].n2 XThC.Tn[13].n0 241.847
R18825 XThC.Tn[13].n74 XThC.Tn[13].n73 205.28
R18826 XThC.Tn[13].n70 XThC.Tn[13].n68 202.094
R18827 XThC.Tn[13].n2 XThC.Tn[13].n1 185
R18828 XThC.Tn[13].n64 XThC.Tn[13].n62 161.365
R18829 XThC.Tn[13].n60 XThC.Tn[13].n58 161.365
R18830 XThC.Tn[13].n56 XThC.Tn[13].n54 161.365
R18831 XThC.Tn[13].n52 XThC.Tn[13].n50 161.365
R18832 XThC.Tn[13].n48 XThC.Tn[13].n46 161.365
R18833 XThC.Tn[13].n44 XThC.Tn[13].n42 161.365
R18834 XThC.Tn[13].n40 XThC.Tn[13].n38 161.365
R18835 XThC.Tn[13].n36 XThC.Tn[13].n34 161.365
R18836 XThC.Tn[13].n32 XThC.Tn[13].n30 161.365
R18837 XThC.Tn[13].n28 XThC.Tn[13].n26 161.365
R18838 XThC.Tn[13].n24 XThC.Tn[13].n22 161.365
R18839 XThC.Tn[13].n20 XThC.Tn[13].n18 161.365
R18840 XThC.Tn[13].n16 XThC.Tn[13].n14 161.365
R18841 XThC.Tn[13].n12 XThC.Tn[13].n10 161.365
R18842 XThC.Tn[13].n8 XThC.Tn[13].n6 161.365
R18843 XThC.Tn[13].n5 XThC.Tn[13].n3 161.365
R18844 XThC.Tn[13].n62 XThC.Tn[13].t33 161.202
R18845 XThC.Tn[13].n58 XThC.Tn[13].t23 161.202
R18846 XThC.Tn[13].n54 XThC.Tn[13].t42 161.202
R18847 XThC.Tn[13].n50 XThC.Tn[13].t39 161.202
R18848 XThC.Tn[13].n46 XThC.Tn[13].t31 161.202
R18849 XThC.Tn[13].n42 XThC.Tn[13].t18 161.202
R18850 XThC.Tn[13].n38 XThC.Tn[13].t17 161.202
R18851 XThC.Tn[13].n34 XThC.Tn[13].t30 161.202
R18852 XThC.Tn[13].n30 XThC.Tn[13].t28 161.202
R18853 XThC.Tn[13].n26 XThC.Tn[13].t19 161.202
R18854 XThC.Tn[13].n22 XThC.Tn[13].t38 161.202
R18855 XThC.Tn[13].n18 XThC.Tn[13].t37 161.202
R18856 XThC.Tn[13].n14 XThC.Tn[13].t16 161.202
R18857 XThC.Tn[13].n10 XThC.Tn[13].t14 161.202
R18858 XThC.Tn[13].n6 XThC.Tn[13].t12 161.202
R18859 XThC.Tn[13].n3 XThC.Tn[13].t27 161.202
R18860 XThC.Tn[13].n62 XThC.Tn[13].t36 145.137
R18861 XThC.Tn[13].n58 XThC.Tn[13].t26 145.137
R18862 XThC.Tn[13].n54 XThC.Tn[13].t13 145.137
R18863 XThC.Tn[13].n50 XThC.Tn[13].t43 145.137
R18864 XThC.Tn[13].n46 XThC.Tn[13].t35 145.137
R18865 XThC.Tn[13].n42 XThC.Tn[13].t24 145.137
R18866 XThC.Tn[13].n38 XThC.Tn[13].t22 145.137
R18867 XThC.Tn[13].n34 XThC.Tn[13].t34 145.137
R18868 XThC.Tn[13].n30 XThC.Tn[13].t32 145.137
R18869 XThC.Tn[13].n26 XThC.Tn[13].t25 145.137
R18870 XThC.Tn[13].n22 XThC.Tn[13].t41 145.137
R18871 XThC.Tn[13].n18 XThC.Tn[13].t40 145.137
R18872 XThC.Tn[13].n14 XThC.Tn[13].t21 145.137
R18873 XThC.Tn[13].n10 XThC.Tn[13].t20 145.137
R18874 XThC.Tn[13].n6 XThC.Tn[13].t15 145.137
R18875 XThC.Tn[13].n3 XThC.Tn[13].t29 145.137
R18876 XThC.Tn[13].n68 XThC.Tn[13].t2 26.5955
R18877 XThC.Tn[13].n68 XThC.Tn[13].t1 26.5955
R18878 XThC.Tn[13].n72 XThC.Tn[13].t9 26.5955
R18879 XThC.Tn[13].n72 XThC.Tn[13].t8 26.5955
R18880 XThC.Tn[13].n73 XThC.Tn[13].t11 26.5955
R18881 XThC.Tn[13].n73 XThC.Tn[13].t10 26.5955
R18882 XThC.Tn[13].n69 XThC.Tn[13].t0 26.5955
R18883 XThC.Tn[13].n69 XThC.Tn[13].t3 26.5955
R18884 XThC.Tn[13].n1 XThC.Tn[13].t4 24.9236
R18885 XThC.Tn[13].n1 XThC.Tn[13].t6 24.9236
R18886 XThC.Tn[13].n0 XThC.Tn[13].t7 24.9236
R18887 XThC.Tn[13].n0 XThC.Tn[13].t5 24.9236
R18888 XThC.Tn[13] XThC.Tn[13].n74 22.9652
R18889 XThC.Tn[13] XThC.Tn[13].n2 18.8943
R18890 XThC.Tn[13].n71 XThC.Tn[13].n70 13.9299
R18891 XThC.Tn[13] XThC.Tn[13].n71 13.9299
R18892 XThC.Tn[13] XThC.Tn[13].n5 8.0245
R18893 XThC.Tn[13].n65 XThC.Tn[13].n64 7.9105
R18894 XThC.Tn[13].n61 XThC.Tn[13].n60 7.9105
R18895 XThC.Tn[13].n57 XThC.Tn[13].n56 7.9105
R18896 XThC.Tn[13].n53 XThC.Tn[13].n52 7.9105
R18897 XThC.Tn[13].n49 XThC.Tn[13].n48 7.9105
R18898 XThC.Tn[13].n45 XThC.Tn[13].n44 7.9105
R18899 XThC.Tn[13].n41 XThC.Tn[13].n40 7.9105
R18900 XThC.Tn[13].n37 XThC.Tn[13].n36 7.9105
R18901 XThC.Tn[13].n33 XThC.Tn[13].n32 7.9105
R18902 XThC.Tn[13].n29 XThC.Tn[13].n28 7.9105
R18903 XThC.Tn[13].n25 XThC.Tn[13].n24 7.9105
R18904 XThC.Tn[13].n21 XThC.Tn[13].n20 7.9105
R18905 XThC.Tn[13].n17 XThC.Tn[13].n16 7.9105
R18906 XThC.Tn[13].n13 XThC.Tn[13].n12 7.9105
R18907 XThC.Tn[13].n9 XThC.Tn[13].n8 7.9105
R18908 XThC.Tn[13].n67 XThC.Tn[13].n66 7.46054
R18909 XThC.Tn[13].n67 XThC.Tn[13] 6.34069
R18910 XThC.Tn[13].n66 XThC.Tn[13] 4.78838
R18911 XThC.Tn[13] XThC.Tn[13].n67 1.79489
R18912 XThC.Tn[13].n66 XThC.Tn[13] 1.51436
R18913 XThC.Tn[13].n71 XThC.Tn[13] 1.19676
R18914 XThC.Tn[13].n9 XThC.Tn[13] 0.235138
R18915 XThC.Tn[13].n13 XThC.Tn[13] 0.235138
R18916 XThC.Tn[13].n17 XThC.Tn[13] 0.235138
R18917 XThC.Tn[13].n21 XThC.Tn[13] 0.235138
R18918 XThC.Tn[13].n25 XThC.Tn[13] 0.235138
R18919 XThC.Tn[13].n29 XThC.Tn[13] 0.235138
R18920 XThC.Tn[13].n33 XThC.Tn[13] 0.235138
R18921 XThC.Tn[13].n37 XThC.Tn[13] 0.235138
R18922 XThC.Tn[13].n41 XThC.Tn[13] 0.235138
R18923 XThC.Tn[13].n45 XThC.Tn[13] 0.235138
R18924 XThC.Tn[13].n49 XThC.Tn[13] 0.235138
R18925 XThC.Tn[13].n53 XThC.Tn[13] 0.235138
R18926 XThC.Tn[13].n57 XThC.Tn[13] 0.235138
R18927 XThC.Tn[13].n61 XThC.Tn[13] 0.235138
R18928 XThC.Tn[13].n65 XThC.Tn[13] 0.235138
R18929 XThC.Tn[13] XThC.Tn[13].n9 0.114505
R18930 XThC.Tn[13] XThC.Tn[13].n13 0.114505
R18931 XThC.Tn[13] XThC.Tn[13].n17 0.114505
R18932 XThC.Tn[13] XThC.Tn[13].n21 0.114505
R18933 XThC.Tn[13] XThC.Tn[13].n25 0.114505
R18934 XThC.Tn[13] XThC.Tn[13].n29 0.114505
R18935 XThC.Tn[13] XThC.Tn[13].n33 0.114505
R18936 XThC.Tn[13] XThC.Tn[13].n37 0.114505
R18937 XThC.Tn[13] XThC.Tn[13].n41 0.114505
R18938 XThC.Tn[13] XThC.Tn[13].n45 0.114505
R18939 XThC.Tn[13] XThC.Tn[13].n49 0.114505
R18940 XThC.Tn[13] XThC.Tn[13].n53 0.114505
R18941 XThC.Tn[13] XThC.Tn[13].n57 0.114505
R18942 XThC.Tn[13] XThC.Tn[13].n61 0.114505
R18943 XThC.Tn[13] XThC.Tn[13].n65 0.114505
R18944 XThC.Tn[13].n64 XThC.Tn[13].n63 0.0599512
R18945 XThC.Tn[13].n60 XThC.Tn[13].n59 0.0599512
R18946 XThC.Tn[13].n56 XThC.Tn[13].n55 0.0599512
R18947 XThC.Tn[13].n52 XThC.Tn[13].n51 0.0599512
R18948 XThC.Tn[13].n48 XThC.Tn[13].n47 0.0599512
R18949 XThC.Tn[13].n44 XThC.Tn[13].n43 0.0599512
R18950 XThC.Tn[13].n40 XThC.Tn[13].n39 0.0599512
R18951 XThC.Tn[13].n36 XThC.Tn[13].n35 0.0599512
R18952 XThC.Tn[13].n32 XThC.Tn[13].n31 0.0599512
R18953 XThC.Tn[13].n28 XThC.Tn[13].n27 0.0599512
R18954 XThC.Tn[13].n24 XThC.Tn[13].n23 0.0599512
R18955 XThC.Tn[13].n20 XThC.Tn[13].n19 0.0599512
R18956 XThC.Tn[13].n16 XThC.Tn[13].n15 0.0599512
R18957 XThC.Tn[13].n12 XThC.Tn[13].n11 0.0599512
R18958 XThC.Tn[13].n8 XThC.Tn[13].n7 0.0599512
R18959 XThC.Tn[13].n5 XThC.Tn[13].n4 0.0599512
R18960 XThC.Tn[13].n63 XThC.Tn[13] 0.0469286
R18961 XThC.Tn[13].n59 XThC.Tn[13] 0.0469286
R18962 XThC.Tn[13].n55 XThC.Tn[13] 0.0469286
R18963 XThC.Tn[13].n51 XThC.Tn[13] 0.0469286
R18964 XThC.Tn[13].n47 XThC.Tn[13] 0.0469286
R18965 XThC.Tn[13].n43 XThC.Tn[13] 0.0469286
R18966 XThC.Tn[13].n39 XThC.Tn[13] 0.0469286
R18967 XThC.Tn[13].n35 XThC.Tn[13] 0.0469286
R18968 XThC.Tn[13].n31 XThC.Tn[13] 0.0469286
R18969 XThC.Tn[13].n27 XThC.Tn[13] 0.0469286
R18970 XThC.Tn[13].n23 XThC.Tn[13] 0.0469286
R18971 XThC.Tn[13].n19 XThC.Tn[13] 0.0469286
R18972 XThC.Tn[13].n15 XThC.Tn[13] 0.0469286
R18973 XThC.Tn[13].n11 XThC.Tn[13] 0.0469286
R18974 XThC.Tn[13].n7 XThC.Tn[13] 0.0469286
R18975 XThC.Tn[13].n4 XThC.Tn[13] 0.0469286
R18976 XThC.Tn[13].n63 XThC.Tn[13] 0.0401341
R18977 XThC.Tn[13].n59 XThC.Tn[13] 0.0401341
R18978 XThC.Tn[13].n55 XThC.Tn[13] 0.0401341
R18979 XThC.Tn[13].n51 XThC.Tn[13] 0.0401341
R18980 XThC.Tn[13].n47 XThC.Tn[13] 0.0401341
R18981 XThC.Tn[13].n43 XThC.Tn[13] 0.0401341
R18982 XThC.Tn[13].n39 XThC.Tn[13] 0.0401341
R18983 XThC.Tn[13].n35 XThC.Tn[13] 0.0401341
R18984 XThC.Tn[13].n31 XThC.Tn[13] 0.0401341
R18985 XThC.Tn[13].n27 XThC.Tn[13] 0.0401341
R18986 XThC.Tn[13].n23 XThC.Tn[13] 0.0401341
R18987 XThC.Tn[13].n19 XThC.Tn[13] 0.0401341
R18988 XThC.Tn[13].n15 XThC.Tn[13] 0.0401341
R18989 XThC.Tn[13].n11 XThC.Tn[13] 0.0401341
R18990 XThC.Tn[13].n7 XThC.Tn[13] 0.0401341
R18991 XThC.Tn[13].n4 XThC.Tn[13] 0.0401341
R18992 XThC.Tn[0].n74 XThC.Tn[0].n73 332.332
R18993 XThC.Tn[0].n74 XThC.Tn[0].n72 296.493
R18994 XThC.Tn[0].n68 XThC.Tn[0].n66 161.365
R18995 XThC.Tn[0].n64 XThC.Tn[0].n62 161.365
R18996 XThC.Tn[0].n60 XThC.Tn[0].n58 161.365
R18997 XThC.Tn[0].n56 XThC.Tn[0].n54 161.365
R18998 XThC.Tn[0].n52 XThC.Tn[0].n50 161.365
R18999 XThC.Tn[0].n48 XThC.Tn[0].n46 161.365
R19000 XThC.Tn[0].n44 XThC.Tn[0].n42 161.365
R19001 XThC.Tn[0].n40 XThC.Tn[0].n38 161.365
R19002 XThC.Tn[0].n36 XThC.Tn[0].n34 161.365
R19003 XThC.Tn[0].n32 XThC.Tn[0].n30 161.365
R19004 XThC.Tn[0].n28 XThC.Tn[0].n26 161.365
R19005 XThC.Tn[0].n24 XThC.Tn[0].n22 161.365
R19006 XThC.Tn[0].n20 XThC.Tn[0].n18 161.365
R19007 XThC.Tn[0].n16 XThC.Tn[0].n14 161.365
R19008 XThC.Tn[0].n12 XThC.Tn[0].n10 161.365
R19009 XThC.Tn[0].n9 XThC.Tn[0].n7 161.365
R19010 XThC.Tn[0].n66 XThC.Tn[0].t29 161.202
R19011 XThC.Tn[0].n62 XThC.Tn[0].t19 161.202
R19012 XThC.Tn[0].n58 XThC.Tn[0].t38 161.202
R19013 XThC.Tn[0].n54 XThC.Tn[0].t36 161.202
R19014 XThC.Tn[0].n50 XThC.Tn[0].t27 161.202
R19015 XThC.Tn[0].n46 XThC.Tn[0].t16 161.202
R19016 XThC.Tn[0].n42 XThC.Tn[0].t15 161.202
R19017 XThC.Tn[0].n38 XThC.Tn[0].t26 161.202
R19018 XThC.Tn[0].n34 XThC.Tn[0].t25 161.202
R19019 XThC.Tn[0].n30 XThC.Tn[0].t17 161.202
R19020 XThC.Tn[0].n26 XThC.Tn[0].t34 161.202
R19021 XThC.Tn[0].n22 XThC.Tn[0].t32 161.202
R19022 XThC.Tn[0].n18 XThC.Tn[0].t13 161.202
R19023 XThC.Tn[0].n14 XThC.Tn[0].t12 161.202
R19024 XThC.Tn[0].n10 XThC.Tn[0].t41 161.202
R19025 XThC.Tn[0].n7 XThC.Tn[0].t22 161.202
R19026 XThC.Tn[0].n66 XThC.Tn[0].t24 145.137
R19027 XThC.Tn[0].n62 XThC.Tn[0].t14 145.137
R19028 XThC.Tn[0].n58 XThC.Tn[0].t33 145.137
R19029 XThC.Tn[0].n54 XThC.Tn[0].t31 145.137
R19030 XThC.Tn[0].n50 XThC.Tn[0].t23 145.137
R19031 XThC.Tn[0].n46 XThC.Tn[0].t42 145.137
R19032 XThC.Tn[0].n42 XThC.Tn[0].t40 145.137
R19033 XThC.Tn[0].n38 XThC.Tn[0].t21 145.137
R19034 XThC.Tn[0].n34 XThC.Tn[0].t20 145.137
R19035 XThC.Tn[0].n30 XThC.Tn[0].t43 145.137
R19036 XThC.Tn[0].n26 XThC.Tn[0].t30 145.137
R19037 XThC.Tn[0].n22 XThC.Tn[0].t28 145.137
R19038 XThC.Tn[0].n18 XThC.Tn[0].t39 145.137
R19039 XThC.Tn[0].n14 XThC.Tn[0].t37 145.137
R19040 XThC.Tn[0].n10 XThC.Tn[0].t35 145.137
R19041 XThC.Tn[0].n7 XThC.Tn[0].t18 145.137
R19042 XThC.Tn[0].n2 XThC.Tn[0].n0 135.248
R19043 XThC.Tn[0].n2 XThC.Tn[0].n1 98.982
R19044 XThC.Tn[0].n4 XThC.Tn[0].n3 98.982
R19045 XThC.Tn[0].n6 XThC.Tn[0].n5 98.982
R19046 XThC.Tn[0].n4 XThC.Tn[0].n2 36.2672
R19047 XThC.Tn[0].n6 XThC.Tn[0].n4 36.2672
R19048 XThC.Tn[0].n71 XThC.Tn[0].n6 32.6405
R19049 XThC.Tn[0].n72 XThC.Tn[0].t1 26.5955
R19050 XThC.Tn[0].n72 XThC.Tn[0].t0 26.5955
R19051 XThC.Tn[0].n73 XThC.Tn[0].t3 26.5955
R19052 XThC.Tn[0].n73 XThC.Tn[0].t2 26.5955
R19053 XThC.Tn[0].n0 XThC.Tn[0].t11 24.9236
R19054 XThC.Tn[0].n0 XThC.Tn[0].t8 24.9236
R19055 XThC.Tn[0].n1 XThC.Tn[0].t9 24.9236
R19056 XThC.Tn[0].n1 XThC.Tn[0].t10 24.9236
R19057 XThC.Tn[0].n3 XThC.Tn[0].t7 24.9236
R19058 XThC.Tn[0].n3 XThC.Tn[0].t6 24.9236
R19059 XThC.Tn[0].n5 XThC.Tn[0].t5 24.9236
R19060 XThC.Tn[0].n5 XThC.Tn[0].t4 24.9236
R19061 XThC.Tn[0].n75 XThC.Tn[0].n74 18.5605
R19062 XThC.Tn[0].n75 XThC.Tn[0].n71 11.5205
R19063 XThC.Tn[0] XThC.Tn[0].n9 8.0245
R19064 XThC.Tn[0].n69 XThC.Tn[0].n68 7.9105
R19065 XThC.Tn[0].n65 XThC.Tn[0].n64 7.9105
R19066 XThC.Tn[0].n61 XThC.Tn[0].n60 7.9105
R19067 XThC.Tn[0].n57 XThC.Tn[0].n56 7.9105
R19068 XThC.Tn[0].n53 XThC.Tn[0].n52 7.9105
R19069 XThC.Tn[0].n49 XThC.Tn[0].n48 7.9105
R19070 XThC.Tn[0].n45 XThC.Tn[0].n44 7.9105
R19071 XThC.Tn[0].n41 XThC.Tn[0].n40 7.9105
R19072 XThC.Tn[0].n37 XThC.Tn[0].n36 7.9105
R19073 XThC.Tn[0].n33 XThC.Tn[0].n32 7.9105
R19074 XThC.Tn[0].n29 XThC.Tn[0].n28 7.9105
R19075 XThC.Tn[0].n25 XThC.Tn[0].n24 7.9105
R19076 XThC.Tn[0].n21 XThC.Tn[0].n20 7.9105
R19077 XThC.Tn[0].n17 XThC.Tn[0].n16 7.9105
R19078 XThC.Tn[0].n13 XThC.Tn[0].n12 7.9105
R19079 XThC.Tn[0].n70 XThC.Tn[0] 5.95611
R19080 XThC.Tn[0].n71 XThC.Tn[0].n70 4.6005
R19081 XThC.Tn[0].n70 XThC.Tn[0] 1.89022
R19082 XThC.Tn[0] XThC.Tn[0].n75 0.6405
R19083 XThC.Tn[0].n13 XThC.Tn[0] 0.235138
R19084 XThC.Tn[0].n17 XThC.Tn[0] 0.235138
R19085 XThC.Tn[0].n21 XThC.Tn[0] 0.235138
R19086 XThC.Tn[0].n25 XThC.Tn[0] 0.235138
R19087 XThC.Tn[0].n29 XThC.Tn[0] 0.235138
R19088 XThC.Tn[0].n33 XThC.Tn[0] 0.235138
R19089 XThC.Tn[0].n37 XThC.Tn[0] 0.235138
R19090 XThC.Tn[0].n41 XThC.Tn[0] 0.235138
R19091 XThC.Tn[0].n45 XThC.Tn[0] 0.235138
R19092 XThC.Tn[0].n49 XThC.Tn[0] 0.235138
R19093 XThC.Tn[0].n53 XThC.Tn[0] 0.235138
R19094 XThC.Tn[0].n57 XThC.Tn[0] 0.235138
R19095 XThC.Tn[0].n61 XThC.Tn[0] 0.235138
R19096 XThC.Tn[0].n65 XThC.Tn[0] 0.235138
R19097 XThC.Tn[0].n69 XThC.Tn[0] 0.235138
R19098 XThC.Tn[0] XThC.Tn[0].n13 0.114505
R19099 XThC.Tn[0] XThC.Tn[0].n17 0.114505
R19100 XThC.Tn[0] XThC.Tn[0].n21 0.114505
R19101 XThC.Tn[0] XThC.Tn[0].n25 0.114505
R19102 XThC.Tn[0] XThC.Tn[0].n29 0.114505
R19103 XThC.Tn[0] XThC.Tn[0].n33 0.114505
R19104 XThC.Tn[0] XThC.Tn[0].n37 0.114505
R19105 XThC.Tn[0] XThC.Tn[0].n41 0.114505
R19106 XThC.Tn[0] XThC.Tn[0].n45 0.114505
R19107 XThC.Tn[0] XThC.Tn[0].n49 0.114505
R19108 XThC.Tn[0] XThC.Tn[0].n53 0.114505
R19109 XThC.Tn[0] XThC.Tn[0].n57 0.114505
R19110 XThC.Tn[0] XThC.Tn[0].n61 0.114505
R19111 XThC.Tn[0] XThC.Tn[0].n65 0.114505
R19112 XThC.Tn[0] XThC.Tn[0].n69 0.114505
R19113 XThC.Tn[0].n68 XThC.Tn[0].n67 0.0599512
R19114 XThC.Tn[0].n64 XThC.Tn[0].n63 0.0599512
R19115 XThC.Tn[0].n60 XThC.Tn[0].n59 0.0599512
R19116 XThC.Tn[0].n56 XThC.Tn[0].n55 0.0599512
R19117 XThC.Tn[0].n52 XThC.Tn[0].n51 0.0599512
R19118 XThC.Tn[0].n48 XThC.Tn[0].n47 0.0599512
R19119 XThC.Tn[0].n44 XThC.Tn[0].n43 0.0599512
R19120 XThC.Tn[0].n40 XThC.Tn[0].n39 0.0599512
R19121 XThC.Tn[0].n36 XThC.Tn[0].n35 0.0599512
R19122 XThC.Tn[0].n32 XThC.Tn[0].n31 0.0599512
R19123 XThC.Tn[0].n28 XThC.Tn[0].n27 0.0599512
R19124 XThC.Tn[0].n24 XThC.Tn[0].n23 0.0599512
R19125 XThC.Tn[0].n20 XThC.Tn[0].n19 0.0599512
R19126 XThC.Tn[0].n16 XThC.Tn[0].n15 0.0599512
R19127 XThC.Tn[0].n12 XThC.Tn[0].n11 0.0599512
R19128 XThC.Tn[0].n9 XThC.Tn[0].n8 0.0599512
R19129 XThC.Tn[0].n67 XThC.Tn[0] 0.0469286
R19130 XThC.Tn[0].n63 XThC.Tn[0] 0.0469286
R19131 XThC.Tn[0].n59 XThC.Tn[0] 0.0469286
R19132 XThC.Tn[0].n55 XThC.Tn[0] 0.0469286
R19133 XThC.Tn[0].n51 XThC.Tn[0] 0.0469286
R19134 XThC.Tn[0].n47 XThC.Tn[0] 0.0469286
R19135 XThC.Tn[0].n43 XThC.Tn[0] 0.0469286
R19136 XThC.Tn[0].n39 XThC.Tn[0] 0.0469286
R19137 XThC.Tn[0].n35 XThC.Tn[0] 0.0469286
R19138 XThC.Tn[0].n31 XThC.Tn[0] 0.0469286
R19139 XThC.Tn[0].n27 XThC.Tn[0] 0.0469286
R19140 XThC.Tn[0].n23 XThC.Tn[0] 0.0469286
R19141 XThC.Tn[0].n19 XThC.Tn[0] 0.0469286
R19142 XThC.Tn[0].n15 XThC.Tn[0] 0.0469286
R19143 XThC.Tn[0].n11 XThC.Tn[0] 0.0469286
R19144 XThC.Tn[0].n8 XThC.Tn[0] 0.0469286
R19145 XThC.Tn[0].n67 XThC.Tn[0] 0.0401341
R19146 XThC.Tn[0].n63 XThC.Tn[0] 0.0401341
R19147 XThC.Tn[0].n59 XThC.Tn[0] 0.0401341
R19148 XThC.Tn[0].n55 XThC.Tn[0] 0.0401341
R19149 XThC.Tn[0].n51 XThC.Tn[0] 0.0401341
R19150 XThC.Tn[0].n47 XThC.Tn[0] 0.0401341
R19151 XThC.Tn[0].n43 XThC.Tn[0] 0.0401341
R19152 XThC.Tn[0].n39 XThC.Tn[0] 0.0401341
R19153 XThC.Tn[0].n35 XThC.Tn[0] 0.0401341
R19154 XThC.Tn[0].n31 XThC.Tn[0] 0.0401341
R19155 XThC.Tn[0].n27 XThC.Tn[0] 0.0401341
R19156 XThC.Tn[0].n23 XThC.Tn[0] 0.0401341
R19157 XThC.Tn[0].n19 XThC.Tn[0] 0.0401341
R19158 XThC.Tn[0].n15 XThC.Tn[0] 0.0401341
R19159 XThC.Tn[0].n11 XThC.Tn[0] 0.0401341
R19160 XThC.Tn[0].n8 XThC.Tn[0] 0.0401341
R19161 XThC.XTB4.Y.n21 XThC.XTB4.Y.t0 235.56
R19162 XThC.XTB4.Y.n3 XThC.XTB4.Y.t3 212.081
R19163 XThC.XTB4.Y.n2 XThC.XTB4.Y.t2 212.081
R19164 XThC.XTB4.Y.n8 XThC.XTB4.Y.t17 212.081
R19165 XThC.XTB4.Y.n0 XThC.XTB4.Y.t13 212.081
R19166 XThC.XTB4.Y.n12 XThC.XTB4.Y.t8 212.081
R19167 XThC.XTB4.Y.n13 XThC.XTB4.Y.t12 212.081
R19168 XThC.XTB4.Y.n15 XThC.XTB4.Y.t6 212.081
R19169 XThC.XTB4.Y.n11 XThC.XTB4.Y.t16 212.081
R19170 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 173.761
R19171 XThC.XTB4.Y.n14 XThC.XTB4.Y 158.656
R19172 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 152
R19173 XThC.XTB4.Y.n5 XThC.XTB4.Y.n1 152
R19174 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 152
R19175 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 152
R19176 XThC.XTB4.Y.n3 XThC.XTB4.Y.t14 139.78
R19177 XThC.XTB4.Y.n2 XThC.XTB4.Y.t10 139.78
R19178 XThC.XTB4.Y.n8 XThC.XTB4.Y.t7 139.78
R19179 XThC.XTB4.Y.n0 XThC.XTB4.Y.t4 139.78
R19180 XThC.XTB4.Y.n12 XThC.XTB4.Y.t11 139.78
R19181 XThC.XTB4.Y.n13 XThC.XTB4.Y.t15 139.78
R19182 XThC.XTB4.Y.n15 XThC.XTB4.Y.t9 139.78
R19183 XThC.XTB4.Y.n11 XThC.XTB4.Y.t5 139.78
R19184 XThC.XTB4.Y.n20 XThC.XTB4.Y.t1 133.386
R19185 XThC.XTB4.Y.n19 XThC.XTB4.Y.n10 72.9296
R19186 XThC.XTB4.Y.n13 XThC.XTB4.Y.n12 61.346
R19187 XThC.XTB4.Y.n7 XThC.XTB4.Y.n1 49.6611
R19188 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 45.2793
R19189 XThC.XTB4.Y.n4 XThC.XTB4.Y.n2 42.3581
R19190 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 38.1854
R19191 XThC.XTB4.Y.n16 XThC.XTB4.Y.n11 30.6732
R19192 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R19193 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R19194 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 30.6732
R19195 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 21.7605
R19196 XThC.XTB4.Y XThC.XTB4.Y.n20 19.5051
R19197 XThC.XTB4.Y.n4 XThC.XTB4.Y.n3 18.9884
R19198 XThC.XTB4.Y.n9 XThC.XTB4.Y.n0 16.0672
R19199 XThC.XTB4.Y.n17 XThC.XTB4.Y 14.7905
R19200 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 11.994
R19201 XThC.XTB4.Y.n10 XThC.XTB4.Y 11.5205
R19202 XThC.XTB4.Y.n6 XThC.XTB4.Y 10.2405
R19203 XThC.XTB4.Y.n2 XThC.XTB4.Y.n1 7.30353
R19204 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 7.24578
R19205 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 4.38232
R19206 XThC.XTB4.Y.n21 XThC.XTB4.Y 2.22659
R19207 XThC.XTB4.Y XThC.XTB4.Y.n21 1.55202
R19208 XThC.XTB4.Y.n18 XThC.XTB4.Y 0.966538
R19209 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19210 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19211 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19212 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19213 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19214 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19215 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19216 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19217 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19218 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19219 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19220 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19221 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19222 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19223 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19224 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19225 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19226 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19227 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19228 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19229 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19230 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19231 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19232 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19233 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19234 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19235 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19236 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19237 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19238 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19239 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19240 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19241 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19242 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19243 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19244 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19245 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19246 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19247 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19248 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19249 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19250 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19251 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19252 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19253 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19254 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19255 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19256 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19257 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19258 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19259 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19260 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19261 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19262 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19263 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19264 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19265 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19266 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19267 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19268 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19269 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19270 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19271 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19272 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19273 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19274 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19275 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19276 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19277 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19278 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19279 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19280 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19281 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19282 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19283 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19284 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19285 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19286 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19287 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19288 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19289 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19290 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19291 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19292 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19293 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19294 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19295 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19296 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19297 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19298 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19299 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19300 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19301 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19302 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19303 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19304 XThR.Tn[3].n7 XThR.Tn[3].n6 135.249
R19305 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19306 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19307 XThR.Tn[3].n7 XThR.Tn[3].n5 98.981
R19308 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19309 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19310 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19311 XThR.Tn[3].n1 XThR.Tn[3].t7 26.5955
R19312 XThR.Tn[3].n1 XThR.Tn[3].t10 26.5955
R19313 XThR.Tn[3].n0 XThR.Tn[3].t8 26.5955
R19314 XThR.Tn[3].n0 XThR.Tn[3].t9 26.5955
R19315 XThR.Tn[3].n3 XThR.Tn[3].t6 24.9236
R19316 XThR.Tn[3].n3 XThR.Tn[3].t3 24.9236
R19317 XThR.Tn[3].n4 XThR.Tn[3].t5 24.9236
R19318 XThR.Tn[3].n4 XThR.Tn[3].t4 24.9236
R19319 XThR.Tn[3].n5 XThR.Tn[3].t11 24.9236
R19320 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19321 XThR.Tn[3].n6 XThR.Tn[3].t0 24.9236
R19322 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19323 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19324 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19325 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19326 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19327 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19328 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19329 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19330 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19331 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19332 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19333 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19334 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19335 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19336 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19337 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19338 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19339 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19340 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19341 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19342 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19343 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19344 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19345 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19346 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19347 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19348 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19349 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19350 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19351 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19352 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19353 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19354 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19355 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19356 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19357 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19358 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19359 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19360 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19361 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19362 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19363 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19364 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19365 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19366 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19367 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19368 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19369 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19370 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19371 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19372 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19373 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19374 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19375 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19376 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19377 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19378 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19379 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19380 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19381 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19382 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19383 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19384 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19385 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19386 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19387 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19388 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19389 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19390 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19391 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19392 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19393 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19394 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19395 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19396 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19397 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19398 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19399 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19400 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19401 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19402 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19403 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19404 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19405 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19406 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19407 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19408 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19409 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19410 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19411 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19412 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19413 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19414 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19415 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19416 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19417 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19418 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19419 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19420 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19421 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19422 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19423 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19424 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19425 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19426 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19427 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19428 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19429 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19430 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19431 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19432 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19433 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19434 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19435 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19436 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19437 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19438 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19439 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19440 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19441 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19442 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19443 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19444 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19445 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19446 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19447 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19448 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19449 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19450 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19451 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19452 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19453 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19454 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19455 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19456 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19457 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19458 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19459 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19460 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19461 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19462 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19463 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19464 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19465 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19466 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19467 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19468 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19469 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19470 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19471 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19472 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19473 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19474 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19475 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19476 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19477 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19478 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19479 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19480 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19481 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19482 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19483 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19484 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19485 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19486 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19487 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19488 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19489 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19490 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19491 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19492 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19493 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19494 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19495 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19496 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19497 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19498 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19499 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19500 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19501 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19502 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19503 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19504 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19505 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19506 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19507 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19508 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19509 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19510 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19511 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19512 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19513 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19514 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19515 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19516 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19517 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19518 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19519 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19520 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19521 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19522 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19523 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19524 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19525 XThR.Tn[5].n1 XThR.Tn[5].t5 26.5955
R19526 XThR.Tn[5].n1 XThR.Tn[5].t4 26.5955
R19527 XThR.Tn[5].n0 XThR.Tn[5].t6 26.5955
R19528 XThR.Tn[5].n0 XThR.Tn[5].t7 26.5955
R19529 XThR.Tn[5].n3 XThR.Tn[5].t11 24.9236
R19530 XThR.Tn[5].n3 XThR.Tn[5].t8 24.9236
R19531 XThR.Tn[5].n4 XThR.Tn[5].t10 24.9236
R19532 XThR.Tn[5].n4 XThR.Tn[5].t9 24.9236
R19533 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19534 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19535 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19536 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19537 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19538 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19539 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19540 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19541 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19542 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19543 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19544 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19545 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19546 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19547 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19548 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19549 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19550 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19551 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19552 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19553 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19554 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19555 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19556 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19557 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19558 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19559 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19560 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19561 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19562 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19563 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19564 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19565 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19566 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19567 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19568 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19569 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19570 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19571 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19572 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19573 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19574 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19575 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19576 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19577 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19578 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19579 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19580 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19581 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19582 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19583 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19584 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19585 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19586 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19587 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19588 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19589 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19590 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19591 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19592 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R19593 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R19594 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R19595 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R19596 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R19597 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R19598 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R19599 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R19600 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R19601 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R19602 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19603 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R19604 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R19605 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R19606 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R19607 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R19608 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R19609 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R19610 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R19611 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R19612 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R19613 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R19614 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R19615 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R19616 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R19617 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R19618 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R19619 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R19620 XThR.Tn[5] XThR.Tn[5].n87 0.038
R19621 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R19622 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R19623 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R19624 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R19625 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R19626 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R19627 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R19628 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R19629 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R19630 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R19631 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R19632 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R19633 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R19634 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R19635 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R19636 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R19637 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R19638 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R19639 XThC.Tn[4].n71 XThC.Tn[4].n69 161.365
R19640 XThC.Tn[4].n67 XThC.Tn[4].n65 161.365
R19641 XThC.Tn[4].n63 XThC.Tn[4].n61 161.365
R19642 XThC.Tn[4].n59 XThC.Tn[4].n57 161.365
R19643 XThC.Tn[4].n55 XThC.Tn[4].n53 161.365
R19644 XThC.Tn[4].n51 XThC.Tn[4].n49 161.365
R19645 XThC.Tn[4].n47 XThC.Tn[4].n45 161.365
R19646 XThC.Tn[4].n43 XThC.Tn[4].n41 161.365
R19647 XThC.Tn[4].n39 XThC.Tn[4].n37 161.365
R19648 XThC.Tn[4].n35 XThC.Tn[4].n33 161.365
R19649 XThC.Tn[4].n31 XThC.Tn[4].n29 161.365
R19650 XThC.Tn[4].n27 XThC.Tn[4].n25 161.365
R19651 XThC.Tn[4].n23 XThC.Tn[4].n21 161.365
R19652 XThC.Tn[4].n19 XThC.Tn[4].n17 161.365
R19653 XThC.Tn[4].n15 XThC.Tn[4].n13 161.365
R19654 XThC.Tn[4].n12 XThC.Tn[4].n10 161.365
R19655 XThC.Tn[4].n69 XThC.Tn[4].t32 161.202
R19656 XThC.Tn[4].n65 XThC.Tn[4].t22 161.202
R19657 XThC.Tn[4].n61 XThC.Tn[4].t41 161.202
R19658 XThC.Tn[4].n57 XThC.Tn[4].t38 161.202
R19659 XThC.Tn[4].n53 XThC.Tn[4].t30 161.202
R19660 XThC.Tn[4].n49 XThC.Tn[4].t17 161.202
R19661 XThC.Tn[4].n45 XThC.Tn[4].t16 161.202
R19662 XThC.Tn[4].n41 XThC.Tn[4].t29 161.202
R19663 XThC.Tn[4].n37 XThC.Tn[4].t27 161.202
R19664 XThC.Tn[4].n33 XThC.Tn[4].t18 161.202
R19665 XThC.Tn[4].n29 XThC.Tn[4].t37 161.202
R19666 XThC.Tn[4].n25 XThC.Tn[4].t36 161.202
R19667 XThC.Tn[4].n21 XThC.Tn[4].t15 161.202
R19668 XThC.Tn[4].n17 XThC.Tn[4].t13 161.202
R19669 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R19670 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R19671 XThC.Tn[4].n69 XThC.Tn[4].t35 145.137
R19672 XThC.Tn[4].n65 XThC.Tn[4].t25 145.137
R19673 XThC.Tn[4].n61 XThC.Tn[4].t12 145.137
R19674 XThC.Tn[4].n57 XThC.Tn[4].t42 145.137
R19675 XThC.Tn[4].n53 XThC.Tn[4].t34 145.137
R19676 XThC.Tn[4].n49 XThC.Tn[4].t23 145.137
R19677 XThC.Tn[4].n45 XThC.Tn[4].t21 145.137
R19678 XThC.Tn[4].n41 XThC.Tn[4].t33 145.137
R19679 XThC.Tn[4].n37 XThC.Tn[4].t31 145.137
R19680 XThC.Tn[4].n33 XThC.Tn[4].t24 145.137
R19681 XThC.Tn[4].n29 XThC.Tn[4].t40 145.137
R19682 XThC.Tn[4].n25 XThC.Tn[4].t39 145.137
R19683 XThC.Tn[4].n21 XThC.Tn[4].t20 145.137
R19684 XThC.Tn[4].n17 XThC.Tn[4].t19 145.137
R19685 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R19686 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R19687 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R19688 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R19689 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R19690 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R19691 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R19692 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R19693 XThC.Tn[4].n73 XThC.Tn[4].n9 32.6405
R19694 XThC.Tn[4].n1 XThC.Tn[4].t7 26.5955
R19695 XThC.Tn[4].n1 XThC.Tn[4].t6 26.5955
R19696 XThC.Tn[4].n0 XThC.Tn[4].t5 26.5955
R19697 XThC.Tn[4].n0 XThC.Tn[4].t4 26.5955
R19698 XThC.Tn[4].n3 XThC.Tn[4].t9 24.9236
R19699 XThC.Tn[4].n3 XThC.Tn[4].t8 24.9236
R19700 XThC.Tn[4].n4 XThC.Tn[4].t11 24.9236
R19701 XThC.Tn[4].n4 XThC.Tn[4].t10 24.9236
R19702 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R19703 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R19704 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R19705 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R19706 XThC.Tn[4].n74 XThC.Tn[4].n2 18.5605
R19707 XThC.Tn[4].n74 XThC.Tn[4].n73 11.5205
R19708 XThC.Tn[4] XThC.Tn[4].n12 8.0245
R19709 XThC.Tn[4].n72 XThC.Tn[4].n71 7.9105
R19710 XThC.Tn[4].n68 XThC.Tn[4].n67 7.9105
R19711 XThC.Tn[4].n64 XThC.Tn[4].n63 7.9105
R19712 XThC.Tn[4].n60 XThC.Tn[4].n59 7.9105
R19713 XThC.Tn[4].n56 XThC.Tn[4].n55 7.9105
R19714 XThC.Tn[4].n52 XThC.Tn[4].n51 7.9105
R19715 XThC.Tn[4].n48 XThC.Tn[4].n47 7.9105
R19716 XThC.Tn[4].n44 XThC.Tn[4].n43 7.9105
R19717 XThC.Tn[4].n40 XThC.Tn[4].n39 7.9105
R19718 XThC.Tn[4].n36 XThC.Tn[4].n35 7.9105
R19719 XThC.Tn[4].n32 XThC.Tn[4].n31 7.9105
R19720 XThC.Tn[4].n28 XThC.Tn[4].n27 7.9105
R19721 XThC.Tn[4].n24 XThC.Tn[4].n23 7.9105
R19722 XThC.Tn[4].n20 XThC.Tn[4].n19 7.9105
R19723 XThC.Tn[4].n16 XThC.Tn[4].n15 7.9105
R19724 XThC.Tn[4].n73 XThC.Tn[4] 5.77342
R19725 XThC.Tn[4] XThC.Tn[4].n74 0.6405
R19726 XThC.Tn[4].n16 XThC.Tn[4] 0.235138
R19727 XThC.Tn[4].n20 XThC.Tn[4] 0.235138
R19728 XThC.Tn[4].n24 XThC.Tn[4] 0.235138
R19729 XThC.Tn[4].n28 XThC.Tn[4] 0.235138
R19730 XThC.Tn[4].n32 XThC.Tn[4] 0.235138
R19731 XThC.Tn[4].n36 XThC.Tn[4] 0.235138
R19732 XThC.Tn[4].n40 XThC.Tn[4] 0.235138
R19733 XThC.Tn[4].n44 XThC.Tn[4] 0.235138
R19734 XThC.Tn[4].n48 XThC.Tn[4] 0.235138
R19735 XThC.Tn[4].n52 XThC.Tn[4] 0.235138
R19736 XThC.Tn[4].n56 XThC.Tn[4] 0.235138
R19737 XThC.Tn[4].n60 XThC.Tn[4] 0.235138
R19738 XThC.Tn[4].n64 XThC.Tn[4] 0.235138
R19739 XThC.Tn[4].n68 XThC.Tn[4] 0.235138
R19740 XThC.Tn[4].n72 XThC.Tn[4] 0.235138
R19741 XThC.Tn[4] XThC.Tn[4].n16 0.114505
R19742 XThC.Tn[4] XThC.Tn[4].n20 0.114505
R19743 XThC.Tn[4] XThC.Tn[4].n24 0.114505
R19744 XThC.Tn[4] XThC.Tn[4].n28 0.114505
R19745 XThC.Tn[4] XThC.Tn[4].n32 0.114505
R19746 XThC.Tn[4] XThC.Tn[4].n36 0.114505
R19747 XThC.Tn[4] XThC.Tn[4].n40 0.114505
R19748 XThC.Tn[4] XThC.Tn[4].n44 0.114505
R19749 XThC.Tn[4] XThC.Tn[4].n48 0.114505
R19750 XThC.Tn[4] XThC.Tn[4].n52 0.114505
R19751 XThC.Tn[4] XThC.Tn[4].n56 0.114505
R19752 XThC.Tn[4] XThC.Tn[4].n60 0.114505
R19753 XThC.Tn[4] XThC.Tn[4].n64 0.114505
R19754 XThC.Tn[4] XThC.Tn[4].n68 0.114505
R19755 XThC.Tn[4] XThC.Tn[4].n72 0.114505
R19756 XThC.Tn[4].n71 XThC.Tn[4].n70 0.0599512
R19757 XThC.Tn[4].n67 XThC.Tn[4].n66 0.0599512
R19758 XThC.Tn[4].n63 XThC.Tn[4].n62 0.0599512
R19759 XThC.Tn[4].n59 XThC.Tn[4].n58 0.0599512
R19760 XThC.Tn[4].n55 XThC.Tn[4].n54 0.0599512
R19761 XThC.Tn[4].n51 XThC.Tn[4].n50 0.0599512
R19762 XThC.Tn[4].n47 XThC.Tn[4].n46 0.0599512
R19763 XThC.Tn[4].n43 XThC.Tn[4].n42 0.0599512
R19764 XThC.Tn[4].n39 XThC.Tn[4].n38 0.0599512
R19765 XThC.Tn[4].n35 XThC.Tn[4].n34 0.0599512
R19766 XThC.Tn[4].n31 XThC.Tn[4].n30 0.0599512
R19767 XThC.Tn[4].n27 XThC.Tn[4].n26 0.0599512
R19768 XThC.Tn[4].n23 XThC.Tn[4].n22 0.0599512
R19769 XThC.Tn[4].n19 XThC.Tn[4].n18 0.0599512
R19770 XThC.Tn[4].n15 XThC.Tn[4].n14 0.0599512
R19771 XThC.Tn[4].n12 XThC.Tn[4].n11 0.0599512
R19772 XThC.Tn[4].n70 XThC.Tn[4] 0.0469286
R19773 XThC.Tn[4].n66 XThC.Tn[4] 0.0469286
R19774 XThC.Tn[4].n62 XThC.Tn[4] 0.0469286
R19775 XThC.Tn[4].n58 XThC.Tn[4] 0.0469286
R19776 XThC.Tn[4].n54 XThC.Tn[4] 0.0469286
R19777 XThC.Tn[4].n50 XThC.Tn[4] 0.0469286
R19778 XThC.Tn[4].n46 XThC.Tn[4] 0.0469286
R19779 XThC.Tn[4].n42 XThC.Tn[4] 0.0469286
R19780 XThC.Tn[4].n38 XThC.Tn[4] 0.0469286
R19781 XThC.Tn[4].n34 XThC.Tn[4] 0.0469286
R19782 XThC.Tn[4].n30 XThC.Tn[4] 0.0469286
R19783 XThC.Tn[4].n26 XThC.Tn[4] 0.0469286
R19784 XThC.Tn[4].n22 XThC.Tn[4] 0.0469286
R19785 XThC.Tn[4].n18 XThC.Tn[4] 0.0469286
R19786 XThC.Tn[4].n14 XThC.Tn[4] 0.0469286
R19787 XThC.Tn[4].n11 XThC.Tn[4] 0.0469286
R19788 XThC.Tn[4].n70 XThC.Tn[4] 0.0401341
R19789 XThC.Tn[4].n66 XThC.Tn[4] 0.0401341
R19790 XThC.Tn[4].n62 XThC.Tn[4] 0.0401341
R19791 XThC.Tn[4].n58 XThC.Tn[4] 0.0401341
R19792 XThC.Tn[4].n54 XThC.Tn[4] 0.0401341
R19793 XThC.Tn[4].n50 XThC.Tn[4] 0.0401341
R19794 XThC.Tn[4].n46 XThC.Tn[4] 0.0401341
R19795 XThC.Tn[4].n42 XThC.Tn[4] 0.0401341
R19796 XThC.Tn[4].n38 XThC.Tn[4] 0.0401341
R19797 XThC.Tn[4].n34 XThC.Tn[4] 0.0401341
R19798 XThC.Tn[4].n30 XThC.Tn[4] 0.0401341
R19799 XThC.Tn[4].n26 XThC.Tn[4] 0.0401341
R19800 XThC.Tn[4].n22 XThC.Tn[4] 0.0401341
R19801 XThC.Tn[4].n18 XThC.Tn[4] 0.0401341
R19802 XThC.Tn[4].n14 XThC.Tn[4] 0.0401341
R19803 XThC.Tn[4].n11 XThC.Tn[4] 0.0401341
R19804 XThC.Tn[2].n74 XThC.Tn[2].n72 332.332
R19805 XThC.Tn[2].n74 XThC.Tn[2].n73 296.493
R19806 XThC.Tn[2].n68 XThC.Tn[2].n66 161.365
R19807 XThC.Tn[2].n64 XThC.Tn[2].n62 161.365
R19808 XThC.Tn[2].n60 XThC.Tn[2].n58 161.365
R19809 XThC.Tn[2].n56 XThC.Tn[2].n54 161.365
R19810 XThC.Tn[2].n52 XThC.Tn[2].n50 161.365
R19811 XThC.Tn[2].n48 XThC.Tn[2].n46 161.365
R19812 XThC.Tn[2].n44 XThC.Tn[2].n42 161.365
R19813 XThC.Tn[2].n40 XThC.Tn[2].n38 161.365
R19814 XThC.Tn[2].n36 XThC.Tn[2].n34 161.365
R19815 XThC.Tn[2].n32 XThC.Tn[2].n30 161.365
R19816 XThC.Tn[2].n28 XThC.Tn[2].n26 161.365
R19817 XThC.Tn[2].n24 XThC.Tn[2].n22 161.365
R19818 XThC.Tn[2].n20 XThC.Tn[2].n18 161.365
R19819 XThC.Tn[2].n16 XThC.Tn[2].n14 161.365
R19820 XThC.Tn[2].n12 XThC.Tn[2].n10 161.365
R19821 XThC.Tn[2].n9 XThC.Tn[2].n7 161.365
R19822 XThC.Tn[2].n66 XThC.Tn[2].t24 161.202
R19823 XThC.Tn[2].n62 XThC.Tn[2].t14 161.202
R19824 XThC.Tn[2].n58 XThC.Tn[2].t33 161.202
R19825 XThC.Tn[2].n54 XThC.Tn[2].t30 161.202
R19826 XThC.Tn[2].n50 XThC.Tn[2].t22 161.202
R19827 XThC.Tn[2].n46 XThC.Tn[2].t41 161.202
R19828 XThC.Tn[2].n42 XThC.Tn[2].t40 161.202
R19829 XThC.Tn[2].n38 XThC.Tn[2].t21 161.202
R19830 XThC.Tn[2].n34 XThC.Tn[2].t19 161.202
R19831 XThC.Tn[2].n30 XThC.Tn[2].t42 161.202
R19832 XThC.Tn[2].n26 XThC.Tn[2].t29 161.202
R19833 XThC.Tn[2].n22 XThC.Tn[2].t28 161.202
R19834 XThC.Tn[2].n18 XThC.Tn[2].t39 161.202
R19835 XThC.Tn[2].n14 XThC.Tn[2].t37 161.202
R19836 XThC.Tn[2].n10 XThC.Tn[2].t35 161.202
R19837 XThC.Tn[2].n7 XThC.Tn[2].t18 161.202
R19838 XThC.Tn[2].n66 XThC.Tn[2].t27 145.137
R19839 XThC.Tn[2].n62 XThC.Tn[2].t17 145.137
R19840 XThC.Tn[2].n58 XThC.Tn[2].t36 145.137
R19841 XThC.Tn[2].n54 XThC.Tn[2].t34 145.137
R19842 XThC.Tn[2].n50 XThC.Tn[2].t26 145.137
R19843 XThC.Tn[2].n46 XThC.Tn[2].t15 145.137
R19844 XThC.Tn[2].n42 XThC.Tn[2].t13 145.137
R19845 XThC.Tn[2].n38 XThC.Tn[2].t25 145.137
R19846 XThC.Tn[2].n34 XThC.Tn[2].t23 145.137
R19847 XThC.Tn[2].n30 XThC.Tn[2].t16 145.137
R19848 XThC.Tn[2].n26 XThC.Tn[2].t32 145.137
R19849 XThC.Tn[2].n22 XThC.Tn[2].t31 145.137
R19850 XThC.Tn[2].n18 XThC.Tn[2].t12 145.137
R19851 XThC.Tn[2].n14 XThC.Tn[2].t43 145.137
R19852 XThC.Tn[2].n10 XThC.Tn[2].t38 145.137
R19853 XThC.Tn[2].n7 XThC.Tn[2].t20 145.137
R19854 XThC.Tn[2].n2 XThC.Tn[2].n0 135.248
R19855 XThC.Tn[2].n2 XThC.Tn[2].n1 98.982
R19856 XThC.Tn[2].n4 XThC.Tn[2].n3 98.982
R19857 XThC.Tn[2].n6 XThC.Tn[2].n5 98.982
R19858 XThC.Tn[2].n4 XThC.Tn[2].n2 36.2672
R19859 XThC.Tn[2].n6 XThC.Tn[2].n4 36.2672
R19860 XThC.Tn[2].n71 XThC.Tn[2].n6 32.6405
R19861 XThC.Tn[2].n72 XThC.Tn[2].t1 26.5955
R19862 XThC.Tn[2].n72 XThC.Tn[2].t0 26.5955
R19863 XThC.Tn[2].n73 XThC.Tn[2].t3 26.5955
R19864 XThC.Tn[2].n73 XThC.Tn[2].t2 26.5955
R19865 XThC.Tn[2].n0 XThC.Tn[2].t8 24.9236
R19866 XThC.Tn[2].n0 XThC.Tn[2].t10 24.9236
R19867 XThC.Tn[2].n1 XThC.Tn[2].t11 24.9236
R19868 XThC.Tn[2].n1 XThC.Tn[2].t9 24.9236
R19869 XThC.Tn[2].n3 XThC.Tn[2].t5 24.9236
R19870 XThC.Tn[2].n3 XThC.Tn[2].t4 24.9236
R19871 XThC.Tn[2].n5 XThC.Tn[2].t7 24.9236
R19872 XThC.Tn[2].n5 XThC.Tn[2].t6 24.9236
R19873 XThC.Tn[2].n75 XThC.Tn[2].n74 18.5605
R19874 XThC.Tn[2].n75 XThC.Tn[2].n71 11.5205
R19875 XThC.Tn[2] XThC.Tn[2].n9 8.0245
R19876 XThC.Tn[2].n69 XThC.Tn[2].n68 7.9105
R19877 XThC.Tn[2].n65 XThC.Tn[2].n64 7.9105
R19878 XThC.Tn[2].n61 XThC.Tn[2].n60 7.9105
R19879 XThC.Tn[2].n57 XThC.Tn[2].n56 7.9105
R19880 XThC.Tn[2].n53 XThC.Tn[2].n52 7.9105
R19881 XThC.Tn[2].n49 XThC.Tn[2].n48 7.9105
R19882 XThC.Tn[2].n45 XThC.Tn[2].n44 7.9105
R19883 XThC.Tn[2].n41 XThC.Tn[2].n40 7.9105
R19884 XThC.Tn[2].n37 XThC.Tn[2].n36 7.9105
R19885 XThC.Tn[2].n33 XThC.Tn[2].n32 7.9105
R19886 XThC.Tn[2].n29 XThC.Tn[2].n28 7.9105
R19887 XThC.Tn[2].n25 XThC.Tn[2].n24 7.9105
R19888 XThC.Tn[2].n21 XThC.Tn[2].n20 7.9105
R19889 XThC.Tn[2].n17 XThC.Tn[2].n16 7.9105
R19890 XThC.Tn[2].n13 XThC.Tn[2].n12 7.9105
R19891 XThC.Tn[2].n70 XThC.Tn[2] 5.58686
R19892 XThC.Tn[2].n71 XThC.Tn[2].n70 4.6005
R19893 XThC.Tn[2].n70 XThC.Tn[2] 1.83383
R19894 XThC.Tn[2] XThC.Tn[2].n75 0.6405
R19895 XThC.Tn[2].n13 XThC.Tn[2] 0.235138
R19896 XThC.Tn[2].n17 XThC.Tn[2] 0.235138
R19897 XThC.Tn[2].n21 XThC.Tn[2] 0.235138
R19898 XThC.Tn[2].n25 XThC.Tn[2] 0.235138
R19899 XThC.Tn[2].n29 XThC.Tn[2] 0.235138
R19900 XThC.Tn[2].n33 XThC.Tn[2] 0.235138
R19901 XThC.Tn[2].n37 XThC.Tn[2] 0.235138
R19902 XThC.Tn[2].n41 XThC.Tn[2] 0.235138
R19903 XThC.Tn[2].n45 XThC.Tn[2] 0.235138
R19904 XThC.Tn[2].n49 XThC.Tn[2] 0.235138
R19905 XThC.Tn[2].n53 XThC.Tn[2] 0.235138
R19906 XThC.Tn[2].n57 XThC.Tn[2] 0.235138
R19907 XThC.Tn[2].n61 XThC.Tn[2] 0.235138
R19908 XThC.Tn[2].n65 XThC.Tn[2] 0.235138
R19909 XThC.Tn[2].n69 XThC.Tn[2] 0.235138
R19910 XThC.Tn[2] XThC.Tn[2].n13 0.114505
R19911 XThC.Tn[2] XThC.Tn[2].n17 0.114505
R19912 XThC.Tn[2] XThC.Tn[2].n21 0.114505
R19913 XThC.Tn[2] XThC.Tn[2].n25 0.114505
R19914 XThC.Tn[2] XThC.Tn[2].n29 0.114505
R19915 XThC.Tn[2] XThC.Tn[2].n33 0.114505
R19916 XThC.Tn[2] XThC.Tn[2].n37 0.114505
R19917 XThC.Tn[2] XThC.Tn[2].n41 0.114505
R19918 XThC.Tn[2] XThC.Tn[2].n45 0.114505
R19919 XThC.Tn[2] XThC.Tn[2].n49 0.114505
R19920 XThC.Tn[2] XThC.Tn[2].n53 0.114505
R19921 XThC.Tn[2] XThC.Tn[2].n57 0.114505
R19922 XThC.Tn[2] XThC.Tn[2].n61 0.114505
R19923 XThC.Tn[2] XThC.Tn[2].n65 0.114505
R19924 XThC.Tn[2] XThC.Tn[2].n69 0.114505
R19925 XThC.Tn[2].n68 XThC.Tn[2].n67 0.0599512
R19926 XThC.Tn[2].n64 XThC.Tn[2].n63 0.0599512
R19927 XThC.Tn[2].n60 XThC.Tn[2].n59 0.0599512
R19928 XThC.Tn[2].n56 XThC.Tn[2].n55 0.0599512
R19929 XThC.Tn[2].n52 XThC.Tn[2].n51 0.0599512
R19930 XThC.Tn[2].n48 XThC.Tn[2].n47 0.0599512
R19931 XThC.Tn[2].n44 XThC.Tn[2].n43 0.0599512
R19932 XThC.Tn[2].n40 XThC.Tn[2].n39 0.0599512
R19933 XThC.Tn[2].n36 XThC.Tn[2].n35 0.0599512
R19934 XThC.Tn[2].n32 XThC.Tn[2].n31 0.0599512
R19935 XThC.Tn[2].n28 XThC.Tn[2].n27 0.0599512
R19936 XThC.Tn[2].n24 XThC.Tn[2].n23 0.0599512
R19937 XThC.Tn[2].n20 XThC.Tn[2].n19 0.0599512
R19938 XThC.Tn[2].n16 XThC.Tn[2].n15 0.0599512
R19939 XThC.Tn[2].n12 XThC.Tn[2].n11 0.0599512
R19940 XThC.Tn[2].n9 XThC.Tn[2].n8 0.0599512
R19941 XThC.Tn[2].n67 XThC.Tn[2] 0.0469286
R19942 XThC.Tn[2].n63 XThC.Tn[2] 0.0469286
R19943 XThC.Tn[2].n59 XThC.Tn[2] 0.0469286
R19944 XThC.Tn[2].n55 XThC.Tn[2] 0.0469286
R19945 XThC.Tn[2].n51 XThC.Tn[2] 0.0469286
R19946 XThC.Tn[2].n47 XThC.Tn[2] 0.0469286
R19947 XThC.Tn[2].n43 XThC.Tn[2] 0.0469286
R19948 XThC.Tn[2].n39 XThC.Tn[2] 0.0469286
R19949 XThC.Tn[2].n35 XThC.Tn[2] 0.0469286
R19950 XThC.Tn[2].n31 XThC.Tn[2] 0.0469286
R19951 XThC.Tn[2].n27 XThC.Tn[2] 0.0469286
R19952 XThC.Tn[2].n23 XThC.Tn[2] 0.0469286
R19953 XThC.Tn[2].n19 XThC.Tn[2] 0.0469286
R19954 XThC.Tn[2].n15 XThC.Tn[2] 0.0469286
R19955 XThC.Tn[2].n11 XThC.Tn[2] 0.0469286
R19956 XThC.Tn[2].n8 XThC.Tn[2] 0.0469286
R19957 XThC.Tn[2].n67 XThC.Tn[2] 0.0401341
R19958 XThC.Tn[2].n63 XThC.Tn[2] 0.0401341
R19959 XThC.Tn[2].n59 XThC.Tn[2] 0.0401341
R19960 XThC.Tn[2].n55 XThC.Tn[2] 0.0401341
R19961 XThC.Tn[2].n51 XThC.Tn[2] 0.0401341
R19962 XThC.Tn[2].n47 XThC.Tn[2] 0.0401341
R19963 XThC.Tn[2].n43 XThC.Tn[2] 0.0401341
R19964 XThC.Tn[2].n39 XThC.Tn[2] 0.0401341
R19965 XThC.Tn[2].n35 XThC.Tn[2] 0.0401341
R19966 XThC.Tn[2].n31 XThC.Tn[2] 0.0401341
R19967 XThC.Tn[2].n27 XThC.Tn[2] 0.0401341
R19968 XThC.Tn[2].n23 XThC.Tn[2] 0.0401341
R19969 XThC.Tn[2].n19 XThC.Tn[2] 0.0401341
R19970 XThC.Tn[2].n15 XThC.Tn[2] 0.0401341
R19971 XThC.Tn[2].n11 XThC.Tn[2] 0.0401341
R19972 XThC.Tn[2].n8 XThC.Tn[2] 0.0401341
R19973 Vbias.n1 Vbias.t3 651.571
R19974 Vbias.n1 Vbias.t4 651.571
R19975 Vbias.n2 Vbias.t0 651.571
R19976 Vbias.n2 Vbias.t5 651.571
R19977 Vbias.n337 Vbias.t260 119.309
R19978 Vbias.n383 Vbias.t194 119.309
R19979 Vbias.n384 Vbias.t61 119.309
R19980 Vbias.n334 Vbias.t215 119.309
R19981 Vbias.n292 Vbias.t86 119.309
R19982 Vbias.n284 Vbias.t186 119.309
R19983 Vbias.n288 Vbias.t109 119.309
R19984 Vbias.n280 Vbias.t189 119.309
R19985 Vbias.n194 Vbias.t64 119.309
R19986 Vbias.n149 Vbias.t82 119.309
R19987 Vbias.n189 Vbias.t105 119.309
R19988 Vbias.n145 Vbias.t121 119.309
R19989 Vbias.n678 Vbias.t255 119.309
R19990 Vbias.n102 Vbias.t16 119.309
R19991 Vbias.n10 Vbias.t146 119.309
R19992 Vbias.n57 Vbias.t57 119.309
R19993 Vbias.n58 Vbias.t129 119.309
R19994 Vbias.n54 Vbias.t201 119.309
R19995 Vbias.n440 Vbias.t79 119.309
R19996 Vbias.n343 Vbias.t216 119.309
R19997 Vbias.n333 Vbias.t31 119.309
R19998 Vbias.n331 Vbias.t100 119.309
R19999 Vbias.n577 Vbias.t6 119.309
R20000 Vbias.n278 Vbias.t128 119.309
R20001 Vbias.n276 Vbias.t10 119.309
R20002 Vbias.n197 Vbias.t83 119.309
R20003 Vbias.n150 Vbias.t154 119.309
R20004 Vbias.n152 Vbias.t122 119.309
R20005 Vbias.n789 Vbias.t195 119.309
R20006 Vbias.n105 Vbias.t17 119.309
R20007 Vbias.n103 Vbias.t88 119.309
R20008 Vbias.n97 Vbias.t160 119.309
R20009 Vbias.n56 Vbias.t130 119.309
R20010 Vbias.n53 Vbias.t41 119.309
R20011 Vbias.n437 Vbias.t174 119.309
R20012 Vbias.n346 Vbias.t59 119.309
R20013 Vbias.n326 Vbias.t132 119.309
R20014 Vbias.n328 Vbias.t203 119.309
R20015 Vbias.n574 Vbias.t103 119.309
R20016 Vbias.n273 Vbias.t226 119.309
R20017 Vbias.n275 Vbias.t108 119.309
R20018 Vbias.n200 Vbias.t180 119.309
R20019 Vbias.n155 Vbias.t257 119.309
R20020 Vbias.n153 Vbias.t222 119.309
R20021 Vbias.n792 Vbias.t37 119.309
R20022 Vbias.n106 Vbias.t113 119.309
R20023 Vbias.n108 Vbias.t185 119.309
R20024 Vbias.n94 Vbias.t261 119.309
R20025 Vbias.n51 Vbias.t229 119.309
R20026 Vbias.n48 Vbias.t56 119.309
R20027 Vbias.n434 Vbias.t182 119.309
R20028 Vbias.n349 Vbias.t67 119.309
R20029 Vbias.n325 Vbias.t139 119.309
R20030 Vbias.n323 Vbias.t214 119.309
R20031 Vbias.n571 Vbias.t115 119.309
R20032 Vbias.n272 Vbias.t241 119.309
R20033 Vbias.n270 Vbias.t117 119.309
R20034 Vbias.n203 Vbias.t188 119.309
R20035 Vbias.n156 Vbias.t8 119.309
R20036 Vbias.n158 Vbias.t235 119.309
R20037 Vbias.n795 Vbias.t48 119.309
R20038 Vbias.n111 Vbias.t124 119.309
R20039 Vbias.n109 Vbias.t196 119.309
R20040 Vbias.n91 Vbias.t14 119.309
R20041 Vbias.n50 Vbias.t242 119.309
R20042 Vbias.n47 Vbias.t141 119.309
R20043 Vbias.n431 Vbias.t15 119.309
R20044 Vbias.n352 Vbias.t152 119.309
R20045 Vbias.n320 Vbias.t224 119.309
R20046 Vbias.n322 Vbias.t38 119.309
R20047 Vbias.n568 Vbias.t206 119.309
R20048 Vbias.n267 Vbias.t66 119.309
R20049 Vbias.n269 Vbias.t208 119.309
R20050 Vbias.n206 Vbias.t23 119.309
R20051 Vbias.n161 Vbias.t93 119.309
R20052 Vbias.n159 Vbias.t63 119.309
R20053 Vbias.n798 Vbias.t135 119.309
R20054 Vbias.n112 Vbias.t213 119.309
R20055 Vbias.n114 Vbias.t29 119.309
R20056 Vbias.n88 Vbias.t99 119.309
R20057 Vbias.n45 Vbias.t69 119.309
R20058 Vbias.n42 Vbias.t227 119.309
R20059 Vbias.n428 Vbias.t101 119.309
R20060 Vbias.n355 Vbias.t245 119.309
R20061 Vbias.n319 Vbias.t58 119.309
R20062 Vbias.n317 Vbias.t131 119.309
R20063 Vbias.n565 Vbias.t34 119.309
R20064 Vbias.n266 Vbias.t155 119.309
R20065 Vbias.n264 Vbias.t36 119.309
R20066 Vbias.n209 Vbias.t107 119.309
R20067 Vbias.n162 Vbias.t179 119.309
R20068 Vbias.n164 Vbias.t150 119.309
R20069 Vbias.n801 Vbias.t221 119.309
R20070 Vbias.n117 Vbias.t40 119.309
R20071 Vbias.n115 Vbias.t112 119.309
R20072 Vbias.n85 Vbias.t183 119.309
R20073 Vbias.n44 Vbias.t156 119.309
R20074 Vbias.n41 Vbias.t60 119.309
R20075 Vbias.n425 Vbias.t184 119.309
R20076 Vbias.n358 Vbias.t72 119.309
R20077 Vbias.n314 Vbias.t145 119.309
R20078 Vbias.n316 Vbias.t218 119.309
R20079 Vbias.n562 Vbias.t116 119.309
R20080 Vbias.n261 Vbias.t244 119.309
R20081 Vbias.n263 Vbias.t120 119.309
R20082 Vbias.n212 Vbias.t192 119.309
R20083 Vbias.n167 Vbias.t11 119.309
R20084 Vbias.n165 Vbias.t237 119.309
R20085 Vbias.n804 Vbias.t50 119.309
R20086 Vbias.n118 Vbias.t127 119.309
R20087 Vbias.n120 Vbias.t200 119.309
R20088 Vbias.n82 Vbias.t18 119.309
R20089 Vbias.n39 Vbias.t247 119.309
R20090 Vbias.n36 Vbias.t147 119.309
R20091 Vbias.n422 Vbias.t19 119.309
R20092 Vbias.n361 Vbias.t158 119.309
R20093 Vbias.n313 Vbias.t230 119.309
R20094 Vbias.n311 Vbias.t42 119.309
R20095 Vbias.n559 Vbias.t209 119.309
R20096 Vbias.n260 Vbias.t74 119.309
R20097 Vbias.n258 Vbias.t212 119.309
R20098 Vbias.n215 Vbias.t28 119.309
R20099 Vbias.n168 Vbias.t98 119.309
R20100 Vbias.n170 Vbias.t68 119.309
R20101 Vbias.n807 Vbias.t138 119.309
R20102 Vbias.n123 Vbias.t219 119.309
R20103 Vbias.n121 Vbias.t33 119.309
R20104 Vbias.n79 Vbias.t102 119.309
R20105 Vbias.n38 Vbias.t76 119.309
R20106 Vbias.n35 Vbias.t169 119.309
R20107 Vbias.n419 Vbias.t39 119.309
R20108 Vbias.n364 Vbias.t178 119.309
R20109 Vbias.n308 Vbias.t253 119.309
R20110 Vbias.n310 Vbias.t70 119.309
R20111 Vbias.n556 Vbias.t231 119.309
R20112 Vbias.n255 Vbias.t94 119.309
R20113 Vbias.n257 Vbias.t234 119.309
R20114 Vbias.n218 Vbias.t45 119.309
R20115 Vbias.n173 Vbias.t118 119.309
R20116 Vbias.n171 Vbias.t91 119.309
R20117 Vbias.n810 Vbias.t163 119.309
R20118 Vbias.n124 Vbias.t240 119.309
R20119 Vbias.n126 Vbias.t53 119.309
R20120 Vbias.n76 Vbias.t125 119.309
R20121 Vbias.n33 Vbias.t96 119.309
R20122 Vbias.n30 Vbias.t246 119.309
R20123 Vbias.n416 Vbias.t111 119.309
R20124 Vbias.n367 Vbias.t254 119.309
R20125 Vbias.n307 Vbias.t71 119.309
R20126 Vbias.n305 Vbias.t143 119.309
R20127 Vbias.n553 Vbias.t43 119.309
R20128 Vbias.n254 Vbias.t167 119.309
R20129 Vbias.n252 Vbias.t46 119.309
R20130 Vbias.n221 Vbias.t119 119.309
R20131 Vbias.n174 Vbias.t190 119.309
R20132 Vbias.n176 Vbias.t164 119.309
R20133 Vbias.n813 Vbias.t236 119.309
R20134 Vbias.n129 Vbias.t54 119.309
R20135 Vbias.n127 Vbias.t126 119.309
R20136 Vbias.n73 Vbias.t199 119.309
R20137 Vbias.n32 Vbias.t171 119.309
R20138 Vbias.n29 Vbias.t75 119.309
R20139 Vbias.n413 Vbias.t202 119.309
R20140 Vbias.n370 Vbias.t84 119.309
R20141 Vbias.n302 Vbias.t157 119.309
R20142 Vbias.n304 Vbias.t228 119.309
R20143 Vbias.n550 Vbias.t134 119.309
R20144 Vbias.n249 Vbias.t256 119.309
R20145 Vbias.n251 Vbias.t136 119.309
R20146 Vbias.n224 Vbias.t211 119.309
R20147 Vbias.n179 Vbias.t27 119.309
R20148 Vbias.n177 Vbias.t251 119.309
R20149 Vbias.n816 Vbias.t65 119.309
R20150 Vbias.n130 Vbias.t144 119.309
R20151 Vbias.n132 Vbias.t217 119.309
R20152 Vbias.n70 Vbias.t32 119.309
R20153 Vbias.n27 Vbias.t258 119.309
R20154 Vbias.n24 Vbias.t95 119.309
R20155 Vbias.n410 Vbias.t223 119.309
R20156 Vbias.n373 Vbias.t106 119.309
R20157 Vbias.n301 Vbias.t177 119.309
R20158 Vbias.n299 Vbias.t252 119.309
R20159 Vbias.n547 Vbias.t159 119.309
R20160 Vbias.n248 Vbias.t22 119.309
R20161 Vbias.n246 Vbias.t162 119.309
R20162 Vbias.n227 Vbias.t233 119.309
R20163 Vbias.n180 Vbias.t44 119.309
R20164 Vbias.n182 Vbias.t21 119.309
R20165 Vbias.n819 Vbias.t90 119.309
R20166 Vbias.n135 Vbias.t166 119.309
R20167 Vbias.n133 Vbias.t239 119.309
R20168 Vbias.n67 Vbias.t52 119.309
R20169 Vbias.n26 Vbias.t25 119.309
R20170 Vbias.n23 Vbias.t248 119.309
R20171 Vbias.n407 Vbias.t114 119.309
R20172 Vbias.n376 Vbias.t259 119.309
R20173 Vbias.n296 Vbias.t77 119.309
R20174 Vbias.n298 Vbias.t148 119.309
R20175 Vbias.n544 Vbias.t47 119.309
R20176 Vbias.n243 Vbias.t172 119.309
R20177 Vbias.n245 Vbias.t51 119.309
R20178 Vbias.n230 Vbias.t123 119.309
R20179 Vbias.n185 Vbias.t197 119.309
R20180 Vbias.n183 Vbias.t168 119.309
R20181 Vbias.n822 Vbias.t243 119.309
R20182 Vbias.n136 Vbias.t62 119.309
R20183 Vbias.n138 Vbias.t133 119.309
R20184 Vbias.n64 Vbias.t205 119.309
R20185 Vbias.n21 Vbias.t173 119.309
R20186 Vbias.n16 Vbias.t12 119.309
R20187 Vbias.n404 Vbias.t142 119.309
R20188 Vbias.n379 Vbias.t26 119.309
R20189 Vbias.n295 Vbias.t97 119.309
R20190 Vbias.n293 Vbias.t170 119.309
R20191 Vbias.n541 Vbias.t78 119.309
R20192 Vbias.n242 Vbias.t191 119.309
R20193 Vbias.n240 Vbias.t80 119.309
R20194 Vbias.n233 Vbias.t149 119.309
R20195 Vbias.n186 Vbias.t220 119.309
R20196 Vbias.n188 Vbias.t187 119.309
R20197 Vbias.n825 Vbias.t7 119.309
R20198 Vbias.n141 Vbias.t81 119.309
R20199 Vbias.n139 Vbias.t153 119.309
R20200 Vbias.n61 Vbias.t225 119.309
R20201 Vbias.n18 Vbias.t193 119.309
R20202 Vbias.n15 Vbias.t24 119.309
R20203 Vbias.n338 Vbias.t151 119.309
R20204 Vbias.n339 Vbias.t35 119.309
R20205 Vbias.n341 Vbias.t104 119.309
R20206 Vbias.n525 Vbias.t175 119.309
R20207 Vbias.n285 Vbias.t85 119.309
R20208 Vbias.n287 Vbias.t207 119.309
R20209 Vbias.n662 Vbias.t89 119.309
R20210 Vbias.n236 Vbias.t161 119.309
R20211 Vbias.n238 Vbias.t232 119.309
R20212 Vbias.n703 Vbias.t204 119.309
R20213 Vbias.n144 Vbias.t20 119.309
R20214 Vbias.n142 Vbias.t92 119.309
R20215 Vbias.n671 Vbias.t165 119.309
R20216 Vbias.n11 Vbias.t238 119.309
R20217 Vbias.n13 Vbias.t210 119.309
R20218 Vbias.n6 Vbias.t181 119.309
R20219 Vbias.n7 Vbias.t110 119.309
R20220 Vbias.n60 Vbias.t87 119.309
R20221 Vbias.n674 Vbias.t73 119.309
R20222 Vbias.n906 Vbias.t198 119.309
R20223 Vbias.n683 Vbias.t176 119.309
R20224 Vbias.n146 Vbias.t49 119.309
R20225 Vbias.n191 Vbias.t137 119.309
R20226 Vbias.n195 Vbias.t9 119.309
R20227 Vbias.n665 Vbias.t250 119.309
R20228 Vbias.n279 Vbias.t55 119.309
R20229 Vbias.n289 Vbias.t249 119.309
R20230 Vbias.n329 Vbias.t30 119.309
R20231 Vbias.n395 Vbias.t13 119.309
R20232 Vbias.n335 Vbias.t140 119.309
R20233 Vbias.n0 Vbias.t1 77.1834
R20234 Vbias.n0 Vbias.t2 34.3787
R20235 Vbias.n3 Vbias.n1 4.78773
R20236 Vbias.n3 Vbias.n2 4.78773
R20237 Vbias.n386 Vbias.n384 4.5005
R20238 Vbias.n441 Vbias.n440 4.5005
R20239 Vbias.n344 Vbias.n343 4.5005
R20240 Vbias.n448 Vbias.n333 4.5005
R20241 Vbias.n451 Vbias.n331 4.5005
R20242 Vbias.n578 Vbias.n577 4.5005
R20243 Vbias.n585 Vbias.n278 4.5005
R20244 Vbias.n588 Vbias.n276 4.5005
R20245 Vbias.n198 Vbias.n197 4.5005
R20246 Vbias.n782 Vbias.n150 4.5005
R20247 Vbias.n779 Vbias.n152 4.5005
R20248 Vbias.n790 Vbias.n789 4.5005
R20249 Vbias.n909 Vbias.n105 4.5005
R20250 Vbias.n912 Vbias.n103 4.5005
R20251 Vbias.n98 Vbias.n97 4.5005
R20252 Vbias.n920 Vbias.n56 4.5005
R20253 Vbias.n922 Vbias.n54 4.5005
R20254 Vbias.n438 Vbias.n437 4.5005
R20255 Vbias.n347 Vbias.n346 4.5005
R20256 Vbias.n457 Vbias.n326 4.5005
R20257 Vbias.n454 Vbias.n328 4.5005
R20258 Vbias.n575 Vbias.n574 4.5005
R20259 Vbias.n594 Vbias.n273 4.5005
R20260 Vbias.n591 Vbias.n275 4.5005
R20261 Vbias.n201 Vbias.n200 4.5005
R20262 Vbias.n773 Vbias.n155 4.5005
R20263 Vbias.n776 Vbias.n153 4.5005
R20264 Vbias.n793 Vbias.n792 4.5005
R20265 Vbias.n904 Vbias.n106 4.5005
R20266 Vbias.n901 Vbias.n108 4.5005
R20267 Vbias.n95 Vbias.n94 4.5005
R20268 Vbias.n927 Vbias.n51 4.5005
R20269 Vbias.n925 Vbias.n53 4.5005
R20270 Vbias.n435 Vbias.n434 4.5005
R20271 Vbias.n350 Vbias.n349 4.5005
R20272 Vbias.n460 Vbias.n325 4.5005
R20273 Vbias.n463 Vbias.n323 4.5005
R20274 Vbias.n572 Vbias.n571 4.5005
R20275 Vbias.n597 Vbias.n272 4.5005
R20276 Vbias.n600 Vbias.n270 4.5005
R20277 Vbias.n204 Vbias.n203 4.5005
R20278 Vbias.n770 Vbias.n156 4.5005
R20279 Vbias.n767 Vbias.n158 4.5005
R20280 Vbias.n796 Vbias.n795 4.5005
R20281 Vbias.n895 Vbias.n111 4.5005
R20282 Vbias.n898 Vbias.n109 4.5005
R20283 Vbias.n92 Vbias.n91 4.5005
R20284 Vbias.n930 Vbias.n50 4.5005
R20285 Vbias.n932 Vbias.n48 4.5005
R20286 Vbias.n432 Vbias.n431 4.5005
R20287 Vbias.n353 Vbias.n352 4.5005
R20288 Vbias.n469 Vbias.n320 4.5005
R20289 Vbias.n466 Vbias.n322 4.5005
R20290 Vbias.n569 Vbias.n568 4.5005
R20291 Vbias.n606 Vbias.n267 4.5005
R20292 Vbias.n603 Vbias.n269 4.5005
R20293 Vbias.n207 Vbias.n206 4.5005
R20294 Vbias.n761 Vbias.n161 4.5005
R20295 Vbias.n764 Vbias.n159 4.5005
R20296 Vbias.n799 Vbias.n798 4.5005
R20297 Vbias.n892 Vbias.n112 4.5005
R20298 Vbias.n889 Vbias.n114 4.5005
R20299 Vbias.n89 Vbias.n88 4.5005
R20300 Vbias.n937 Vbias.n45 4.5005
R20301 Vbias.n935 Vbias.n47 4.5005
R20302 Vbias.n429 Vbias.n428 4.5005
R20303 Vbias.n356 Vbias.n355 4.5005
R20304 Vbias.n472 Vbias.n319 4.5005
R20305 Vbias.n475 Vbias.n317 4.5005
R20306 Vbias.n566 Vbias.n565 4.5005
R20307 Vbias.n609 Vbias.n266 4.5005
R20308 Vbias.n612 Vbias.n264 4.5005
R20309 Vbias.n210 Vbias.n209 4.5005
R20310 Vbias.n758 Vbias.n162 4.5005
R20311 Vbias.n755 Vbias.n164 4.5005
R20312 Vbias.n802 Vbias.n801 4.5005
R20313 Vbias.n883 Vbias.n117 4.5005
R20314 Vbias.n886 Vbias.n115 4.5005
R20315 Vbias.n86 Vbias.n85 4.5005
R20316 Vbias.n940 Vbias.n44 4.5005
R20317 Vbias.n942 Vbias.n42 4.5005
R20318 Vbias.n426 Vbias.n425 4.5005
R20319 Vbias.n359 Vbias.n358 4.5005
R20320 Vbias.n481 Vbias.n314 4.5005
R20321 Vbias.n478 Vbias.n316 4.5005
R20322 Vbias.n563 Vbias.n562 4.5005
R20323 Vbias.n618 Vbias.n261 4.5005
R20324 Vbias.n615 Vbias.n263 4.5005
R20325 Vbias.n213 Vbias.n212 4.5005
R20326 Vbias.n749 Vbias.n167 4.5005
R20327 Vbias.n752 Vbias.n165 4.5005
R20328 Vbias.n805 Vbias.n804 4.5005
R20329 Vbias.n880 Vbias.n118 4.5005
R20330 Vbias.n877 Vbias.n120 4.5005
R20331 Vbias.n83 Vbias.n82 4.5005
R20332 Vbias.n947 Vbias.n39 4.5005
R20333 Vbias.n945 Vbias.n41 4.5005
R20334 Vbias.n423 Vbias.n422 4.5005
R20335 Vbias.n362 Vbias.n361 4.5005
R20336 Vbias.n484 Vbias.n313 4.5005
R20337 Vbias.n487 Vbias.n311 4.5005
R20338 Vbias.n560 Vbias.n559 4.5005
R20339 Vbias.n621 Vbias.n260 4.5005
R20340 Vbias.n624 Vbias.n258 4.5005
R20341 Vbias.n216 Vbias.n215 4.5005
R20342 Vbias.n746 Vbias.n168 4.5005
R20343 Vbias.n743 Vbias.n170 4.5005
R20344 Vbias.n808 Vbias.n807 4.5005
R20345 Vbias.n871 Vbias.n123 4.5005
R20346 Vbias.n874 Vbias.n121 4.5005
R20347 Vbias.n80 Vbias.n79 4.5005
R20348 Vbias.n950 Vbias.n38 4.5005
R20349 Vbias.n952 Vbias.n36 4.5005
R20350 Vbias.n420 Vbias.n419 4.5005
R20351 Vbias.n365 Vbias.n364 4.5005
R20352 Vbias.n493 Vbias.n308 4.5005
R20353 Vbias.n490 Vbias.n310 4.5005
R20354 Vbias.n557 Vbias.n556 4.5005
R20355 Vbias.n630 Vbias.n255 4.5005
R20356 Vbias.n627 Vbias.n257 4.5005
R20357 Vbias.n219 Vbias.n218 4.5005
R20358 Vbias.n737 Vbias.n173 4.5005
R20359 Vbias.n740 Vbias.n171 4.5005
R20360 Vbias.n811 Vbias.n810 4.5005
R20361 Vbias.n868 Vbias.n124 4.5005
R20362 Vbias.n865 Vbias.n126 4.5005
R20363 Vbias.n77 Vbias.n76 4.5005
R20364 Vbias.n957 Vbias.n33 4.5005
R20365 Vbias.n955 Vbias.n35 4.5005
R20366 Vbias.n417 Vbias.n416 4.5005
R20367 Vbias.n368 Vbias.n367 4.5005
R20368 Vbias.n496 Vbias.n307 4.5005
R20369 Vbias.n499 Vbias.n305 4.5005
R20370 Vbias.n554 Vbias.n553 4.5005
R20371 Vbias.n633 Vbias.n254 4.5005
R20372 Vbias.n636 Vbias.n252 4.5005
R20373 Vbias.n222 Vbias.n221 4.5005
R20374 Vbias.n734 Vbias.n174 4.5005
R20375 Vbias.n731 Vbias.n176 4.5005
R20376 Vbias.n814 Vbias.n813 4.5005
R20377 Vbias.n859 Vbias.n129 4.5005
R20378 Vbias.n862 Vbias.n127 4.5005
R20379 Vbias.n74 Vbias.n73 4.5005
R20380 Vbias.n960 Vbias.n32 4.5005
R20381 Vbias.n962 Vbias.n30 4.5005
R20382 Vbias.n414 Vbias.n413 4.5005
R20383 Vbias.n371 Vbias.n370 4.5005
R20384 Vbias.n505 Vbias.n302 4.5005
R20385 Vbias.n502 Vbias.n304 4.5005
R20386 Vbias.n551 Vbias.n550 4.5005
R20387 Vbias.n642 Vbias.n249 4.5005
R20388 Vbias.n639 Vbias.n251 4.5005
R20389 Vbias.n225 Vbias.n224 4.5005
R20390 Vbias.n725 Vbias.n179 4.5005
R20391 Vbias.n728 Vbias.n177 4.5005
R20392 Vbias.n817 Vbias.n816 4.5005
R20393 Vbias.n856 Vbias.n130 4.5005
R20394 Vbias.n853 Vbias.n132 4.5005
R20395 Vbias.n71 Vbias.n70 4.5005
R20396 Vbias.n967 Vbias.n27 4.5005
R20397 Vbias.n965 Vbias.n29 4.5005
R20398 Vbias.n411 Vbias.n410 4.5005
R20399 Vbias.n374 Vbias.n373 4.5005
R20400 Vbias.n508 Vbias.n301 4.5005
R20401 Vbias.n511 Vbias.n299 4.5005
R20402 Vbias.n548 Vbias.n547 4.5005
R20403 Vbias.n645 Vbias.n248 4.5005
R20404 Vbias.n648 Vbias.n246 4.5005
R20405 Vbias.n228 Vbias.n227 4.5005
R20406 Vbias.n722 Vbias.n180 4.5005
R20407 Vbias.n719 Vbias.n182 4.5005
R20408 Vbias.n820 Vbias.n819 4.5005
R20409 Vbias.n847 Vbias.n135 4.5005
R20410 Vbias.n850 Vbias.n133 4.5005
R20411 Vbias.n68 Vbias.n67 4.5005
R20412 Vbias.n970 Vbias.n26 4.5005
R20413 Vbias.n972 Vbias.n24 4.5005
R20414 Vbias.n408 Vbias.n407 4.5005
R20415 Vbias.n377 Vbias.n376 4.5005
R20416 Vbias.n517 Vbias.n296 4.5005
R20417 Vbias.n514 Vbias.n298 4.5005
R20418 Vbias.n545 Vbias.n544 4.5005
R20419 Vbias.n654 Vbias.n243 4.5005
R20420 Vbias.n651 Vbias.n245 4.5005
R20421 Vbias.n231 Vbias.n230 4.5005
R20422 Vbias.n713 Vbias.n185 4.5005
R20423 Vbias.n716 Vbias.n183 4.5005
R20424 Vbias.n823 Vbias.n822 4.5005
R20425 Vbias.n844 Vbias.n136 4.5005
R20426 Vbias.n841 Vbias.n138 4.5005
R20427 Vbias.n65 Vbias.n64 4.5005
R20428 Vbias.n977 Vbias.n21 4.5005
R20429 Vbias.n975 Vbias.n23 4.5005
R20430 Vbias.n405 Vbias.n404 4.5005
R20431 Vbias.n380 Vbias.n379 4.5005
R20432 Vbias.n520 Vbias.n295 4.5005
R20433 Vbias.n523 Vbias.n293 4.5005
R20434 Vbias.n542 Vbias.n541 4.5005
R20435 Vbias.n657 Vbias.n242 4.5005
R20436 Vbias.n660 Vbias.n240 4.5005
R20437 Vbias.n234 Vbias.n233 4.5005
R20438 Vbias.n710 Vbias.n186 4.5005
R20439 Vbias.n707 Vbias.n188 4.5005
R20440 Vbias.n826 Vbias.n825 4.5005
R20441 Vbias.n835 Vbias.n141 4.5005
R20442 Vbias.n838 Vbias.n139 4.5005
R20443 Vbias.n62 Vbias.n61 4.5005
R20444 Vbias.n980 Vbias.n18 4.5005
R20445 Vbias.n982 Vbias.n16 4.5005
R20446 Vbias.n402 Vbias.n338 4.5005
R20447 Vbias.n340 Vbias.n339 4.5005
R20448 Vbias.n399 Vbias.n341 4.5005
R20449 Vbias.n526 Vbias.n525 4.5005
R20450 Vbias.n539 Vbias.n285 4.5005
R20451 Vbias.n536 Vbias.n287 4.5005
R20452 Vbias.n663 Vbias.n662 4.5005
R20453 Vbias.n694 Vbias.n236 4.5005
R20454 Vbias.n691 Vbias.n238 4.5005
R20455 Vbias.n704 Vbias.n703 4.5005
R20456 Vbias.n829 Vbias.n144 4.5005
R20457 Vbias.n832 Vbias.n142 4.5005
R20458 Vbias.n672 Vbias.n671 4.5005
R20459 Vbias.n988 Vbias.n11 4.5005
R20460 Vbias.n14 Vbias.n13 4.5005
R20461 Vbias.n985 Vbias.n15 4.5005
R20462 Vbias.n994 Vbias.n6 4.5005
R20463 Vbias.n59 Vbias.n58 4.5005
R20464 Vbias.n918 Vbias.n57 4.5005
R20465 Vbias.n8 Vbias.n7 4.5005
R20466 Vbias.n991 Vbias.n10 4.5005
R20467 Vbias.n100 Vbias.n60 4.5005
R20468 Vbias.n914 Vbias.n102 4.5005
R20469 Vbias.n675 Vbias.n674 4.5005
R20470 Vbias.n680 Vbias.n678 4.5005
R20471 Vbias.n907 Vbias.n906 4.5005
R20472 Vbias.n788 Vbias.n145 4.5005
R20473 Vbias.n684 Vbias.n683 4.5005
R20474 Vbias.n701 Vbias.n189 4.5005
R20475 Vbias.n147 Vbias.n146 4.5005
R20476 Vbias.n784 Vbias.n149 4.5005
R20477 Vbias.n192 Vbias.n191 4.5005
R20478 Vbias.n697 Vbias.n194 4.5005
R20479 Vbias.n196 Vbias.n195 4.5005
R20480 Vbias.n281 Vbias.n280 4.5005
R20481 Vbias.n666 Vbias.n665 4.5005
R20482 Vbias.n533 Vbias.n288 4.5005
R20483 Vbias.n583 Vbias.n279 4.5005
R20484 Vbias.n580 Vbias.n284 4.5005
R20485 Vbias.n290 Vbias.n289 4.5005
R20486 Vbias.n529 Vbias.n292 4.5005
R20487 Vbias.n330 Vbias.n329 4.5005
R20488 Vbias.n446 Vbias.n334 4.5005
R20489 Vbias.n396 Vbias.n395 4.5005
R20490 Vbias.n388 Vbias.n383 4.5005
R20491 Vbias.n336 Vbias.n335 4.5005
R20492 Vbias.n443 Vbias.n337 4.5005
R20493 Vbias.n59 Vbias 3.50727
R20494 Vbias Vbias.n918 3.50727
R20495 Vbias.n100 Vbias 3.50727
R20496 Vbias.n914 Vbias 3.50727
R20497 Vbias Vbias.n907 3.50727
R20498 Vbias Vbias.n788 3.50727
R20499 Vbias Vbias.n147 3.50727
R20500 Vbias.n784 Vbias 3.50727
R20501 Vbias Vbias.n196 3.50727
R20502 Vbias.n281 Vbias 3.50727
R20503 Vbias Vbias.n583 3.50727
R20504 Vbias.n580 Vbias 3.50727
R20505 Vbias Vbias.n330 3.50727
R20506 Vbias Vbias.n446 3.50727
R20507 Vbias Vbias.n336 3.50727
R20508 Vbias.n443 Vbias 3.50727
R20509 Vbias.n995 Vbias.n994 3.4105
R20510 Vbias.n985 Vbias.n984 3.4105
R20511 Vbias.n983 Vbias.n982 3.4105
R20512 Vbias.n975 Vbias.n974 3.4105
R20513 Vbias.n973 Vbias.n972 3.4105
R20514 Vbias.n965 Vbias.n964 3.4105
R20515 Vbias.n963 Vbias.n962 3.4105
R20516 Vbias.n955 Vbias.n954 3.4105
R20517 Vbias.n953 Vbias.n952 3.4105
R20518 Vbias.n945 Vbias.n944 3.4105
R20519 Vbias.n943 Vbias.n942 3.4105
R20520 Vbias.n935 Vbias.n934 3.4105
R20521 Vbias.n933 Vbias.n932 3.4105
R20522 Vbias.n925 Vbias.n924 3.4105
R20523 Vbias.n923 Vbias.n922 3.4105
R20524 Vbias.n920 Vbias.n919 3.4105
R20525 Vbias.n928 Vbias.n927 3.4105
R20526 Vbias.n930 Vbias.n929 3.4105
R20527 Vbias.n938 Vbias.n937 3.4105
R20528 Vbias.n940 Vbias.n939 3.4105
R20529 Vbias.n948 Vbias.n947 3.4105
R20530 Vbias.n950 Vbias.n949 3.4105
R20531 Vbias.n958 Vbias.n957 3.4105
R20532 Vbias.n960 Vbias.n959 3.4105
R20533 Vbias.n968 Vbias.n967 3.4105
R20534 Vbias.n970 Vbias.n969 3.4105
R20535 Vbias.n978 Vbias.n977 3.4105
R20536 Vbias.n980 Vbias.n979 3.4105
R20537 Vbias.n20 Vbias.n14 3.4105
R20538 Vbias.n19 Vbias.n8 3.4105
R20539 Vbias.n991 Vbias.n990 3.4105
R20540 Vbias.n989 Vbias.n988 3.4105
R20541 Vbias.n63 Vbias.n62 3.4105
R20542 Vbias.n66 Vbias.n65 3.4105
R20543 Vbias.n69 Vbias.n68 3.4105
R20544 Vbias.n72 Vbias.n71 3.4105
R20545 Vbias.n75 Vbias.n74 3.4105
R20546 Vbias.n78 Vbias.n77 3.4105
R20547 Vbias.n81 Vbias.n80 3.4105
R20548 Vbias.n84 Vbias.n83 3.4105
R20549 Vbias.n87 Vbias.n86 3.4105
R20550 Vbias.n90 Vbias.n89 3.4105
R20551 Vbias.n93 Vbias.n92 3.4105
R20552 Vbias.n96 Vbias.n95 3.4105
R20553 Vbias.n99 Vbias.n98 3.4105
R20554 Vbias.n913 Vbias.n912 3.4105
R20555 Vbias.n901 Vbias.n900 3.4105
R20556 Vbias.n899 Vbias.n898 3.4105
R20557 Vbias.n889 Vbias.n888 3.4105
R20558 Vbias.n887 Vbias.n886 3.4105
R20559 Vbias.n877 Vbias.n876 3.4105
R20560 Vbias.n875 Vbias.n874 3.4105
R20561 Vbias.n865 Vbias.n864 3.4105
R20562 Vbias.n863 Vbias.n862 3.4105
R20563 Vbias.n853 Vbias.n852 3.4105
R20564 Vbias.n851 Vbias.n850 3.4105
R20565 Vbias.n841 Vbias.n840 3.4105
R20566 Vbias.n839 Vbias.n838 3.4105
R20567 Vbias.n673 Vbias.n672 3.4105
R20568 Vbias.n676 Vbias.n675 3.4105
R20569 Vbias.n681 Vbias.n680 3.4105
R20570 Vbias.n833 Vbias.n832 3.4105
R20571 Vbias.n835 Vbias.n834 3.4105
R20572 Vbias.n845 Vbias.n844 3.4105
R20573 Vbias.n847 Vbias.n846 3.4105
R20574 Vbias.n857 Vbias.n856 3.4105
R20575 Vbias.n859 Vbias.n858 3.4105
R20576 Vbias.n869 Vbias.n868 3.4105
R20577 Vbias.n871 Vbias.n870 3.4105
R20578 Vbias.n881 Vbias.n880 3.4105
R20579 Vbias.n883 Vbias.n882 3.4105
R20580 Vbias.n893 Vbias.n892 3.4105
R20581 Vbias.n895 Vbias.n894 3.4105
R20582 Vbias.n905 Vbias.n904 3.4105
R20583 Vbias.n909 Vbias.n908 3.4105
R20584 Vbias.n791 Vbias.n790 3.4105
R20585 Vbias.n794 Vbias.n793 3.4105
R20586 Vbias.n797 Vbias.n796 3.4105
R20587 Vbias.n800 Vbias.n799 3.4105
R20588 Vbias.n803 Vbias.n802 3.4105
R20589 Vbias.n806 Vbias.n805 3.4105
R20590 Vbias.n809 Vbias.n808 3.4105
R20591 Vbias.n812 Vbias.n811 3.4105
R20592 Vbias.n815 Vbias.n814 3.4105
R20593 Vbias.n818 Vbias.n817 3.4105
R20594 Vbias.n821 Vbias.n820 3.4105
R20595 Vbias.n824 Vbias.n823 3.4105
R20596 Vbias.n827 Vbias.n826 3.4105
R20597 Vbias.n829 Vbias.n828 3.4105
R20598 Vbias.n685 Vbias.n684 3.4105
R20599 Vbias.n702 Vbias.n701 3.4105
R20600 Vbias.n705 Vbias.n704 3.4105
R20601 Vbias.n707 Vbias.n706 3.4105
R20602 Vbias.n717 Vbias.n716 3.4105
R20603 Vbias.n719 Vbias.n718 3.4105
R20604 Vbias.n729 Vbias.n728 3.4105
R20605 Vbias.n731 Vbias.n730 3.4105
R20606 Vbias.n741 Vbias.n740 3.4105
R20607 Vbias.n743 Vbias.n742 3.4105
R20608 Vbias.n753 Vbias.n752 3.4105
R20609 Vbias.n755 Vbias.n754 3.4105
R20610 Vbias.n765 Vbias.n764 3.4105
R20611 Vbias.n767 Vbias.n766 3.4105
R20612 Vbias.n777 Vbias.n776 3.4105
R20613 Vbias.n779 Vbias.n778 3.4105
R20614 Vbias.n783 Vbias.n782 3.4105
R20615 Vbias.n773 Vbias.n772 3.4105
R20616 Vbias.n771 Vbias.n770 3.4105
R20617 Vbias.n761 Vbias.n760 3.4105
R20618 Vbias.n759 Vbias.n758 3.4105
R20619 Vbias.n749 Vbias.n748 3.4105
R20620 Vbias.n747 Vbias.n746 3.4105
R20621 Vbias.n737 Vbias.n736 3.4105
R20622 Vbias.n735 Vbias.n734 3.4105
R20623 Vbias.n725 Vbias.n724 3.4105
R20624 Vbias.n723 Vbias.n722 3.4105
R20625 Vbias.n713 Vbias.n712 3.4105
R20626 Vbias.n711 Vbias.n710 3.4105
R20627 Vbias.n691 Vbias.n690 3.4105
R20628 Vbias.n689 Vbias.n192 3.4105
R20629 Vbias.n697 Vbias.n696 3.4105
R20630 Vbias.n695 Vbias.n694 3.4105
R20631 Vbias.n235 Vbias.n234 3.4105
R20632 Vbias.n232 Vbias.n231 3.4105
R20633 Vbias.n229 Vbias.n228 3.4105
R20634 Vbias.n226 Vbias.n225 3.4105
R20635 Vbias.n223 Vbias.n222 3.4105
R20636 Vbias.n220 Vbias.n219 3.4105
R20637 Vbias.n217 Vbias.n216 3.4105
R20638 Vbias.n214 Vbias.n213 3.4105
R20639 Vbias.n211 Vbias.n210 3.4105
R20640 Vbias.n208 Vbias.n207 3.4105
R20641 Vbias.n205 Vbias.n204 3.4105
R20642 Vbias.n202 Vbias.n201 3.4105
R20643 Vbias.n199 Vbias.n198 3.4105
R20644 Vbias.n589 Vbias.n588 3.4105
R20645 Vbias.n591 Vbias.n590 3.4105
R20646 Vbias.n601 Vbias.n600 3.4105
R20647 Vbias.n603 Vbias.n602 3.4105
R20648 Vbias.n613 Vbias.n612 3.4105
R20649 Vbias.n615 Vbias.n614 3.4105
R20650 Vbias.n625 Vbias.n624 3.4105
R20651 Vbias.n627 Vbias.n626 3.4105
R20652 Vbias.n637 Vbias.n636 3.4105
R20653 Vbias.n639 Vbias.n638 3.4105
R20654 Vbias.n649 Vbias.n648 3.4105
R20655 Vbias.n651 Vbias.n650 3.4105
R20656 Vbias.n661 Vbias.n660 3.4105
R20657 Vbias.n664 Vbias.n663 3.4105
R20658 Vbias.n667 Vbias.n666 3.4105
R20659 Vbias.n534 Vbias.n533 3.4105
R20660 Vbias.n536 Vbias.n535 3.4105
R20661 Vbias.n657 Vbias.n656 3.4105
R20662 Vbias.n655 Vbias.n654 3.4105
R20663 Vbias.n645 Vbias.n644 3.4105
R20664 Vbias.n643 Vbias.n642 3.4105
R20665 Vbias.n633 Vbias.n632 3.4105
R20666 Vbias.n631 Vbias.n630 3.4105
R20667 Vbias.n621 Vbias.n620 3.4105
R20668 Vbias.n619 Vbias.n618 3.4105
R20669 Vbias.n609 Vbias.n608 3.4105
R20670 Vbias.n607 Vbias.n606 3.4105
R20671 Vbias.n597 Vbias.n596 3.4105
R20672 Vbias.n595 Vbias.n594 3.4105
R20673 Vbias.n585 Vbias.n584 3.4105
R20674 Vbias.n579 Vbias.n578 3.4105
R20675 Vbias.n576 Vbias.n575 3.4105
R20676 Vbias.n573 Vbias.n572 3.4105
R20677 Vbias.n570 Vbias.n569 3.4105
R20678 Vbias.n567 Vbias.n566 3.4105
R20679 Vbias.n564 Vbias.n563 3.4105
R20680 Vbias.n561 Vbias.n560 3.4105
R20681 Vbias.n558 Vbias.n557 3.4105
R20682 Vbias.n555 Vbias.n554 3.4105
R20683 Vbias.n552 Vbias.n551 3.4105
R20684 Vbias.n549 Vbias.n548 3.4105
R20685 Vbias.n546 Vbias.n545 3.4105
R20686 Vbias.n543 Vbias.n542 3.4105
R20687 Vbias.n540 Vbias.n539 3.4105
R20688 Vbias.n391 Vbias.n290 3.4105
R20689 Vbias.n529 Vbias.n528 3.4105
R20690 Vbias.n527 Vbias.n526 3.4105
R20691 Vbias.n524 Vbias.n523 3.4105
R20692 Vbias.n514 Vbias.n513 3.4105
R20693 Vbias.n512 Vbias.n511 3.4105
R20694 Vbias.n502 Vbias.n501 3.4105
R20695 Vbias.n500 Vbias.n499 3.4105
R20696 Vbias.n490 Vbias.n489 3.4105
R20697 Vbias.n488 Vbias.n487 3.4105
R20698 Vbias.n478 Vbias.n477 3.4105
R20699 Vbias.n476 Vbias.n475 3.4105
R20700 Vbias.n466 Vbias.n465 3.4105
R20701 Vbias.n464 Vbias.n463 3.4105
R20702 Vbias.n454 Vbias.n453 3.4105
R20703 Vbias.n452 Vbias.n451 3.4105
R20704 Vbias.n448 Vbias.n447 3.4105
R20705 Vbias.n458 Vbias.n457 3.4105
R20706 Vbias.n460 Vbias.n459 3.4105
R20707 Vbias.n470 Vbias.n469 3.4105
R20708 Vbias.n472 Vbias.n471 3.4105
R20709 Vbias.n482 Vbias.n481 3.4105
R20710 Vbias.n484 Vbias.n483 3.4105
R20711 Vbias.n494 Vbias.n493 3.4105
R20712 Vbias.n496 Vbias.n495 3.4105
R20713 Vbias.n506 Vbias.n505 3.4105
R20714 Vbias.n508 Vbias.n507 3.4105
R20715 Vbias.n518 Vbias.n517 3.4105
R20716 Vbias.n520 Vbias.n519 3.4105
R20717 Vbias.n399 Vbias.n398 3.4105
R20718 Vbias.n397 Vbias.n396 3.4105
R20719 Vbias.n389 Vbias.n388 3.4105
R20720 Vbias.n382 Vbias.n340 3.4105
R20721 Vbias.n381 Vbias.n380 3.4105
R20722 Vbias.n378 Vbias.n377 3.4105
R20723 Vbias.n375 Vbias.n374 3.4105
R20724 Vbias.n372 Vbias.n371 3.4105
R20725 Vbias.n369 Vbias.n368 3.4105
R20726 Vbias.n366 Vbias.n365 3.4105
R20727 Vbias.n363 Vbias.n362 3.4105
R20728 Vbias.n360 Vbias.n359 3.4105
R20729 Vbias.n357 Vbias.n356 3.4105
R20730 Vbias.n354 Vbias.n353 3.4105
R20731 Vbias.n351 Vbias.n350 3.4105
R20732 Vbias.n348 Vbias.n347 3.4105
R20733 Vbias.n345 Vbias.n344 3.4105
R20734 Vbias.n442 Vbias.n441 3.4105
R20735 Vbias.n439 Vbias.n438 3.4105
R20736 Vbias.n436 Vbias.n435 3.4105
R20737 Vbias.n433 Vbias.n432 3.4105
R20738 Vbias.n430 Vbias.n429 3.4105
R20739 Vbias.n427 Vbias.n426 3.4105
R20740 Vbias.n424 Vbias.n423 3.4105
R20741 Vbias.n421 Vbias.n420 3.4105
R20742 Vbias.n418 Vbias.n417 3.4105
R20743 Vbias.n415 Vbias.n414 3.4105
R20744 Vbias.n412 Vbias.n411 3.4105
R20745 Vbias.n409 Vbias.n408 3.4105
R20746 Vbias.n406 Vbias.n405 3.4105
R20747 Vbias.n403 Vbias.n402 3.4105
R20748 Vbias.n386 Vbias.n385 3.4105
R20749 Vbias.n387 Vbias.n386 2.9408
R20750 Vbias.n441 Vbias.n332 2.9408
R20751 Vbias.n922 Vbias.n921 2.9408
R20752 Vbias.n438 Vbias.n327 2.9408
R20753 Vbias.n926 Vbias.n925 2.9408
R20754 Vbias.n435 Vbias.n324 2.9408
R20755 Vbias.n932 Vbias.n931 2.9408
R20756 Vbias.n432 Vbias.n321 2.9408
R20757 Vbias.n936 Vbias.n935 2.9408
R20758 Vbias.n429 Vbias.n318 2.9408
R20759 Vbias.n942 Vbias.n941 2.9408
R20760 Vbias.n426 Vbias.n315 2.9408
R20761 Vbias.n946 Vbias.n945 2.9408
R20762 Vbias.n423 Vbias.n312 2.9408
R20763 Vbias.n952 Vbias.n951 2.9408
R20764 Vbias.n420 Vbias.n309 2.9408
R20765 Vbias.n956 Vbias.n955 2.9408
R20766 Vbias.n417 Vbias.n306 2.9408
R20767 Vbias.n962 Vbias.n961 2.9408
R20768 Vbias.n414 Vbias.n303 2.9408
R20769 Vbias.n966 Vbias.n965 2.9408
R20770 Vbias.n411 Vbias.n300 2.9408
R20771 Vbias.n972 Vbias.n971 2.9408
R20772 Vbias.n408 Vbias.n297 2.9408
R20773 Vbias.n976 Vbias.n975 2.9408
R20774 Vbias.n405 Vbias.n294 2.9408
R20775 Vbias.n982 Vbias.n981 2.9408
R20776 Vbias.n402 Vbias.n401 2.9408
R20777 Vbias.n986 Vbias.n985 2.9408
R20778 Vbias.n994 Vbias.n993 2.9408
R20779 Vbias.n917 Vbias.n59 2.9408
R20780 Vbias.n444 Vbias.n443 2.9408
R20781 Vbias.n449 Vbias.n332 2.76612
R20782 Vbias.n450 Vbias.n449 2.76612
R20783 Vbias.n450 Vbias.n277 2.76612
R20784 Vbias.n586 Vbias.n277 2.76612
R20785 Vbias.n587 Vbias.n586 2.76612
R20786 Vbias.n587 Vbias.n151 2.76612
R20787 Vbias.n781 Vbias.n151 2.76612
R20788 Vbias.n781 Vbias.n780 2.76612
R20789 Vbias.n780 Vbias.n104 2.76612
R20790 Vbias.n910 Vbias.n104 2.76612
R20791 Vbias.n911 Vbias.n910 2.76612
R20792 Vbias.n911 Vbias.n55 2.76612
R20793 Vbias.n921 Vbias.n55 2.76612
R20794 Vbias.n456 Vbias.n327 2.76612
R20795 Vbias.n456 Vbias.n455 2.76612
R20796 Vbias.n455 Vbias.n274 2.76612
R20797 Vbias.n593 Vbias.n274 2.76612
R20798 Vbias.n593 Vbias.n592 2.76612
R20799 Vbias.n592 Vbias.n154 2.76612
R20800 Vbias.n774 Vbias.n154 2.76612
R20801 Vbias.n775 Vbias.n774 2.76612
R20802 Vbias.n775 Vbias.n107 2.76612
R20803 Vbias.n903 Vbias.n107 2.76612
R20804 Vbias.n903 Vbias.n902 2.76612
R20805 Vbias.n902 Vbias.n52 2.76612
R20806 Vbias.n926 Vbias.n52 2.76612
R20807 Vbias.n461 Vbias.n324 2.76612
R20808 Vbias.n462 Vbias.n461 2.76612
R20809 Vbias.n462 Vbias.n271 2.76612
R20810 Vbias.n598 Vbias.n271 2.76612
R20811 Vbias.n599 Vbias.n598 2.76612
R20812 Vbias.n599 Vbias.n157 2.76612
R20813 Vbias.n769 Vbias.n157 2.76612
R20814 Vbias.n769 Vbias.n768 2.76612
R20815 Vbias.n768 Vbias.n110 2.76612
R20816 Vbias.n896 Vbias.n110 2.76612
R20817 Vbias.n897 Vbias.n896 2.76612
R20818 Vbias.n897 Vbias.n49 2.76612
R20819 Vbias.n931 Vbias.n49 2.76612
R20820 Vbias.n468 Vbias.n321 2.76612
R20821 Vbias.n468 Vbias.n467 2.76612
R20822 Vbias.n467 Vbias.n268 2.76612
R20823 Vbias.n605 Vbias.n268 2.76612
R20824 Vbias.n605 Vbias.n604 2.76612
R20825 Vbias.n604 Vbias.n160 2.76612
R20826 Vbias.n762 Vbias.n160 2.76612
R20827 Vbias.n763 Vbias.n762 2.76612
R20828 Vbias.n763 Vbias.n113 2.76612
R20829 Vbias.n891 Vbias.n113 2.76612
R20830 Vbias.n891 Vbias.n890 2.76612
R20831 Vbias.n890 Vbias.n46 2.76612
R20832 Vbias.n936 Vbias.n46 2.76612
R20833 Vbias.n473 Vbias.n318 2.76612
R20834 Vbias.n474 Vbias.n473 2.76612
R20835 Vbias.n474 Vbias.n265 2.76612
R20836 Vbias.n610 Vbias.n265 2.76612
R20837 Vbias.n611 Vbias.n610 2.76612
R20838 Vbias.n611 Vbias.n163 2.76612
R20839 Vbias.n757 Vbias.n163 2.76612
R20840 Vbias.n757 Vbias.n756 2.76612
R20841 Vbias.n756 Vbias.n116 2.76612
R20842 Vbias.n884 Vbias.n116 2.76612
R20843 Vbias.n885 Vbias.n884 2.76612
R20844 Vbias.n885 Vbias.n43 2.76612
R20845 Vbias.n941 Vbias.n43 2.76612
R20846 Vbias.n480 Vbias.n315 2.76612
R20847 Vbias.n480 Vbias.n479 2.76612
R20848 Vbias.n479 Vbias.n262 2.76612
R20849 Vbias.n617 Vbias.n262 2.76612
R20850 Vbias.n617 Vbias.n616 2.76612
R20851 Vbias.n616 Vbias.n166 2.76612
R20852 Vbias.n750 Vbias.n166 2.76612
R20853 Vbias.n751 Vbias.n750 2.76612
R20854 Vbias.n751 Vbias.n119 2.76612
R20855 Vbias.n879 Vbias.n119 2.76612
R20856 Vbias.n879 Vbias.n878 2.76612
R20857 Vbias.n878 Vbias.n40 2.76612
R20858 Vbias.n946 Vbias.n40 2.76612
R20859 Vbias.n485 Vbias.n312 2.76612
R20860 Vbias.n486 Vbias.n485 2.76612
R20861 Vbias.n486 Vbias.n259 2.76612
R20862 Vbias.n622 Vbias.n259 2.76612
R20863 Vbias.n623 Vbias.n622 2.76612
R20864 Vbias.n623 Vbias.n169 2.76612
R20865 Vbias.n745 Vbias.n169 2.76612
R20866 Vbias.n745 Vbias.n744 2.76612
R20867 Vbias.n744 Vbias.n122 2.76612
R20868 Vbias.n872 Vbias.n122 2.76612
R20869 Vbias.n873 Vbias.n872 2.76612
R20870 Vbias.n873 Vbias.n37 2.76612
R20871 Vbias.n951 Vbias.n37 2.76612
R20872 Vbias.n492 Vbias.n309 2.76612
R20873 Vbias.n492 Vbias.n491 2.76612
R20874 Vbias.n491 Vbias.n256 2.76612
R20875 Vbias.n629 Vbias.n256 2.76612
R20876 Vbias.n629 Vbias.n628 2.76612
R20877 Vbias.n628 Vbias.n172 2.76612
R20878 Vbias.n738 Vbias.n172 2.76612
R20879 Vbias.n739 Vbias.n738 2.76612
R20880 Vbias.n739 Vbias.n125 2.76612
R20881 Vbias.n867 Vbias.n125 2.76612
R20882 Vbias.n867 Vbias.n866 2.76612
R20883 Vbias.n866 Vbias.n34 2.76612
R20884 Vbias.n956 Vbias.n34 2.76612
R20885 Vbias.n497 Vbias.n306 2.76612
R20886 Vbias.n498 Vbias.n497 2.76612
R20887 Vbias.n498 Vbias.n253 2.76612
R20888 Vbias.n634 Vbias.n253 2.76612
R20889 Vbias.n635 Vbias.n634 2.76612
R20890 Vbias.n635 Vbias.n175 2.76612
R20891 Vbias.n733 Vbias.n175 2.76612
R20892 Vbias.n733 Vbias.n732 2.76612
R20893 Vbias.n732 Vbias.n128 2.76612
R20894 Vbias.n860 Vbias.n128 2.76612
R20895 Vbias.n861 Vbias.n860 2.76612
R20896 Vbias.n861 Vbias.n31 2.76612
R20897 Vbias.n961 Vbias.n31 2.76612
R20898 Vbias.n504 Vbias.n303 2.76612
R20899 Vbias.n504 Vbias.n503 2.76612
R20900 Vbias.n503 Vbias.n250 2.76612
R20901 Vbias.n641 Vbias.n250 2.76612
R20902 Vbias.n641 Vbias.n640 2.76612
R20903 Vbias.n640 Vbias.n178 2.76612
R20904 Vbias.n726 Vbias.n178 2.76612
R20905 Vbias.n727 Vbias.n726 2.76612
R20906 Vbias.n727 Vbias.n131 2.76612
R20907 Vbias.n855 Vbias.n131 2.76612
R20908 Vbias.n855 Vbias.n854 2.76612
R20909 Vbias.n854 Vbias.n28 2.76612
R20910 Vbias.n966 Vbias.n28 2.76612
R20911 Vbias.n509 Vbias.n300 2.76612
R20912 Vbias.n510 Vbias.n509 2.76612
R20913 Vbias.n510 Vbias.n247 2.76612
R20914 Vbias.n646 Vbias.n247 2.76612
R20915 Vbias.n647 Vbias.n646 2.76612
R20916 Vbias.n647 Vbias.n181 2.76612
R20917 Vbias.n721 Vbias.n181 2.76612
R20918 Vbias.n721 Vbias.n720 2.76612
R20919 Vbias.n720 Vbias.n134 2.76612
R20920 Vbias.n848 Vbias.n134 2.76612
R20921 Vbias.n849 Vbias.n848 2.76612
R20922 Vbias.n849 Vbias.n25 2.76612
R20923 Vbias.n971 Vbias.n25 2.76612
R20924 Vbias.n516 Vbias.n297 2.76612
R20925 Vbias.n516 Vbias.n515 2.76612
R20926 Vbias.n515 Vbias.n244 2.76612
R20927 Vbias.n653 Vbias.n244 2.76612
R20928 Vbias.n653 Vbias.n652 2.76612
R20929 Vbias.n652 Vbias.n184 2.76612
R20930 Vbias.n714 Vbias.n184 2.76612
R20931 Vbias.n715 Vbias.n714 2.76612
R20932 Vbias.n715 Vbias.n137 2.76612
R20933 Vbias.n843 Vbias.n137 2.76612
R20934 Vbias.n843 Vbias.n842 2.76612
R20935 Vbias.n842 Vbias.n22 2.76612
R20936 Vbias.n976 Vbias.n22 2.76612
R20937 Vbias.n521 Vbias.n294 2.76612
R20938 Vbias.n522 Vbias.n521 2.76612
R20939 Vbias.n522 Vbias.n241 2.76612
R20940 Vbias.n658 Vbias.n241 2.76612
R20941 Vbias.n659 Vbias.n658 2.76612
R20942 Vbias.n659 Vbias.n187 2.76612
R20943 Vbias.n709 Vbias.n187 2.76612
R20944 Vbias.n709 Vbias.n708 2.76612
R20945 Vbias.n708 Vbias.n140 2.76612
R20946 Vbias.n836 Vbias.n140 2.76612
R20947 Vbias.n837 Vbias.n836 2.76612
R20948 Vbias.n837 Vbias.n17 2.76612
R20949 Vbias.n981 Vbias.n17 2.76612
R20950 Vbias.n401 Vbias.n400 2.76612
R20951 Vbias.n400 Vbias.n286 2.76612
R20952 Vbias.n538 Vbias.n286 2.76612
R20953 Vbias.n538 Vbias.n537 2.76612
R20954 Vbias.n537 Vbias.n237 2.76612
R20955 Vbias.n693 Vbias.n237 2.76612
R20956 Vbias.n693 Vbias.n692 2.76612
R20957 Vbias.n692 Vbias.n143 2.76612
R20958 Vbias.n830 Vbias.n143 2.76612
R20959 Vbias.n831 Vbias.n830 2.76612
R20960 Vbias.n831 Vbias.n12 2.76612
R20961 Vbias.n987 Vbias.n12 2.76612
R20962 Vbias.n987 Vbias.n986 2.76612
R20963 Vbias.n917 Vbias.n916 2.76612
R20964 Vbias.n993 Vbias.n992 2.76612
R20965 Vbias.n992 Vbias.n9 2.76612
R20966 Vbias.n916 Vbias.n915 2.76612
R20967 Vbias.n915 Vbias.n101 2.76612
R20968 Vbias.n679 Vbias.n9 2.76612
R20969 Vbias.n679 Vbias.n190 2.76612
R20970 Vbias.n787 Vbias.n101 2.76612
R20971 Vbias.n787 Vbias.n786 2.76612
R20972 Vbias.n700 Vbias.n190 2.76612
R20973 Vbias.n700 Vbias.n699 2.76612
R20974 Vbias.n786 Vbias.n785 2.76612
R20975 Vbias.n785 Vbias.n148 2.76612
R20976 Vbias.n699 Vbias.n698 2.76612
R20977 Vbias.n698 Vbias.n193 2.76612
R20978 Vbias.n282 Vbias.n148 2.76612
R20979 Vbias.n582 Vbias.n282 2.76612
R20980 Vbias.n532 Vbias.n193 2.76612
R20981 Vbias.n532 Vbias.n531 2.76612
R20982 Vbias.n582 Vbias.n581 2.76612
R20983 Vbias.n581 Vbias.n283 2.76612
R20984 Vbias.n531 Vbias.n530 2.76612
R20985 Vbias.n530 Vbias.n291 2.76612
R20986 Vbias.n445 Vbias.n283 2.76612
R20987 Vbias.n445 Vbias.n444 2.76612
R20988 Vbias.n387 Vbias.n291 2.76612
R20989 Vbias.n4 Vbias.n3 2.06591
R20990 Vbias Vbias.n342 1.6647
R20991 Vbias Vbias.n394 1.6647
R20992 Vbias.n392 Vbias 1.6647
R20993 Vbias.n668 Vbias 1.6647
R20994 Vbias Vbias.n688 1.6647
R20995 Vbias.n686 Vbias 1.6647
R20996 Vbias.n677 Vbias 1.6647
R20997 Vbias Vbias.n5 1.6647
R20998 Vbias.n996 Vbias 1.6647
R20999 Vbias.n670 Vbias 1.6647
R21000 Vbias.n682 Vbias 1.6647
R21001 Vbias.n687 Vbias 1.6647
R21002 Vbias.n669 Vbias 1.6647
R21003 Vbias Vbias.n239 1.6647
R21004 Vbias.n393 Vbias 1.6647
R21005 Vbias.n390 Vbias 1.6647
R21006 Vbias Vbias.n997 1.57836
R21007 Vbias.n4 Vbias.n0 1.13456
R21008 Vbias Vbias.n4 0.782551
R21009 Vbias.n997 Vbias 0.412011
R21010 Vbias.n390 Vbias.n342 0.410967
R21011 Vbias.n394 Vbias.n390 0.410967
R21012 Vbias.n394 Vbias.n393 0.410967
R21013 Vbias.n393 Vbias.n392 0.410967
R21014 Vbias.n392 Vbias.n239 0.410967
R21015 Vbias.n668 Vbias.n239 0.410967
R21016 Vbias.n669 Vbias.n668 0.410967
R21017 Vbias.n688 Vbias.n669 0.410967
R21018 Vbias.n688 Vbias.n687 0.410967
R21019 Vbias.n687 Vbias.n686 0.410967
R21020 Vbias.n686 Vbias.n682 0.410967
R21021 Vbias.n682 Vbias.n677 0.410967
R21022 Vbias.n677 Vbias.n670 0.410967
R21023 Vbias.n670 Vbias.n5 0.410967
R21024 Vbias.n996 Vbias.n5 0.410967
R21025 Vbias.n342 Vbias 0.383811
R21026 Vbias.n997 Vbias.n996 0.332633
R21027 Vbias.n995 Vbias 0.252372
R21028 Vbias.n984 Vbias 0.252372
R21029 Vbias.n983 Vbias 0.252372
R21030 Vbias.n974 Vbias 0.252372
R21031 Vbias.n973 Vbias 0.252372
R21032 Vbias.n964 Vbias 0.252372
R21033 Vbias.n963 Vbias 0.252372
R21034 Vbias.n954 Vbias 0.252372
R21035 Vbias.n953 Vbias 0.252372
R21036 Vbias.n944 Vbias 0.252372
R21037 Vbias.n943 Vbias 0.252372
R21038 Vbias.n934 Vbias 0.252372
R21039 Vbias.n933 Vbias 0.252372
R21040 Vbias.n924 Vbias 0.252372
R21041 Vbias.n923 Vbias 0.252372
R21042 Vbias.n919 Vbias 0.252372
R21043 Vbias.n928 Vbias 0.252372
R21044 Vbias.n929 Vbias 0.252372
R21045 Vbias.n938 Vbias 0.252372
R21046 Vbias.n939 Vbias 0.252372
R21047 Vbias.n948 Vbias 0.252372
R21048 Vbias.n949 Vbias 0.252372
R21049 Vbias.n958 Vbias 0.252372
R21050 Vbias.n959 Vbias 0.252372
R21051 Vbias.n968 Vbias 0.252372
R21052 Vbias.n969 Vbias 0.252372
R21053 Vbias.n978 Vbias 0.252372
R21054 Vbias.n979 Vbias 0.252372
R21055 Vbias Vbias.n20 0.252372
R21056 Vbias Vbias.n19 0.252372
R21057 Vbias.n990 Vbias 0.252372
R21058 Vbias.n989 Vbias 0.252372
R21059 Vbias Vbias.n63 0.252372
R21060 Vbias Vbias.n66 0.252372
R21061 Vbias Vbias.n69 0.252372
R21062 Vbias Vbias.n72 0.252372
R21063 Vbias Vbias.n75 0.252372
R21064 Vbias Vbias.n78 0.252372
R21065 Vbias Vbias.n81 0.252372
R21066 Vbias Vbias.n84 0.252372
R21067 Vbias Vbias.n87 0.252372
R21068 Vbias Vbias.n90 0.252372
R21069 Vbias Vbias.n93 0.252372
R21070 Vbias Vbias.n96 0.252372
R21071 Vbias Vbias.n99 0.252372
R21072 Vbias Vbias.n913 0.252372
R21073 Vbias.n900 Vbias 0.252372
R21074 Vbias Vbias.n899 0.252372
R21075 Vbias.n888 Vbias 0.252372
R21076 Vbias Vbias.n887 0.252372
R21077 Vbias.n876 Vbias 0.252372
R21078 Vbias Vbias.n875 0.252372
R21079 Vbias.n864 Vbias 0.252372
R21080 Vbias Vbias.n863 0.252372
R21081 Vbias.n852 Vbias 0.252372
R21082 Vbias Vbias.n851 0.252372
R21083 Vbias.n840 Vbias 0.252372
R21084 Vbias Vbias.n839 0.252372
R21085 Vbias.n673 Vbias 0.252372
R21086 Vbias.n676 Vbias 0.252372
R21087 Vbias.n681 Vbias 0.252372
R21088 Vbias Vbias.n833 0.252372
R21089 Vbias.n834 Vbias 0.252372
R21090 Vbias Vbias.n845 0.252372
R21091 Vbias.n846 Vbias 0.252372
R21092 Vbias Vbias.n857 0.252372
R21093 Vbias.n858 Vbias 0.252372
R21094 Vbias Vbias.n869 0.252372
R21095 Vbias.n870 Vbias 0.252372
R21096 Vbias Vbias.n881 0.252372
R21097 Vbias.n882 Vbias 0.252372
R21098 Vbias Vbias.n893 0.252372
R21099 Vbias.n894 Vbias 0.252372
R21100 Vbias Vbias.n905 0.252372
R21101 Vbias.n908 Vbias 0.252372
R21102 Vbias.n791 Vbias 0.252372
R21103 Vbias.n794 Vbias 0.252372
R21104 Vbias.n797 Vbias 0.252372
R21105 Vbias.n800 Vbias 0.252372
R21106 Vbias.n803 Vbias 0.252372
R21107 Vbias.n806 Vbias 0.252372
R21108 Vbias.n809 Vbias 0.252372
R21109 Vbias.n812 Vbias 0.252372
R21110 Vbias.n815 Vbias 0.252372
R21111 Vbias.n818 Vbias 0.252372
R21112 Vbias.n821 Vbias 0.252372
R21113 Vbias.n824 Vbias 0.252372
R21114 Vbias.n827 Vbias 0.252372
R21115 Vbias.n828 Vbias 0.252372
R21116 Vbias.n685 Vbias 0.252372
R21117 Vbias Vbias.n702 0.252372
R21118 Vbias Vbias.n705 0.252372
R21119 Vbias.n706 Vbias 0.252372
R21120 Vbias Vbias.n717 0.252372
R21121 Vbias.n718 Vbias 0.252372
R21122 Vbias Vbias.n729 0.252372
R21123 Vbias.n730 Vbias 0.252372
R21124 Vbias Vbias.n741 0.252372
R21125 Vbias.n742 Vbias 0.252372
R21126 Vbias Vbias.n753 0.252372
R21127 Vbias.n754 Vbias 0.252372
R21128 Vbias Vbias.n765 0.252372
R21129 Vbias.n766 Vbias 0.252372
R21130 Vbias Vbias.n777 0.252372
R21131 Vbias.n778 Vbias 0.252372
R21132 Vbias Vbias.n783 0.252372
R21133 Vbias.n772 Vbias 0.252372
R21134 Vbias Vbias.n771 0.252372
R21135 Vbias.n760 Vbias 0.252372
R21136 Vbias Vbias.n759 0.252372
R21137 Vbias.n748 Vbias 0.252372
R21138 Vbias Vbias.n747 0.252372
R21139 Vbias.n736 Vbias 0.252372
R21140 Vbias Vbias.n735 0.252372
R21141 Vbias.n724 Vbias 0.252372
R21142 Vbias Vbias.n723 0.252372
R21143 Vbias.n712 Vbias 0.252372
R21144 Vbias Vbias.n711 0.252372
R21145 Vbias.n690 Vbias 0.252372
R21146 Vbias Vbias.n689 0.252372
R21147 Vbias.n696 Vbias 0.252372
R21148 Vbias.n695 Vbias 0.252372
R21149 Vbias.n235 Vbias 0.252372
R21150 Vbias.n232 Vbias 0.252372
R21151 Vbias.n229 Vbias 0.252372
R21152 Vbias.n226 Vbias 0.252372
R21153 Vbias.n223 Vbias 0.252372
R21154 Vbias.n220 Vbias 0.252372
R21155 Vbias.n217 Vbias 0.252372
R21156 Vbias.n214 Vbias 0.252372
R21157 Vbias.n211 Vbias 0.252372
R21158 Vbias.n208 Vbias 0.252372
R21159 Vbias.n205 Vbias 0.252372
R21160 Vbias.n202 Vbias 0.252372
R21161 Vbias.n199 Vbias 0.252372
R21162 Vbias.n589 Vbias 0.252372
R21163 Vbias.n590 Vbias 0.252372
R21164 Vbias.n601 Vbias 0.252372
R21165 Vbias.n602 Vbias 0.252372
R21166 Vbias.n613 Vbias 0.252372
R21167 Vbias.n614 Vbias 0.252372
R21168 Vbias.n625 Vbias 0.252372
R21169 Vbias.n626 Vbias 0.252372
R21170 Vbias.n637 Vbias 0.252372
R21171 Vbias.n638 Vbias 0.252372
R21172 Vbias.n649 Vbias 0.252372
R21173 Vbias.n650 Vbias 0.252372
R21174 Vbias.n661 Vbias 0.252372
R21175 Vbias.n664 Vbias 0.252372
R21176 Vbias.n667 Vbias 0.252372
R21177 Vbias Vbias.n534 0.252372
R21178 Vbias.n535 Vbias 0.252372
R21179 Vbias.n656 Vbias 0.252372
R21180 Vbias.n655 Vbias 0.252372
R21181 Vbias.n644 Vbias 0.252372
R21182 Vbias.n643 Vbias 0.252372
R21183 Vbias.n632 Vbias 0.252372
R21184 Vbias.n631 Vbias 0.252372
R21185 Vbias.n620 Vbias 0.252372
R21186 Vbias.n619 Vbias 0.252372
R21187 Vbias.n608 Vbias 0.252372
R21188 Vbias.n607 Vbias 0.252372
R21189 Vbias.n596 Vbias 0.252372
R21190 Vbias.n595 Vbias 0.252372
R21191 Vbias.n584 Vbias 0.252372
R21192 Vbias Vbias.n579 0.252372
R21193 Vbias Vbias.n576 0.252372
R21194 Vbias Vbias.n573 0.252372
R21195 Vbias Vbias.n570 0.252372
R21196 Vbias Vbias.n567 0.252372
R21197 Vbias Vbias.n564 0.252372
R21198 Vbias Vbias.n561 0.252372
R21199 Vbias Vbias.n558 0.252372
R21200 Vbias Vbias.n555 0.252372
R21201 Vbias Vbias.n552 0.252372
R21202 Vbias Vbias.n549 0.252372
R21203 Vbias Vbias.n546 0.252372
R21204 Vbias Vbias.n543 0.252372
R21205 Vbias Vbias.n540 0.252372
R21206 Vbias.n391 Vbias 0.252372
R21207 Vbias.n528 Vbias 0.252372
R21208 Vbias.n527 Vbias 0.252372
R21209 Vbias.n524 Vbias 0.252372
R21210 Vbias.n513 Vbias 0.252372
R21211 Vbias.n512 Vbias 0.252372
R21212 Vbias.n501 Vbias 0.252372
R21213 Vbias.n500 Vbias 0.252372
R21214 Vbias.n489 Vbias 0.252372
R21215 Vbias.n488 Vbias 0.252372
R21216 Vbias.n477 Vbias 0.252372
R21217 Vbias.n476 Vbias 0.252372
R21218 Vbias.n465 Vbias 0.252372
R21219 Vbias.n464 Vbias 0.252372
R21220 Vbias.n453 Vbias 0.252372
R21221 Vbias.n452 Vbias 0.252372
R21222 Vbias.n447 Vbias 0.252372
R21223 Vbias.n458 Vbias 0.252372
R21224 Vbias.n459 Vbias 0.252372
R21225 Vbias.n470 Vbias 0.252372
R21226 Vbias.n471 Vbias 0.252372
R21227 Vbias.n482 Vbias 0.252372
R21228 Vbias.n483 Vbias 0.252372
R21229 Vbias.n494 Vbias 0.252372
R21230 Vbias.n495 Vbias 0.252372
R21231 Vbias.n506 Vbias 0.252372
R21232 Vbias.n507 Vbias 0.252372
R21233 Vbias.n518 Vbias 0.252372
R21234 Vbias.n519 Vbias 0.252372
R21235 Vbias.n398 Vbias 0.252372
R21236 Vbias Vbias.n397 0.252372
R21237 Vbias.n389 Vbias 0.252372
R21238 Vbias.n382 Vbias 0.252372
R21239 Vbias.n381 Vbias 0.252372
R21240 Vbias.n378 Vbias 0.252372
R21241 Vbias.n375 Vbias 0.252372
R21242 Vbias.n372 Vbias 0.252372
R21243 Vbias.n369 Vbias 0.252372
R21244 Vbias.n366 Vbias 0.252372
R21245 Vbias.n363 Vbias 0.252372
R21246 Vbias.n360 Vbias 0.252372
R21247 Vbias.n357 Vbias 0.252372
R21248 Vbias.n354 Vbias 0.252372
R21249 Vbias.n351 Vbias 0.252372
R21250 Vbias.n348 Vbias 0.252372
R21251 Vbias.n345 Vbias 0.252372
R21252 Vbias Vbias.n442 0.252372
R21253 Vbias Vbias.n439 0.252372
R21254 Vbias Vbias.n436 0.252372
R21255 Vbias Vbias.n433 0.252372
R21256 Vbias Vbias.n430 0.252372
R21257 Vbias Vbias.n427 0.252372
R21258 Vbias Vbias.n424 0.252372
R21259 Vbias Vbias.n421 0.252372
R21260 Vbias Vbias.n418 0.252372
R21261 Vbias Vbias.n415 0.252372
R21262 Vbias Vbias.n412 0.252372
R21263 Vbias Vbias.n409 0.252372
R21264 Vbias Vbias.n406 0.252372
R21265 Vbias Vbias.n403 0.252372
R21266 Vbias.n385 Vbias 0.252372
R21267 Vbias.n344 Vbias.n332 0.175179
R21268 Vbias.n449 Vbias.n448 0.175179
R21269 Vbias.n451 Vbias.n450 0.175179
R21270 Vbias.n578 Vbias.n277 0.175179
R21271 Vbias.n586 Vbias.n585 0.175179
R21272 Vbias.n588 Vbias.n587 0.175179
R21273 Vbias.n198 Vbias.n151 0.175179
R21274 Vbias.n782 Vbias.n781 0.175179
R21275 Vbias.n780 Vbias.n779 0.175179
R21276 Vbias.n790 Vbias.n104 0.175179
R21277 Vbias.n910 Vbias.n909 0.175179
R21278 Vbias.n912 Vbias.n911 0.175179
R21279 Vbias.n98 Vbias.n55 0.175179
R21280 Vbias.n921 Vbias.n920 0.175179
R21281 Vbias.n347 Vbias.n327 0.175179
R21282 Vbias.n457 Vbias.n456 0.175179
R21283 Vbias.n455 Vbias.n454 0.175179
R21284 Vbias.n575 Vbias.n274 0.175179
R21285 Vbias.n594 Vbias.n593 0.175179
R21286 Vbias.n592 Vbias.n591 0.175179
R21287 Vbias.n201 Vbias.n154 0.175179
R21288 Vbias.n774 Vbias.n773 0.175179
R21289 Vbias.n776 Vbias.n775 0.175179
R21290 Vbias.n793 Vbias.n107 0.175179
R21291 Vbias.n904 Vbias.n903 0.175179
R21292 Vbias.n902 Vbias.n901 0.175179
R21293 Vbias.n95 Vbias.n52 0.175179
R21294 Vbias.n927 Vbias.n926 0.175179
R21295 Vbias.n350 Vbias.n324 0.175179
R21296 Vbias.n461 Vbias.n460 0.175179
R21297 Vbias.n463 Vbias.n462 0.175179
R21298 Vbias.n572 Vbias.n271 0.175179
R21299 Vbias.n598 Vbias.n597 0.175179
R21300 Vbias.n600 Vbias.n599 0.175179
R21301 Vbias.n204 Vbias.n157 0.175179
R21302 Vbias.n770 Vbias.n769 0.175179
R21303 Vbias.n768 Vbias.n767 0.175179
R21304 Vbias.n796 Vbias.n110 0.175179
R21305 Vbias.n896 Vbias.n895 0.175179
R21306 Vbias.n898 Vbias.n897 0.175179
R21307 Vbias.n92 Vbias.n49 0.175179
R21308 Vbias.n931 Vbias.n930 0.175179
R21309 Vbias.n353 Vbias.n321 0.175179
R21310 Vbias.n469 Vbias.n468 0.175179
R21311 Vbias.n467 Vbias.n466 0.175179
R21312 Vbias.n569 Vbias.n268 0.175179
R21313 Vbias.n606 Vbias.n605 0.175179
R21314 Vbias.n604 Vbias.n603 0.175179
R21315 Vbias.n207 Vbias.n160 0.175179
R21316 Vbias.n762 Vbias.n761 0.175179
R21317 Vbias.n764 Vbias.n763 0.175179
R21318 Vbias.n799 Vbias.n113 0.175179
R21319 Vbias.n892 Vbias.n891 0.175179
R21320 Vbias.n890 Vbias.n889 0.175179
R21321 Vbias.n89 Vbias.n46 0.175179
R21322 Vbias.n937 Vbias.n936 0.175179
R21323 Vbias.n356 Vbias.n318 0.175179
R21324 Vbias.n473 Vbias.n472 0.175179
R21325 Vbias.n475 Vbias.n474 0.175179
R21326 Vbias.n566 Vbias.n265 0.175179
R21327 Vbias.n610 Vbias.n609 0.175179
R21328 Vbias.n612 Vbias.n611 0.175179
R21329 Vbias.n210 Vbias.n163 0.175179
R21330 Vbias.n758 Vbias.n757 0.175179
R21331 Vbias.n756 Vbias.n755 0.175179
R21332 Vbias.n802 Vbias.n116 0.175179
R21333 Vbias.n884 Vbias.n883 0.175179
R21334 Vbias.n886 Vbias.n885 0.175179
R21335 Vbias.n86 Vbias.n43 0.175179
R21336 Vbias.n941 Vbias.n940 0.175179
R21337 Vbias.n359 Vbias.n315 0.175179
R21338 Vbias.n481 Vbias.n480 0.175179
R21339 Vbias.n479 Vbias.n478 0.175179
R21340 Vbias.n563 Vbias.n262 0.175179
R21341 Vbias.n618 Vbias.n617 0.175179
R21342 Vbias.n616 Vbias.n615 0.175179
R21343 Vbias.n213 Vbias.n166 0.175179
R21344 Vbias.n750 Vbias.n749 0.175179
R21345 Vbias.n752 Vbias.n751 0.175179
R21346 Vbias.n805 Vbias.n119 0.175179
R21347 Vbias.n880 Vbias.n879 0.175179
R21348 Vbias.n878 Vbias.n877 0.175179
R21349 Vbias.n83 Vbias.n40 0.175179
R21350 Vbias.n947 Vbias.n946 0.175179
R21351 Vbias.n362 Vbias.n312 0.175179
R21352 Vbias.n485 Vbias.n484 0.175179
R21353 Vbias.n487 Vbias.n486 0.175179
R21354 Vbias.n560 Vbias.n259 0.175179
R21355 Vbias.n622 Vbias.n621 0.175179
R21356 Vbias.n624 Vbias.n623 0.175179
R21357 Vbias.n216 Vbias.n169 0.175179
R21358 Vbias.n746 Vbias.n745 0.175179
R21359 Vbias.n744 Vbias.n743 0.175179
R21360 Vbias.n808 Vbias.n122 0.175179
R21361 Vbias.n872 Vbias.n871 0.175179
R21362 Vbias.n874 Vbias.n873 0.175179
R21363 Vbias.n80 Vbias.n37 0.175179
R21364 Vbias.n951 Vbias.n950 0.175179
R21365 Vbias.n365 Vbias.n309 0.175179
R21366 Vbias.n493 Vbias.n492 0.175179
R21367 Vbias.n491 Vbias.n490 0.175179
R21368 Vbias.n557 Vbias.n256 0.175179
R21369 Vbias.n630 Vbias.n629 0.175179
R21370 Vbias.n628 Vbias.n627 0.175179
R21371 Vbias.n219 Vbias.n172 0.175179
R21372 Vbias.n738 Vbias.n737 0.175179
R21373 Vbias.n740 Vbias.n739 0.175179
R21374 Vbias.n811 Vbias.n125 0.175179
R21375 Vbias.n868 Vbias.n867 0.175179
R21376 Vbias.n866 Vbias.n865 0.175179
R21377 Vbias.n77 Vbias.n34 0.175179
R21378 Vbias.n957 Vbias.n956 0.175179
R21379 Vbias.n368 Vbias.n306 0.175179
R21380 Vbias.n497 Vbias.n496 0.175179
R21381 Vbias.n499 Vbias.n498 0.175179
R21382 Vbias.n554 Vbias.n253 0.175179
R21383 Vbias.n634 Vbias.n633 0.175179
R21384 Vbias.n636 Vbias.n635 0.175179
R21385 Vbias.n222 Vbias.n175 0.175179
R21386 Vbias.n734 Vbias.n733 0.175179
R21387 Vbias.n732 Vbias.n731 0.175179
R21388 Vbias.n814 Vbias.n128 0.175179
R21389 Vbias.n860 Vbias.n859 0.175179
R21390 Vbias.n862 Vbias.n861 0.175179
R21391 Vbias.n74 Vbias.n31 0.175179
R21392 Vbias.n961 Vbias.n960 0.175179
R21393 Vbias.n371 Vbias.n303 0.175179
R21394 Vbias.n505 Vbias.n504 0.175179
R21395 Vbias.n503 Vbias.n502 0.175179
R21396 Vbias.n551 Vbias.n250 0.175179
R21397 Vbias.n642 Vbias.n641 0.175179
R21398 Vbias.n640 Vbias.n639 0.175179
R21399 Vbias.n225 Vbias.n178 0.175179
R21400 Vbias.n726 Vbias.n725 0.175179
R21401 Vbias.n728 Vbias.n727 0.175179
R21402 Vbias.n817 Vbias.n131 0.175179
R21403 Vbias.n856 Vbias.n855 0.175179
R21404 Vbias.n854 Vbias.n853 0.175179
R21405 Vbias.n71 Vbias.n28 0.175179
R21406 Vbias.n967 Vbias.n966 0.175179
R21407 Vbias.n374 Vbias.n300 0.175179
R21408 Vbias.n509 Vbias.n508 0.175179
R21409 Vbias.n511 Vbias.n510 0.175179
R21410 Vbias.n548 Vbias.n247 0.175179
R21411 Vbias.n646 Vbias.n645 0.175179
R21412 Vbias.n648 Vbias.n647 0.175179
R21413 Vbias.n228 Vbias.n181 0.175179
R21414 Vbias.n722 Vbias.n721 0.175179
R21415 Vbias.n720 Vbias.n719 0.175179
R21416 Vbias.n820 Vbias.n134 0.175179
R21417 Vbias.n848 Vbias.n847 0.175179
R21418 Vbias.n850 Vbias.n849 0.175179
R21419 Vbias.n68 Vbias.n25 0.175179
R21420 Vbias.n971 Vbias.n970 0.175179
R21421 Vbias.n377 Vbias.n297 0.175179
R21422 Vbias.n517 Vbias.n516 0.175179
R21423 Vbias.n515 Vbias.n514 0.175179
R21424 Vbias.n545 Vbias.n244 0.175179
R21425 Vbias.n654 Vbias.n653 0.175179
R21426 Vbias.n652 Vbias.n651 0.175179
R21427 Vbias.n231 Vbias.n184 0.175179
R21428 Vbias.n714 Vbias.n713 0.175179
R21429 Vbias.n716 Vbias.n715 0.175179
R21430 Vbias.n823 Vbias.n137 0.175179
R21431 Vbias.n844 Vbias.n843 0.175179
R21432 Vbias.n842 Vbias.n841 0.175179
R21433 Vbias.n65 Vbias.n22 0.175179
R21434 Vbias.n977 Vbias.n976 0.175179
R21435 Vbias.n380 Vbias.n294 0.175179
R21436 Vbias.n521 Vbias.n520 0.175179
R21437 Vbias.n523 Vbias.n522 0.175179
R21438 Vbias.n542 Vbias.n241 0.175179
R21439 Vbias.n658 Vbias.n657 0.175179
R21440 Vbias.n660 Vbias.n659 0.175179
R21441 Vbias.n234 Vbias.n187 0.175179
R21442 Vbias.n710 Vbias.n709 0.175179
R21443 Vbias.n708 Vbias.n707 0.175179
R21444 Vbias.n826 Vbias.n140 0.175179
R21445 Vbias.n836 Vbias.n835 0.175179
R21446 Vbias.n838 Vbias.n837 0.175179
R21447 Vbias.n62 Vbias.n17 0.175179
R21448 Vbias.n981 Vbias.n980 0.175179
R21449 Vbias.n401 Vbias.n340 0.175179
R21450 Vbias.n400 Vbias.n399 0.175179
R21451 Vbias.n526 Vbias.n286 0.175179
R21452 Vbias.n539 Vbias.n538 0.175179
R21453 Vbias.n537 Vbias.n536 0.175179
R21454 Vbias.n663 Vbias.n237 0.175179
R21455 Vbias.n694 Vbias.n693 0.175179
R21456 Vbias.n692 Vbias.n691 0.175179
R21457 Vbias.n704 Vbias.n143 0.175179
R21458 Vbias.n830 Vbias.n829 0.175179
R21459 Vbias.n832 Vbias.n831 0.175179
R21460 Vbias.n672 Vbias.n12 0.175179
R21461 Vbias.n988 Vbias.n987 0.175179
R21462 Vbias.n986 Vbias.n14 0.175179
R21463 Vbias.n918 Vbias.n917 0.175179
R21464 Vbias.n993 Vbias.n8 0.175179
R21465 Vbias.n992 Vbias.n991 0.175179
R21466 Vbias.n916 Vbias.n100 0.175179
R21467 Vbias.n915 Vbias.n914 0.175179
R21468 Vbias.n675 Vbias.n9 0.175179
R21469 Vbias.n680 Vbias.n679 0.175179
R21470 Vbias.n907 Vbias.n101 0.175179
R21471 Vbias.n788 Vbias.n787 0.175179
R21472 Vbias.n684 Vbias.n190 0.175179
R21473 Vbias.n701 Vbias.n700 0.175179
R21474 Vbias.n786 Vbias.n147 0.175179
R21475 Vbias.n785 Vbias.n784 0.175179
R21476 Vbias.n699 Vbias.n192 0.175179
R21477 Vbias.n698 Vbias.n697 0.175179
R21478 Vbias.n196 Vbias.n148 0.175179
R21479 Vbias.n282 Vbias.n281 0.175179
R21480 Vbias.n666 Vbias.n193 0.175179
R21481 Vbias.n533 Vbias.n532 0.175179
R21482 Vbias.n583 Vbias.n582 0.175179
R21483 Vbias.n581 Vbias.n580 0.175179
R21484 Vbias.n531 Vbias.n290 0.175179
R21485 Vbias.n530 Vbias.n529 0.175179
R21486 Vbias.n330 Vbias.n283 0.175179
R21487 Vbias.n446 Vbias.n445 0.175179
R21488 Vbias.n396 Vbias.n291 0.175179
R21489 Vbias.n388 Vbias.n387 0.175179
R21490 Vbias.n444 Vbias.n336 0.175179
R21491 Vbias.n397 Vbias 0.0972718
R21492 Vbias Vbias.n391 0.0972718
R21493 Vbias Vbias.n667 0.0972718
R21494 Vbias.n689 Vbias 0.0972718
R21495 Vbias Vbias.n685 0.0972718
R21496 Vbias Vbias.n676 0.0972718
R21497 Vbias.n19 Vbias 0.0972718
R21498 Vbias Vbias.n995 0.0972718
R21499 Vbias.n984 Vbias 0.0972718
R21500 Vbias Vbias.n983 0.0972718
R21501 Vbias.n974 Vbias 0.0972718
R21502 Vbias Vbias.n973 0.0972718
R21503 Vbias.n964 Vbias 0.0972718
R21504 Vbias Vbias.n963 0.0972718
R21505 Vbias.n954 Vbias 0.0972718
R21506 Vbias Vbias.n953 0.0972718
R21507 Vbias.n944 Vbias 0.0972718
R21508 Vbias Vbias.n943 0.0972718
R21509 Vbias.n934 Vbias 0.0972718
R21510 Vbias Vbias.n933 0.0972718
R21511 Vbias.n924 Vbias 0.0972718
R21512 Vbias Vbias.n923 0.0972718
R21513 Vbias.n919 Vbias 0.0972718
R21514 Vbias Vbias.n928 0.0972718
R21515 Vbias.n929 Vbias 0.0972718
R21516 Vbias Vbias.n938 0.0972718
R21517 Vbias.n939 Vbias 0.0972718
R21518 Vbias Vbias.n948 0.0972718
R21519 Vbias.n949 Vbias 0.0972718
R21520 Vbias Vbias.n958 0.0972718
R21521 Vbias.n959 Vbias 0.0972718
R21522 Vbias Vbias.n968 0.0972718
R21523 Vbias.n969 Vbias 0.0972718
R21524 Vbias Vbias.n978 0.0972718
R21525 Vbias.n979 Vbias 0.0972718
R21526 Vbias.n20 Vbias 0.0972718
R21527 Vbias.n990 Vbias 0.0972718
R21528 Vbias Vbias.n989 0.0972718
R21529 Vbias.n63 Vbias 0.0972718
R21530 Vbias.n66 Vbias 0.0972718
R21531 Vbias.n69 Vbias 0.0972718
R21532 Vbias.n72 Vbias 0.0972718
R21533 Vbias.n75 Vbias 0.0972718
R21534 Vbias.n78 Vbias 0.0972718
R21535 Vbias.n81 Vbias 0.0972718
R21536 Vbias.n84 Vbias 0.0972718
R21537 Vbias.n87 Vbias 0.0972718
R21538 Vbias.n90 Vbias 0.0972718
R21539 Vbias.n93 Vbias 0.0972718
R21540 Vbias.n96 Vbias 0.0972718
R21541 Vbias.n99 Vbias 0.0972718
R21542 Vbias.n913 Vbias 0.0972718
R21543 Vbias.n900 Vbias 0.0972718
R21544 Vbias.n899 Vbias 0.0972718
R21545 Vbias.n888 Vbias 0.0972718
R21546 Vbias.n887 Vbias 0.0972718
R21547 Vbias.n876 Vbias 0.0972718
R21548 Vbias.n875 Vbias 0.0972718
R21549 Vbias.n864 Vbias 0.0972718
R21550 Vbias.n863 Vbias 0.0972718
R21551 Vbias.n852 Vbias 0.0972718
R21552 Vbias.n851 Vbias 0.0972718
R21553 Vbias.n840 Vbias 0.0972718
R21554 Vbias.n839 Vbias 0.0972718
R21555 Vbias Vbias.n673 0.0972718
R21556 Vbias Vbias.n681 0.0972718
R21557 Vbias.n833 Vbias 0.0972718
R21558 Vbias.n834 Vbias 0.0972718
R21559 Vbias.n845 Vbias 0.0972718
R21560 Vbias.n846 Vbias 0.0972718
R21561 Vbias.n857 Vbias 0.0972718
R21562 Vbias.n858 Vbias 0.0972718
R21563 Vbias.n869 Vbias 0.0972718
R21564 Vbias.n870 Vbias 0.0972718
R21565 Vbias.n881 Vbias 0.0972718
R21566 Vbias.n882 Vbias 0.0972718
R21567 Vbias.n893 Vbias 0.0972718
R21568 Vbias.n894 Vbias 0.0972718
R21569 Vbias.n905 Vbias 0.0972718
R21570 Vbias.n908 Vbias 0.0972718
R21571 Vbias Vbias.n791 0.0972718
R21572 Vbias Vbias.n794 0.0972718
R21573 Vbias Vbias.n797 0.0972718
R21574 Vbias Vbias.n800 0.0972718
R21575 Vbias Vbias.n803 0.0972718
R21576 Vbias Vbias.n806 0.0972718
R21577 Vbias Vbias.n809 0.0972718
R21578 Vbias Vbias.n812 0.0972718
R21579 Vbias Vbias.n815 0.0972718
R21580 Vbias Vbias.n818 0.0972718
R21581 Vbias Vbias.n821 0.0972718
R21582 Vbias Vbias.n824 0.0972718
R21583 Vbias Vbias.n827 0.0972718
R21584 Vbias.n828 Vbias 0.0972718
R21585 Vbias.n702 Vbias 0.0972718
R21586 Vbias.n705 Vbias 0.0972718
R21587 Vbias.n706 Vbias 0.0972718
R21588 Vbias.n717 Vbias 0.0972718
R21589 Vbias.n718 Vbias 0.0972718
R21590 Vbias.n729 Vbias 0.0972718
R21591 Vbias.n730 Vbias 0.0972718
R21592 Vbias.n741 Vbias 0.0972718
R21593 Vbias.n742 Vbias 0.0972718
R21594 Vbias.n753 Vbias 0.0972718
R21595 Vbias.n754 Vbias 0.0972718
R21596 Vbias.n765 Vbias 0.0972718
R21597 Vbias.n766 Vbias 0.0972718
R21598 Vbias.n777 Vbias 0.0972718
R21599 Vbias.n778 Vbias 0.0972718
R21600 Vbias.n783 Vbias 0.0972718
R21601 Vbias.n772 Vbias 0.0972718
R21602 Vbias.n771 Vbias 0.0972718
R21603 Vbias.n760 Vbias 0.0972718
R21604 Vbias.n759 Vbias 0.0972718
R21605 Vbias.n748 Vbias 0.0972718
R21606 Vbias.n747 Vbias 0.0972718
R21607 Vbias.n736 Vbias 0.0972718
R21608 Vbias.n735 Vbias 0.0972718
R21609 Vbias.n724 Vbias 0.0972718
R21610 Vbias.n723 Vbias 0.0972718
R21611 Vbias.n712 Vbias 0.0972718
R21612 Vbias.n711 Vbias 0.0972718
R21613 Vbias.n690 Vbias 0.0972718
R21614 Vbias.n696 Vbias 0.0972718
R21615 Vbias Vbias.n695 0.0972718
R21616 Vbias Vbias.n235 0.0972718
R21617 Vbias Vbias.n232 0.0972718
R21618 Vbias Vbias.n229 0.0972718
R21619 Vbias Vbias.n226 0.0972718
R21620 Vbias Vbias.n223 0.0972718
R21621 Vbias Vbias.n220 0.0972718
R21622 Vbias Vbias.n217 0.0972718
R21623 Vbias Vbias.n214 0.0972718
R21624 Vbias Vbias.n211 0.0972718
R21625 Vbias Vbias.n208 0.0972718
R21626 Vbias Vbias.n205 0.0972718
R21627 Vbias Vbias.n202 0.0972718
R21628 Vbias Vbias.n199 0.0972718
R21629 Vbias Vbias.n589 0.0972718
R21630 Vbias.n590 Vbias 0.0972718
R21631 Vbias Vbias.n601 0.0972718
R21632 Vbias.n602 Vbias 0.0972718
R21633 Vbias Vbias.n613 0.0972718
R21634 Vbias.n614 Vbias 0.0972718
R21635 Vbias Vbias.n625 0.0972718
R21636 Vbias.n626 Vbias 0.0972718
R21637 Vbias Vbias.n637 0.0972718
R21638 Vbias.n638 Vbias 0.0972718
R21639 Vbias Vbias.n649 0.0972718
R21640 Vbias.n650 Vbias 0.0972718
R21641 Vbias Vbias.n661 0.0972718
R21642 Vbias Vbias.n664 0.0972718
R21643 Vbias.n534 Vbias 0.0972718
R21644 Vbias.n535 Vbias 0.0972718
R21645 Vbias.n656 Vbias 0.0972718
R21646 Vbias Vbias.n655 0.0972718
R21647 Vbias.n644 Vbias 0.0972718
R21648 Vbias Vbias.n643 0.0972718
R21649 Vbias.n632 Vbias 0.0972718
R21650 Vbias Vbias.n631 0.0972718
R21651 Vbias.n620 Vbias 0.0972718
R21652 Vbias Vbias.n619 0.0972718
R21653 Vbias.n608 Vbias 0.0972718
R21654 Vbias Vbias.n607 0.0972718
R21655 Vbias.n596 Vbias 0.0972718
R21656 Vbias Vbias.n595 0.0972718
R21657 Vbias.n584 Vbias 0.0972718
R21658 Vbias.n579 Vbias 0.0972718
R21659 Vbias.n576 Vbias 0.0972718
R21660 Vbias.n573 Vbias 0.0972718
R21661 Vbias.n570 Vbias 0.0972718
R21662 Vbias.n567 Vbias 0.0972718
R21663 Vbias.n564 Vbias 0.0972718
R21664 Vbias.n561 Vbias 0.0972718
R21665 Vbias.n558 Vbias 0.0972718
R21666 Vbias.n555 Vbias 0.0972718
R21667 Vbias.n552 Vbias 0.0972718
R21668 Vbias.n549 Vbias 0.0972718
R21669 Vbias.n546 Vbias 0.0972718
R21670 Vbias.n543 Vbias 0.0972718
R21671 Vbias.n540 Vbias 0.0972718
R21672 Vbias.n528 Vbias 0.0972718
R21673 Vbias Vbias.n527 0.0972718
R21674 Vbias Vbias.n524 0.0972718
R21675 Vbias.n513 Vbias 0.0972718
R21676 Vbias Vbias.n512 0.0972718
R21677 Vbias.n501 Vbias 0.0972718
R21678 Vbias Vbias.n500 0.0972718
R21679 Vbias.n489 Vbias 0.0972718
R21680 Vbias Vbias.n488 0.0972718
R21681 Vbias.n477 Vbias 0.0972718
R21682 Vbias Vbias.n476 0.0972718
R21683 Vbias.n465 Vbias 0.0972718
R21684 Vbias Vbias.n464 0.0972718
R21685 Vbias.n453 Vbias 0.0972718
R21686 Vbias Vbias.n452 0.0972718
R21687 Vbias.n447 Vbias 0.0972718
R21688 Vbias Vbias.n458 0.0972718
R21689 Vbias.n459 Vbias 0.0972718
R21690 Vbias Vbias.n470 0.0972718
R21691 Vbias.n471 Vbias 0.0972718
R21692 Vbias Vbias.n482 0.0972718
R21693 Vbias.n483 Vbias 0.0972718
R21694 Vbias Vbias.n494 0.0972718
R21695 Vbias.n495 Vbias 0.0972718
R21696 Vbias Vbias.n506 0.0972718
R21697 Vbias.n507 Vbias 0.0972718
R21698 Vbias Vbias.n518 0.0972718
R21699 Vbias.n519 Vbias 0.0972718
R21700 Vbias.n398 Vbias 0.0972718
R21701 Vbias Vbias.n389 0.0972718
R21702 Vbias Vbias.n382 0.0972718
R21703 Vbias Vbias.n381 0.0972718
R21704 Vbias Vbias.n378 0.0972718
R21705 Vbias Vbias.n375 0.0972718
R21706 Vbias Vbias.n372 0.0972718
R21707 Vbias Vbias.n369 0.0972718
R21708 Vbias Vbias.n366 0.0972718
R21709 Vbias Vbias.n363 0.0972718
R21710 Vbias Vbias.n360 0.0972718
R21711 Vbias Vbias.n357 0.0972718
R21712 Vbias Vbias.n354 0.0972718
R21713 Vbias Vbias.n351 0.0972718
R21714 Vbias Vbias.n348 0.0972718
R21715 Vbias Vbias.n345 0.0972718
R21716 Vbias.n442 Vbias 0.0972718
R21717 Vbias.n439 Vbias 0.0972718
R21718 Vbias.n436 Vbias 0.0972718
R21719 Vbias.n433 Vbias 0.0972718
R21720 Vbias.n430 Vbias 0.0972718
R21721 Vbias.n427 Vbias 0.0972718
R21722 Vbias.n424 Vbias 0.0972718
R21723 Vbias.n421 Vbias 0.0972718
R21724 Vbias.n418 Vbias 0.0972718
R21725 Vbias.n415 Vbias 0.0972718
R21726 Vbias.n412 Vbias 0.0972718
R21727 Vbias.n409 Vbias 0.0972718
R21728 Vbias.n406 Vbias 0.0972718
R21729 Vbias.n403 Vbias 0.0972718
R21730 Vbias.n385 Vbias 0.0972718
R21731 Vbias.n337 Vbias 0.0489375
R21732 Vbias.n383 Vbias 0.0489375
R21733 Vbias.n384 Vbias 0.0489375
R21734 Vbias.n334 Vbias 0.0489375
R21735 Vbias.n292 Vbias 0.0489375
R21736 Vbias.n284 Vbias 0.0489375
R21737 Vbias.n288 Vbias 0.0489375
R21738 Vbias.n280 Vbias 0.0489375
R21739 Vbias.n194 Vbias 0.0489375
R21740 Vbias.n149 Vbias 0.0489375
R21741 Vbias.n189 Vbias 0.0489375
R21742 Vbias.n145 Vbias 0.0489375
R21743 Vbias.n678 Vbias 0.0489375
R21744 Vbias.n102 Vbias 0.0489375
R21745 Vbias.n10 Vbias 0.0489375
R21746 Vbias.n57 Vbias 0.0489375
R21747 Vbias.n58 Vbias 0.0489375
R21748 Vbias.n54 Vbias 0.0489375
R21749 Vbias.n440 Vbias 0.0489375
R21750 Vbias.n343 Vbias 0.0489375
R21751 Vbias.n333 Vbias 0.0489375
R21752 Vbias.n331 Vbias 0.0489375
R21753 Vbias.n577 Vbias 0.0489375
R21754 Vbias.n278 Vbias 0.0489375
R21755 Vbias.n276 Vbias 0.0489375
R21756 Vbias.n197 Vbias 0.0489375
R21757 Vbias.n150 Vbias 0.0489375
R21758 Vbias.n152 Vbias 0.0489375
R21759 Vbias.n789 Vbias 0.0489375
R21760 Vbias.n105 Vbias 0.0489375
R21761 Vbias.n103 Vbias 0.0489375
R21762 Vbias.n97 Vbias 0.0489375
R21763 Vbias.n56 Vbias 0.0489375
R21764 Vbias.n53 Vbias 0.0489375
R21765 Vbias.n437 Vbias 0.0489375
R21766 Vbias.n346 Vbias 0.0489375
R21767 Vbias.n326 Vbias 0.0489375
R21768 Vbias.n328 Vbias 0.0489375
R21769 Vbias.n574 Vbias 0.0489375
R21770 Vbias.n273 Vbias 0.0489375
R21771 Vbias.n275 Vbias 0.0489375
R21772 Vbias.n200 Vbias 0.0489375
R21773 Vbias.n155 Vbias 0.0489375
R21774 Vbias.n153 Vbias 0.0489375
R21775 Vbias.n792 Vbias 0.0489375
R21776 Vbias.n106 Vbias 0.0489375
R21777 Vbias.n108 Vbias 0.0489375
R21778 Vbias.n94 Vbias 0.0489375
R21779 Vbias.n51 Vbias 0.0489375
R21780 Vbias.n48 Vbias 0.0489375
R21781 Vbias.n434 Vbias 0.0489375
R21782 Vbias.n349 Vbias 0.0489375
R21783 Vbias.n325 Vbias 0.0489375
R21784 Vbias.n323 Vbias 0.0489375
R21785 Vbias.n571 Vbias 0.0489375
R21786 Vbias.n272 Vbias 0.0489375
R21787 Vbias.n270 Vbias 0.0489375
R21788 Vbias.n203 Vbias 0.0489375
R21789 Vbias.n156 Vbias 0.0489375
R21790 Vbias.n158 Vbias 0.0489375
R21791 Vbias.n795 Vbias 0.0489375
R21792 Vbias.n111 Vbias 0.0489375
R21793 Vbias.n109 Vbias 0.0489375
R21794 Vbias.n91 Vbias 0.0489375
R21795 Vbias.n50 Vbias 0.0489375
R21796 Vbias.n47 Vbias 0.0489375
R21797 Vbias.n431 Vbias 0.0489375
R21798 Vbias.n352 Vbias 0.0489375
R21799 Vbias.n320 Vbias 0.0489375
R21800 Vbias.n322 Vbias 0.0489375
R21801 Vbias.n568 Vbias 0.0489375
R21802 Vbias.n267 Vbias 0.0489375
R21803 Vbias.n269 Vbias 0.0489375
R21804 Vbias.n206 Vbias 0.0489375
R21805 Vbias.n161 Vbias 0.0489375
R21806 Vbias.n159 Vbias 0.0489375
R21807 Vbias.n798 Vbias 0.0489375
R21808 Vbias.n112 Vbias 0.0489375
R21809 Vbias.n114 Vbias 0.0489375
R21810 Vbias.n88 Vbias 0.0489375
R21811 Vbias.n45 Vbias 0.0489375
R21812 Vbias.n42 Vbias 0.0489375
R21813 Vbias.n428 Vbias 0.0489375
R21814 Vbias.n355 Vbias 0.0489375
R21815 Vbias.n319 Vbias 0.0489375
R21816 Vbias.n317 Vbias 0.0489375
R21817 Vbias.n565 Vbias 0.0489375
R21818 Vbias.n266 Vbias 0.0489375
R21819 Vbias.n264 Vbias 0.0489375
R21820 Vbias.n209 Vbias 0.0489375
R21821 Vbias.n162 Vbias 0.0489375
R21822 Vbias.n164 Vbias 0.0489375
R21823 Vbias.n801 Vbias 0.0489375
R21824 Vbias.n117 Vbias 0.0489375
R21825 Vbias.n115 Vbias 0.0489375
R21826 Vbias.n85 Vbias 0.0489375
R21827 Vbias.n44 Vbias 0.0489375
R21828 Vbias.n41 Vbias 0.0489375
R21829 Vbias.n425 Vbias 0.0489375
R21830 Vbias.n358 Vbias 0.0489375
R21831 Vbias.n314 Vbias 0.0489375
R21832 Vbias.n316 Vbias 0.0489375
R21833 Vbias.n562 Vbias 0.0489375
R21834 Vbias.n261 Vbias 0.0489375
R21835 Vbias.n263 Vbias 0.0489375
R21836 Vbias.n212 Vbias 0.0489375
R21837 Vbias.n167 Vbias 0.0489375
R21838 Vbias.n165 Vbias 0.0489375
R21839 Vbias.n804 Vbias 0.0489375
R21840 Vbias.n118 Vbias 0.0489375
R21841 Vbias.n120 Vbias 0.0489375
R21842 Vbias.n82 Vbias 0.0489375
R21843 Vbias.n39 Vbias 0.0489375
R21844 Vbias.n36 Vbias 0.0489375
R21845 Vbias.n422 Vbias 0.0489375
R21846 Vbias.n361 Vbias 0.0489375
R21847 Vbias.n313 Vbias 0.0489375
R21848 Vbias.n311 Vbias 0.0489375
R21849 Vbias.n559 Vbias 0.0489375
R21850 Vbias.n260 Vbias 0.0489375
R21851 Vbias.n258 Vbias 0.0489375
R21852 Vbias.n215 Vbias 0.0489375
R21853 Vbias.n168 Vbias 0.0489375
R21854 Vbias.n170 Vbias 0.0489375
R21855 Vbias.n807 Vbias 0.0489375
R21856 Vbias.n123 Vbias 0.0489375
R21857 Vbias.n121 Vbias 0.0489375
R21858 Vbias.n79 Vbias 0.0489375
R21859 Vbias.n38 Vbias 0.0489375
R21860 Vbias.n35 Vbias 0.0489375
R21861 Vbias.n419 Vbias 0.0489375
R21862 Vbias.n364 Vbias 0.0489375
R21863 Vbias.n308 Vbias 0.0489375
R21864 Vbias.n310 Vbias 0.0489375
R21865 Vbias.n556 Vbias 0.0489375
R21866 Vbias.n255 Vbias 0.0489375
R21867 Vbias.n257 Vbias 0.0489375
R21868 Vbias.n218 Vbias 0.0489375
R21869 Vbias.n173 Vbias 0.0489375
R21870 Vbias.n171 Vbias 0.0489375
R21871 Vbias.n810 Vbias 0.0489375
R21872 Vbias.n124 Vbias 0.0489375
R21873 Vbias.n126 Vbias 0.0489375
R21874 Vbias.n76 Vbias 0.0489375
R21875 Vbias.n33 Vbias 0.0489375
R21876 Vbias.n30 Vbias 0.0489375
R21877 Vbias.n416 Vbias 0.0489375
R21878 Vbias.n367 Vbias 0.0489375
R21879 Vbias.n307 Vbias 0.0489375
R21880 Vbias.n305 Vbias 0.0489375
R21881 Vbias.n553 Vbias 0.0489375
R21882 Vbias.n254 Vbias 0.0489375
R21883 Vbias.n252 Vbias 0.0489375
R21884 Vbias.n221 Vbias 0.0489375
R21885 Vbias.n174 Vbias 0.0489375
R21886 Vbias.n176 Vbias 0.0489375
R21887 Vbias.n813 Vbias 0.0489375
R21888 Vbias.n129 Vbias 0.0489375
R21889 Vbias.n127 Vbias 0.0489375
R21890 Vbias.n73 Vbias 0.0489375
R21891 Vbias.n32 Vbias 0.0489375
R21892 Vbias.n29 Vbias 0.0489375
R21893 Vbias.n413 Vbias 0.0489375
R21894 Vbias.n370 Vbias 0.0489375
R21895 Vbias.n302 Vbias 0.0489375
R21896 Vbias.n304 Vbias 0.0489375
R21897 Vbias.n550 Vbias 0.0489375
R21898 Vbias.n249 Vbias 0.0489375
R21899 Vbias.n251 Vbias 0.0489375
R21900 Vbias.n224 Vbias 0.0489375
R21901 Vbias.n179 Vbias 0.0489375
R21902 Vbias.n177 Vbias 0.0489375
R21903 Vbias.n816 Vbias 0.0489375
R21904 Vbias.n130 Vbias 0.0489375
R21905 Vbias.n132 Vbias 0.0489375
R21906 Vbias.n70 Vbias 0.0489375
R21907 Vbias.n27 Vbias 0.0489375
R21908 Vbias.n24 Vbias 0.0489375
R21909 Vbias.n410 Vbias 0.0489375
R21910 Vbias.n373 Vbias 0.0489375
R21911 Vbias.n301 Vbias 0.0489375
R21912 Vbias.n299 Vbias 0.0489375
R21913 Vbias.n547 Vbias 0.0489375
R21914 Vbias.n248 Vbias 0.0489375
R21915 Vbias.n246 Vbias 0.0489375
R21916 Vbias.n227 Vbias 0.0489375
R21917 Vbias.n180 Vbias 0.0489375
R21918 Vbias.n182 Vbias 0.0489375
R21919 Vbias.n819 Vbias 0.0489375
R21920 Vbias.n135 Vbias 0.0489375
R21921 Vbias.n133 Vbias 0.0489375
R21922 Vbias.n67 Vbias 0.0489375
R21923 Vbias.n26 Vbias 0.0489375
R21924 Vbias.n23 Vbias 0.0489375
R21925 Vbias.n407 Vbias 0.0489375
R21926 Vbias.n376 Vbias 0.0489375
R21927 Vbias.n296 Vbias 0.0489375
R21928 Vbias.n298 Vbias 0.0489375
R21929 Vbias.n544 Vbias 0.0489375
R21930 Vbias.n243 Vbias 0.0489375
R21931 Vbias.n245 Vbias 0.0489375
R21932 Vbias.n230 Vbias 0.0489375
R21933 Vbias.n185 Vbias 0.0489375
R21934 Vbias.n183 Vbias 0.0489375
R21935 Vbias.n822 Vbias 0.0489375
R21936 Vbias.n136 Vbias 0.0489375
R21937 Vbias.n138 Vbias 0.0489375
R21938 Vbias.n64 Vbias 0.0489375
R21939 Vbias.n21 Vbias 0.0489375
R21940 Vbias.n16 Vbias 0.0489375
R21941 Vbias.n404 Vbias 0.0489375
R21942 Vbias.n379 Vbias 0.0489375
R21943 Vbias.n295 Vbias 0.0489375
R21944 Vbias.n293 Vbias 0.0489375
R21945 Vbias.n541 Vbias 0.0489375
R21946 Vbias.n242 Vbias 0.0489375
R21947 Vbias.n240 Vbias 0.0489375
R21948 Vbias.n233 Vbias 0.0489375
R21949 Vbias.n186 Vbias 0.0489375
R21950 Vbias.n188 Vbias 0.0489375
R21951 Vbias.n825 Vbias 0.0489375
R21952 Vbias.n141 Vbias 0.0489375
R21953 Vbias.n139 Vbias 0.0489375
R21954 Vbias.n61 Vbias 0.0489375
R21955 Vbias.n18 Vbias 0.0489375
R21956 Vbias.n15 Vbias 0.0489375
R21957 Vbias.n338 Vbias 0.0489375
R21958 Vbias.n339 Vbias 0.0489375
R21959 Vbias.n341 Vbias 0.0489375
R21960 Vbias.n525 Vbias 0.0489375
R21961 Vbias.n285 Vbias 0.0489375
R21962 Vbias.n287 Vbias 0.0489375
R21963 Vbias.n662 Vbias 0.0489375
R21964 Vbias.n236 Vbias 0.0489375
R21965 Vbias.n238 Vbias 0.0489375
R21966 Vbias.n703 Vbias 0.0489375
R21967 Vbias.n144 Vbias 0.0489375
R21968 Vbias.n142 Vbias 0.0489375
R21969 Vbias.n671 Vbias 0.0489375
R21970 Vbias.n11 Vbias 0.0489375
R21971 Vbias.n13 Vbias 0.0489375
R21972 Vbias.n6 Vbias 0.0489375
R21973 Vbias.n7 Vbias 0.0489375
R21974 Vbias.n60 Vbias 0.0489375
R21975 Vbias.n674 Vbias 0.0489375
R21976 Vbias.n906 Vbias 0.0489375
R21977 Vbias.n683 Vbias 0.0489375
R21978 Vbias.n146 Vbias 0.0489375
R21979 Vbias.n191 Vbias 0.0489375
R21980 Vbias.n195 Vbias 0.0489375
R21981 Vbias.n665 Vbias 0.0489375
R21982 Vbias.n279 Vbias 0.0489375
R21983 Vbias.n289 Vbias 0.0489375
R21984 Vbias.n329 Vbias 0.0489375
R21985 Vbias.n395 Vbias 0.0489375
R21986 Vbias.n335 Vbias 0.0489375
R21987 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R21988 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R21989 XThC.Tn[1].n71 XThC.Tn[1].n69 161.365
R21990 XThC.Tn[1].n67 XThC.Tn[1].n65 161.365
R21991 XThC.Tn[1].n63 XThC.Tn[1].n61 161.365
R21992 XThC.Tn[1].n59 XThC.Tn[1].n57 161.365
R21993 XThC.Tn[1].n55 XThC.Tn[1].n53 161.365
R21994 XThC.Tn[1].n51 XThC.Tn[1].n49 161.365
R21995 XThC.Tn[1].n47 XThC.Tn[1].n45 161.365
R21996 XThC.Tn[1].n43 XThC.Tn[1].n41 161.365
R21997 XThC.Tn[1].n39 XThC.Tn[1].n37 161.365
R21998 XThC.Tn[1].n35 XThC.Tn[1].n33 161.365
R21999 XThC.Tn[1].n31 XThC.Tn[1].n29 161.365
R22000 XThC.Tn[1].n27 XThC.Tn[1].n25 161.365
R22001 XThC.Tn[1].n23 XThC.Tn[1].n21 161.365
R22002 XThC.Tn[1].n19 XThC.Tn[1].n17 161.365
R22003 XThC.Tn[1].n15 XThC.Tn[1].n13 161.365
R22004 XThC.Tn[1].n12 XThC.Tn[1].n10 161.365
R22005 XThC.Tn[1].n69 XThC.Tn[1].t35 161.202
R22006 XThC.Tn[1].n65 XThC.Tn[1].t25 161.202
R22007 XThC.Tn[1].n61 XThC.Tn[1].t12 161.202
R22008 XThC.Tn[1].n57 XThC.Tn[1].t41 161.202
R22009 XThC.Tn[1].n53 XThC.Tn[1].t33 161.202
R22010 XThC.Tn[1].n49 XThC.Tn[1].t20 161.202
R22011 XThC.Tn[1].n45 XThC.Tn[1].t19 161.202
R22012 XThC.Tn[1].n41 XThC.Tn[1].t32 161.202
R22013 XThC.Tn[1].n37 XThC.Tn[1].t30 161.202
R22014 XThC.Tn[1].n33 XThC.Tn[1].t21 161.202
R22015 XThC.Tn[1].n29 XThC.Tn[1].t40 161.202
R22016 XThC.Tn[1].n25 XThC.Tn[1].t39 161.202
R22017 XThC.Tn[1].n21 XThC.Tn[1].t18 161.202
R22018 XThC.Tn[1].n17 XThC.Tn[1].t16 161.202
R22019 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R22020 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R22021 XThC.Tn[1].n69 XThC.Tn[1].t38 145.137
R22022 XThC.Tn[1].n65 XThC.Tn[1].t28 145.137
R22023 XThC.Tn[1].n61 XThC.Tn[1].t15 145.137
R22024 XThC.Tn[1].n57 XThC.Tn[1].t13 145.137
R22025 XThC.Tn[1].n53 XThC.Tn[1].t37 145.137
R22026 XThC.Tn[1].n49 XThC.Tn[1].t26 145.137
R22027 XThC.Tn[1].n45 XThC.Tn[1].t24 145.137
R22028 XThC.Tn[1].n41 XThC.Tn[1].t36 145.137
R22029 XThC.Tn[1].n37 XThC.Tn[1].t34 145.137
R22030 XThC.Tn[1].n33 XThC.Tn[1].t27 145.137
R22031 XThC.Tn[1].n29 XThC.Tn[1].t43 145.137
R22032 XThC.Tn[1].n25 XThC.Tn[1].t42 145.137
R22033 XThC.Tn[1].n21 XThC.Tn[1].t23 145.137
R22034 XThC.Tn[1].n17 XThC.Tn[1].t22 145.137
R22035 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R22036 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R22037 XThC.Tn[1].n5 XThC.Tn[1].n3 135.249
R22038 XThC.Tn[1].n5 XThC.Tn[1].n4 98.981
R22039 XThC.Tn[1].n7 XThC.Tn[1].n6 98.981
R22040 XThC.Tn[1].n9 XThC.Tn[1].n8 98.981
R22041 XThC.Tn[1].n7 XThC.Tn[1].n5 36.2672
R22042 XThC.Tn[1].n9 XThC.Tn[1].n7 36.2672
R22043 XThC.Tn[1].n74 XThC.Tn[1].n9 32.6405
R22044 XThC.Tn[1].n1 XThC.Tn[1].t1 26.5955
R22045 XThC.Tn[1].n1 XThC.Tn[1].t0 26.5955
R22046 XThC.Tn[1].n0 XThC.Tn[1].t3 26.5955
R22047 XThC.Tn[1].n0 XThC.Tn[1].t2 26.5955
R22048 XThC.Tn[1].n3 XThC.Tn[1].t11 24.9236
R22049 XThC.Tn[1].n3 XThC.Tn[1].t10 24.9236
R22050 XThC.Tn[1].n4 XThC.Tn[1].t9 24.9236
R22051 XThC.Tn[1].n4 XThC.Tn[1].t8 24.9236
R22052 XThC.Tn[1].n6 XThC.Tn[1].t7 24.9236
R22053 XThC.Tn[1].n6 XThC.Tn[1].t6 24.9236
R22054 XThC.Tn[1].n8 XThC.Tn[1].t5 24.9236
R22055 XThC.Tn[1].n8 XThC.Tn[1].t4 24.9236
R22056 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R22057 XThC.Tn[1] XThC.Tn[1].n12 8.0245
R22058 XThC.Tn[1].n72 XThC.Tn[1].n71 7.9105
R22059 XThC.Tn[1].n68 XThC.Tn[1].n67 7.9105
R22060 XThC.Tn[1].n64 XThC.Tn[1].n63 7.9105
R22061 XThC.Tn[1].n60 XThC.Tn[1].n59 7.9105
R22062 XThC.Tn[1].n56 XThC.Tn[1].n55 7.9105
R22063 XThC.Tn[1].n52 XThC.Tn[1].n51 7.9105
R22064 XThC.Tn[1].n48 XThC.Tn[1].n47 7.9105
R22065 XThC.Tn[1].n44 XThC.Tn[1].n43 7.9105
R22066 XThC.Tn[1].n40 XThC.Tn[1].n39 7.9105
R22067 XThC.Tn[1].n36 XThC.Tn[1].n35 7.9105
R22068 XThC.Tn[1].n32 XThC.Tn[1].n31 7.9105
R22069 XThC.Tn[1].n28 XThC.Tn[1].n27 7.9105
R22070 XThC.Tn[1].n24 XThC.Tn[1].n23 7.9105
R22071 XThC.Tn[1].n20 XThC.Tn[1].n19 7.9105
R22072 XThC.Tn[1].n16 XThC.Tn[1].n15 7.9105
R22073 XThC.Tn[1] XThC.Tn[1].n74 6.7205
R22074 XThC.Tn[1].n73 XThC.Tn[1] 6.08068
R22075 XThC.Tn[1].n74 XThC.Tn[1].n73 4.65249
R22076 XThC.Tn[1].n73 XThC.Tn[1] 1.8942
R22077 XThC.Tn[1].n16 XThC.Tn[1] 0.235138
R22078 XThC.Tn[1].n20 XThC.Tn[1] 0.235138
R22079 XThC.Tn[1].n24 XThC.Tn[1] 0.235138
R22080 XThC.Tn[1].n28 XThC.Tn[1] 0.235138
R22081 XThC.Tn[1].n32 XThC.Tn[1] 0.235138
R22082 XThC.Tn[1].n36 XThC.Tn[1] 0.235138
R22083 XThC.Tn[1].n40 XThC.Tn[1] 0.235138
R22084 XThC.Tn[1].n44 XThC.Tn[1] 0.235138
R22085 XThC.Tn[1].n48 XThC.Tn[1] 0.235138
R22086 XThC.Tn[1].n52 XThC.Tn[1] 0.235138
R22087 XThC.Tn[1].n56 XThC.Tn[1] 0.235138
R22088 XThC.Tn[1].n60 XThC.Tn[1] 0.235138
R22089 XThC.Tn[1].n64 XThC.Tn[1] 0.235138
R22090 XThC.Tn[1].n68 XThC.Tn[1] 0.235138
R22091 XThC.Tn[1].n72 XThC.Tn[1] 0.235138
R22092 XThC.Tn[1] XThC.Tn[1].n16 0.114505
R22093 XThC.Tn[1] XThC.Tn[1].n20 0.114505
R22094 XThC.Tn[1] XThC.Tn[1].n24 0.114505
R22095 XThC.Tn[1] XThC.Tn[1].n28 0.114505
R22096 XThC.Tn[1] XThC.Tn[1].n32 0.114505
R22097 XThC.Tn[1] XThC.Tn[1].n36 0.114505
R22098 XThC.Tn[1] XThC.Tn[1].n40 0.114505
R22099 XThC.Tn[1] XThC.Tn[1].n44 0.114505
R22100 XThC.Tn[1] XThC.Tn[1].n48 0.114505
R22101 XThC.Tn[1] XThC.Tn[1].n52 0.114505
R22102 XThC.Tn[1] XThC.Tn[1].n56 0.114505
R22103 XThC.Tn[1] XThC.Tn[1].n60 0.114505
R22104 XThC.Tn[1] XThC.Tn[1].n64 0.114505
R22105 XThC.Tn[1] XThC.Tn[1].n68 0.114505
R22106 XThC.Tn[1] XThC.Tn[1].n72 0.114505
R22107 XThC.Tn[1].n71 XThC.Tn[1].n70 0.0599512
R22108 XThC.Tn[1].n67 XThC.Tn[1].n66 0.0599512
R22109 XThC.Tn[1].n63 XThC.Tn[1].n62 0.0599512
R22110 XThC.Tn[1].n59 XThC.Tn[1].n58 0.0599512
R22111 XThC.Tn[1].n55 XThC.Tn[1].n54 0.0599512
R22112 XThC.Tn[1].n51 XThC.Tn[1].n50 0.0599512
R22113 XThC.Tn[1].n47 XThC.Tn[1].n46 0.0599512
R22114 XThC.Tn[1].n43 XThC.Tn[1].n42 0.0599512
R22115 XThC.Tn[1].n39 XThC.Tn[1].n38 0.0599512
R22116 XThC.Tn[1].n35 XThC.Tn[1].n34 0.0599512
R22117 XThC.Tn[1].n31 XThC.Tn[1].n30 0.0599512
R22118 XThC.Tn[1].n27 XThC.Tn[1].n26 0.0599512
R22119 XThC.Tn[1].n23 XThC.Tn[1].n22 0.0599512
R22120 XThC.Tn[1].n19 XThC.Tn[1].n18 0.0599512
R22121 XThC.Tn[1].n15 XThC.Tn[1].n14 0.0599512
R22122 XThC.Tn[1].n12 XThC.Tn[1].n11 0.0599512
R22123 XThC.Tn[1].n70 XThC.Tn[1] 0.0469286
R22124 XThC.Tn[1].n66 XThC.Tn[1] 0.0469286
R22125 XThC.Tn[1].n62 XThC.Tn[1] 0.0469286
R22126 XThC.Tn[1].n58 XThC.Tn[1] 0.0469286
R22127 XThC.Tn[1].n54 XThC.Tn[1] 0.0469286
R22128 XThC.Tn[1].n50 XThC.Tn[1] 0.0469286
R22129 XThC.Tn[1].n46 XThC.Tn[1] 0.0469286
R22130 XThC.Tn[1].n42 XThC.Tn[1] 0.0469286
R22131 XThC.Tn[1].n38 XThC.Tn[1] 0.0469286
R22132 XThC.Tn[1].n34 XThC.Tn[1] 0.0469286
R22133 XThC.Tn[1].n30 XThC.Tn[1] 0.0469286
R22134 XThC.Tn[1].n26 XThC.Tn[1] 0.0469286
R22135 XThC.Tn[1].n22 XThC.Tn[1] 0.0469286
R22136 XThC.Tn[1].n18 XThC.Tn[1] 0.0469286
R22137 XThC.Tn[1].n14 XThC.Tn[1] 0.0469286
R22138 XThC.Tn[1].n11 XThC.Tn[1] 0.0469286
R22139 XThC.Tn[1].n70 XThC.Tn[1] 0.0401341
R22140 XThC.Tn[1].n66 XThC.Tn[1] 0.0401341
R22141 XThC.Tn[1].n62 XThC.Tn[1] 0.0401341
R22142 XThC.Tn[1].n58 XThC.Tn[1] 0.0401341
R22143 XThC.Tn[1].n54 XThC.Tn[1] 0.0401341
R22144 XThC.Tn[1].n50 XThC.Tn[1] 0.0401341
R22145 XThC.Tn[1].n46 XThC.Tn[1] 0.0401341
R22146 XThC.Tn[1].n42 XThC.Tn[1] 0.0401341
R22147 XThC.Tn[1].n38 XThC.Tn[1] 0.0401341
R22148 XThC.Tn[1].n34 XThC.Tn[1] 0.0401341
R22149 XThC.Tn[1].n30 XThC.Tn[1] 0.0401341
R22150 XThC.Tn[1].n26 XThC.Tn[1] 0.0401341
R22151 XThC.Tn[1].n22 XThC.Tn[1] 0.0401341
R22152 XThC.Tn[1].n18 XThC.Tn[1] 0.0401341
R22153 XThC.Tn[1].n14 XThC.Tn[1] 0.0401341
R22154 XThC.Tn[1].n11 XThC.Tn[1] 0.0401341
R22155 XThC.Tn[3].n2 XThC.Tn[3].n1 332.334
R22156 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R22157 XThC.Tn[3].n71 XThC.Tn[3].n69 161.365
R22158 XThC.Tn[3].n67 XThC.Tn[3].n65 161.365
R22159 XThC.Tn[3].n63 XThC.Tn[3].n61 161.365
R22160 XThC.Tn[3].n59 XThC.Tn[3].n57 161.365
R22161 XThC.Tn[3].n55 XThC.Tn[3].n53 161.365
R22162 XThC.Tn[3].n51 XThC.Tn[3].n49 161.365
R22163 XThC.Tn[3].n47 XThC.Tn[3].n45 161.365
R22164 XThC.Tn[3].n43 XThC.Tn[3].n41 161.365
R22165 XThC.Tn[3].n39 XThC.Tn[3].n37 161.365
R22166 XThC.Tn[3].n35 XThC.Tn[3].n33 161.365
R22167 XThC.Tn[3].n31 XThC.Tn[3].n29 161.365
R22168 XThC.Tn[3].n27 XThC.Tn[3].n25 161.365
R22169 XThC.Tn[3].n23 XThC.Tn[3].n21 161.365
R22170 XThC.Tn[3].n19 XThC.Tn[3].n17 161.365
R22171 XThC.Tn[3].n15 XThC.Tn[3].n13 161.365
R22172 XThC.Tn[3].n12 XThC.Tn[3].n10 161.365
R22173 XThC.Tn[3].n69 XThC.Tn[3].t16 161.202
R22174 XThC.Tn[3].n65 XThC.Tn[3].t38 161.202
R22175 XThC.Tn[3].n61 XThC.Tn[3].t25 161.202
R22176 XThC.Tn[3].n57 XThC.Tn[3].t22 161.202
R22177 XThC.Tn[3].n53 XThC.Tn[3].t14 161.202
R22178 XThC.Tn[3].n49 XThC.Tn[3].t33 161.202
R22179 XThC.Tn[3].n45 XThC.Tn[3].t32 161.202
R22180 XThC.Tn[3].n41 XThC.Tn[3].t13 161.202
R22181 XThC.Tn[3].n37 XThC.Tn[3].t43 161.202
R22182 XThC.Tn[3].n33 XThC.Tn[3].t34 161.202
R22183 XThC.Tn[3].n29 XThC.Tn[3].t21 161.202
R22184 XThC.Tn[3].n25 XThC.Tn[3].t20 161.202
R22185 XThC.Tn[3].n21 XThC.Tn[3].t31 161.202
R22186 XThC.Tn[3].n17 XThC.Tn[3].t29 161.202
R22187 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R22188 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R22189 XThC.Tn[3].n69 XThC.Tn[3].t19 145.137
R22190 XThC.Tn[3].n65 XThC.Tn[3].t41 145.137
R22191 XThC.Tn[3].n61 XThC.Tn[3].t28 145.137
R22192 XThC.Tn[3].n57 XThC.Tn[3].t26 145.137
R22193 XThC.Tn[3].n53 XThC.Tn[3].t18 145.137
R22194 XThC.Tn[3].n49 XThC.Tn[3].t39 145.137
R22195 XThC.Tn[3].n45 XThC.Tn[3].t37 145.137
R22196 XThC.Tn[3].n41 XThC.Tn[3].t17 145.137
R22197 XThC.Tn[3].n37 XThC.Tn[3].t15 145.137
R22198 XThC.Tn[3].n33 XThC.Tn[3].t40 145.137
R22199 XThC.Tn[3].n29 XThC.Tn[3].t24 145.137
R22200 XThC.Tn[3].n25 XThC.Tn[3].t23 145.137
R22201 XThC.Tn[3].n21 XThC.Tn[3].t36 145.137
R22202 XThC.Tn[3].n17 XThC.Tn[3].t35 145.137
R22203 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R22204 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R22205 XThC.Tn[3].n5 XThC.Tn[3].n3 135.249
R22206 XThC.Tn[3].n5 XThC.Tn[3].n4 98.981
R22207 XThC.Tn[3].n7 XThC.Tn[3].n6 98.981
R22208 XThC.Tn[3].n9 XThC.Tn[3].n8 98.981
R22209 XThC.Tn[3].n7 XThC.Tn[3].n5 36.2672
R22210 XThC.Tn[3].n9 XThC.Tn[3].n7 36.2672
R22211 XThC.Tn[3].n74 XThC.Tn[3].n9 32.6405
R22212 XThC.Tn[3].n0 XThC.Tn[3].t1 26.5955
R22213 XThC.Tn[3].n0 XThC.Tn[3].t0 26.5955
R22214 XThC.Tn[3].n1 XThC.Tn[3].t3 26.5955
R22215 XThC.Tn[3].n1 XThC.Tn[3].t2 26.5955
R22216 XThC.Tn[3].n3 XThC.Tn[3].t11 24.9236
R22217 XThC.Tn[3].n3 XThC.Tn[3].t10 24.9236
R22218 XThC.Tn[3].n4 XThC.Tn[3].t9 24.9236
R22219 XThC.Tn[3].n4 XThC.Tn[3].t8 24.9236
R22220 XThC.Tn[3].n6 XThC.Tn[3].t7 24.9236
R22221 XThC.Tn[3].n6 XThC.Tn[3].t6 24.9236
R22222 XThC.Tn[3].n8 XThC.Tn[3].t5 24.9236
R22223 XThC.Tn[3].n8 XThC.Tn[3].t4 24.9236
R22224 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R22225 XThC.Tn[3] XThC.Tn[3].n12 8.0245
R22226 XThC.Tn[3].n72 XThC.Tn[3].n71 7.9105
R22227 XThC.Tn[3].n68 XThC.Tn[3].n67 7.9105
R22228 XThC.Tn[3].n64 XThC.Tn[3].n63 7.9105
R22229 XThC.Tn[3].n60 XThC.Tn[3].n59 7.9105
R22230 XThC.Tn[3].n56 XThC.Tn[3].n55 7.9105
R22231 XThC.Tn[3].n52 XThC.Tn[3].n51 7.9105
R22232 XThC.Tn[3].n48 XThC.Tn[3].n47 7.9105
R22233 XThC.Tn[3].n44 XThC.Tn[3].n43 7.9105
R22234 XThC.Tn[3].n40 XThC.Tn[3].n39 7.9105
R22235 XThC.Tn[3].n36 XThC.Tn[3].n35 7.9105
R22236 XThC.Tn[3].n32 XThC.Tn[3].n31 7.9105
R22237 XThC.Tn[3].n28 XThC.Tn[3].n27 7.9105
R22238 XThC.Tn[3].n24 XThC.Tn[3].n23 7.9105
R22239 XThC.Tn[3].n20 XThC.Tn[3].n19 7.9105
R22240 XThC.Tn[3].n16 XThC.Tn[3].n15 7.9105
R22241 XThC.Tn[3].n73 XThC.Tn[3] 7.48718
R22242 XThC.Tn[3] XThC.Tn[3].n74 6.7205
R22243 XThC.Tn[3].n74 XThC.Tn[3].n73 5.06464
R22244 XThC.Tn[3].n73 XThC.Tn[3] 1.18175
R22245 XThC.Tn[3].n16 XThC.Tn[3] 0.235138
R22246 XThC.Tn[3].n20 XThC.Tn[3] 0.235138
R22247 XThC.Tn[3].n24 XThC.Tn[3] 0.235138
R22248 XThC.Tn[3].n28 XThC.Tn[3] 0.235138
R22249 XThC.Tn[3].n32 XThC.Tn[3] 0.235138
R22250 XThC.Tn[3].n36 XThC.Tn[3] 0.235138
R22251 XThC.Tn[3].n40 XThC.Tn[3] 0.235138
R22252 XThC.Tn[3].n44 XThC.Tn[3] 0.235138
R22253 XThC.Tn[3].n48 XThC.Tn[3] 0.235138
R22254 XThC.Tn[3].n52 XThC.Tn[3] 0.235138
R22255 XThC.Tn[3].n56 XThC.Tn[3] 0.235138
R22256 XThC.Tn[3].n60 XThC.Tn[3] 0.235138
R22257 XThC.Tn[3].n64 XThC.Tn[3] 0.235138
R22258 XThC.Tn[3].n68 XThC.Tn[3] 0.235138
R22259 XThC.Tn[3].n72 XThC.Tn[3] 0.235138
R22260 XThC.Tn[3] XThC.Tn[3].n16 0.114505
R22261 XThC.Tn[3] XThC.Tn[3].n20 0.114505
R22262 XThC.Tn[3] XThC.Tn[3].n24 0.114505
R22263 XThC.Tn[3] XThC.Tn[3].n28 0.114505
R22264 XThC.Tn[3] XThC.Tn[3].n32 0.114505
R22265 XThC.Tn[3] XThC.Tn[3].n36 0.114505
R22266 XThC.Tn[3] XThC.Tn[3].n40 0.114505
R22267 XThC.Tn[3] XThC.Tn[3].n44 0.114505
R22268 XThC.Tn[3] XThC.Tn[3].n48 0.114505
R22269 XThC.Tn[3] XThC.Tn[3].n52 0.114505
R22270 XThC.Tn[3] XThC.Tn[3].n56 0.114505
R22271 XThC.Tn[3] XThC.Tn[3].n60 0.114505
R22272 XThC.Tn[3] XThC.Tn[3].n64 0.114505
R22273 XThC.Tn[3] XThC.Tn[3].n68 0.114505
R22274 XThC.Tn[3] XThC.Tn[3].n72 0.114505
R22275 XThC.Tn[3].n71 XThC.Tn[3].n70 0.0599512
R22276 XThC.Tn[3].n67 XThC.Tn[3].n66 0.0599512
R22277 XThC.Tn[3].n63 XThC.Tn[3].n62 0.0599512
R22278 XThC.Tn[3].n59 XThC.Tn[3].n58 0.0599512
R22279 XThC.Tn[3].n55 XThC.Tn[3].n54 0.0599512
R22280 XThC.Tn[3].n51 XThC.Tn[3].n50 0.0599512
R22281 XThC.Tn[3].n47 XThC.Tn[3].n46 0.0599512
R22282 XThC.Tn[3].n43 XThC.Tn[3].n42 0.0599512
R22283 XThC.Tn[3].n39 XThC.Tn[3].n38 0.0599512
R22284 XThC.Tn[3].n35 XThC.Tn[3].n34 0.0599512
R22285 XThC.Tn[3].n31 XThC.Tn[3].n30 0.0599512
R22286 XThC.Tn[3].n27 XThC.Tn[3].n26 0.0599512
R22287 XThC.Tn[3].n23 XThC.Tn[3].n22 0.0599512
R22288 XThC.Tn[3].n19 XThC.Tn[3].n18 0.0599512
R22289 XThC.Tn[3].n15 XThC.Tn[3].n14 0.0599512
R22290 XThC.Tn[3].n12 XThC.Tn[3].n11 0.0599512
R22291 XThC.Tn[3].n70 XThC.Tn[3] 0.0469286
R22292 XThC.Tn[3].n66 XThC.Tn[3] 0.0469286
R22293 XThC.Tn[3].n62 XThC.Tn[3] 0.0469286
R22294 XThC.Tn[3].n58 XThC.Tn[3] 0.0469286
R22295 XThC.Tn[3].n54 XThC.Tn[3] 0.0469286
R22296 XThC.Tn[3].n50 XThC.Tn[3] 0.0469286
R22297 XThC.Tn[3].n46 XThC.Tn[3] 0.0469286
R22298 XThC.Tn[3].n42 XThC.Tn[3] 0.0469286
R22299 XThC.Tn[3].n38 XThC.Tn[3] 0.0469286
R22300 XThC.Tn[3].n34 XThC.Tn[3] 0.0469286
R22301 XThC.Tn[3].n30 XThC.Tn[3] 0.0469286
R22302 XThC.Tn[3].n26 XThC.Tn[3] 0.0469286
R22303 XThC.Tn[3].n22 XThC.Tn[3] 0.0469286
R22304 XThC.Tn[3].n18 XThC.Tn[3] 0.0469286
R22305 XThC.Tn[3].n14 XThC.Tn[3] 0.0469286
R22306 XThC.Tn[3].n11 XThC.Tn[3] 0.0469286
R22307 XThC.Tn[3].n70 XThC.Tn[3] 0.0401341
R22308 XThC.Tn[3].n66 XThC.Tn[3] 0.0401341
R22309 XThC.Tn[3].n62 XThC.Tn[3] 0.0401341
R22310 XThC.Tn[3].n58 XThC.Tn[3] 0.0401341
R22311 XThC.Tn[3].n54 XThC.Tn[3] 0.0401341
R22312 XThC.Tn[3].n50 XThC.Tn[3] 0.0401341
R22313 XThC.Tn[3].n46 XThC.Tn[3] 0.0401341
R22314 XThC.Tn[3].n42 XThC.Tn[3] 0.0401341
R22315 XThC.Tn[3].n38 XThC.Tn[3] 0.0401341
R22316 XThC.Tn[3].n34 XThC.Tn[3] 0.0401341
R22317 XThC.Tn[3].n30 XThC.Tn[3] 0.0401341
R22318 XThC.Tn[3].n26 XThC.Tn[3] 0.0401341
R22319 XThC.Tn[3].n22 XThC.Tn[3] 0.0401341
R22320 XThC.Tn[3].n18 XThC.Tn[3] 0.0401341
R22321 XThC.Tn[3].n14 XThC.Tn[3] 0.0401341
R22322 XThC.Tn[3].n11 XThC.Tn[3] 0.0401341
R22323 XThR.Tn[10].n87 XThR.Tn[10].n86 256.103
R22324 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R22325 XThR.Tn[10].n5 XThR.Tn[10].n3 241.847
R22326 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R22327 XThR.Tn[10].n87 XThR.Tn[10].n85 202.094
R22328 XThR.Tn[10].n5 XThR.Tn[10].n4 185
R22329 XThR.Tn[10] XThR.Tn[10].n78 161.363
R22330 XThR.Tn[10] XThR.Tn[10].n73 161.363
R22331 XThR.Tn[10] XThR.Tn[10].n68 161.363
R22332 XThR.Tn[10] XThR.Tn[10].n63 161.363
R22333 XThR.Tn[10] XThR.Tn[10].n58 161.363
R22334 XThR.Tn[10] XThR.Tn[10].n53 161.363
R22335 XThR.Tn[10] XThR.Tn[10].n48 161.363
R22336 XThR.Tn[10] XThR.Tn[10].n43 161.363
R22337 XThR.Tn[10] XThR.Tn[10].n38 161.363
R22338 XThR.Tn[10] XThR.Tn[10].n33 161.363
R22339 XThR.Tn[10] XThR.Tn[10].n28 161.363
R22340 XThR.Tn[10] XThR.Tn[10].n23 161.363
R22341 XThR.Tn[10] XThR.Tn[10].n18 161.363
R22342 XThR.Tn[10] XThR.Tn[10].n13 161.363
R22343 XThR.Tn[10] XThR.Tn[10].n8 161.363
R22344 XThR.Tn[10] XThR.Tn[10].n6 161.363
R22345 XThR.Tn[10].n80 XThR.Tn[10].n79 161.3
R22346 XThR.Tn[10].n75 XThR.Tn[10].n74 161.3
R22347 XThR.Tn[10].n70 XThR.Tn[10].n69 161.3
R22348 XThR.Tn[10].n65 XThR.Tn[10].n64 161.3
R22349 XThR.Tn[10].n60 XThR.Tn[10].n59 161.3
R22350 XThR.Tn[10].n55 XThR.Tn[10].n54 161.3
R22351 XThR.Tn[10].n50 XThR.Tn[10].n49 161.3
R22352 XThR.Tn[10].n45 XThR.Tn[10].n44 161.3
R22353 XThR.Tn[10].n40 XThR.Tn[10].n39 161.3
R22354 XThR.Tn[10].n35 XThR.Tn[10].n34 161.3
R22355 XThR.Tn[10].n30 XThR.Tn[10].n29 161.3
R22356 XThR.Tn[10].n25 XThR.Tn[10].n24 161.3
R22357 XThR.Tn[10].n20 XThR.Tn[10].n19 161.3
R22358 XThR.Tn[10].n15 XThR.Tn[10].n14 161.3
R22359 XThR.Tn[10].n10 XThR.Tn[10].n9 161.3
R22360 XThR.Tn[10].n78 XThR.Tn[10].t37 161.106
R22361 XThR.Tn[10].n73 XThR.Tn[10].t45 161.106
R22362 XThR.Tn[10].n68 XThR.Tn[10].t27 161.106
R22363 XThR.Tn[10].n63 XThR.Tn[10].t72 161.106
R22364 XThR.Tn[10].n58 XThR.Tn[10].t35 161.106
R22365 XThR.Tn[10].n53 XThR.Tn[10].t61 161.106
R22366 XThR.Tn[10].n48 XThR.Tn[10].t43 161.106
R22367 XThR.Tn[10].n43 XThR.Tn[10].t24 161.106
R22368 XThR.Tn[10].n38 XThR.Tn[10].t69 161.106
R22369 XThR.Tn[10].n33 XThR.Tn[10].t15 161.106
R22370 XThR.Tn[10].n28 XThR.Tn[10].t59 161.106
R22371 XThR.Tn[10].n23 XThR.Tn[10].t26 161.106
R22372 XThR.Tn[10].n18 XThR.Tn[10].t58 161.106
R22373 XThR.Tn[10].n13 XThR.Tn[10].t41 161.106
R22374 XThR.Tn[10].n8 XThR.Tn[10].t63 161.106
R22375 XThR.Tn[10].n6 XThR.Tn[10].t47 161.106
R22376 XThR.Tn[10].n79 XThR.Tn[10].t34 159.978
R22377 XThR.Tn[10].n74 XThR.Tn[10].t39 159.978
R22378 XThR.Tn[10].n69 XThR.Tn[10].t22 159.978
R22379 XThR.Tn[10].n64 XThR.Tn[10].t68 159.978
R22380 XThR.Tn[10].n59 XThR.Tn[10].t32 159.978
R22381 XThR.Tn[10].n54 XThR.Tn[10].t57 159.978
R22382 XThR.Tn[10].n49 XThR.Tn[10].t38 159.978
R22383 XThR.Tn[10].n44 XThR.Tn[10].t20 159.978
R22384 XThR.Tn[10].n39 XThR.Tn[10].t66 159.978
R22385 XThR.Tn[10].n34 XThR.Tn[10].t12 159.978
R22386 XThR.Tn[10].n29 XThR.Tn[10].t56 159.978
R22387 XThR.Tn[10].n24 XThR.Tn[10].t21 159.978
R22388 XThR.Tn[10].n19 XThR.Tn[10].t55 159.978
R22389 XThR.Tn[10].n14 XThR.Tn[10].t36 159.978
R22390 XThR.Tn[10].n9 XThR.Tn[10].t60 159.978
R22391 XThR.Tn[10].n78 XThR.Tn[10].t29 145.038
R22392 XThR.Tn[10].n73 XThR.Tn[10].t49 145.038
R22393 XThR.Tn[10].n68 XThR.Tn[10].t31 145.038
R22394 XThR.Tn[10].n63 XThR.Tn[10].t16 145.038
R22395 XThR.Tn[10].n58 XThR.Tn[10].t46 145.038
R22396 XThR.Tn[10].n53 XThR.Tn[10].t28 145.038
R22397 XThR.Tn[10].n48 XThR.Tn[10].t33 145.038
R22398 XThR.Tn[10].n43 XThR.Tn[10].t17 145.038
R22399 XThR.Tn[10].n38 XThR.Tn[10].t14 145.038
R22400 XThR.Tn[10].n33 XThR.Tn[10].t44 145.038
R22401 XThR.Tn[10].n28 XThR.Tn[10].t67 145.038
R22402 XThR.Tn[10].n23 XThR.Tn[10].t30 145.038
R22403 XThR.Tn[10].n18 XThR.Tn[10].t65 145.038
R22404 XThR.Tn[10].n13 XThR.Tn[10].t48 145.038
R22405 XThR.Tn[10].n8 XThR.Tn[10].t13 145.038
R22406 XThR.Tn[10].n6 XThR.Tn[10].t54 145.038
R22407 XThR.Tn[10].n79 XThR.Tn[10].t64 143.911
R22408 XThR.Tn[10].n74 XThR.Tn[10].t25 143.911
R22409 XThR.Tn[10].n69 XThR.Tn[10].t71 143.911
R22410 XThR.Tn[10].n64 XThR.Tn[10].t52 143.911
R22411 XThR.Tn[10].n59 XThR.Tn[10].t19 143.911
R22412 XThR.Tn[10].n54 XThR.Tn[10].t62 143.911
R22413 XThR.Tn[10].n49 XThR.Tn[10].t73 143.911
R22414 XThR.Tn[10].n44 XThR.Tn[10].t53 143.911
R22415 XThR.Tn[10].n39 XThR.Tn[10].t51 143.911
R22416 XThR.Tn[10].n34 XThR.Tn[10].t18 143.911
R22417 XThR.Tn[10].n29 XThR.Tn[10].t42 143.911
R22418 XThR.Tn[10].n24 XThR.Tn[10].t70 143.911
R22419 XThR.Tn[10].n19 XThR.Tn[10].t40 143.911
R22420 XThR.Tn[10].n14 XThR.Tn[10].t23 143.911
R22421 XThR.Tn[10].n9 XThR.Tn[10].t50 143.911
R22422 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R22423 XThR.Tn[10].n86 XThR.Tn[10].t1 26.5955
R22424 XThR.Tn[10].n86 XThR.Tn[10].t5 26.5955
R22425 XThR.Tn[10].n0 XThR.Tn[10].t9 26.5955
R22426 XThR.Tn[10].n0 XThR.Tn[10].t7 26.5955
R22427 XThR.Tn[10].n1 XThR.Tn[10].t10 26.5955
R22428 XThR.Tn[10].n1 XThR.Tn[10].t8 26.5955
R22429 XThR.Tn[10].n85 XThR.Tn[10].t3 26.5955
R22430 XThR.Tn[10].n85 XThR.Tn[10].t0 26.5955
R22431 XThR.Tn[10].n4 XThR.Tn[10].t4 24.9236
R22432 XThR.Tn[10].n4 XThR.Tn[10].t11 24.9236
R22433 XThR.Tn[10].n3 XThR.Tn[10].t2 24.9236
R22434 XThR.Tn[10].n3 XThR.Tn[10].t6 24.9236
R22435 XThR.Tn[10] XThR.Tn[10].n5 18.8943
R22436 XThR.Tn[10].n88 XThR.Tn[10].n87 13.5534
R22437 XThR.Tn[10].n84 XThR.Tn[10] 7.84567
R22438 XThR.Tn[10].n84 XThR.Tn[10] 6.34069
R22439 XThR.Tn[10] XThR.Tn[10].n7 5.34038
R22440 XThR.Tn[10].n12 XThR.Tn[10].n11 4.5005
R22441 XThR.Tn[10].n17 XThR.Tn[10].n16 4.5005
R22442 XThR.Tn[10].n22 XThR.Tn[10].n21 4.5005
R22443 XThR.Tn[10].n27 XThR.Tn[10].n26 4.5005
R22444 XThR.Tn[10].n32 XThR.Tn[10].n31 4.5005
R22445 XThR.Tn[10].n37 XThR.Tn[10].n36 4.5005
R22446 XThR.Tn[10].n42 XThR.Tn[10].n41 4.5005
R22447 XThR.Tn[10].n47 XThR.Tn[10].n46 4.5005
R22448 XThR.Tn[10].n52 XThR.Tn[10].n51 4.5005
R22449 XThR.Tn[10].n57 XThR.Tn[10].n56 4.5005
R22450 XThR.Tn[10].n62 XThR.Tn[10].n61 4.5005
R22451 XThR.Tn[10].n67 XThR.Tn[10].n66 4.5005
R22452 XThR.Tn[10].n72 XThR.Tn[10].n71 4.5005
R22453 XThR.Tn[10].n77 XThR.Tn[10].n76 4.5005
R22454 XThR.Tn[10].n82 XThR.Tn[10].n81 4.5005
R22455 XThR.Tn[10].n83 XThR.Tn[10] 3.70586
R22456 XThR.Tn[10].n12 XThR.Tn[10] 2.52282
R22457 XThR.Tn[10].n17 XThR.Tn[10] 2.52282
R22458 XThR.Tn[10].n22 XThR.Tn[10] 2.52282
R22459 XThR.Tn[10].n27 XThR.Tn[10] 2.52282
R22460 XThR.Tn[10].n32 XThR.Tn[10] 2.52282
R22461 XThR.Tn[10].n37 XThR.Tn[10] 2.52282
R22462 XThR.Tn[10].n42 XThR.Tn[10] 2.52282
R22463 XThR.Tn[10].n47 XThR.Tn[10] 2.52282
R22464 XThR.Tn[10].n52 XThR.Tn[10] 2.52282
R22465 XThR.Tn[10].n57 XThR.Tn[10] 2.52282
R22466 XThR.Tn[10].n62 XThR.Tn[10] 2.52282
R22467 XThR.Tn[10].n67 XThR.Tn[10] 2.52282
R22468 XThR.Tn[10].n72 XThR.Tn[10] 2.52282
R22469 XThR.Tn[10].n77 XThR.Tn[10] 2.52282
R22470 XThR.Tn[10].n82 XThR.Tn[10] 2.52282
R22471 XThR.Tn[10] XThR.Tn[10].n84 1.79489
R22472 XThR.Tn[10] XThR.Tn[10].n88 1.50638
R22473 XThR.Tn[10].n88 XThR.Tn[10] 1.19676
R22474 XThR.Tn[10].n80 XThR.Tn[10] 1.08677
R22475 XThR.Tn[10].n75 XThR.Tn[10] 1.08677
R22476 XThR.Tn[10].n70 XThR.Tn[10] 1.08677
R22477 XThR.Tn[10].n65 XThR.Tn[10] 1.08677
R22478 XThR.Tn[10].n60 XThR.Tn[10] 1.08677
R22479 XThR.Tn[10].n55 XThR.Tn[10] 1.08677
R22480 XThR.Tn[10].n50 XThR.Tn[10] 1.08677
R22481 XThR.Tn[10].n45 XThR.Tn[10] 1.08677
R22482 XThR.Tn[10].n40 XThR.Tn[10] 1.08677
R22483 XThR.Tn[10].n35 XThR.Tn[10] 1.08677
R22484 XThR.Tn[10].n30 XThR.Tn[10] 1.08677
R22485 XThR.Tn[10].n25 XThR.Tn[10] 1.08677
R22486 XThR.Tn[10].n20 XThR.Tn[10] 1.08677
R22487 XThR.Tn[10].n15 XThR.Tn[10] 1.08677
R22488 XThR.Tn[10].n10 XThR.Tn[10] 1.08677
R22489 XThR.Tn[10] XThR.Tn[10].n12 0.839786
R22490 XThR.Tn[10] XThR.Tn[10].n17 0.839786
R22491 XThR.Tn[10] XThR.Tn[10].n22 0.839786
R22492 XThR.Tn[10] XThR.Tn[10].n27 0.839786
R22493 XThR.Tn[10] XThR.Tn[10].n32 0.839786
R22494 XThR.Tn[10] XThR.Tn[10].n37 0.839786
R22495 XThR.Tn[10] XThR.Tn[10].n42 0.839786
R22496 XThR.Tn[10] XThR.Tn[10].n47 0.839786
R22497 XThR.Tn[10] XThR.Tn[10].n52 0.839786
R22498 XThR.Tn[10] XThR.Tn[10].n57 0.839786
R22499 XThR.Tn[10] XThR.Tn[10].n62 0.839786
R22500 XThR.Tn[10] XThR.Tn[10].n67 0.839786
R22501 XThR.Tn[10] XThR.Tn[10].n72 0.839786
R22502 XThR.Tn[10] XThR.Tn[10].n77 0.839786
R22503 XThR.Tn[10] XThR.Tn[10].n82 0.839786
R22504 XThR.Tn[10].n7 XThR.Tn[10] 0.499542
R22505 XThR.Tn[10].n81 XThR.Tn[10] 0.063
R22506 XThR.Tn[10].n76 XThR.Tn[10] 0.063
R22507 XThR.Tn[10].n71 XThR.Tn[10] 0.063
R22508 XThR.Tn[10].n66 XThR.Tn[10] 0.063
R22509 XThR.Tn[10].n61 XThR.Tn[10] 0.063
R22510 XThR.Tn[10].n56 XThR.Tn[10] 0.063
R22511 XThR.Tn[10].n51 XThR.Tn[10] 0.063
R22512 XThR.Tn[10].n46 XThR.Tn[10] 0.063
R22513 XThR.Tn[10].n41 XThR.Tn[10] 0.063
R22514 XThR.Tn[10].n36 XThR.Tn[10] 0.063
R22515 XThR.Tn[10].n31 XThR.Tn[10] 0.063
R22516 XThR.Tn[10].n26 XThR.Tn[10] 0.063
R22517 XThR.Tn[10].n21 XThR.Tn[10] 0.063
R22518 XThR.Tn[10].n16 XThR.Tn[10] 0.063
R22519 XThR.Tn[10].n11 XThR.Tn[10] 0.063
R22520 XThR.Tn[10].n83 XThR.Tn[10] 0.0540714
R22521 XThR.Tn[10] XThR.Tn[10].n83 0.038
R22522 XThR.Tn[10].n7 XThR.Tn[10] 0.0143889
R22523 XThR.Tn[10].n81 XThR.Tn[10].n80 0.00771154
R22524 XThR.Tn[10].n76 XThR.Tn[10].n75 0.00771154
R22525 XThR.Tn[10].n71 XThR.Tn[10].n70 0.00771154
R22526 XThR.Tn[10].n66 XThR.Tn[10].n65 0.00771154
R22527 XThR.Tn[10].n61 XThR.Tn[10].n60 0.00771154
R22528 XThR.Tn[10].n56 XThR.Tn[10].n55 0.00771154
R22529 XThR.Tn[10].n51 XThR.Tn[10].n50 0.00771154
R22530 XThR.Tn[10].n46 XThR.Tn[10].n45 0.00771154
R22531 XThR.Tn[10].n41 XThR.Tn[10].n40 0.00771154
R22532 XThR.Tn[10].n36 XThR.Tn[10].n35 0.00771154
R22533 XThR.Tn[10].n31 XThR.Tn[10].n30 0.00771154
R22534 XThR.Tn[10].n26 XThR.Tn[10].n25 0.00771154
R22535 XThR.Tn[10].n21 XThR.Tn[10].n20 0.00771154
R22536 XThR.Tn[10].n16 XThR.Tn[10].n15 0.00771154
R22537 XThR.Tn[10].n11 XThR.Tn[10].n10 0.00771154
R22538 XThC.Tn[14].n70 XThC.Tn[14].n69 256.103
R22539 XThC.Tn[14].n74 XThC.Tn[14].n72 243.68
R22540 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22541 XThC.Tn[14].n74 XThC.Tn[14].n73 205.28
R22542 XThC.Tn[14].n70 XThC.Tn[14].n68 202.095
R22543 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22544 XThC.Tn[14].n64 XThC.Tn[14].n62 161.365
R22545 XThC.Tn[14].n60 XThC.Tn[14].n58 161.365
R22546 XThC.Tn[14].n56 XThC.Tn[14].n54 161.365
R22547 XThC.Tn[14].n52 XThC.Tn[14].n50 161.365
R22548 XThC.Tn[14].n48 XThC.Tn[14].n46 161.365
R22549 XThC.Tn[14].n44 XThC.Tn[14].n42 161.365
R22550 XThC.Tn[14].n40 XThC.Tn[14].n38 161.365
R22551 XThC.Tn[14].n36 XThC.Tn[14].n34 161.365
R22552 XThC.Tn[14].n32 XThC.Tn[14].n30 161.365
R22553 XThC.Tn[14].n28 XThC.Tn[14].n26 161.365
R22554 XThC.Tn[14].n24 XThC.Tn[14].n22 161.365
R22555 XThC.Tn[14].n20 XThC.Tn[14].n18 161.365
R22556 XThC.Tn[14].n16 XThC.Tn[14].n14 161.365
R22557 XThC.Tn[14].n12 XThC.Tn[14].n10 161.365
R22558 XThC.Tn[14].n8 XThC.Tn[14].n6 161.365
R22559 XThC.Tn[14].n5 XThC.Tn[14].n3 161.365
R22560 XThC.Tn[14].n62 XThC.Tn[14].t12 161.202
R22561 XThC.Tn[14].n58 XThC.Tn[14].t33 161.202
R22562 XThC.Tn[14].n54 XThC.Tn[14].t21 161.202
R22563 XThC.Tn[14].n50 XThC.Tn[14].t19 161.202
R22564 XThC.Tn[14].n46 XThC.Tn[14].t42 161.202
R22565 XThC.Tn[14].n42 XThC.Tn[14].t30 161.202
R22566 XThC.Tn[14].n38 XThC.Tn[14].t27 161.202
R22567 XThC.Tn[14].n34 XThC.Tn[14].t41 161.202
R22568 XThC.Tn[14].n30 XThC.Tn[14].t39 161.202
R22569 XThC.Tn[14].n26 XThC.Tn[14].t31 161.202
R22570 XThC.Tn[14].n22 XThC.Tn[14].t17 161.202
R22571 XThC.Tn[14].n18 XThC.Tn[14].t14 161.202
R22572 XThC.Tn[14].n14 XThC.Tn[14].t26 161.202
R22573 XThC.Tn[14].n10 XThC.Tn[14].t25 161.202
R22574 XThC.Tn[14].n6 XThC.Tn[14].t22 161.202
R22575 XThC.Tn[14].n3 XThC.Tn[14].t38 161.202
R22576 XThC.Tn[14].n62 XThC.Tn[14].t18 145.137
R22577 XThC.Tn[14].n58 XThC.Tn[14].t40 145.137
R22578 XThC.Tn[14].n54 XThC.Tn[14].t28 145.137
R22579 XThC.Tn[14].n50 XThC.Tn[14].t24 145.137
R22580 XThC.Tn[14].n46 XThC.Tn[14].t16 145.137
R22581 XThC.Tn[14].n42 XThC.Tn[14].t36 145.137
R22582 XThC.Tn[14].n38 XThC.Tn[14].t35 145.137
R22583 XThC.Tn[14].n34 XThC.Tn[14].t15 145.137
R22584 XThC.Tn[14].n30 XThC.Tn[14].t13 145.137
R22585 XThC.Tn[14].n26 XThC.Tn[14].t37 145.137
R22586 XThC.Tn[14].n22 XThC.Tn[14].t23 145.137
R22587 XThC.Tn[14].n18 XThC.Tn[14].t20 145.137
R22588 XThC.Tn[14].n14 XThC.Tn[14].t34 145.137
R22589 XThC.Tn[14].n10 XThC.Tn[14].t32 145.137
R22590 XThC.Tn[14].n6 XThC.Tn[14].t29 145.137
R22591 XThC.Tn[14].n3 XThC.Tn[14].t43 145.137
R22592 XThC.Tn[14].n68 XThC.Tn[14].t0 26.5955
R22593 XThC.Tn[14].n68 XThC.Tn[14].t1 26.5955
R22594 XThC.Tn[14].n72 XThC.Tn[14].t11 26.5955
R22595 XThC.Tn[14].n72 XThC.Tn[14].t10 26.5955
R22596 XThC.Tn[14].n73 XThC.Tn[14].t9 26.5955
R22597 XThC.Tn[14].n73 XThC.Tn[14].t8 26.5955
R22598 XThC.Tn[14].n69 XThC.Tn[14].t3 26.5955
R22599 XThC.Tn[14].n69 XThC.Tn[14].t2 26.5955
R22600 XThC.Tn[14].n1 XThC.Tn[14].t5 24.9236
R22601 XThC.Tn[14].n1 XThC.Tn[14].t7 24.9236
R22602 XThC.Tn[14].n0 XThC.Tn[14].t4 24.9236
R22603 XThC.Tn[14].n0 XThC.Tn[14].t6 24.9236
R22604 XThC.Tn[14] XThC.Tn[14].n74 22.9652
R22605 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22606 XThC.Tn[14].n71 XThC.Tn[14].n70 13.9299
R22607 XThC.Tn[14] XThC.Tn[14].n71 13.9299
R22608 XThC.Tn[14] XThC.Tn[14].n5 8.0245
R22609 XThC.Tn[14].n65 XThC.Tn[14].n64 7.9105
R22610 XThC.Tn[14].n61 XThC.Tn[14].n60 7.9105
R22611 XThC.Tn[14].n57 XThC.Tn[14].n56 7.9105
R22612 XThC.Tn[14].n53 XThC.Tn[14].n52 7.9105
R22613 XThC.Tn[14].n49 XThC.Tn[14].n48 7.9105
R22614 XThC.Tn[14].n45 XThC.Tn[14].n44 7.9105
R22615 XThC.Tn[14].n41 XThC.Tn[14].n40 7.9105
R22616 XThC.Tn[14].n37 XThC.Tn[14].n36 7.9105
R22617 XThC.Tn[14].n33 XThC.Tn[14].n32 7.9105
R22618 XThC.Tn[14].n29 XThC.Tn[14].n28 7.9105
R22619 XThC.Tn[14].n25 XThC.Tn[14].n24 7.9105
R22620 XThC.Tn[14].n21 XThC.Tn[14].n20 7.9105
R22621 XThC.Tn[14].n17 XThC.Tn[14].n16 7.9105
R22622 XThC.Tn[14].n13 XThC.Tn[14].n12 7.9105
R22623 XThC.Tn[14].n9 XThC.Tn[14].n8 7.9105
R22624 XThC.Tn[14].n67 XThC.Tn[14].n66 7.51947
R22625 XThC.Tn[14].n66 XThC.Tn[14] 5.85107
R22626 XThC.Tn[14].n71 XThC.Tn[14].n67 2.99115
R22627 XThC.Tn[14].n71 XThC.Tn[14] 2.87153
R22628 XThC.Tn[14].n67 XThC.Tn[14] 2.2734
R22629 XThC.Tn[14].n66 XThC.Tn[14] 1.06164
R22630 XThC.Tn[14].n9 XThC.Tn[14] 0.235138
R22631 XThC.Tn[14].n13 XThC.Tn[14] 0.235138
R22632 XThC.Tn[14].n17 XThC.Tn[14] 0.235138
R22633 XThC.Tn[14].n21 XThC.Tn[14] 0.235138
R22634 XThC.Tn[14].n25 XThC.Tn[14] 0.235138
R22635 XThC.Tn[14].n29 XThC.Tn[14] 0.235138
R22636 XThC.Tn[14].n33 XThC.Tn[14] 0.235138
R22637 XThC.Tn[14].n37 XThC.Tn[14] 0.235138
R22638 XThC.Tn[14].n41 XThC.Tn[14] 0.235138
R22639 XThC.Tn[14].n45 XThC.Tn[14] 0.235138
R22640 XThC.Tn[14].n49 XThC.Tn[14] 0.235138
R22641 XThC.Tn[14].n53 XThC.Tn[14] 0.235138
R22642 XThC.Tn[14].n57 XThC.Tn[14] 0.235138
R22643 XThC.Tn[14].n61 XThC.Tn[14] 0.235138
R22644 XThC.Tn[14].n65 XThC.Tn[14] 0.235138
R22645 XThC.Tn[14] XThC.Tn[14].n9 0.114505
R22646 XThC.Tn[14] XThC.Tn[14].n13 0.114505
R22647 XThC.Tn[14] XThC.Tn[14].n17 0.114505
R22648 XThC.Tn[14] XThC.Tn[14].n21 0.114505
R22649 XThC.Tn[14] XThC.Tn[14].n25 0.114505
R22650 XThC.Tn[14] XThC.Tn[14].n29 0.114505
R22651 XThC.Tn[14] XThC.Tn[14].n33 0.114505
R22652 XThC.Tn[14] XThC.Tn[14].n37 0.114505
R22653 XThC.Tn[14] XThC.Tn[14].n41 0.114505
R22654 XThC.Tn[14] XThC.Tn[14].n45 0.114505
R22655 XThC.Tn[14] XThC.Tn[14].n49 0.114505
R22656 XThC.Tn[14] XThC.Tn[14].n53 0.114505
R22657 XThC.Tn[14] XThC.Tn[14].n57 0.114505
R22658 XThC.Tn[14] XThC.Tn[14].n61 0.114505
R22659 XThC.Tn[14] XThC.Tn[14].n65 0.114505
R22660 XThC.Tn[14].n64 XThC.Tn[14].n63 0.0599512
R22661 XThC.Tn[14].n60 XThC.Tn[14].n59 0.0599512
R22662 XThC.Tn[14].n56 XThC.Tn[14].n55 0.0599512
R22663 XThC.Tn[14].n52 XThC.Tn[14].n51 0.0599512
R22664 XThC.Tn[14].n48 XThC.Tn[14].n47 0.0599512
R22665 XThC.Tn[14].n44 XThC.Tn[14].n43 0.0599512
R22666 XThC.Tn[14].n40 XThC.Tn[14].n39 0.0599512
R22667 XThC.Tn[14].n36 XThC.Tn[14].n35 0.0599512
R22668 XThC.Tn[14].n32 XThC.Tn[14].n31 0.0599512
R22669 XThC.Tn[14].n28 XThC.Tn[14].n27 0.0599512
R22670 XThC.Tn[14].n24 XThC.Tn[14].n23 0.0599512
R22671 XThC.Tn[14].n20 XThC.Tn[14].n19 0.0599512
R22672 XThC.Tn[14].n16 XThC.Tn[14].n15 0.0599512
R22673 XThC.Tn[14].n12 XThC.Tn[14].n11 0.0599512
R22674 XThC.Tn[14].n8 XThC.Tn[14].n7 0.0599512
R22675 XThC.Tn[14].n5 XThC.Tn[14].n4 0.0599512
R22676 XThC.Tn[14].n63 XThC.Tn[14] 0.0469286
R22677 XThC.Tn[14].n59 XThC.Tn[14] 0.0469286
R22678 XThC.Tn[14].n55 XThC.Tn[14] 0.0469286
R22679 XThC.Tn[14].n51 XThC.Tn[14] 0.0469286
R22680 XThC.Tn[14].n47 XThC.Tn[14] 0.0469286
R22681 XThC.Tn[14].n43 XThC.Tn[14] 0.0469286
R22682 XThC.Tn[14].n39 XThC.Tn[14] 0.0469286
R22683 XThC.Tn[14].n35 XThC.Tn[14] 0.0469286
R22684 XThC.Tn[14].n31 XThC.Tn[14] 0.0469286
R22685 XThC.Tn[14].n27 XThC.Tn[14] 0.0469286
R22686 XThC.Tn[14].n23 XThC.Tn[14] 0.0469286
R22687 XThC.Tn[14].n19 XThC.Tn[14] 0.0469286
R22688 XThC.Tn[14].n15 XThC.Tn[14] 0.0469286
R22689 XThC.Tn[14].n11 XThC.Tn[14] 0.0469286
R22690 XThC.Tn[14].n7 XThC.Tn[14] 0.0469286
R22691 XThC.Tn[14].n4 XThC.Tn[14] 0.0469286
R22692 XThC.Tn[14].n63 XThC.Tn[14] 0.0401341
R22693 XThC.Tn[14].n59 XThC.Tn[14] 0.0401341
R22694 XThC.Tn[14].n55 XThC.Tn[14] 0.0401341
R22695 XThC.Tn[14].n51 XThC.Tn[14] 0.0401341
R22696 XThC.Tn[14].n47 XThC.Tn[14] 0.0401341
R22697 XThC.Tn[14].n43 XThC.Tn[14] 0.0401341
R22698 XThC.Tn[14].n39 XThC.Tn[14] 0.0401341
R22699 XThC.Tn[14].n35 XThC.Tn[14] 0.0401341
R22700 XThC.Tn[14].n31 XThC.Tn[14] 0.0401341
R22701 XThC.Tn[14].n27 XThC.Tn[14] 0.0401341
R22702 XThC.Tn[14].n23 XThC.Tn[14] 0.0401341
R22703 XThC.Tn[14].n19 XThC.Tn[14] 0.0401341
R22704 XThC.Tn[14].n15 XThC.Tn[14] 0.0401341
R22705 XThC.Tn[14].n11 XThC.Tn[14] 0.0401341
R22706 XThC.Tn[14].n7 XThC.Tn[14] 0.0401341
R22707 XThC.Tn[14].n4 XThC.Tn[14] 0.0401341
R22708 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R22709 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R22710 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R22711 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R22712 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R22713 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R22714 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R22715 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R22716 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R22717 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22718 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22719 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22720 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22721 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22722 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22723 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22724 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22725 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22726 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22727 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22728 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22729 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22730 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22731 XThC.XTB1.Y.n0 XThC.XTB1.Y.t2 132.067
R22732 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22733 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22734 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22735 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22736 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22737 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22738 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22739 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22740 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22741 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22742 XThC.XTB1.Y.n2 XThC.XTB1.Y.t1 26.5955
R22743 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22744 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22745 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22746 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22747 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22748 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22749 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22750 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22751 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22752 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22753 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22754 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22755 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22756 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22757 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22758 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22759 XThC.Tn[8].n71 XThC.Tn[8].n70 256.104
R22760 XThC.Tn[8].n75 XThC.Tn[8].n74 243.679
R22761 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22762 XThC.Tn[8].n75 XThC.Tn[8].n73 205.28
R22763 XThC.Tn[8].n71 XThC.Tn[8].n69 202.095
R22764 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22765 XThC.Tn[8].n65 XThC.Tn[8].n63 161.365
R22766 XThC.Tn[8].n61 XThC.Tn[8].n59 161.365
R22767 XThC.Tn[8].n57 XThC.Tn[8].n55 161.365
R22768 XThC.Tn[8].n53 XThC.Tn[8].n51 161.365
R22769 XThC.Tn[8].n49 XThC.Tn[8].n47 161.365
R22770 XThC.Tn[8].n45 XThC.Tn[8].n43 161.365
R22771 XThC.Tn[8].n41 XThC.Tn[8].n39 161.365
R22772 XThC.Tn[8].n37 XThC.Tn[8].n35 161.365
R22773 XThC.Tn[8].n33 XThC.Tn[8].n31 161.365
R22774 XThC.Tn[8].n29 XThC.Tn[8].n27 161.365
R22775 XThC.Tn[8].n25 XThC.Tn[8].n23 161.365
R22776 XThC.Tn[8].n21 XThC.Tn[8].n19 161.365
R22777 XThC.Tn[8].n17 XThC.Tn[8].n15 161.365
R22778 XThC.Tn[8].n13 XThC.Tn[8].n11 161.365
R22779 XThC.Tn[8].n9 XThC.Tn[8].n7 161.365
R22780 XThC.Tn[8].n6 XThC.Tn[8].n4 161.365
R22781 XThC.Tn[8].n63 XThC.Tn[8].t15 161.202
R22782 XThC.Tn[8].n59 XThC.Tn[8].t37 161.202
R22783 XThC.Tn[8].n55 XThC.Tn[8].t24 161.202
R22784 XThC.Tn[8].n51 XThC.Tn[8].t21 161.202
R22785 XThC.Tn[8].n47 XThC.Tn[8].t13 161.202
R22786 XThC.Tn[8].n43 XThC.Tn[8].t32 161.202
R22787 XThC.Tn[8].n39 XThC.Tn[8].t31 161.202
R22788 XThC.Tn[8].n35 XThC.Tn[8].t12 161.202
R22789 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R22790 XThC.Tn[8].n27 XThC.Tn[8].t33 161.202
R22791 XThC.Tn[8].n23 XThC.Tn[8].t20 161.202
R22792 XThC.Tn[8].n19 XThC.Tn[8].t19 161.202
R22793 XThC.Tn[8].n15 XThC.Tn[8].t30 161.202
R22794 XThC.Tn[8].n11 XThC.Tn[8].t28 161.202
R22795 XThC.Tn[8].n7 XThC.Tn[8].t26 161.202
R22796 XThC.Tn[8].n4 XThC.Tn[8].t41 161.202
R22797 XThC.Tn[8].n63 XThC.Tn[8].t18 145.137
R22798 XThC.Tn[8].n59 XThC.Tn[8].t40 145.137
R22799 XThC.Tn[8].n55 XThC.Tn[8].t27 145.137
R22800 XThC.Tn[8].n51 XThC.Tn[8].t25 145.137
R22801 XThC.Tn[8].n47 XThC.Tn[8].t17 145.137
R22802 XThC.Tn[8].n43 XThC.Tn[8].t38 145.137
R22803 XThC.Tn[8].n39 XThC.Tn[8].t36 145.137
R22804 XThC.Tn[8].n35 XThC.Tn[8].t16 145.137
R22805 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R22806 XThC.Tn[8].n27 XThC.Tn[8].t39 145.137
R22807 XThC.Tn[8].n23 XThC.Tn[8].t23 145.137
R22808 XThC.Tn[8].n19 XThC.Tn[8].t22 145.137
R22809 XThC.Tn[8].n15 XThC.Tn[8].t35 145.137
R22810 XThC.Tn[8].n11 XThC.Tn[8].t34 145.137
R22811 XThC.Tn[8].n7 XThC.Tn[8].t29 145.137
R22812 XThC.Tn[8].n4 XThC.Tn[8].t43 145.137
R22813 XThC.Tn[8].n69 XThC.Tn[8].t5 26.5955
R22814 XThC.Tn[8].n69 XThC.Tn[8].t6 26.5955
R22815 XThC.Tn[8].n70 XThC.Tn[8].t4 26.5955
R22816 XThC.Tn[8].n70 XThC.Tn[8].t7 26.5955
R22817 XThC.Tn[8].n73 XThC.Tn[8].t2 26.5955
R22818 XThC.Tn[8].n73 XThC.Tn[8].t1 26.5955
R22819 XThC.Tn[8].n74 XThC.Tn[8].t0 26.5955
R22820 XThC.Tn[8].n74 XThC.Tn[8].t3 26.5955
R22821 XThC.Tn[8].n1 XThC.Tn[8].t11 24.9236
R22822 XThC.Tn[8].n1 XThC.Tn[8].t10 24.9236
R22823 XThC.Tn[8].n0 XThC.Tn[8].t9 24.9236
R22824 XThC.Tn[8].n0 XThC.Tn[8].t8 24.9236
R22825 XThC.Tn[8] XThC.Tn[8].n75 22.9652
R22826 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22827 XThC.Tn[8].n72 XThC.Tn[8].n71 13.9299
R22828 XThC.Tn[8] XThC.Tn[8].n72 13.9299
R22829 XThC.Tn[8] XThC.Tn[8].n6 8.0245
R22830 XThC.Tn[8].n66 XThC.Tn[8].n65 7.9105
R22831 XThC.Tn[8].n62 XThC.Tn[8].n61 7.9105
R22832 XThC.Tn[8].n58 XThC.Tn[8].n57 7.9105
R22833 XThC.Tn[8].n54 XThC.Tn[8].n53 7.9105
R22834 XThC.Tn[8].n50 XThC.Tn[8].n49 7.9105
R22835 XThC.Tn[8].n46 XThC.Tn[8].n45 7.9105
R22836 XThC.Tn[8].n42 XThC.Tn[8].n41 7.9105
R22837 XThC.Tn[8].n38 XThC.Tn[8].n37 7.9105
R22838 XThC.Tn[8].n34 XThC.Tn[8].n33 7.9105
R22839 XThC.Tn[8].n30 XThC.Tn[8].n29 7.9105
R22840 XThC.Tn[8].n26 XThC.Tn[8].n25 7.9105
R22841 XThC.Tn[8].n22 XThC.Tn[8].n21 7.9105
R22842 XThC.Tn[8].n18 XThC.Tn[8].n17 7.9105
R22843 XThC.Tn[8].n14 XThC.Tn[8].n13 7.9105
R22844 XThC.Tn[8].n10 XThC.Tn[8].n9 7.9105
R22845 XThC.Tn[8].n68 XThC.Tn[8].n67 7.42331
R22846 XThC.Tn[8].n67 XThC.Tn[8] 4.24005
R22847 XThC.Tn[8].n72 XThC.Tn[8].n68 2.99115
R22848 XThC.Tn[8].n72 XThC.Tn[8] 2.87153
R22849 XThC.Tn[8].n68 XThC.Tn[8] 2.2734
R22850 XThC.Tn[8].n3 XThC.Tn[8] 0.672375
R22851 XThC.Tn[8].n10 XThC.Tn[8] 0.235138
R22852 XThC.Tn[8].n14 XThC.Tn[8] 0.235138
R22853 XThC.Tn[8].n18 XThC.Tn[8] 0.235138
R22854 XThC.Tn[8].n22 XThC.Tn[8] 0.235138
R22855 XThC.Tn[8].n26 XThC.Tn[8] 0.235138
R22856 XThC.Tn[8].n30 XThC.Tn[8] 0.235138
R22857 XThC.Tn[8].n34 XThC.Tn[8] 0.235138
R22858 XThC.Tn[8].n38 XThC.Tn[8] 0.235138
R22859 XThC.Tn[8].n42 XThC.Tn[8] 0.235138
R22860 XThC.Tn[8].n46 XThC.Tn[8] 0.235138
R22861 XThC.Tn[8].n50 XThC.Tn[8] 0.235138
R22862 XThC.Tn[8].n54 XThC.Tn[8] 0.235138
R22863 XThC.Tn[8].n58 XThC.Tn[8] 0.235138
R22864 XThC.Tn[8].n62 XThC.Tn[8] 0.235138
R22865 XThC.Tn[8].n66 XThC.Tn[8] 0.235138
R22866 XThC.Tn[8].n67 XThC.Tn[8].n3 0.220435
R22867 XThC.Tn[8].n3 XThC.Tn[8] 0.168469
R22868 XThC.Tn[8] XThC.Tn[8].n10 0.114505
R22869 XThC.Tn[8] XThC.Tn[8].n14 0.114505
R22870 XThC.Tn[8] XThC.Tn[8].n18 0.114505
R22871 XThC.Tn[8] XThC.Tn[8].n22 0.114505
R22872 XThC.Tn[8] XThC.Tn[8].n26 0.114505
R22873 XThC.Tn[8] XThC.Tn[8].n30 0.114505
R22874 XThC.Tn[8] XThC.Tn[8].n34 0.114505
R22875 XThC.Tn[8] XThC.Tn[8].n38 0.114505
R22876 XThC.Tn[8] XThC.Tn[8].n42 0.114505
R22877 XThC.Tn[8] XThC.Tn[8].n46 0.114505
R22878 XThC.Tn[8] XThC.Tn[8].n50 0.114505
R22879 XThC.Tn[8] XThC.Tn[8].n54 0.114505
R22880 XThC.Tn[8] XThC.Tn[8].n58 0.114505
R22881 XThC.Tn[8] XThC.Tn[8].n62 0.114505
R22882 XThC.Tn[8] XThC.Tn[8].n66 0.114505
R22883 XThC.Tn[8].n65 XThC.Tn[8].n64 0.0599512
R22884 XThC.Tn[8].n61 XThC.Tn[8].n60 0.0599512
R22885 XThC.Tn[8].n57 XThC.Tn[8].n56 0.0599512
R22886 XThC.Tn[8].n53 XThC.Tn[8].n52 0.0599512
R22887 XThC.Tn[8].n49 XThC.Tn[8].n48 0.0599512
R22888 XThC.Tn[8].n45 XThC.Tn[8].n44 0.0599512
R22889 XThC.Tn[8].n41 XThC.Tn[8].n40 0.0599512
R22890 XThC.Tn[8].n37 XThC.Tn[8].n36 0.0599512
R22891 XThC.Tn[8].n33 XThC.Tn[8].n32 0.0599512
R22892 XThC.Tn[8].n29 XThC.Tn[8].n28 0.0599512
R22893 XThC.Tn[8].n25 XThC.Tn[8].n24 0.0599512
R22894 XThC.Tn[8].n21 XThC.Tn[8].n20 0.0599512
R22895 XThC.Tn[8].n17 XThC.Tn[8].n16 0.0599512
R22896 XThC.Tn[8].n13 XThC.Tn[8].n12 0.0599512
R22897 XThC.Tn[8].n9 XThC.Tn[8].n8 0.0599512
R22898 XThC.Tn[8].n6 XThC.Tn[8].n5 0.0599512
R22899 XThC.Tn[8].n64 XThC.Tn[8] 0.0469286
R22900 XThC.Tn[8].n60 XThC.Tn[8] 0.0469286
R22901 XThC.Tn[8].n56 XThC.Tn[8] 0.0469286
R22902 XThC.Tn[8].n52 XThC.Tn[8] 0.0469286
R22903 XThC.Tn[8].n48 XThC.Tn[8] 0.0469286
R22904 XThC.Tn[8].n44 XThC.Tn[8] 0.0469286
R22905 XThC.Tn[8].n40 XThC.Tn[8] 0.0469286
R22906 XThC.Tn[8].n36 XThC.Tn[8] 0.0469286
R22907 XThC.Tn[8].n32 XThC.Tn[8] 0.0469286
R22908 XThC.Tn[8].n28 XThC.Tn[8] 0.0469286
R22909 XThC.Tn[8].n24 XThC.Tn[8] 0.0469286
R22910 XThC.Tn[8].n20 XThC.Tn[8] 0.0469286
R22911 XThC.Tn[8].n16 XThC.Tn[8] 0.0469286
R22912 XThC.Tn[8].n12 XThC.Tn[8] 0.0469286
R22913 XThC.Tn[8].n8 XThC.Tn[8] 0.0469286
R22914 XThC.Tn[8].n5 XThC.Tn[8] 0.0469286
R22915 XThC.Tn[8].n64 XThC.Tn[8] 0.0401341
R22916 XThC.Tn[8].n60 XThC.Tn[8] 0.0401341
R22917 XThC.Tn[8].n56 XThC.Tn[8] 0.0401341
R22918 XThC.Tn[8].n52 XThC.Tn[8] 0.0401341
R22919 XThC.Tn[8].n48 XThC.Tn[8] 0.0401341
R22920 XThC.Tn[8].n44 XThC.Tn[8] 0.0401341
R22921 XThC.Tn[8].n40 XThC.Tn[8] 0.0401341
R22922 XThC.Tn[8].n36 XThC.Tn[8] 0.0401341
R22923 XThC.Tn[8].n32 XThC.Tn[8] 0.0401341
R22924 XThC.Tn[8].n28 XThC.Tn[8] 0.0401341
R22925 XThC.Tn[8].n24 XThC.Tn[8] 0.0401341
R22926 XThC.Tn[8].n20 XThC.Tn[8] 0.0401341
R22927 XThC.Tn[8].n16 XThC.Tn[8] 0.0401341
R22928 XThC.Tn[8].n12 XThC.Tn[8] 0.0401341
R22929 XThC.Tn[8].n8 XThC.Tn[8] 0.0401341
R22930 XThC.Tn[8].n5 XThC.Tn[8] 0.0401341
R22931 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R22932 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R22933 XThR.Tn[1] XThR.Tn[1].n82 161.363
R22934 XThR.Tn[1] XThR.Tn[1].n77 161.363
R22935 XThR.Tn[1] XThR.Tn[1].n72 161.363
R22936 XThR.Tn[1] XThR.Tn[1].n67 161.363
R22937 XThR.Tn[1] XThR.Tn[1].n62 161.363
R22938 XThR.Tn[1] XThR.Tn[1].n57 161.363
R22939 XThR.Tn[1] XThR.Tn[1].n52 161.363
R22940 XThR.Tn[1] XThR.Tn[1].n47 161.363
R22941 XThR.Tn[1] XThR.Tn[1].n42 161.363
R22942 XThR.Tn[1] XThR.Tn[1].n37 161.363
R22943 XThR.Tn[1] XThR.Tn[1].n32 161.363
R22944 XThR.Tn[1] XThR.Tn[1].n27 161.363
R22945 XThR.Tn[1] XThR.Tn[1].n22 161.363
R22946 XThR.Tn[1] XThR.Tn[1].n17 161.363
R22947 XThR.Tn[1] XThR.Tn[1].n12 161.363
R22948 XThR.Tn[1] XThR.Tn[1].n10 161.363
R22949 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R22950 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R22951 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R22952 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R22953 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R22954 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R22955 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R22956 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R22957 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R22958 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R22959 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R22960 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R22961 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R22962 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R22963 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R22964 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R22965 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R22966 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R22967 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R22968 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R22969 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R22970 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R22971 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R22972 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R22973 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R22974 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R22975 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R22976 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R22977 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R22978 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R22979 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R22980 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R22981 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R22982 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R22983 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R22984 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R22985 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R22986 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R22987 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R22988 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R22989 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R22990 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R22991 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R22992 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R22993 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R22994 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R22995 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R22996 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R22997 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R22998 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R22999 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R23000 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R23001 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R23002 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R23003 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R23004 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R23005 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R23006 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R23007 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R23008 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R23009 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R23010 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R23011 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R23012 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R23013 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R23014 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R23015 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R23016 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R23017 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R23018 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R23019 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R23020 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R23021 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R23022 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R23023 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R23024 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R23025 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R23026 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R23027 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R23028 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R23029 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R23030 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R23031 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R23032 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R23033 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R23034 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R23035 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R23036 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R23037 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R23038 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R23039 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R23040 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R23041 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R23042 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R23043 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R23044 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R23045 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R23046 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R23047 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R23048 XThR.Tn[1] XThR.Tn[1].n11 5.34038
R23049 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R23050 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R23051 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R23052 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R23053 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R23054 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R23055 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R23056 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R23057 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R23058 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R23059 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R23060 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R23061 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R23062 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R23063 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R23064 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R23065 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R23066 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R23067 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R23068 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R23069 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R23070 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R23071 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R23072 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R23073 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R23074 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R23075 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R23076 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R23077 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R23078 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R23079 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R23080 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R23081 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R23082 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R23083 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R23084 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R23085 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R23086 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R23087 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R23088 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R23089 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R23090 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R23091 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R23092 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R23093 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R23094 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R23095 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R23096 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R23097 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R23098 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R23099 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R23100 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R23101 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R23102 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R23103 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R23104 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R23105 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R23106 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R23107 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R23108 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R23109 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R23110 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R23111 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R23112 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R23113 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R23114 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R23115 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R23116 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R23117 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R23118 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R23119 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R23120 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R23121 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R23122 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R23123 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R23124 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R23125 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R23126 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R23127 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R23128 XThR.Tn[1] XThR.Tn[1].n87 0.038
R23129 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R23130 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R23131 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R23132 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R23133 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R23134 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R23135 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R23136 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R23137 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R23138 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R23139 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R23140 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R23141 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R23142 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R23143 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R23144 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R23145 XThC.Tn[7].n5 XThC.Tn[7].n4 255.096
R23146 XThC.Tn[7].n2 XThC.Tn[7].n0 236.589
R23147 XThC.Tn[7].n5 XThC.Tn[7].n3 201.845
R23148 XThC.Tn[7].n2 XThC.Tn[7].n1 200.321
R23149 XThC.Tn[7].n67 XThC.Tn[7].n65 161.365
R23150 XThC.Tn[7].n63 XThC.Tn[7].n61 161.365
R23151 XThC.Tn[7].n59 XThC.Tn[7].n57 161.365
R23152 XThC.Tn[7].n55 XThC.Tn[7].n53 161.365
R23153 XThC.Tn[7].n51 XThC.Tn[7].n49 161.365
R23154 XThC.Tn[7].n47 XThC.Tn[7].n45 161.365
R23155 XThC.Tn[7].n43 XThC.Tn[7].n41 161.365
R23156 XThC.Tn[7].n39 XThC.Tn[7].n37 161.365
R23157 XThC.Tn[7].n35 XThC.Tn[7].n33 161.365
R23158 XThC.Tn[7].n31 XThC.Tn[7].n29 161.365
R23159 XThC.Tn[7].n27 XThC.Tn[7].n25 161.365
R23160 XThC.Tn[7].n23 XThC.Tn[7].n21 161.365
R23161 XThC.Tn[7].n19 XThC.Tn[7].n17 161.365
R23162 XThC.Tn[7].n15 XThC.Tn[7].n13 161.365
R23163 XThC.Tn[7].n11 XThC.Tn[7].n9 161.365
R23164 XThC.Tn[7].n8 XThC.Tn[7].n6 161.365
R23165 XThC.Tn[7].n65 XThC.Tn[7].t19 161.202
R23166 XThC.Tn[7].n61 XThC.Tn[7].t9 161.202
R23167 XThC.Tn[7].n57 XThC.Tn[7].t28 161.202
R23168 XThC.Tn[7].n53 XThC.Tn[7].t26 161.202
R23169 XThC.Tn[7].n49 XThC.Tn[7].t17 161.202
R23170 XThC.Tn[7].n45 XThC.Tn[7].t38 161.202
R23171 XThC.Tn[7].n41 XThC.Tn[7].t36 161.202
R23172 XThC.Tn[7].n37 XThC.Tn[7].t16 161.202
R23173 XThC.Tn[7].n33 XThC.Tn[7].t14 161.202
R23174 XThC.Tn[7].n29 XThC.Tn[7].t39 161.202
R23175 XThC.Tn[7].n25 XThC.Tn[7].t23 161.202
R23176 XThC.Tn[7].n21 XThC.Tn[7].t22 161.202
R23177 XThC.Tn[7].n17 XThC.Tn[7].t35 161.202
R23178 XThC.Tn[7].n13 XThC.Tn[7].t34 161.202
R23179 XThC.Tn[7].n9 XThC.Tn[7].t30 161.202
R23180 XThC.Tn[7].n6 XThC.Tn[7].t11 161.202
R23181 XThC.Tn[7].n65 XThC.Tn[7].t15 145.137
R23182 XThC.Tn[7].n61 XThC.Tn[7].t37 145.137
R23183 XThC.Tn[7].n57 XThC.Tn[7].t24 145.137
R23184 XThC.Tn[7].n53 XThC.Tn[7].t21 145.137
R23185 XThC.Tn[7].n49 XThC.Tn[7].t13 145.137
R23186 XThC.Tn[7].n45 XThC.Tn[7].t32 145.137
R23187 XThC.Tn[7].n41 XThC.Tn[7].t31 145.137
R23188 XThC.Tn[7].n37 XThC.Tn[7].t12 145.137
R23189 XThC.Tn[7].n33 XThC.Tn[7].t10 145.137
R23190 XThC.Tn[7].n29 XThC.Tn[7].t33 145.137
R23191 XThC.Tn[7].n25 XThC.Tn[7].t20 145.137
R23192 XThC.Tn[7].n21 XThC.Tn[7].t18 145.137
R23193 XThC.Tn[7].n17 XThC.Tn[7].t29 145.137
R23194 XThC.Tn[7].n13 XThC.Tn[7].t27 145.137
R23195 XThC.Tn[7].n9 XThC.Tn[7].t25 145.137
R23196 XThC.Tn[7].n6 XThC.Tn[7].t8 145.137
R23197 XThC.Tn[7].n4 XThC.Tn[7].t2 26.5955
R23198 XThC.Tn[7].n4 XThC.Tn[7].t1 26.5955
R23199 XThC.Tn[7].n3 XThC.Tn[7].t0 26.5955
R23200 XThC.Tn[7].n3 XThC.Tn[7].t3 26.5955
R23201 XThC.Tn[7] XThC.Tn[7].n5 26.4992
R23202 XThC.Tn[7].n0 XThC.Tn[7].t6 24.9236
R23203 XThC.Tn[7].n0 XThC.Tn[7].t5 24.9236
R23204 XThC.Tn[7].n1 XThC.Tn[7].t4 24.9236
R23205 XThC.Tn[7].n1 XThC.Tn[7].t7 24.9236
R23206 XThC.Tn[7].n70 XThC.Tn[7].n2 12.0894
R23207 XThC.Tn[7].n70 XThC.Tn[7] 9.64206
R23208 XThC.Tn[7].n69 XThC.Tn[7] 8.14595
R23209 XThC.Tn[7] XThC.Tn[7].n8 8.0245
R23210 XThC.Tn[7].n68 XThC.Tn[7].n67 7.9105
R23211 XThC.Tn[7].n64 XThC.Tn[7].n63 7.9105
R23212 XThC.Tn[7].n60 XThC.Tn[7].n59 7.9105
R23213 XThC.Tn[7].n56 XThC.Tn[7].n55 7.9105
R23214 XThC.Tn[7].n52 XThC.Tn[7].n51 7.9105
R23215 XThC.Tn[7].n48 XThC.Tn[7].n47 7.9105
R23216 XThC.Tn[7].n44 XThC.Tn[7].n43 7.9105
R23217 XThC.Tn[7].n40 XThC.Tn[7].n39 7.9105
R23218 XThC.Tn[7].n36 XThC.Tn[7].n35 7.9105
R23219 XThC.Tn[7].n32 XThC.Tn[7].n31 7.9105
R23220 XThC.Tn[7].n28 XThC.Tn[7].n27 7.9105
R23221 XThC.Tn[7].n24 XThC.Tn[7].n23 7.9105
R23222 XThC.Tn[7].n20 XThC.Tn[7].n19 7.9105
R23223 XThC.Tn[7].n16 XThC.Tn[7].n15 7.9105
R23224 XThC.Tn[7].n12 XThC.Tn[7].n11 7.9105
R23225 XThC.Tn[7].n69 XThC.Tn[7] 5.30358
R23226 XThC.Tn[7] XThC.Tn[7].n69 3.15894
R23227 XThC.Tn[7] XThC.Tn[7].n70 1.66284
R23228 XThC.Tn[7].n12 XThC.Tn[7] 0.235138
R23229 XThC.Tn[7].n16 XThC.Tn[7] 0.235138
R23230 XThC.Tn[7].n20 XThC.Tn[7] 0.235138
R23231 XThC.Tn[7].n24 XThC.Tn[7] 0.235138
R23232 XThC.Tn[7].n28 XThC.Tn[7] 0.235138
R23233 XThC.Tn[7].n32 XThC.Tn[7] 0.235138
R23234 XThC.Tn[7].n36 XThC.Tn[7] 0.235138
R23235 XThC.Tn[7].n40 XThC.Tn[7] 0.235138
R23236 XThC.Tn[7].n44 XThC.Tn[7] 0.235138
R23237 XThC.Tn[7].n48 XThC.Tn[7] 0.235138
R23238 XThC.Tn[7].n52 XThC.Tn[7] 0.235138
R23239 XThC.Tn[7].n56 XThC.Tn[7] 0.235138
R23240 XThC.Tn[7].n60 XThC.Tn[7] 0.235138
R23241 XThC.Tn[7].n64 XThC.Tn[7] 0.235138
R23242 XThC.Tn[7].n68 XThC.Tn[7] 0.235138
R23243 XThC.Tn[7] XThC.Tn[7].n12 0.114505
R23244 XThC.Tn[7] XThC.Tn[7].n16 0.114505
R23245 XThC.Tn[7] XThC.Tn[7].n20 0.114505
R23246 XThC.Tn[7] XThC.Tn[7].n24 0.114505
R23247 XThC.Tn[7] XThC.Tn[7].n28 0.114505
R23248 XThC.Tn[7] XThC.Tn[7].n32 0.114505
R23249 XThC.Tn[7] XThC.Tn[7].n36 0.114505
R23250 XThC.Tn[7] XThC.Tn[7].n40 0.114505
R23251 XThC.Tn[7] XThC.Tn[7].n44 0.114505
R23252 XThC.Tn[7] XThC.Tn[7].n48 0.114505
R23253 XThC.Tn[7] XThC.Tn[7].n52 0.114505
R23254 XThC.Tn[7] XThC.Tn[7].n56 0.114505
R23255 XThC.Tn[7] XThC.Tn[7].n60 0.114505
R23256 XThC.Tn[7] XThC.Tn[7].n64 0.114505
R23257 XThC.Tn[7] XThC.Tn[7].n68 0.114505
R23258 XThC.Tn[7].n67 XThC.Tn[7].n66 0.0599512
R23259 XThC.Tn[7].n63 XThC.Tn[7].n62 0.0599512
R23260 XThC.Tn[7].n59 XThC.Tn[7].n58 0.0599512
R23261 XThC.Tn[7].n55 XThC.Tn[7].n54 0.0599512
R23262 XThC.Tn[7].n51 XThC.Tn[7].n50 0.0599512
R23263 XThC.Tn[7].n47 XThC.Tn[7].n46 0.0599512
R23264 XThC.Tn[7].n43 XThC.Tn[7].n42 0.0599512
R23265 XThC.Tn[7].n39 XThC.Tn[7].n38 0.0599512
R23266 XThC.Tn[7].n35 XThC.Tn[7].n34 0.0599512
R23267 XThC.Tn[7].n31 XThC.Tn[7].n30 0.0599512
R23268 XThC.Tn[7].n27 XThC.Tn[7].n26 0.0599512
R23269 XThC.Tn[7].n23 XThC.Tn[7].n22 0.0599512
R23270 XThC.Tn[7].n19 XThC.Tn[7].n18 0.0599512
R23271 XThC.Tn[7].n15 XThC.Tn[7].n14 0.0599512
R23272 XThC.Tn[7].n11 XThC.Tn[7].n10 0.0599512
R23273 XThC.Tn[7].n8 XThC.Tn[7].n7 0.0599512
R23274 XThC.Tn[7].n66 XThC.Tn[7] 0.0469286
R23275 XThC.Tn[7].n62 XThC.Tn[7] 0.0469286
R23276 XThC.Tn[7].n58 XThC.Tn[7] 0.0469286
R23277 XThC.Tn[7].n54 XThC.Tn[7] 0.0469286
R23278 XThC.Tn[7].n50 XThC.Tn[7] 0.0469286
R23279 XThC.Tn[7].n46 XThC.Tn[7] 0.0469286
R23280 XThC.Tn[7].n42 XThC.Tn[7] 0.0469286
R23281 XThC.Tn[7].n38 XThC.Tn[7] 0.0469286
R23282 XThC.Tn[7].n34 XThC.Tn[7] 0.0469286
R23283 XThC.Tn[7].n30 XThC.Tn[7] 0.0469286
R23284 XThC.Tn[7].n26 XThC.Tn[7] 0.0469286
R23285 XThC.Tn[7].n22 XThC.Tn[7] 0.0469286
R23286 XThC.Tn[7].n18 XThC.Tn[7] 0.0469286
R23287 XThC.Tn[7].n14 XThC.Tn[7] 0.0469286
R23288 XThC.Tn[7].n10 XThC.Tn[7] 0.0469286
R23289 XThC.Tn[7].n7 XThC.Tn[7] 0.0469286
R23290 XThC.Tn[7].n66 XThC.Tn[7] 0.0401341
R23291 XThC.Tn[7].n62 XThC.Tn[7] 0.0401341
R23292 XThC.Tn[7].n58 XThC.Tn[7] 0.0401341
R23293 XThC.Tn[7].n54 XThC.Tn[7] 0.0401341
R23294 XThC.Tn[7].n50 XThC.Tn[7] 0.0401341
R23295 XThC.Tn[7].n46 XThC.Tn[7] 0.0401341
R23296 XThC.Tn[7].n42 XThC.Tn[7] 0.0401341
R23297 XThC.Tn[7].n38 XThC.Tn[7] 0.0401341
R23298 XThC.Tn[7].n34 XThC.Tn[7] 0.0401341
R23299 XThC.Tn[7].n30 XThC.Tn[7] 0.0401341
R23300 XThC.Tn[7].n26 XThC.Tn[7] 0.0401341
R23301 XThC.Tn[7].n22 XThC.Tn[7] 0.0401341
R23302 XThC.Tn[7].n18 XThC.Tn[7] 0.0401341
R23303 XThC.Tn[7].n14 XThC.Tn[7] 0.0401341
R23304 XThC.Tn[7].n10 XThC.Tn[7] 0.0401341
R23305 XThC.Tn[7].n7 XThC.Tn[7] 0.0401341
R23306 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R23307 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R23308 XThR.Tn[4] XThR.Tn[4].n82 161.363
R23309 XThR.Tn[4] XThR.Tn[4].n77 161.363
R23310 XThR.Tn[4] XThR.Tn[4].n72 161.363
R23311 XThR.Tn[4] XThR.Tn[4].n67 161.363
R23312 XThR.Tn[4] XThR.Tn[4].n62 161.363
R23313 XThR.Tn[4] XThR.Tn[4].n57 161.363
R23314 XThR.Tn[4] XThR.Tn[4].n52 161.363
R23315 XThR.Tn[4] XThR.Tn[4].n47 161.363
R23316 XThR.Tn[4] XThR.Tn[4].n42 161.363
R23317 XThR.Tn[4] XThR.Tn[4].n37 161.363
R23318 XThR.Tn[4] XThR.Tn[4].n32 161.363
R23319 XThR.Tn[4] XThR.Tn[4].n27 161.363
R23320 XThR.Tn[4] XThR.Tn[4].n22 161.363
R23321 XThR.Tn[4] XThR.Tn[4].n17 161.363
R23322 XThR.Tn[4] XThR.Tn[4].n12 161.363
R23323 XThR.Tn[4] XThR.Tn[4].n10 161.363
R23324 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R23325 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R23326 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R23327 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R23328 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R23329 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R23330 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R23331 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R23332 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R23333 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R23334 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R23335 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R23336 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R23337 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R23338 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R23339 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R23340 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R23341 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R23342 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R23343 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R23344 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R23345 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R23346 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R23347 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R23348 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R23349 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R23350 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R23351 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R23352 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R23353 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R23354 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R23355 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R23356 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R23357 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R23358 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R23359 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R23360 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R23361 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R23362 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R23363 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R23364 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R23365 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R23366 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R23367 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R23368 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R23369 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R23370 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R23371 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R23372 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R23373 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R23374 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R23375 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R23376 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R23377 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R23378 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R23379 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R23380 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R23381 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R23382 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R23383 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R23384 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R23385 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R23386 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R23387 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R23388 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R23389 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R23390 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R23391 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R23392 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R23393 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R23394 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R23395 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R23396 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R23397 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R23398 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R23399 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R23400 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R23401 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R23402 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R23403 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R23404 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R23405 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R23406 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R23407 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R23408 XThR.Tn[4].n1 XThR.Tn[4].t8 26.5955
R23409 XThR.Tn[4].n1 XThR.Tn[4].t11 26.5955
R23410 XThR.Tn[4].n0 XThR.Tn[4].t9 26.5955
R23411 XThR.Tn[4].n0 XThR.Tn[4].t10 26.5955
R23412 XThR.Tn[4].n3 XThR.Tn[4].t7 24.9236
R23413 XThR.Tn[4].n3 XThR.Tn[4].t4 24.9236
R23414 XThR.Tn[4].n4 XThR.Tn[4].t6 24.9236
R23415 XThR.Tn[4].n4 XThR.Tn[4].t5 24.9236
R23416 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R23417 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R23418 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R23419 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R23420 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R23421 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R23422 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R23423 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R23424 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R23425 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R23426 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R23427 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R23428 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R23429 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R23430 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R23431 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R23432 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R23433 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R23434 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R23435 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R23436 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R23437 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R23438 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R23439 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R23440 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R23441 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R23442 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R23443 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R23444 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R23445 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R23446 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R23447 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R23448 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R23449 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R23450 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R23451 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R23452 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R23453 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R23454 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R23455 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R23456 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R23457 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R23458 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R23459 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R23460 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R23461 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R23462 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R23463 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R23464 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R23465 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R23466 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R23467 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R23468 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R23469 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R23470 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R23471 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R23472 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R23473 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R23474 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R23475 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R23476 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R23477 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R23478 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R23479 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R23480 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R23481 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R23482 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R23483 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R23484 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R23485 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R23486 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R23487 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R23488 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R23489 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R23490 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R23491 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R23492 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R23493 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R23494 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R23495 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R23496 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R23497 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R23498 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R23499 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R23500 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R23501 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R23502 XThR.Tn[4] XThR.Tn[4].n87 0.038
R23503 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R23504 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R23505 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R23506 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R23507 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R23508 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R23509 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R23510 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R23511 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R23512 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R23513 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R23514 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R23515 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R23516 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R23517 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R23518 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R23519 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R23520 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R23521 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R23522 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R23523 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R23524 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R23525 XThR.Tn[11] XThR.Tn[11].n82 161.363
R23526 XThR.Tn[11] XThR.Tn[11].n77 161.363
R23527 XThR.Tn[11] XThR.Tn[11].n72 161.363
R23528 XThR.Tn[11] XThR.Tn[11].n67 161.363
R23529 XThR.Tn[11] XThR.Tn[11].n62 161.363
R23530 XThR.Tn[11] XThR.Tn[11].n57 161.363
R23531 XThR.Tn[11] XThR.Tn[11].n52 161.363
R23532 XThR.Tn[11] XThR.Tn[11].n47 161.363
R23533 XThR.Tn[11] XThR.Tn[11].n42 161.363
R23534 XThR.Tn[11] XThR.Tn[11].n37 161.363
R23535 XThR.Tn[11] XThR.Tn[11].n32 161.363
R23536 XThR.Tn[11] XThR.Tn[11].n27 161.363
R23537 XThR.Tn[11] XThR.Tn[11].n22 161.363
R23538 XThR.Tn[11] XThR.Tn[11].n17 161.363
R23539 XThR.Tn[11] XThR.Tn[11].n12 161.363
R23540 XThR.Tn[11] XThR.Tn[11].n10 161.363
R23541 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R23542 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R23543 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R23544 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R23545 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R23546 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R23547 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R23548 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R23549 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R23550 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R23551 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R23552 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R23553 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R23554 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R23555 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R23556 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R23557 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R23558 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R23559 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R23560 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R23561 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R23562 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R23563 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R23564 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R23565 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R23566 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R23567 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R23568 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R23569 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R23570 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R23571 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R23572 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R23573 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R23574 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R23575 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R23576 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R23577 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R23578 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R23579 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R23580 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R23581 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R23582 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R23583 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R23584 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R23585 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R23586 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R23587 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R23588 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R23589 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R23590 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R23591 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R23592 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R23593 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R23594 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R23595 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R23596 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R23597 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R23598 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R23599 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R23600 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R23601 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R23602 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R23603 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R23604 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R23605 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R23606 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R23607 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R23608 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R23609 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R23610 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R23611 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R23612 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R23613 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R23614 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R23615 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R23616 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R23617 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R23618 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R23619 XThR.Tn[11].n6 XThR.Tn[11].t3 26.5955
R23620 XThR.Tn[11].n6 XThR.Tn[11].t11 26.5955
R23621 XThR.Tn[11].n7 XThR.Tn[11].t1 26.5955
R23622 XThR.Tn[11].n7 XThR.Tn[11].t10 26.5955
R23623 XThR.Tn[11].n3 XThR.Tn[11].t6 26.5955
R23624 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R23625 XThR.Tn[11].n4 XThR.Tn[11].t7 26.5955
R23626 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R23627 XThR.Tn[11].n0 XThR.Tn[11].t5 24.9236
R23628 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R23629 XThR.Tn[11].n1 XThR.Tn[11].t4 24.9236
R23630 XThR.Tn[11].n1 XThR.Tn[11].t0 24.9236
R23631 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R23632 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R23633 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R23634 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R23635 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R23636 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R23637 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R23638 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R23639 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R23640 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R23641 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R23642 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R23643 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R23644 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R23645 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R23646 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R23647 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R23648 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R23649 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R23650 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R23651 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R23652 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R23653 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R23654 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R23655 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R23656 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R23657 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R23658 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R23659 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R23660 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R23661 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R23662 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R23663 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R23664 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R23665 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R23666 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R23667 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R23668 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R23669 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R23670 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R23671 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R23672 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R23673 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R23674 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R23675 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R23676 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R23677 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R23678 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R23679 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R23680 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R23681 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R23682 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R23683 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R23684 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R23685 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R23686 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R23687 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R23688 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R23689 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R23690 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R23691 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R23692 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R23693 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R23694 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R23695 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R23696 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R23697 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R23698 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R23699 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R23700 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R23701 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R23702 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R23703 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R23704 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R23705 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R23706 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R23707 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R23708 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R23709 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R23710 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R23711 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R23712 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R23713 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R23714 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R23715 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R23716 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R23717 XThR.Tn[11] XThR.Tn[11].n87 0.038
R23718 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R23719 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R23720 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R23721 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R23722 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R23723 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R23724 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R23725 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R23726 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R23727 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R23728 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R23729 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R23730 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R23731 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R23732 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R23733 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R23734 XThR.Tn[7].n5 XThR.Tn[7].n3 244.067
R23735 XThR.Tn[7].n2 XThR.Tn[7].n0 236.589
R23736 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23737 XThR.Tn[7].n2 XThR.Tn[7].n1 200.321
R23738 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23739 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23740 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23741 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23742 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23743 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23744 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23745 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23746 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23747 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23748 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23749 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23750 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23751 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23752 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23753 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23754 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23755 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23756 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23757 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23758 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23759 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23760 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23761 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23762 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23763 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23764 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23765 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23766 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23767 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23768 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23769 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23770 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23771 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23772 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23773 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23774 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23775 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23776 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23777 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23778 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23779 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23780 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23781 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23782 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23783 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23784 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23785 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23786 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23787 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23788 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23789 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23790 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23791 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23792 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23793 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23794 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23795 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23796 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23797 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23798 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23799 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23800 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23801 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23802 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23803 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23804 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23805 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23806 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23807 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23808 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23809 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23810 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23811 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23812 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23813 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23814 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23815 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23816 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23817 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23818 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23819 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23820 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23821 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23822 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23823 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23824 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23825 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23826 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23827 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23828 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23829 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23830 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23831 XThR.Tn[7].n4 XThR.Tn[7].t1 26.5955
R23832 XThR.Tn[7].n4 XThR.Tn[7].t0 26.5955
R23833 XThR.Tn[7].n3 XThR.Tn[7].t2 26.5955
R23834 XThR.Tn[7].n3 XThR.Tn[7].t3 26.5955
R23835 XThR.Tn[7].n0 XThR.Tn[7].t7 24.9236
R23836 XThR.Tn[7].n0 XThR.Tn[7].t4 24.9236
R23837 XThR.Tn[7].n1 XThR.Tn[7].t6 24.9236
R23838 XThR.Tn[7].n1 XThR.Tn[7].t5 24.9236
R23839 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23840 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23841 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23842 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23843 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R23844 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23845 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23846 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23847 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23848 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23849 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23850 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23851 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23852 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23853 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23854 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23855 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23856 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23857 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23858 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23859 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23860 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23861 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23862 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23863 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23864 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23865 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23866 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23867 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23868 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23869 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23870 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23871 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23872 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23873 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23874 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23875 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23876 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23877 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23878 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23879 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23880 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23881 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23882 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23883 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23884 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23885 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23886 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23887 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23888 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23889 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23890 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23891 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23892 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23893 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23894 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23895 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23896 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23897 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23898 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23899 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23900 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23901 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23902 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23903 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23904 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23905 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23906 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23907 XThR.Tn[7].n6 XThR.Tn[7] 0.830612
R23908 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23909 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23910 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23911 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23912 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23913 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23914 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23915 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23916 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23917 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23918 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23919 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23920 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23921 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23922 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23923 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23924 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R23925 XThR.Tn[7] XThR.Tn[7].n84 0.038
R23926 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R23927 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R23928 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R23929 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R23930 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R23931 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R23932 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R23933 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R23934 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R23935 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R23936 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R23937 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R23938 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R23939 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R23940 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R23941 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R23942 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23943 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23944 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23945 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23946 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23947 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23948 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23949 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23950 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23951 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23952 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23953 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23954 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23955 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23956 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23957 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23958 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23959 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23960 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23961 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23962 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23963 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23964 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23965 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23966 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23967 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23968 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23969 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23970 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23971 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23972 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23973 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23974 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23975 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23976 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23977 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23978 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23979 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23980 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23981 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23982 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23983 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23984 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23985 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23986 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23987 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23988 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23989 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23990 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23991 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23992 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23993 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23994 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23995 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23996 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23997 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R23998 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R23999 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R24000 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R24001 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R24002 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R24003 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R24004 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R24005 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R24006 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R24007 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R24008 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R24009 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R24010 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R24011 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R24012 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R24013 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R24014 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R24015 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R24016 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R24017 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R24018 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R24019 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R24020 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R24021 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R24022 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R24023 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R24024 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R24025 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R24026 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R24027 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R24028 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R24029 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R24030 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R24031 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R24032 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R24033 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R24034 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R24035 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R24036 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R24037 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R24038 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R24039 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R24040 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R24041 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R24042 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R24043 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R24044 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R24045 XThR.Tn[0].n1 XThR.Tn[0].t3 26.5955
R24046 XThR.Tn[0].n0 XThR.Tn[0].t5 26.5955
R24047 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R24048 XThR.Tn[0].n3 XThR.Tn[0].t8 24.9236
R24049 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R24050 XThR.Tn[0].n4 XThR.Tn[0].t7 24.9236
R24051 XThR.Tn[0].n4 XThR.Tn[0].t10 24.9236
R24052 XThR.Tn[0].n5 XThR.Tn[0].t11 24.9236
R24053 XThR.Tn[0].n5 XThR.Tn[0].t1 24.9236
R24054 XThR.Tn[0].n6 XThR.Tn[0].t2 24.9236
R24055 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R24056 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R24057 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R24058 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R24059 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R24060 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R24061 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R24062 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R24063 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R24064 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R24065 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R24066 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R24067 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R24068 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R24069 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R24070 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R24071 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R24072 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R24073 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R24074 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R24075 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R24076 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R24077 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R24078 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R24079 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R24080 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R24081 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R24082 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R24083 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R24084 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R24085 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R24086 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R24087 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R24088 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R24089 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R24090 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R24091 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R24092 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R24093 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R24094 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R24095 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R24096 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R24097 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R24098 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R24099 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R24100 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R24101 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R24102 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R24103 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R24104 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R24105 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R24106 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R24107 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R24108 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R24109 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R24110 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R24111 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R24112 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R24113 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R24114 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R24115 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R24116 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R24117 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R24118 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R24119 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R24120 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R24121 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R24122 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R24123 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R24124 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R24125 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R24126 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R24127 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R24128 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R24129 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R24130 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R24131 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R24132 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R24133 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R24134 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R24135 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R24136 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R24137 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R24138 XThR.Tn[0] XThR.Tn[0].n87 0.038
R24139 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R24140 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R24141 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R24142 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R24143 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R24144 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R24145 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R24146 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R24147 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R24148 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R24149 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R24150 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R24151 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R24152 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R24153 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R24154 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R24155 XThR.Tn[8].n5 XThR.Tn[8].n4 256.103
R24156 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R24157 XThR.Tn[8].n88 XThR.Tn[8].n86 241.847
R24158 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R24159 XThR.Tn[8].n5 XThR.Tn[8].n3 202.095
R24160 XThR.Tn[8].n88 XThR.Tn[8].n87 185
R24161 XThR.Tn[8] XThR.Tn[8].n79 161.363
R24162 XThR.Tn[8] XThR.Tn[8].n74 161.363
R24163 XThR.Tn[8] XThR.Tn[8].n69 161.363
R24164 XThR.Tn[8] XThR.Tn[8].n64 161.363
R24165 XThR.Tn[8] XThR.Tn[8].n59 161.363
R24166 XThR.Tn[8] XThR.Tn[8].n54 161.363
R24167 XThR.Tn[8] XThR.Tn[8].n49 161.363
R24168 XThR.Tn[8] XThR.Tn[8].n44 161.363
R24169 XThR.Tn[8] XThR.Tn[8].n39 161.363
R24170 XThR.Tn[8] XThR.Tn[8].n34 161.363
R24171 XThR.Tn[8] XThR.Tn[8].n29 161.363
R24172 XThR.Tn[8] XThR.Tn[8].n24 161.363
R24173 XThR.Tn[8] XThR.Tn[8].n19 161.363
R24174 XThR.Tn[8] XThR.Tn[8].n14 161.363
R24175 XThR.Tn[8] XThR.Tn[8].n9 161.363
R24176 XThR.Tn[8] XThR.Tn[8].n7 161.363
R24177 XThR.Tn[8].n81 XThR.Tn[8].n80 161.3
R24178 XThR.Tn[8].n76 XThR.Tn[8].n75 161.3
R24179 XThR.Tn[8].n71 XThR.Tn[8].n70 161.3
R24180 XThR.Tn[8].n66 XThR.Tn[8].n65 161.3
R24181 XThR.Tn[8].n61 XThR.Tn[8].n60 161.3
R24182 XThR.Tn[8].n56 XThR.Tn[8].n55 161.3
R24183 XThR.Tn[8].n51 XThR.Tn[8].n50 161.3
R24184 XThR.Tn[8].n46 XThR.Tn[8].n45 161.3
R24185 XThR.Tn[8].n41 XThR.Tn[8].n40 161.3
R24186 XThR.Tn[8].n36 XThR.Tn[8].n35 161.3
R24187 XThR.Tn[8].n31 XThR.Tn[8].n30 161.3
R24188 XThR.Tn[8].n26 XThR.Tn[8].n25 161.3
R24189 XThR.Tn[8].n21 XThR.Tn[8].n20 161.3
R24190 XThR.Tn[8].n16 XThR.Tn[8].n15 161.3
R24191 XThR.Tn[8].n11 XThR.Tn[8].n10 161.3
R24192 XThR.Tn[8].n79 XThR.Tn[8].t23 161.106
R24193 XThR.Tn[8].n74 XThR.Tn[8].t29 161.106
R24194 XThR.Tn[8].n69 XThR.Tn[8].t71 161.106
R24195 XThR.Tn[8].n64 XThR.Tn[8].t57 161.106
R24196 XThR.Tn[8].n59 XThR.Tn[8].t21 161.106
R24197 XThR.Tn[8].n54 XThR.Tn[8].t46 161.106
R24198 XThR.Tn[8].n49 XThR.Tn[8].t27 161.106
R24199 XThR.Tn[8].n44 XThR.Tn[8].t69 161.106
R24200 XThR.Tn[8].n39 XThR.Tn[8].t56 161.106
R24201 XThR.Tn[8].n34 XThR.Tn[8].t61 161.106
R24202 XThR.Tn[8].n29 XThR.Tn[8].t44 161.106
R24203 XThR.Tn[8].n24 XThR.Tn[8].t70 161.106
R24204 XThR.Tn[8].n19 XThR.Tn[8].t43 161.106
R24205 XThR.Tn[8].n14 XThR.Tn[8].t26 161.106
R24206 XThR.Tn[8].n9 XThR.Tn[8].t49 161.106
R24207 XThR.Tn[8].n7 XThR.Tn[8].t33 161.106
R24208 XThR.Tn[8].n80 XThR.Tn[8].t19 159.978
R24209 XThR.Tn[8].n75 XThR.Tn[8].t25 159.978
R24210 XThR.Tn[8].n70 XThR.Tn[8].t67 159.978
R24211 XThR.Tn[8].n65 XThR.Tn[8].t54 159.978
R24212 XThR.Tn[8].n60 XThR.Tn[8].t16 159.978
R24213 XThR.Tn[8].n55 XThR.Tn[8].t42 159.978
R24214 XThR.Tn[8].n50 XThR.Tn[8].t24 159.978
R24215 XThR.Tn[8].n45 XThR.Tn[8].t64 159.978
R24216 XThR.Tn[8].n40 XThR.Tn[8].t51 159.978
R24217 XThR.Tn[8].n35 XThR.Tn[8].t58 159.978
R24218 XThR.Tn[8].n30 XThR.Tn[8].t41 159.978
R24219 XThR.Tn[8].n25 XThR.Tn[8].t66 159.978
R24220 XThR.Tn[8].n20 XThR.Tn[8].t40 159.978
R24221 XThR.Tn[8].n15 XThR.Tn[8].t22 159.978
R24222 XThR.Tn[8].n10 XThR.Tn[8].t45 159.978
R24223 XThR.Tn[8].n79 XThR.Tn[8].t73 145.038
R24224 XThR.Tn[8].n74 XThR.Tn[8].t35 145.038
R24225 XThR.Tn[8].n69 XThR.Tn[8].t15 145.038
R24226 XThR.Tn[8].n64 XThR.Tn[8].t62 145.038
R24227 XThR.Tn[8].n59 XThR.Tn[8].t30 145.038
R24228 XThR.Tn[8].n54 XThR.Tn[8].t72 145.038
R24229 XThR.Tn[8].n49 XThR.Tn[8].t17 145.038
R24230 XThR.Tn[8].n44 XThR.Tn[8].t63 145.038
R24231 XThR.Tn[8].n39 XThR.Tn[8].t60 145.038
R24232 XThR.Tn[8].n34 XThR.Tn[8].t28 145.038
R24233 XThR.Tn[8].n29 XThR.Tn[8].t52 145.038
R24234 XThR.Tn[8].n24 XThR.Tn[8].t12 145.038
R24235 XThR.Tn[8].n19 XThR.Tn[8].t50 145.038
R24236 XThR.Tn[8].n14 XThR.Tn[8].t34 145.038
R24237 XThR.Tn[8].n9 XThR.Tn[8].t59 145.038
R24238 XThR.Tn[8].n7 XThR.Tn[8].t39 145.038
R24239 XThR.Tn[8].n80 XThR.Tn[8].t32 143.911
R24240 XThR.Tn[8].n75 XThR.Tn[8].t55 143.911
R24241 XThR.Tn[8].n70 XThR.Tn[8].t37 143.911
R24242 XThR.Tn[8].n65 XThR.Tn[8].t18 143.911
R24243 XThR.Tn[8].n60 XThR.Tn[8].t48 143.911
R24244 XThR.Tn[8].n55 XThR.Tn[8].t31 143.911
R24245 XThR.Tn[8].n50 XThR.Tn[8].t38 143.911
R24246 XThR.Tn[8].n45 XThR.Tn[8].t20 143.911
R24247 XThR.Tn[8].n40 XThR.Tn[8].t14 143.911
R24248 XThR.Tn[8].n35 XThR.Tn[8].t47 143.911
R24249 XThR.Tn[8].n30 XThR.Tn[8].t68 143.911
R24250 XThR.Tn[8].n25 XThR.Tn[8].t36 143.911
R24251 XThR.Tn[8].n20 XThR.Tn[8].t65 143.911
R24252 XThR.Tn[8].n15 XThR.Tn[8].t53 143.911
R24253 XThR.Tn[8].n10 XThR.Tn[8].t13 143.911
R24254 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R24255 XThR.Tn[8].n3 XThR.Tn[8].t8 26.5955
R24256 XThR.Tn[8].n3 XThR.Tn[8].t10 26.5955
R24257 XThR.Tn[8].n4 XThR.Tn[8].t1 26.5955
R24258 XThR.Tn[8].n4 XThR.Tn[8].t9 26.5955
R24259 XThR.Tn[8].n0 XThR.Tn[8].t6 26.5955
R24260 XThR.Tn[8].n0 XThR.Tn[8].t4 26.5955
R24261 XThR.Tn[8].n1 XThR.Tn[8].t7 26.5955
R24262 XThR.Tn[8].n1 XThR.Tn[8].t5 26.5955
R24263 XThR.Tn[8].n86 XThR.Tn[8].t11 24.9236
R24264 XThR.Tn[8].n86 XThR.Tn[8].t3 24.9236
R24265 XThR.Tn[8].n87 XThR.Tn[8].t2 24.9236
R24266 XThR.Tn[8].n87 XThR.Tn[8].t0 24.9236
R24267 XThR.Tn[8] XThR.Tn[8].n88 18.8943
R24268 XThR.Tn[8].n6 XThR.Tn[8].n5 13.5534
R24269 XThR.Tn[8].n85 XThR.Tn[8] 7.82692
R24270 XThR.Tn[8] XThR.Tn[8].n85 6.34069
R24271 XThR.Tn[8] XThR.Tn[8].n8 5.34038
R24272 XThR.Tn[8].n13 XThR.Tn[8].n12 4.5005
R24273 XThR.Tn[8].n18 XThR.Tn[8].n17 4.5005
R24274 XThR.Tn[8].n23 XThR.Tn[8].n22 4.5005
R24275 XThR.Tn[8].n28 XThR.Tn[8].n27 4.5005
R24276 XThR.Tn[8].n33 XThR.Tn[8].n32 4.5005
R24277 XThR.Tn[8].n38 XThR.Tn[8].n37 4.5005
R24278 XThR.Tn[8].n43 XThR.Tn[8].n42 4.5005
R24279 XThR.Tn[8].n48 XThR.Tn[8].n47 4.5005
R24280 XThR.Tn[8].n53 XThR.Tn[8].n52 4.5005
R24281 XThR.Tn[8].n58 XThR.Tn[8].n57 4.5005
R24282 XThR.Tn[8].n63 XThR.Tn[8].n62 4.5005
R24283 XThR.Tn[8].n68 XThR.Tn[8].n67 4.5005
R24284 XThR.Tn[8].n73 XThR.Tn[8].n72 4.5005
R24285 XThR.Tn[8].n78 XThR.Tn[8].n77 4.5005
R24286 XThR.Tn[8].n83 XThR.Tn[8].n82 4.5005
R24287 XThR.Tn[8].n84 XThR.Tn[8] 3.70586
R24288 XThR.Tn[8].n13 XThR.Tn[8] 2.52282
R24289 XThR.Tn[8].n18 XThR.Tn[8] 2.52282
R24290 XThR.Tn[8].n23 XThR.Tn[8] 2.52282
R24291 XThR.Tn[8].n28 XThR.Tn[8] 2.52282
R24292 XThR.Tn[8].n33 XThR.Tn[8] 2.52282
R24293 XThR.Tn[8].n38 XThR.Tn[8] 2.52282
R24294 XThR.Tn[8].n43 XThR.Tn[8] 2.52282
R24295 XThR.Tn[8].n48 XThR.Tn[8] 2.52282
R24296 XThR.Tn[8].n53 XThR.Tn[8] 2.52282
R24297 XThR.Tn[8].n58 XThR.Tn[8] 2.52282
R24298 XThR.Tn[8].n63 XThR.Tn[8] 2.52282
R24299 XThR.Tn[8].n68 XThR.Tn[8] 2.52282
R24300 XThR.Tn[8].n73 XThR.Tn[8] 2.52282
R24301 XThR.Tn[8].n78 XThR.Tn[8] 2.52282
R24302 XThR.Tn[8].n83 XThR.Tn[8] 2.52282
R24303 XThR.Tn[8].n85 XThR.Tn[8] 1.79489
R24304 XThR.Tn[8].n6 XThR.Tn[8] 1.50638
R24305 XThR.Tn[8] XThR.Tn[8].n6 1.19676
R24306 XThR.Tn[8].n81 XThR.Tn[8] 1.08677
R24307 XThR.Tn[8].n76 XThR.Tn[8] 1.08677
R24308 XThR.Tn[8].n71 XThR.Tn[8] 1.08677
R24309 XThR.Tn[8].n66 XThR.Tn[8] 1.08677
R24310 XThR.Tn[8].n61 XThR.Tn[8] 1.08677
R24311 XThR.Tn[8].n56 XThR.Tn[8] 1.08677
R24312 XThR.Tn[8].n51 XThR.Tn[8] 1.08677
R24313 XThR.Tn[8].n46 XThR.Tn[8] 1.08677
R24314 XThR.Tn[8].n41 XThR.Tn[8] 1.08677
R24315 XThR.Tn[8].n36 XThR.Tn[8] 1.08677
R24316 XThR.Tn[8].n31 XThR.Tn[8] 1.08677
R24317 XThR.Tn[8].n26 XThR.Tn[8] 1.08677
R24318 XThR.Tn[8].n21 XThR.Tn[8] 1.08677
R24319 XThR.Tn[8].n16 XThR.Tn[8] 1.08677
R24320 XThR.Tn[8].n11 XThR.Tn[8] 1.08677
R24321 XThR.Tn[8] XThR.Tn[8].n13 0.839786
R24322 XThR.Tn[8] XThR.Tn[8].n18 0.839786
R24323 XThR.Tn[8] XThR.Tn[8].n23 0.839786
R24324 XThR.Tn[8] XThR.Tn[8].n28 0.839786
R24325 XThR.Tn[8] XThR.Tn[8].n33 0.839786
R24326 XThR.Tn[8] XThR.Tn[8].n38 0.839786
R24327 XThR.Tn[8] XThR.Tn[8].n43 0.839786
R24328 XThR.Tn[8] XThR.Tn[8].n48 0.839786
R24329 XThR.Tn[8] XThR.Tn[8].n53 0.839786
R24330 XThR.Tn[8] XThR.Tn[8].n58 0.839786
R24331 XThR.Tn[8] XThR.Tn[8].n63 0.839786
R24332 XThR.Tn[8] XThR.Tn[8].n68 0.839786
R24333 XThR.Tn[8] XThR.Tn[8].n73 0.839786
R24334 XThR.Tn[8] XThR.Tn[8].n78 0.839786
R24335 XThR.Tn[8] XThR.Tn[8].n83 0.839786
R24336 XThR.Tn[8].n8 XThR.Tn[8] 0.499542
R24337 XThR.Tn[8].n82 XThR.Tn[8] 0.063
R24338 XThR.Tn[8].n77 XThR.Tn[8] 0.063
R24339 XThR.Tn[8].n72 XThR.Tn[8] 0.063
R24340 XThR.Tn[8].n67 XThR.Tn[8] 0.063
R24341 XThR.Tn[8].n62 XThR.Tn[8] 0.063
R24342 XThR.Tn[8].n57 XThR.Tn[8] 0.063
R24343 XThR.Tn[8].n52 XThR.Tn[8] 0.063
R24344 XThR.Tn[8].n47 XThR.Tn[8] 0.063
R24345 XThR.Tn[8].n42 XThR.Tn[8] 0.063
R24346 XThR.Tn[8].n37 XThR.Tn[8] 0.063
R24347 XThR.Tn[8].n32 XThR.Tn[8] 0.063
R24348 XThR.Tn[8].n27 XThR.Tn[8] 0.063
R24349 XThR.Tn[8].n22 XThR.Tn[8] 0.063
R24350 XThR.Tn[8].n17 XThR.Tn[8] 0.063
R24351 XThR.Tn[8].n12 XThR.Tn[8] 0.063
R24352 XThR.Tn[8].n84 XThR.Tn[8] 0.0540714
R24353 XThR.Tn[8] XThR.Tn[8].n84 0.038
R24354 XThR.Tn[8].n8 XThR.Tn[8] 0.0143889
R24355 XThR.Tn[8].n82 XThR.Tn[8].n81 0.00771154
R24356 XThR.Tn[8].n77 XThR.Tn[8].n76 0.00771154
R24357 XThR.Tn[8].n72 XThR.Tn[8].n71 0.00771154
R24358 XThR.Tn[8].n67 XThR.Tn[8].n66 0.00771154
R24359 XThR.Tn[8].n62 XThR.Tn[8].n61 0.00771154
R24360 XThR.Tn[8].n57 XThR.Tn[8].n56 0.00771154
R24361 XThR.Tn[8].n52 XThR.Tn[8].n51 0.00771154
R24362 XThR.Tn[8].n47 XThR.Tn[8].n46 0.00771154
R24363 XThR.Tn[8].n42 XThR.Tn[8].n41 0.00771154
R24364 XThR.Tn[8].n37 XThR.Tn[8].n36 0.00771154
R24365 XThR.Tn[8].n32 XThR.Tn[8].n31 0.00771154
R24366 XThR.Tn[8].n27 XThR.Tn[8].n26 0.00771154
R24367 XThR.Tn[8].n22 XThR.Tn[8].n21 0.00771154
R24368 XThR.Tn[8].n17 XThR.Tn[8].n16 0.00771154
R24369 XThR.Tn[8].n12 XThR.Tn[8].n11 0.00771154
R24370 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R24371 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R24372 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R24373 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R24374 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R24375 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R24376 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R24377 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R24378 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R24379 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R24380 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R24381 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R24382 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R24383 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R24384 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R24385 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R24386 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R24387 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R24388 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R24389 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R24390 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R24391 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R24392 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R24393 XThC.XTB3.Y.n0 XThC.XTB3.Y.t2 132.067
R24394 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R24395 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R24396 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R24397 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R24398 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R24399 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R24400 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R24401 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R24402 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R24403 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R24404 XThC.XTB3.Y.n2 XThC.XTB3.Y.t1 26.5955
R24405 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R24406 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R24407 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R24408 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R24409 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R24410 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R24411 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R24412 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R24413 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R24414 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R24415 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R24416 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R24417 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R24418 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R24419 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R24420 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R24421 data[4].n3 data[4].t0 231.835
R24422 data[4].n0 data[4].t3 230.155
R24423 data[4].n0 data[4].t1 157.856
R24424 data[4].n3 data[4].t2 157.07
R24425 data[4].n1 data[4].n0 152
R24426 data[4].n4 data[4].n3 152
R24427 data[4].n2 data[4].n1 25.6681
R24428 data[4].n4 data[4].n2 10.7642
R24429 data[4].n2 data[4] 2.763
R24430 data[4].n1 data[4] 2.10199
R24431 data[4] data[4].n4 2.01193
R24432 XThR.Tn[13].n87 XThR.Tn[13].n86 256.103
R24433 XThR.Tn[13].n2 XThR.Tn[13].n0 243.68
R24434 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R24435 XThR.Tn[13].n2 XThR.Tn[13].n1 205.28
R24436 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R24437 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R24438 XThR.Tn[13] XThR.Tn[13].n78 161.363
R24439 XThR.Tn[13] XThR.Tn[13].n73 161.363
R24440 XThR.Tn[13] XThR.Tn[13].n68 161.363
R24441 XThR.Tn[13] XThR.Tn[13].n63 161.363
R24442 XThR.Tn[13] XThR.Tn[13].n58 161.363
R24443 XThR.Tn[13] XThR.Tn[13].n53 161.363
R24444 XThR.Tn[13] XThR.Tn[13].n48 161.363
R24445 XThR.Tn[13] XThR.Tn[13].n43 161.363
R24446 XThR.Tn[13] XThR.Tn[13].n38 161.363
R24447 XThR.Tn[13] XThR.Tn[13].n33 161.363
R24448 XThR.Tn[13] XThR.Tn[13].n28 161.363
R24449 XThR.Tn[13] XThR.Tn[13].n23 161.363
R24450 XThR.Tn[13] XThR.Tn[13].n18 161.363
R24451 XThR.Tn[13] XThR.Tn[13].n13 161.363
R24452 XThR.Tn[13] XThR.Tn[13].n8 161.363
R24453 XThR.Tn[13] XThR.Tn[13].n6 161.363
R24454 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R24455 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R24456 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R24457 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R24458 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R24459 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R24460 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R24461 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R24462 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R24463 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R24464 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R24465 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R24466 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R24467 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R24468 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R24469 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R24470 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R24471 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R24472 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R24473 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R24474 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R24475 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R24476 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R24477 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R24478 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R24479 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R24480 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R24481 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R24482 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R24483 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R24484 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R24485 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R24486 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R24487 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R24488 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R24489 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R24490 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R24491 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R24492 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R24493 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R24494 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R24495 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R24496 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R24497 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R24498 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R24499 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R24500 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R24501 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R24502 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R24503 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R24504 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R24505 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R24506 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R24507 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R24508 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R24509 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R24510 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R24511 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R24512 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R24513 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R24514 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R24515 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R24516 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R24517 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R24518 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R24519 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R24520 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R24521 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R24522 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R24523 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R24524 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R24525 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R24526 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R24527 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R24528 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R24529 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R24530 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R24531 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R24532 XThR.Tn[13].n85 XThR.Tn[13].t2 26.5955
R24533 XThR.Tn[13].n85 XThR.Tn[13].t0 26.5955
R24534 XThR.Tn[13].n0 XThR.Tn[13].t9 26.5955
R24535 XThR.Tn[13].n0 XThR.Tn[13].t11 26.5955
R24536 XThR.Tn[13].n1 XThR.Tn[13].t10 26.5955
R24537 XThR.Tn[13].n1 XThR.Tn[13].t8 26.5955
R24538 XThR.Tn[13].n86 XThR.Tn[13].t3 26.5955
R24539 XThR.Tn[13].n86 XThR.Tn[13].t1 26.5955
R24540 XThR.Tn[13].n4 XThR.Tn[13].t6 24.9236
R24541 XThR.Tn[13].n4 XThR.Tn[13].t4 24.9236
R24542 XThR.Tn[13].n3 XThR.Tn[13].t7 24.9236
R24543 XThR.Tn[13].n3 XThR.Tn[13].t5 24.9236
R24544 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R24545 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R24546 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R24547 XThR.Tn[13] XThR.Tn[13].n7 5.34038
R24548 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R24549 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R24550 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R24551 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R24552 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R24553 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R24554 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R24555 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R24556 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R24557 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R24558 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R24559 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R24560 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R24561 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R24562 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R24563 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R24564 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R24565 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R24566 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R24567 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R24568 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R24569 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R24570 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R24571 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R24572 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R24573 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R24574 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R24575 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R24576 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R24577 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R24578 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R24579 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R24580 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R24581 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R24582 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R24583 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R24584 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R24585 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R24586 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R24587 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R24588 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R24589 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R24590 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R24591 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R24592 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R24593 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R24594 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R24595 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R24596 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R24597 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R24598 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R24599 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R24600 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R24601 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R24602 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R24603 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R24604 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R24605 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R24606 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R24607 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R24608 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R24609 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R24610 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R24611 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R24612 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R24613 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R24614 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R24615 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R24616 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R24617 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R24618 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R24619 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R24620 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R24621 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R24622 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R24623 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R24624 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R24625 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R24626 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R24627 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R24628 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R24629 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R24630 XThR.Tn[13] XThR.Tn[13].n83 0.038
R24631 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R24632 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R24633 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R24634 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R24635 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R24636 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R24637 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R24638 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R24639 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R24640 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R24641 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R24642 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R24643 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R24644 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R24645 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R24646 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R24647 data[0].n1 data[0].t0 230.155
R24648 data[0].n0 data[0].t2 228.463
R24649 data[0].n1 data[0].t1 157.856
R24650 data[0].n0 data[0].t3 157.07
R24651 data[0].n2 data[0].n1 152.768
R24652 data[0].n4 data[0].n0 152.256
R24653 data[0].n3 data[0].n2 24.1398
R24654 data[0].n4 data[0].n3 9.48418
R24655 data[0] data[0].n4 6.1445
R24656 data[0].n2 data[0] 5.6325
R24657 data[0].n3 data[0] 2.638
R24658 XThR.XTB4.Y XThR.XTB4.Y.t0 230.518
R24659 XThR.XTB4.Y.n10 XThR.XTB4.Y.t12 212.081
R24660 XThR.XTB4.Y.n11 XThR.XTB4.Y.t2 212.081
R24661 XThR.XTB4.Y.n16 XThR.XTB4.Y.t7 212.081
R24662 XThR.XTB4.Y.n17 XThR.XTB4.Y.t6 212.081
R24663 XThR.XTB4.Y.n0 XThR.XTB4.Y.t17 212.081
R24664 XThR.XTB4.Y.n1 XThR.XTB4.Y.t5 212.081
R24665 XThR.XTB4.Y.n3 XThR.XTB4.Y.t15 212.081
R24666 XThR.XTB4.Y.n4 XThR.XTB4.Y.t4 212.081
R24667 XThR.XTB4.Y.n13 XThR.XTB4.Y.n12 173.761
R24668 XThR.XTB4.Y.n2 XThR.XTB4.Y 167.361
R24669 XThR.XTB4.Y.n19 XThR.XTB4.Y.n18 152
R24670 XThR.XTB4.Y.n15 XThR.XTB4.Y.n14 152
R24671 XThR.XTB4.Y.n13 XThR.XTB4.Y.n9 152
R24672 XThR.XTB4.Y.n6 XThR.XTB4.Y.n5 152
R24673 XThR.XTB4.Y.n10 XThR.XTB4.Y.t3 139.78
R24674 XThR.XTB4.Y.n11 XThR.XTB4.Y.t9 139.78
R24675 XThR.XTB4.Y.n16 XThR.XTB4.Y.t14 139.78
R24676 XThR.XTB4.Y.n17 XThR.XTB4.Y.t11 139.78
R24677 XThR.XTB4.Y.n0 XThR.XTB4.Y.t10 139.78
R24678 XThR.XTB4.Y.n1 XThR.XTB4.Y.t16 139.78
R24679 XThR.XTB4.Y.n3 XThR.XTB4.Y.t8 139.78
R24680 XThR.XTB4.Y.n4 XThR.XTB4.Y.t13 139.78
R24681 XThR.XTB4.Y.n21 XThR.XTB4.Y.t1 133.386
R24682 XThR.XTB4.Y.n20 XThR.XTB4.Y.n19 72.9296
R24683 XThR.XTB4.Y.n1 XThR.XTB4.Y.n0 61.346
R24684 XThR.XTB4.Y.n15 XThR.XTB4.Y.n9 49.6611
R24685 XThR.XTB4.Y.n18 XThR.XTB4.Y.n16 45.2793
R24686 XThR.XTB4.Y.n12 XThR.XTB4.Y.n11 42.3581
R24687 XThR.XTB4.Y.n20 XThR.XTB4.Y.n8 38.1854
R24688 XThR.XTB4.Y.n2 XThR.XTB4.Y.n1 30.6732
R24689 XThR.XTB4.Y.n3 XThR.XTB4.Y.n2 30.6732
R24690 XThR.XTB4.Y.n5 XThR.XTB4.Y.n3 30.6732
R24691 XThR.XTB4.Y.n5 XThR.XTB4.Y.n4 30.6732
R24692 XThR.XTB4.Y XThR.XTB4.Y.n21 28.966
R24693 XThR.XTB4.Y.n14 XThR.XTB4.Y.n13 21.7605
R24694 XThR.XTB4.Y.n14 XThR.XTB4.Y 21.1205
R24695 XThR.XTB4.Y.n12 XThR.XTB4.Y.n10 18.9884
R24696 XThR.XTB4.Y.n18 XThR.XTB4.Y.n17 16.0672
R24697 XThR.XTB4.Y.n21 XThR.XTB4.Y.n20 11.994
R24698 XThR.XTB4.Y.n22 XThR.XTB4.Y 11.6875
R24699 XThR.XTB4.Y.n8 XThR.XTB4.Y.n7 8.21182
R24700 XThR.XTB4.Y.n11 XThR.XTB4.Y.n9 7.30353
R24701 XThR.XTB4.Y.n8 XThR.XTB4.Y.n6 7.24578
R24702 XThR.XTB4.Y.n22 XThR.XTB4.Y 7.23528
R24703 XThR.XTB4.Y.n6 XThR.XTB4.Y 6.08654
R24704 XThR.XTB4.Y XThR.XTB4.Y.n22 5.04292
R24705 XThR.XTB4.Y.n16 XThR.XTB4.Y.n15 4.38232
R24706 XThR.XTB4.Y.n7 XThR.XTB4.Y 1.79489
R24707 XThR.XTB4.Y.n7 XThR.XTB4.Y 0.966538
R24708 XThR.XTB4.Y.n19 XThR.XTB4.Y 0.6405
R24709 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R24710 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R24711 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R24712 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R24713 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R24714 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R24715 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R24716 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R24717 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24718 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24719 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24720 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24721 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24722 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24723 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24724 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24725 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24726 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24727 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24728 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24729 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24730 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24731 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24732 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24733 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24734 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24735 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24736 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24737 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24738 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24739 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24740 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24741 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24742 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24743 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24744 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24745 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24746 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24747 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24748 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24749 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24750 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24751 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24752 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24753 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24754 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24755 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24756 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24757 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24758 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24759 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24760 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24761 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R24762 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R24763 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R24764 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R24765 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R24766 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R24767 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R24768 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R24769 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R24770 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R24771 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R24772 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R24773 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R24774 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R24775 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R24776 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R24777 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R24778 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R24779 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R24780 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R24781 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R24782 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R24783 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R24784 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R24785 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R24786 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R24787 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R24788 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R24789 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R24790 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R24791 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R24792 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R24793 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R24794 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R24795 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R24796 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R24797 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R24798 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R24799 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R24800 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R24801 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R24802 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R24803 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R24804 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R24805 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R24806 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R24807 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R24808 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R24809 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R24810 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R24811 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R24812 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R24813 data[6].n0 data[6].t0 230.576
R24814 data[6].n0 data[6].t1 158.275
R24815 data[6].n1 data[6].n0 152
R24816 data[6].n1 data[6] 11.9995
R24817 data[6] data[6].n1 6.66717
R24818 data[1].n4 data[1].t2 230.576
R24819 data[1].n1 data[1].t0 230.363
R24820 data[1].n0 data[1].t4 229.369
R24821 data[1].n4 data[1].t5 158.275
R24822 data[1].n1 data[1].t3 158.064
R24823 data[1].n0 data[1].t1 157.07
R24824 data[1].n2 data[1].n1 153.28
R24825 data[1].n7 data[1].n0 153.147
R24826 data[1].n5 data[1].n4 152
R24827 data[1].n7 data[1].n6 16.3874
R24828 data[1].n6 data[1].n5 14.9641
R24829 data[1].n3 data[1].n2 9.3005
R24830 data[1].n6 data[1].n3 6.49639
R24831 data[1] data[1].n7 3.24826
R24832 data[1].n2 data[1] 2.92621
R24833 data[1].n3 data[1] 2.15819
R24834 data[1].n5 data[1] 2.13383
R24835 data[2].n0 data[2].t0 230.576
R24836 data[2].n0 data[2].t1 158.275
R24837 data[2].n1 data[2].n0 152
R24838 data[2].n1 data[2] 12.7714
R24839 data[2] data[2].n1 2.13383
R24840 data[5].n4 data[5].t2 230.576
R24841 data[5].n1 data[5].t0 230.363
R24842 data[5].n0 data[5].t1 229.369
R24843 data[5].n4 data[5].t5 158.275
R24844 data[5].n1 data[5].t3 158.064
R24845 data[5].n0 data[5].t4 157.07
R24846 data[5].n2 data[5].n1 152.256
R24847 data[5].n7 data[5].n0 152.238
R24848 data[5].n5 data[5].n4 152
R24849 data[5].n7 data[5].n6 16.3874
R24850 data[5].n6 data[5].n5 14.6005
R24851 data[5].n3 data[5].n2 9.3005
R24852 data[5].n5 data[5] 6.66717
R24853 data[5].n6 data[5].n3 6.49639
R24854 data[5].n2 data[5] 6.1445
R24855 data[5] data[5].n7 5.68939
R24856 data[5].n3 data[5] 2.28319
R24857 data[3].n0 data[3].t1 230.576
R24858 data[3].n0 data[3].t0 158.275
R24859 data[3].n1 data[3].n0 153.553
R24860 data[3].n1 data[3] 11.6078
R24861 data[3] data[3].n1 2.90959
R24862 data[7].n0 data[7].t0 230.576
R24863 data[7].n0 data[7].t1 158.275
R24864 data[7].n1 data[7].n0 152
R24865 data[7].n1 data[7] 11.9995
R24866 data[7] data[7].n1 6.66717
R24867 bias[1] bias[1].t0 23.8076
R24868 bias[2] bias[2].t0 57.7456
R24869 bias[0] bias[0].t0 12.1467
C0 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.03425f
C1 XA.XIR[6].XIC[10].icell.Ien VPWR 0.1903f
C2 a_7331_10587# data[0] 0.00451f
C3 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.15202f
C4 XA.XIR[3].XIC[1].icell.SM Iout 0.00388f
C5 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PUM 0.00465f
C6 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PDM 0.0059f
C7 XA.XIR[13].XIC[13].icell.PDM VPWR 0.00799f
C8 XA.XIR[5].XIC[13].icell.PUM VPWR 0.00937f
C9 XThR.Tn[4] XA.XIR[5].XIC[1].icell.Ien 0.00338f
C10 XA.XIR[6].XIC[6].icell.Ien Iout 0.06417f
C11 XA.XIR[8].XIC[3].icell.PUM Vbias 0.0031f
C12 XA.XIR[4].XIC[1].icell.PDM VPWR 0.00799f
C13 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7] 0.00341f
C14 XThR.XTBN.Y XA.XIR[14].XIC_dummy_left.icell.Iout 0.00116f
C15 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.SM 0.0039f
C16 XA.XIR[15].XIC[7].icell.SM Iout 0.00388f
C17 XA.XIR[15].XIC_dummy_right.icell.Ien Vbias 0.00288f
C18 XThR.Tn[3] XA.XIR[4].XIC[1].icell.Ien 0.00338f
C19 XA.XIR[3].XIC[9].icell.PDM VPWR 0.00799f
C20 XA.XIR[4].XIC[14].icell.SM VPWR 0.00207f
C21 XA.XIR[8].XIC[11].icell.PDM VPWR 0.00799f
C22 XA.XIR[14].XIC[4].icell.Ien VPWR 0.19084f
C23 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C24 XA.XIR[0].XIC[12].icell.PDM Vbias 0.04282f
C25 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00584f
C26 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13] 0.00341f
C27 XA.XIR[11].XIC[2].icell.SM Vbias 0.00701f
C28 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PUM 0.00465f
C29 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07214f
C30 XA.XIR[4].XIC[10].icell.SM Iout 0.00388f
C31 XThC.XTBN.A a_8739_9569# 0.01719f
C32 XA.XIR[13].XIC[14].icell.Ien Vbias 0.21098f
C33 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C34 XA.XIR[13].XIC[6].icell.Ien VPWR 0.1903f
C35 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.04036f
C36 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.0353f
C37 XA.XIR[9].XIC[12].icell.PUM Vbias 0.0031f
C38 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04031f
C39 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C40 XA.XIR[8].XIC[8].icell.SM VPWR 0.00158f
C41 XA.XIR[10].XIC[4].icell.SM Vbias 0.00701f
C42 XA.XIR[2].XIC[3].icell.PDM Iout 0.00117f
C43 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01577f
C44 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00584f
C45 XA.XIR[12].XIC[8].icell.PUM VPWR 0.00937f
C46 XA.XIR[13].XIC[2].icell.Ien Iout 0.06417f
C47 XThC.Tn[4] XThR.Tn[2] 0.28739f
C48 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C49 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12] 0.00341f
C50 XA.XIR[8].XIC[4].icell.SM Iout 0.00388f
C51 XA.XIR[0].XIC[5].icell.PUM Vbias 0.0031f
C52 XThR.Tn[8] XA.XIR[9].XIC[4].icell.SM 0.00121f
C53 XThR.XTB6.Y XThR.Tn[14] 0.00128f
C54 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C55 XThR.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.00353f
C56 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00584f
C57 XA.XIR[11].XIC[9].icell.Ien VPWR 0.1903f
C58 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.SM 0.00168f
C59 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.SM 0.0039f
C60 XA.XIR[3].XIC[13].icell.SM Vbias 0.00701f
C61 XThC.Tn[13] XThR.Tn[14] 0.2874f
C62 XThR.Tn[4] XA.XIR[5].XIC[6].icell.Ien 0.00338f
C63 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C64 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.SM 0.00168f
C65 XA.XIR[11].XIC[5].icell.Ien Iout 0.06417f
C66 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00214f
C67 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C68 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C69 XThR.Tn[3] XA.XIR[4].XIC[6].icell.Ien 0.00338f
C70 XA.XIR[9].XIC[13].icell.SM Iout 0.00388f
C71 XA.XIR[2].XIC[6].icell.SM Vbias 0.00701f
C72 XA.XIR[7].XIC[8].icell.PUM Vbias 0.0031f
C73 XA.XIR[10].XIC[7].icell.Ien Iout 0.06417f
C74 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C75 a_7875_9569# XThC.Tn[9] 0.19329f
C76 XA.XIR[0].XIC[10].icell.SM VPWR 0.00158f
C77 XThR.Tn[9] XA.XIR[10].XIC[7].icell.Ien 0.00338f
C78 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.SM 0.00168f
C79 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5] 0.00341f
C80 XThC.XTB6.A XThC.Tn[5] 0.00363f
C81 XA.XIR[1].XIC[8].icell.SM Vbias 0.00704f
C82 XA.XIR[0].XIC[6].icell.SM Iout 0.00367f
C83 XThC.XTB2.Y XThC.Tn[9] 0.292f
C84 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.SM 0.0039f
C85 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C86 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.04036f
C87 XA.XIR[10].XIC[10].icell.Ien Vbias 0.21098f
C88 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C89 XA.XIR[2].XIC[0].icell.PUM VPWR 0.00937f
C90 XThR.XTB3.Y XThR.Tn[6] 0.00298f
C91 XA.XIR[3].XIC_dummy_right.icell.SM VPWR 0.00123f
C92 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PUM 0.00465f
C93 XThR.Tn[13] XA.XIR[14].XIC[1].icell.SM 0.00121f
C94 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8] 0.00341f
C95 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04031f
C96 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C97 XA.XIR[2].XIC[13].icell.Ien VPWR 0.1903f
C98 XA.XIR[11].XIC_15.icell.SM Iout 0.0047f
C99 XThR.XTB1.Y XThR.Tn[1] 0.0099f
C100 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PUM 0.00465f
C101 XA.XIR[7].XIC[13].icell.SM VPWR 0.00158f
C102 XThR.XTBN.Y XThR.Tn[9] 0.48048f
C103 XThC.Tn[0] XThR.Tn[6] 0.28741f
C104 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02762f
C105 XA.XIR[1].XIC[1].icell.PUM VPWR 0.00937f
C106 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.SM 0.00168f
C107 XA.XIR[13].XIC[11].icell.PUM Vbias 0.0031f
C108 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6] 0.00341f
C109 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C110 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PUM 0.00465f
C111 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.SM 0.0039f
C112 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C113 XA.XIR[2].XIC[9].icell.Ien Iout 0.06417f
C114 XA.XIR[1].XIC_15.icell.Ien VPWR 0.25566f
C115 XA.XIR[7].XIC[9].icell.SM Iout 0.00388f
C116 XThR.Tn[0] XA.XIR[1].XIC[4].icell.SM 0.00121f
C117 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.15202f
C118 XA.XIR[11].XIC[10].icell.SM VPWR 0.00158f
C119 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.15202f
C120 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C121 XThC.XTBN.A XThC.Tn[11] 0.12129f
C122 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PUM 0.00465f
C123 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02774f
C124 XThR.XTB5.Y a_n1049_5317# 0.00907f
C125 XThR.Tn[12] XA.XIR[13].XIC[5].icell.Ien 0.00338f
C126 XA.XIR[4].XIC[1].icell.PUM VPWR 0.00937f
C127 XA.XIR[1].XIC[11].icell.Ien Iout 0.06417f
C128 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C129 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.SM 0.00168f
C130 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Ien 0.00584f
C131 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PUM 0.00465f
C132 XThC.Tn[2] XThR.Tn[11] 0.28739f
C133 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C134 XA.XIR[13].XIC[0].icell.SM VPWR 0.00158f
C135 XThR.Tn[7] XA.XIR[8].XIC[10].icell.SM 0.00121f
C136 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02762f
C137 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C138 XThC.XTBN.Y a_4067_9615# 0.08456f
C139 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11] 0.00341f
C140 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C141 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.SM 0.0039f
C142 XThC.Tn[0] Vbias 1.91132f
C143 XThR.Tn[5] XA.XIR[6].XIC[6].icell.SM 0.00121f
C144 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PUM 0.00465f
C145 XThR.Tn[11] XA.XIR[12].XIC[8].icell.Ien 0.00338f
C146 XA.XIR[6].XIC[3].icell.PDM Vbias 0.04261f
C147 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C148 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[0].icell.SM 0.0039f
C149 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.SM 0.0039f
C150 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Iout 0.00347f
C151 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.15202f
C152 XA.XIR[5].XIC[10].icell.PDM Vbias 0.04261f
C153 XA.XIR[14].XIC[0].icell.PDM Vbias 0.04207f
C154 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C155 XA.XIR[15].XIC[3].icell.PUM VPWR 0.00937f
C156 XA.XIR[5].XIC[3].icell.Ien VPWR 0.1903f
C157 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07214f
C158 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C159 XThC.XTB3.Y a_8739_9569# 0.07285f
C160 XA.XIR[13].XIC[4].icell.PDM Vbias 0.04261f
C161 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C162 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02762f
C163 XA.XIR[13].XIC[12].icell.Ien Vbias 0.21098f
C164 XThC.XTB6.Y XThC.Tn[7] 0.01462f
C165 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.SM 0.0039f
C166 XA.XIR[4].XIC[6].icell.PUM VPWR 0.00937f
C167 XA.XIR[7].XIC[3].icell.PDM Iout 0.00117f
C168 XThR.Tn[10] Iout 1.16231f
C169 XThR.Tn[1] XA.XIR[2].XIC[12].icell.Ien 0.00338f
C170 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.SM 0.0039f
C171 XThR.Tn[9] XThR.Tn[10] 0.07779f
C172 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C173 XA.XIR[12].XIC[9].icell.PDM Vbias 0.04261f
C174 XA.XIR[11].XIC[13].icell.PUM VPWR 0.00937f
C175 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00214f
C176 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.15202f
C177 XA.XIR[15].XIC[1].icell.PDM Iout 0.00117f
C178 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.03535f
C179 XThC.Tn[5] XThR.Tn[1] 0.2874f
C180 XA.XIR[6].XIC[10].icell.PDM Iout 0.00117f
C181 XA.XIR[10].XIC[11].icell.PDM VPWR 0.00799f
C182 XThR.XTB5.Y data[7] 0.00931f
C183 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00584f
C184 XA.XIR[9].XIC[2].icell.Ien Vbias 0.21098f
C185 XThC.Tn[9] Iout 0.83793f
C186 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.SM 0.00168f
C187 XThC.Tn[9] XThR.Tn[9] 0.28739f
C188 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00584f
C189 XA.XIR[14].XIC[7].icell.PDM Iout 0.00117f
C190 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00256f
C191 XA.XIR[14].XIC[12].icell.SM VPWR 0.00158f
C192 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C193 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00584f
C194 XThC.Tn[5] XThR.Tn[12] 0.28739f
C195 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.03425f
C196 XA.XIR[9].XIC[11].icell.PDM VPWR 0.00799f
C197 XA.XIR[13].XIC[12].icell.PDM VPWR 0.00799f
C198 XThC.Tn[14] XThR.Tn[8] 0.28745f
C199 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00584f
C200 XA.XIR[0].XIC[3].icell.PDM VPWR 0.00774f
C201 XThR.XTB3.Y XThR.Tn[4] 0.00382f
C202 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PUM 0.00465f
C203 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.SM 0.00168f
C204 XThC.XTBN.A data[0] 0.02545f
C205 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C206 XA.XIR[3].XIC[5].icell.PUM Vbias 0.0031f
C207 XThC.XTB6.Y a_5949_10571# 0.01283f
C208 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00584f
C209 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C210 XA.XIR[1].XIC[0].icell.SM VPWR 0.00158f
C211 XThR.XTB3.Y a_n1049_7493# 0.23056f
C212 XA.XIR[6].XIC[8].icell.SM Vbias 0.00701f
C213 XA.XIR[9].XIC[9].icell.PUM VPWR 0.00937f
C214 XThC.Tn[0] XThR.Tn[4] 0.28743f
C215 XA.XIR[10].XIC[1].icell.SM VPWR 0.00158f
C216 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C217 XThC.XTBN.Y XThC.Tn[3] 0.62681f
C218 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C219 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C220 XThR.XTBN.A VPWR 0.90694f
C221 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02762f
C222 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C223 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02762f
C224 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.SM 0.0039f
C225 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.PDM 0.0059f
C226 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00584f
C227 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.15202f
C228 XA.XIR[5].XIC[11].icell.Ien Vbias 0.21098f
C229 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C230 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.SM 0.00168f
C231 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.03425f
C232 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00214f
C233 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.SM 0.00168f
C234 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04031f
C235 XThR.XTB5.Y a_n1049_6405# 0.24821f
C236 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04038f
C237 XA.XIR[11].XIC[14].icell.Ien VPWR 0.19036f
C238 XA.XIR[3].XIC[5].icell.PDM Vbias 0.04261f
C239 XThR.Tn[6] VPWR 6.58002f
C240 XA.XIR[4].XIC[14].icell.PUM Vbias 0.0031f
C241 XA.XIR[3].XIC[10].icell.SM VPWR 0.00158f
C242 XA.XIR[8].XIC[7].icell.PDM Vbias 0.04261f
C243 XA.XIR[14].XIC[2].icell.SM Vbias 0.00701f
C244 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C245 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10] 0.00341f
C246 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C247 XThC.XTB4.Y XThC.Tn[7] 0.01797f
C248 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01721f
C249 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C250 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02762f
C251 XA.XIR[6].XIC_15.icell.Ien VPWR 0.25566f
C252 XThC.Tn[4] XThR.Tn[10] 0.28739f
C253 XA.XIR[2].XIC[11].icell.PDM Vbias 0.04261f
C254 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14] 0.00341f
C255 XA.XIR[3].XIC[6].icell.SM Iout 0.00388f
C256 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02762f
C257 XA.XIR[13].XIC[4].icell.SM Vbias 0.00701f
C258 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C259 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.15202f
C260 XA.XIR[1].XIC[4].icell.PDM Iout 0.00117f
C261 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[5].icell.SM 0.0039f
C262 XA.XIR[6].XIC[11].icell.Ien Iout 0.06417f
C263 XA.XIR[7].XIC[5].icell.PUM VPWR 0.00937f
C264 XA.XIR[2].XIC[3].icell.SM VPWR 0.00158f
C265 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01577f
C266 XA.XIR[8].XIC[8].icell.PUM Vbias 0.0031f
C267 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C268 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.03023f
C269 XA.XIR[12].XIC[6].icell.Ien Vbias 0.21098f
C270 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C271 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PUM 0.00465f
C272 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.SM 0.0039f
C273 XA.XIR[1].XIC[5].icell.SM VPWR 0.00158f
C274 XA.XIR[4].XIC[4].icell.PDM Iout 0.00117f
C275 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00214f
C276 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.SM 0.0039f
C277 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C278 XA.XIR[14].XIC[9].icell.Ien VPWR 0.19084f
C279 XA.XIR[10].XIC_15.icell.Ien Vbias 0.21234f
C280 VPWR Vbias 0.2164p
C281 XA.XIR[11].XIC[7].icell.SM Vbias 0.00701f
C282 XA.XIR[3].XIC[12].icell.PDM Iout 0.00117f
C283 a_4861_9615# XThC.Tn[3] 0.27012f
C284 XA.XIR[1].XIC[1].icell.SM Iout 0.00388f
C285 XA.XIR[8].XIC[14].icell.PDM Iout 0.00117f
C286 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C287 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PDM 0.00172f
C288 XA.XIR[14].XIC[5].icell.Ien Iout 0.06417f
C289 XThC.Tn[0] XA.XIR[10].XIC_dummy_left.icell.Iout 0.00109f
C290 XA.XIR[8].XIC[13].icell.SM VPWR 0.00158f
C291 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.389f
C292 XA.XIR[13].XIC[7].icell.Ien Iout 0.06417f
C293 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C294 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.15202f
C295 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.SM 0.00168f
C296 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C297 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00256f
C298 XA.XIR[8].XIC[9].icell.SM Iout 0.00388f
C299 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C300 XThR.Tn[8] XA.XIR[9].XIC[9].icell.SM 0.00121f
C301 XA.XIR[0].XIC[10].icell.PUM Vbias 0.0031f
C302 XThR.Tn[0] XA.XIR[0].XIC_15.icell.PDM 0.00341f
C303 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C304 XThR.Tn[2] XA.XIR[3].XIC[4].icell.Ien 0.00338f
C305 XA.XIR[13].XIC[10].icell.Ien Vbias 0.21098f
C306 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C307 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.SM 0.0039f
C308 XThR.Tn[4] XA.XIR[5].XIC[11].icell.Ien 0.00338f
C309 XThR.Tn[1] XA.XIR[1].XIC[13].icell.PDM 0.00341f
C310 XA.XIR[11].XIC[11].icell.PUM VPWR 0.00937f
C311 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04031f
C312 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C313 XA.XIR[14].XIC_15.icell.SM Iout 0.0047f
C314 XThR.Tn[3] XA.XIR[4].XIC[11].icell.Ien 0.00338f
C315 XA.XIR[2].XIC[11].icell.SM Vbias 0.00701f
C316 a_7331_10587# VPWR 0.0063f
C317 XA.XIR[7].XIC[13].icell.PUM Vbias 0.0031f
C318 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00584f
C319 XThR.Tn[1] XA.XIR[2].XIC[2].icell.SM 0.00121f
C320 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02762f
C321 XA.XIR[14].XIC[10].icell.SM VPWR 0.00158f
C322 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04031f
C323 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C324 XA.XIR[1].XIC[13].icell.SM Vbias 0.00704f
C325 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11] 0.00341f
C326 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00584f
C327 XA.XIR[0].XIC[11].icell.SM Iout 0.00367f
C328 XA.XIR[5].XIC[1].icell.PDM VPWR 0.00799f
C329 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02762f
C330 XThR.Tn[2] XA.XIR[2].XIC[10].icell.PDM 0.00341f
C331 XThC.Tn[2] XThR.Tn[14] 0.28739f
C332 XThC.XTB3.Y data[0] 0.03253f
C333 XA.XIR[6].XIC[0].icell.SM VPWR 0.00158f
C334 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04031f
C335 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.03425f
C336 XThR.Tn[13] XA.XIR[14].XIC[6].icell.SM 0.00121f
C337 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[13].icell.Ien 0.00214f
C338 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00584f
C339 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02762f
C340 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.SM 0.00168f
C341 XA.XIR[3].XIC[2].icell.PUM Vbias 0.0031f
C342 XThR.Tn[4] VPWR 6.61651f
C343 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C344 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.03425f
C345 XA.XIR[2].XIC[14].icell.Ien Iout 0.06417f
C346 XA.XIR[12].XIC[0].icell.PDM VPWR 0.00799f
C347 XA.XIR[12].XIC[0].icell.SM Vbias 0.00675f
C348 XA.XIR[7].XIC[14].icell.SM Iout 0.00388f
C349 XThR.Tn[0] XA.XIR[1].XIC[9].icell.SM 0.00121f
C350 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00214f
C351 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C352 a_n1049_7493# VPWR 0.72084f
C353 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C354 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PUM 0.00465f
C355 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C356 XA.XIR[11].XIC[6].icell.PDM VPWR 0.00799f
C357 XA.XIR[1].XIC_dummy_right.icell.SM VPWR 0.00123f
C358 XA.XIR[11].XIC[12].icell.Ien VPWR 0.1903f
C359 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C360 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00584f
C361 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02762f
C362 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C363 XA.XIR[14].XIC[0].icell.Ien Iout 0.06411f
C364 XA.XIR[5].XIC[1].icell.SM Vbias 0.00701f
C365 XA.XIR[7].XIC[11].icell.PDM Vbias 0.04261f
C366 XA.XIR[10].XIC[10].icell.PDM VPWR 0.00799f
C367 XThR.Tn[13] Iout 1.16236f
C368 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.15202f
C369 XThR.XTB6.Y VPWR 1.05512f
C370 XThR.Tn[5] XA.XIR[6].XIC[11].icell.SM 0.00121f
C371 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C372 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00214f
C373 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PUM 0.00465f
C374 XA.XIR[15].XIC[9].icell.PDM Vbias 0.04261f
C375 XA.XIR[14].XIC[13].icell.PUM VPWR 0.00937f
C376 XA.XIR[4].XIC[4].icell.Ien Vbias 0.21098f
C377 XThC.Tn[13] VPWR 6.87751f
C378 XA.XIR[6].XIC[5].icell.SM VPWR 0.00158f
C379 XA.XIR[13].XIC[11].icell.PDM VPWR 0.00799f
C380 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.15202f
C381 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C382 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C383 XA.XIR[15].XIC[8].icell.PUM VPWR 0.00937f
C384 XA.XIR[5].XIC[8].icell.Ien VPWR 0.1903f
C385 XA.XIR[6].XIC[1].icell.SM Iout 0.00388f
C386 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PUM 0.00102f
C387 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C388 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11267f
C389 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.03425f
C390 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C391 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.03425f
C392 XA.XIR[5].XIC[4].icell.Ien Iout 0.06417f
C393 XA.XIR[4].XIC[11].icell.PUM VPWR 0.00937f
C394 XA.XIR[9].XIC[7].icell.PDM Vbias 0.04261f
C395 a_9827_9569# Vbias 0.00417f
C396 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00584f
C397 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C398 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00584f
C399 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.SM 0.0039f
C400 XA.XIR[0].XIC[2].icell.PUM VPWR 0.00877f
C401 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C402 XA.XIR[2].XIC[2].icell.PDM VPWR 0.00799f
C403 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02762f
C404 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C405 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PDM 0.00598f
C406 XA.XIR[13].XIC[1].icell.SM VPWR 0.00158f
C407 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.SM 0.0039f
C408 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00214f
C409 XA.XIR[9].XIC[7].icell.Ien Vbias 0.21098f
C410 XA.XIR[8].XIC[5].icell.PUM VPWR 0.00937f
C411 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02762f
C412 XThR.Tn[6] XA.XIR[7].XIC[3].icell.Ien 0.00338f
C413 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02762f
C414 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C415 XThR.Tn[2] XA.XIR[3].XIC[1].icell.Ien 0.00338f
C416 XA.XIR[12].XIC[3].icell.Ien VPWR 0.1903f
C417 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PUM 0.00465f
C418 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.SM 0.00168f
C419 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.SM 0.00168f
C420 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00584f
C421 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.SM 0.0039f
C422 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02812f
C423 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1909f
C424 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C425 XA.XIR[11].XIC[4].icell.SM VPWR 0.00158f
C426 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04031f
C427 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02762f
C428 XA.XIR[9].XIC[14].icell.PDM Iout 0.00117f
C429 XA.XIR[3].XIC[10].icell.PUM Vbias 0.0031f
C430 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9] 0.00341f
C431 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02762f
C432 XA.XIR[1].XIC[12].icell.PDM Vbias 0.04261f
C433 XThR.Tn[4] XA.XIR[5].XIC[1].icell.SM 0.00121f
C434 XThC.Tn[4] XThR.Tn[13] 0.28739f
C435 XA.XIR[9].XIC[14].icell.PUM VPWR 0.00937f
C436 XA.XIR[6].XIC[13].icell.SM Vbias 0.00701f
C437 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11] 0.00341f
C438 XA.XIR[10].XIC[6].icell.SM VPWR 0.00158f
C439 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00584f
C440 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.SM 0.0039f
C441 XA.XIR[4].XIC_15.icell.SM VPWR 0.00275f
C442 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.0353f
C443 XThR.Tn[14] XA.XIR[15].XIC[3].icell.Ien 0.00338f
C444 XThR.Tn[3] XA.XIR[4].XIC[1].icell.SM 0.00121f
C445 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C446 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.15202f
C447 XA.XIR[2].XIC[3].icell.PUM Vbias 0.0031f
C448 XA.XIR[4].XIC[12].icell.PDM Vbias 0.04261f
C449 XA.XIR[7].XIC[3].icell.Ien Vbias 0.21098f
C450 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.SM 0.00168f
C451 XA.XIR[10].XIC[2].icell.SM Iout 0.00388f
C452 XA.XIR[0].XIC[7].icell.PUM VPWR 0.00877f
C453 XThR.Tn[9] XA.XIR[10].XIC[2].icell.SM 0.00121f
C454 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Iout 0.00347f
C455 XThC.XTB2.Y a_3773_9615# 0.2342f
C456 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00584f
C457 XThC.Tn[7] Iout 0.84037f
C458 XThC.XTB1.Y data[0] 0.06453f
C459 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C460 XThC.Tn[7] XThR.Tn[9] 0.28739f
C461 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00584f
C462 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.SM 0.0039f
C463 XA.XIR[1].XIC[5].icell.PUM Vbias 0.0031f
C464 XThC.XTB7.B Vbias 0.09241f
C465 XA.XIR[13].XIC_15.icell.Ien Vbias 0.21234f
C466 XA.XIR[14].XIC[7].icell.SM Vbias 0.00701f
C467 XThC.Tn[3] XThR.Tn[8] 0.28739f
C468 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PUM 0.00465f
C469 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.04036f
C470 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.03425f
C471 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00214f
C472 XA.XIR[3].XIC[11].icell.SM Iout 0.00388f
C473 XThC.Tn[0] XA.XIR[13].XIC_dummy_left.icell.Iout 0.00109f
C474 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C475 XA.XIR[6].XIC_dummy_right.icell.SM VPWR 0.00123f
C476 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.15202f
C477 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8] 0.00341f
C478 XA.XIR[2].XIC[8].icell.SM VPWR 0.00158f
C479 XA.XIR[7].XIC[10].icell.PUM VPWR 0.00937f
C480 XA.XIR[8].XIC[13].icell.PUM Vbias 0.0031f
C481 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Ien 0.00584f
C482 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C483 XA.XIR[11].XIC[10].icell.Ien VPWR 0.1903f
C484 XA.XIR[2].XIC[4].icell.SM Iout 0.00388f
C485 XA.XIR[1].XIC[10].icell.SM VPWR 0.00158f
C486 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04031f
C487 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PUM 0.00465f
C488 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00584f
C489 XA.XIR[1].XIC[6].icell.SM Iout 0.00388f
C490 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PUM 0.00465f
C491 XA.XIR[14].XIC[11].icell.PUM VPWR 0.00937f
C492 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00214f
C493 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00584f
C494 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11] 0.00341f
C495 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.SM 0.00168f
C496 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.15202f
C497 XThC.XTBN.A VPWR 0.88811f
C498 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00584f
C499 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Ien 0.00232f
C500 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.15202f
C501 XThC.Tn[5] XA.XIR[0].XIC[6].icell.Ien 0.0016f
C502 XA.XIR[8].XIC[14].icell.SM Iout 0.00388f
C503 a_9827_9569# XThC.Tn[13] 0.00173f
C504 XThR.Tn[11] XA.XIR[12].XIC[3].icell.SM 0.00121f
C505 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C506 XA.XIR[2].XIC[1].icell.PUM VPWR 0.00937f
C507 XThR.Tn[8] XA.XIR[9].XIC[14].icell.SM 0.00121f
C508 XA.XIR[0].XIC_15.icell.PUM Vbias 0.0031f
C509 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PUM 0.00465f
C510 XThC.Tn[0] XThC.Tn[2] 0.1179f
C511 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C512 XThR.Tn[2] XA.XIR[3].XIC[9].icell.Ien 0.00338f
C513 XA.XIR[11].XIC[0].icell.Ien VPWR 0.1903f
C514 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.SM 0.00168f
C515 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Ien 0.00584f
C516 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02762f
C517 XThR.Tn[4] XA.XIR[4].XIC[12].icell.PDM 0.00341f
C518 XThC.Tn[5] XThC.Tn[6] 0.30991f
C519 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C520 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04031f
C521 XA.XIR[7].XIC[2].icell.PDM VPWR 0.00799f
C522 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C523 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.15202f
C524 XA.XIR[10].XIC[2].icell.PUM VPWR 0.00937f
C525 XThR.Tn[3] XA.XIR[3].XIC[13].icell.PDM 0.00341f
C526 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C527 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14] 0.00341f
C528 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C529 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C530 XThR.Tn[1] XA.XIR[2].XIC[7].icell.SM 0.00121f
C531 XA.XIR[6].XIC[9].icell.PDM VPWR 0.00799f
C532 XA.XIR[15].XIC[1].icell.Ien Vbias 0.17899f
C533 XA.XIR[15].XIC[0].icell.PDM VPWR 0.0114f
C534 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C535 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.SM 0.0039f
C536 XThR.XTB6.A XThR.Tn[1] 0.00411f
C537 XA.XIR[14].XIC[6].icell.PDM VPWR 0.00799f
C538 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C539 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C540 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C541 XA.XIR[14].XIC[12].icell.Ien VPWR 0.19084f
C542 XA.XIR[11].XIC[2].icell.PDM Vbias 0.04261f
C543 XA.XIR[5].XIC[4].icell.PDM Iout 0.00117f
C544 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.03425f
C545 XA.XIR[13].XIC[10].icell.PDM VPWR 0.00799f
C546 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C547 XA.XIR[10].XIC[6].icell.PDM Vbias 0.04261f
C548 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02762f
C549 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.03574f
C550 XThR.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.00338f
C551 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.0353f
C552 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Iout 0.00395f
C553 XThC.XTB7.Y XThC.Tn[8] 0.07806f
C554 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C555 XThC.XTB7.B XThC.Tn[13] 0.00276f
C556 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Ien 0.00595f
C557 XThR.Tn[0] XA.XIR[1].XIC[14].icell.SM 0.00121f
C558 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.SM 0.00168f
C559 XA.XIR[9].XIC[4].icell.Ien VPWR 0.1903f
C560 XA.XIR[6].XIC[5].icell.PUM Vbias 0.0031f
C561 XA.XIR[12].XIC[3].icell.PDM Iout 0.00117f
C562 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00584f
C563 XThR.Tn[0] XThR.Tn[1] 0.22353f
C564 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.03425f
C565 XA.XIR[15].XIC[6].icell.Ien Vbias 0.17899f
C566 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PUM 0.00465f
C567 XA.XIR[11].XIC[9].icell.PDM Iout 0.00117f
C568 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C569 XA.XIR[5].XIC[6].icell.SM Vbias 0.00701f
C570 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.SM 0.00168f
C571 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11153f
C572 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00214f
C573 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.SM 0.0039f
C574 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.15202f
C575 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C576 XA.XIR[4].XIC[9].icell.Ien Vbias 0.21098f
C577 XA.XIR[3].XIC[7].icell.PUM VPWR 0.00937f
C578 XA.XIR[1].XIC[3].icell.PDM VPWR 0.00799f
C579 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02762f
C580 XA.XIR[0].XIC[0].icell.Ien Vbias 0.20983f
C581 XA.XIR[6].XIC[10].icell.SM VPWR 0.00158f
C582 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.03425f
C583 XA.XIR[6].XIC[6].icell.SM Iout 0.00388f
C584 XA.XIR[5].XIC[13].icell.Ien VPWR 0.1903f
C585 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7] 0.00341f
C586 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C587 XA.XIR[8].XIC[3].icell.Ien Vbias 0.21098f
C588 XA.XIR[4].XIC[3].icell.PDM VPWR 0.00799f
C589 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00584f
C590 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00214f
C591 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C592 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Iout 0.00347f
C593 XA.XIR[12].XIC[1].icell.SM Vbias 0.00701f
C594 XThC.XTB3.Y VPWR 1.07065f
C595 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C596 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C597 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02762f
C598 XThC.XTB1.Y XThC.Tn[0] 0.19116f
C599 XA.XIR[5].XIC[9].icell.Ien Iout 0.06417f
C600 XA.XIR[8].XIC[13].icell.PDM VPWR 0.00799f
C601 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.SM 0.0039f
C602 XA.XIR[3].XIC[11].icell.PDM VPWR 0.00799f
C603 XA.XIR[14].XIC[4].icell.SM VPWR 0.00158f
C604 XThC.Tn[14] XThR.Tn[3] 0.28745f
C605 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13] 0.00341f
C606 XA.XIR[0].XIC[14].icell.PDM Vbias 0.04282f
C607 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PUM 0.00465f
C608 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00214f
C609 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.03425f
C610 XA.XIR[11].XIC[4].icell.PUM Vbias 0.0031f
C611 XThC.Tn[2] VPWR 5.93664f
C612 XThC.XTB7.A a_6243_10571# 0.0017f
C613 XA.XIR[8].XIC[1].icell.PDM Iout 0.00117f
C614 XThC.XTBN.A a_9827_9569# 0.09118f
C615 XA.XIR[13].XIC[6].icell.SM VPWR 0.00158f
C616 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04031f
C617 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04031f
C618 XA.XIR[8].XIC[10].icell.PUM VPWR 0.00937f
C619 XA.XIR[9].XIC[12].icell.Ien Vbias 0.21098f
C620 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C621 XA.XIR[10].XIC[6].icell.PUM Vbias 0.0031f
C622 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.PDM 0.00591f
C623 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00256f
C624 XThR.Tn[6] XA.XIR[7].XIC[8].icell.Ien 0.00338f
C625 XA.XIR[2].XIC[5].icell.PDM Iout 0.00117f
C626 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07214f
C627 XA.XIR[11].XIC_15.icell.Ien VPWR 0.25566f
C628 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00584f
C629 XA.XIR[13].XIC[2].icell.SM Iout 0.00388f
C630 XA.XIR[12].XIC[8].icell.Ien VPWR 0.1903f
C631 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00214f
C632 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C633 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C634 XA.XIR[0].XIC[5].icell.Ien Vbias 0.2113f
C635 XThC.Tn[8] XThR.Tn[0] 0.28773f
C636 XThC.Tn[10] XThR.Tn[5] 0.28739f
C637 XA.XIR[12].XIC[4].icell.Ien Iout 0.06417f
C638 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C639 XThR.Tn[0] XA.XIR[0].XIC[2].icell.PDM 0.00341f
C640 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C641 XA.XIR[3].XIC_15.icell.PUM Vbias 0.0031f
C642 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00214f
C643 XThR.Tn[4] XA.XIR[5].XIC[6].icell.SM 0.00121f
C644 XThR.Tn[1] XA.XIR[1].XIC[0].icell.PDM 0.00347f
C645 XA.XIR[11].XIC[5].icell.SM Iout 0.00388f
C646 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C647 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C648 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.15202f
C649 XThR.Tn[3] XA.XIR[4].XIC[6].icell.SM 0.00121f
C650 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.03425f
C651 XThR.Tn[14] XA.XIR[15].XIC[8].icell.Ien 0.00338f
C652 XA.XIR[14].XIC[10].icell.Ien VPWR 0.19084f
C653 XA.XIR[2].XIC[8].icell.PUM Vbias 0.0031f
C654 XA.XIR[10].XIC_dummy_right.icell.Ien Vbias 0.00288f
C655 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11] 0.00341f
C656 XA.XIR[7].XIC[8].icell.Ien Vbias 0.21098f
C657 XThC.XTB5.Y a_5155_9615# 0.24821f
C658 XA.XIR[10].XIC[7].icell.SM Iout 0.00388f
C659 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C660 XThR.Tn[9] XA.XIR[10].XIC[7].icell.SM 0.00121f
C661 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00214f
C662 XA.XIR[0].XIC[12].icell.PUM VPWR 0.00878f
C663 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5] 0.00341f
C664 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C665 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PUM 0.00465f
C666 XA.XIR[1].XIC[10].icell.PUM Vbias 0.0031f
C667 XThC.XTB7.A a_4067_9615# 0.0127f
C668 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C669 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PDM 0.00172f
C670 XThC.XTBN.A XThC.XTB7.B 0.35142f
C671 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04052f
C672 XA.XIR[11].XIC_dummy_left.icell.SM VPWR 0.00269f
C673 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[10].icell.SM 0.0039f
C674 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01577f
C675 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.03425f
C676 XA.XIR[2].XIC[13].icell.SM VPWR 0.00158f
C677 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C678 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.15202f
C679 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00584f
C680 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PUM 0.00465f
C681 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6] 0.00341f
C682 XA.XIR[2].XIC[9].icell.SM Iout 0.00388f
C683 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14] 0.00341f
C684 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.SM 0.00168f
C685 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.SM 0.0039f
C686 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.03425f
C687 XThR.Tn[12] XA.XIR[13].XIC[5].icell.SM 0.00121f
C688 XA.XIR[4].XIC[1].icell.Ien VPWR 0.1903f
C689 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C690 XA.XIR[1].XIC[11].icell.SM Iout 0.00388f
C691 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C692 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.03425f
C693 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.15202f
C694 XA.XIR[13].XIC[2].icell.PUM VPWR 0.00937f
C695 XThC.XTBN.Y a_5155_9615# 0.07602f
C696 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00214f
C697 XA.XIR[10].XIC[0].icell.Ien Vbias 0.20951f
C698 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.15202f
C699 XThR.Tn[11] XA.XIR[12].XIC[8].icell.SM 0.00121f
C700 XA.XIR[6].XIC[5].icell.PDM Vbias 0.04261f
C701 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.SM 0.00168f
C702 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00214f
C703 XThR.Tn[2] XA.XIR[3].XIC[14].icell.Ien 0.00338f
C704 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.SM 0.0039f
C705 Vbias bias[0] 0.17404f
C706 bias[1] bias[2] 0.03172f
C707 XThC.XTB1.Y VPWR 1.1176f
C708 XA.XIR[14].XIC[2].icell.PDM Vbias 0.04261f
C709 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PUM 0.00176f
C710 XA.XIR[5].XIC[12].icell.PDM Vbias 0.04261f
C711 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C712 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02762f
C713 XA.XIR[15].XIC[3].icell.Ien VPWR 0.32895f
C714 XThR.Tn[7] Iout 1.16233f
C715 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C716 XA.XIR[5].XIC[3].icell.SM VPWR 0.00158f
C717 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.15202f
C718 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.SM 0.0039f
C719 XA.XIR[7].XIC_15.icell.SM Iout 0.0047f
C720 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02762f
C721 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02762f
C722 XA.XIR[13].XIC[6].icell.PDM Vbias 0.04261f
C723 XThC.XTB7.A XThC.Tn[3] 0.03065f
C724 XThR.Tn[1] XA.XIR[2].XIC[12].icell.SM 0.00121f
C725 XA.XIR[7].XIC[5].icell.PDM Iout 0.00117f
C726 XA.XIR[4].XIC[6].icell.Ien VPWR 0.1903f
C727 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01432f
C728 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.15235f
C729 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00214f
C730 XA.XIR[15].XIC[3].icell.PDM Iout 0.00117f
C731 XA.XIR[6].XIC[12].icell.PDM Iout 0.00117f
C732 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PUM 0.00465f
C733 XA.XIR[4].XIC[2].icell.Ien Iout 0.06417f
C734 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C735 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.SM 0.0039f
C736 XA.XIR[9].XIC[2].icell.SM Vbias 0.00701f
C737 a_2979_9615# XThC.Tn[0] 0.28426f
C738 XA.XIR[14].XIC[9].icell.PDM Iout 0.00117f
C739 XA.XIR[9].XIC[13].icell.PDM VPWR 0.00799f
C740 XThC.Tn[12] XThR.Tn[6] 0.28739f
C741 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.SM 0.0039f
C742 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.SM 0.0039f
C743 XA.XIR[0].XIC[5].icell.PDM VPWR 0.00908f
C744 XA.XIR[7].XIC[0].icell.Ien VPWR 0.1903f
C745 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C746 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C747 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.03425f
C748 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00214f
C749 XA.XIR[9].XIC[1].icell.PDM Iout 0.00117f
C750 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.SM 0.00168f
C751 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C752 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C753 XA.XIR[3].XIC[5].icell.Ien Vbias 0.21098f
C754 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9] 0.00341f
C755 XA.XIR[1].XIC[2].icell.PUM VPWR 0.00937f
C756 XA.XIR[6].XIC[10].icell.PUM Vbias 0.0031f
C757 XA.XIR[9].XIC[9].icell.Ien VPWR 0.1903f
C758 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00584f
C759 XA.XIR[10].XIC[3].icell.PUM VPWR 0.00937f
C760 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00584f
C761 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.SM 0.00168f
C762 XThC.Tn[14] XThR.Tn[11] 0.28745f
C763 XA.XIR[12].XIC[12].icell.SM Iout 0.00388f
C764 XA.XIR[9].XIC[5].icell.Ien Iout 0.06417f
C765 XA.XIR[5].XIC[11].icell.SM Vbias 0.00701f
C766 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C767 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C768 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18966f
C769 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.15202f
C770 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04031f
C771 XThC.Tn[4] XThR.Tn[7] 0.28739f
C772 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C773 XA.XIR[11].XIC[14].icell.PDM VPWR 0.00809f
C774 XThC.Tn[12] Vbias 2.48601f
C775 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04031f
C776 XA.XIR[8].XIC[9].icell.PDM Vbias 0.04261f
C777 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04031f
C778 XA.XIR[3].XIC[7].icell.PDM Vbias 0.04261f
C779 XA.XIR[4].XIC[14].icell.Ien Vbias 0.21098f
C780 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02771f
C781 XA.XIR[14].XIC[4].icell.PUM Vbias 0.0031f
C782 XThC.XTB7.B XThC.Tn[2] 0.00273f
C783 XA.XIR[3].XIC[12].icell.PUM VPWR 0.00937f
C784 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10] 0.00341f
C785 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.SM 0.00168f
C786 XThC.XTB7.Y XThC.Tn[6] 0.2144f
C787 XA.XIR[2].XIC[13].icell.PDM Vbias 0.04261f
C788 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14] 0.00341f
C789 XA.XIR[1].XIC[6].icell.PDM Iout 0.00117f
C790 XA.XIR[13].XIC[6].icell.PUM Vbias 0.0031f
C791 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.SM 0.00168f
C792 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07214f
C793 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02762f
C794 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C795 XA.XIR[8].XIC[8].icell.Ien Vbias 0.21098f
C796 XThC.XTB6.Y XThC.Tn[10] 0.02461f
C797 XA.XIR[2].XIC[5].icell.PUM VPWR 0.00937f
C798 XA.XIR[14].XIC_15.icell.Ien VPWR 0.25598f
C799 XA.XIR[7].XIC[5].icell.Ien VPWR 0.1903f
C800 XA.XIR[6].XIC[11].icell.SM Iout 0.00388f
C801 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PUM 0.00465f
C802 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.03425f
C803 XA.XIR[12].XIC[6].icell.SM Vbias 0.00701f
C804 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Iout 0.00347f
C805 XA.XIR[5].XIC[14].icell.Ien Iout 0.06417f
C806 XA.XIR[4].XIC[6].icell.PDM Iout 0.00117f
C807 XA.XIR[1].XIC[7].icell.PUM VPWR 0.00937f
C808 XThC.Tn[8] XThR.Tn[1] 0.28739f
C809 XA.XIR[10].XIC_15.icell.PDM Vbias 0.04401f
C810 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PUM 0.00429f
C811 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.SM 0.00168f
C812 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11] 0.00341f
C813 XA.XIR[11].XIC[9].icell.PUM Vbias 0.0031f
C814 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.15202f
C815 XA.XIR[3].XIC[14].icell.PDM Iout 0.00117f
C816 XA.XIR[14].XIC[5].icell.SM Iout 0.00388f
C817 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.SM 0.0039f
C818 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.SM 0.00168f
C819 XA.XIR[0].XIC_dummy_left.icell.Ien Vbias 0.00348f
C820 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.15202f
C821 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01577f
C822 XThR.Tn[7] XA.XIR[8].XIC[2].icell.Ien 0.00338f
C823 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C824 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C825 XThR.Tn[6] XA.XIR[7].XIC[13].icell.Ien 0.00338f
C826 XThC.Tn[8] XThR.Tn[12] 0.28739f
C827 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02762f
C828 XA.XIR[13].XIC_dummy_right.icell.Ien Vbias 0.00288f
C829 XA.XIR[13].XIC[7].icell.SM Iout 0.00388f
C830 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C831 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00584f
C832 XA.XIR[0].XIC[10].icell.Ien Vbias 0.2113f
C833 XA.XIR[11].XIC_dummy_right.icell.SM VPWR 0.00123f
C834 XA.XIR[12].XIC[9].icell.Ien Iout 0.06417f
C835 XThR.Tn[2] XA.XIR[3].XIC[4].icell.SM 0.00121f
C836 XThC.Tn[3] XThR.Tn[3] 0.28739f
C837 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.SM 0.0039f
C838 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C839 XThR.Tn[4] XA.XIR[5].XIC[11].icell.SM 0.00121f
C840 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14] 0.00341f
C841 XThR.Tn[1] XA.XIR[1].XIC_15.icell.PDM 0.00341f
C842 XThC.Tn[12] XThR.Tn[4] 0.28739f
C843 XA.XIR[14].XIC[0].icell.PUM VPWR 0.00937f
C844 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00584f
C845 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C846 XThR.Tn[3] XA.XIR[3].XIC[0].icell.PDM 0.00347f
C847 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04052f
C848 XThR.Tn[10] XA.XIR[11].XIC[3].icell.Ien 0.00338f
C849 XThR.Tn[3] XA.XIR[4].XIC[11].icell.SM 0.00121f
C850 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.03425f
C851 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.15202f
C852 a_2979_9615# VPWR 0.70527f
C853 XA.XIR[7].XIC[13].icell.Ien Vbias 0.21098f
C854 XA.XIR[2].XIC[13].icell.PUM Vbias 0.0031f
C855 XThR.Tn[11] XA.XIR[12].XIC[13].icell.SM 0.00121f
C856 XA.XIR[9].XIC[0].icell.Ien Iout 0.06411f
C857 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.15202f
C858 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.15202f
C859 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04031f
C860 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.15202f
C861 XThC.XTB4.Y XThC.Tn[10] 0.01391f
C862 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.SM 0.00168f
C863 XA.XIR[1].XIC_15.icell.PUM Vbias 0.0031f
C864 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.03425f
C865 XA.XIR[5].XIC[3].icell.PDM VPWR 0.00799f
C866 XThR.Tn[2] XA.XIR[2].XIC[12].icell.PDM 0.00341f
C867 XThC.XTB4.Y a_4861_9615# 0.23756f
C868 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00214f
C869 XThC.Tn[6] XThR.Tn[0] 0.28748f
C870 XA.XIR[8].XIC_15.icell.SM Iout 0.0047f
C871 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02762f
C872 XA.XIR[6].XIC[2].icell.PUM VPWR 0.00937f
C873 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.04036f
C874 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C875 XA.XIR[13].XIC[0].icell.Ien Vbias 0.20951f
C876 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.15202f
C877 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PUM 0.00465f
C878 XThC.XTB5.Y a_7875_9569# 0.00418f
C879 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00214f
C880 XThC.Tn[12] XThC.Tn[13] 0.23689f
C881 XA.XIR[12].XIC[2].icell.PDM VPWR 0.00799f
C882 XA.XIR[2].XIC[14].icell.SM Iout 0.00388f
C883 XA.XIR[12].XIC[2].icell.PUM Vbias 0.0031f
C884 XA.XIR[12].XIC[10].icell.SM Iout 0.00388f
C885 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.03425f
C886 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.SM 0.00168f
C887 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C888 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02762f
C889 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.SM 0.00168f
C890 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C891 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PUM 0.00465f
C892 XA.XIR[11].XIC[8].icell.PDM VPWR 0.00799f
C893 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02762f
C894 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02762f
C895 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.SM 0.00168f
C896 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C897 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00584f
C898 XA.XIR[15].XIC[1].icell.SM Vbias 0.00701f
C899 XA.XIR[5].XIC[3].icell.PUM Vbias 0.0031f
C900 XA.XIR[7].XIC[13].icell.PDM Vbias 0.04261f
C901 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00256f
C902 XA.XIR[10].XIC[0].icell.PDM Iout 0.00117f
C903 XA.XIR[4].XIC[4].icell.SM Vbias 0.00701f
C904 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.03425f
C905 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04037f
C906 XA.XIR[3].XIC[2].icell.Ien VPWR 0.1903f
C907 XA.XIR[6].XIC[7].icell.PUM VPWR 0.00937f
C908 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.03425f
C909 XA.XIR[7].XIC_dummy_left.icell.SM VPWR 0.00269f
C910 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Ien 0.00214f
C911 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.SM 0.00168f
C912 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C913 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00214f
C914 XA.XIR[15].XIC[8].icell.Ien VPWR 0.32895f
C915 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02762f
C916 XA.XIR[5].XIC[8].icell.SM VPWR 0.00158f
C917 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00214f
C918 XThC.XTBN.Y a_7875_9569# 0.229f
C919 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.15202f
C920 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00214f
C921 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00584f
C922 XA.XIR[15].XIC[4].icell.Ien Iout 0.06807f
C923 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.15202f
C924 XA.XIR[5].XIC[4].icell.SM Iout 0.00388f
C925 XA.XIR[9].XIC[9].icell.PDM Vbias 0.04261f
C926 a_10915_9569# Vbias 0.00873f
C927 XA.XIR[8].XIC[0].icell.PDM VPWR 0.00799f
C928 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C929 XA.XIR[4].XIC[11].icell.Ien VPWR 0.1903f
C930 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C931 XA.XIR[0].XIC[1].icell.PDM Vbias 0.04282f
C932 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C933 XThC.Tn[5] XThR.Tn[2] 0.28739f
C934 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.SM 0.0039f
C935 XA.XIR[4].XIC[7].icell.Ien Iout 0.06417f
C936 XA.XIR[11].XIC[13].icell.PDM VPWR 0.00799f
C937 XA.XIR[2].XIC[4].icell.PDM VPWR 0.00799f
C938 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PUM 0.00465f
C939 XA.XIR[13].XIC[3].icell.PUM VPWR 0.00937f
C940 XA.XIR[9].XIC[7].icell.SM Vbias 0.00701f
C941 XThC.Tn[14] XThR.Tn[14] 0.28745f
C942 XA.XIR[8].XIC[5].icell.Ien VPWR 0.1903f
C943 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.SM 0.00168f
C944 XThR.Tn[6] XA.XIR[7].XIC[3].icell.SM 0.00121f
C945 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C946 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PUM 0.00465f
C947 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C948 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.03425f
C949 XA.XIR[12].XIC[3].icell.SM VPWR 0.00158f
C950 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C951 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C952 XA.XIR[14].XIC[14].icell.PDM VPWR 0.00809f
C953 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00584f
C954 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.SM 0.00168f
C955 VPWR bias[2] 1.5142f
C956 XA.XIR[11].XIC[6].icell.PUM VPWR 0.00937f
C957 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Ien 0.00584f
C958 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04031f
C959 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00214f
C960 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.SM 0.0039f
C961 a_n1335_4229# data[4] 0.00451f
C962 XThR.Tn[11] XA.XIR[12].XIC[11].icell.SM 0.00121f
C963 XA.XIR[3].XIC[10].icell.Ien Vbias 0.21098f
C964 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C965 XA.XIR[1].XIC[14].icell.PDM Vbias 0.04261f
C966 XA.XIR[7].XIC[1].icell.Ien Iout 0.06417f
C967 XThC.XTB2.Y XThC.Tn[10] 0.00106f
C968 XA.XIR[6].XIC_15.icell.PUM Vbias 0.0031f
C969 XA.XIR[9].XIC[14].icell.Ien VPWR 0.19036f
C970 XA.XIR[10].XIC[8].icell.PUM VPWR 0.00937f
C971 XA.XIR[10].XIC[14].icell.PDM Vbias 0.04261f
C972 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C973 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00214f
C974 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02762f
C975 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.SM 0.00168f
C976 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11] 0.00341f
C977 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00256f
C978 XThR.Tn[14] XA.XIR[15].XIC[3].icell.SM 0.00121f
C979 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Iout 0.00347f
C980 XA.XIR[2].XIC[3].icell.Ien Vbias 0.21098f
C981 XA.XIR[4].XIC[14].icell.PDM Vbias 0.04261f
C982 XA.XIR[7].XIC[3].icell.SM Vbias 0.00701f
C983 XA.XIR[9].XIC[10].icell.Ien Iout 0.06417f
C984 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C985 XThC.XTB2.Y a_4861_9615# 0.00851f
C986 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.15202f
C987 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C988 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18965f
C989 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00214f
C990 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.SM 0.0039f
C991 XThC.Tn[1] XThR.Tn[6] 0.28739f
C992 XA.XIR[12].XIC[14].icell.Ien Iout 0.06417f
C993 XA.XIR[13].XIC_15.icell.PDM Vbias 0.04401f
C994 XA.XIR[1].XIC[5].icell.Ien Vbias 0.21104f
C995 XA.XIR[14].XIC[9].icell.PUM Vbias 0.0031f
C996 XA.XIR[0].XIC[3].icell.Ien Iout 0.06389f
C997 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.03023f
C998 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04031f
C999 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1000 XThC.XTBN.A XThC.Tn[12] 0.22686f
C1001 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C1002 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00584f
C1003 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.SM 0.00168f
C1004 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8] 0.00341f
C1005 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04031f
C1006 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02762f
C1007 XThR.Tn[5] a_n1049_5611# 0.27042f
C1008 XA.XIR[8].XIC[13].icell.Ien Vbias 0.21098f
C1009 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14] 0.00341f
C1010 XA.XIR[2].XIC[10].icell.PUM VPWR 0.00937f
C1011 XA.XIR[7].XIC[10].icell.Ien VPWR 0.1903f
C1012 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C1013 XThC.Tn[3] XThR.Tn[11] 0.28739f
C1014 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00584f
C1015 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.389f
C1016 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.SM 0.0039f
C1017 XA.XIR[1].XIC[12].icell.PUM VPWR 0.00937f
C1018 XA.XIR[14].XIC_dummy_right.icell.SM VPWR 0.00123f
C1019 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00214f
C1020 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00584f
C1021 XA.XIR[7].XIC[6].icell.Ien Iout 0.06417f
C1022 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04031f
C1023 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.03425f
C1024 XThC.Tn[1] Vbias 2.40656f
C1025 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.SM 0.00168f
C1026 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.03425f
C1027 XThC.XTBN.Y Iout 0.00167f
C1028 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C1029 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.SM 0.0039f
C1030 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C1031 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C1032 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.15202f
C1033 XThR.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.00338f
C1034 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.SM 0.0039f
C1035 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.03425f
C1036 XA.XIR[8].XIC[0].icell.Ien VPWR 0.1903f
C1037 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00584f
C1038 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00214f
C1039 XThC.XTB5.Y XThC.Tn[4] 0.19958f
C1040 a_10915_9569# XThC.Tn[13] 0.01061f
C1041 XThR.Tn[5] XA.XIR[6].XIC[3].icell.Ien 0.00338f
C1042 XA.XIR[0].XIC_15.icell.Ien Vbias 0.21265f
C1043 XThC.XTB6.Y a_7651_9569# 0.0046f
C1044 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Ien 0.00584f
C1045 XThR.Tn[2] XA.XIR[3].XIC[9].icell.SM 0.00121f
C1046 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.03425f
C1047 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.SM 0.0039f
C1048 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C1049 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PUM 0.00465f
C1050 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00214f
C1051 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00584f
C1052 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04031f
C1053 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.15202f
C1054 XThR.Tn[4] XA.XIR[4].XIC[14].icell.PDM 0.00341f
C1055 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02762f
C1056 XA.XIR[7].XIC[4].icell.PDM VPWR 0.00799f
C1057 XThC.Tn[6] XThR.Tn[1] 0.2874f
C1058 XThR.Tn[3] XA.XIR[3].XIC_15.icell.PDM 0.00341f
C1059 XA.XIR[6].XIC[0].icell.Ien Vbias 0.20951f
C1060 XThR.Tn[10] XA.XIR[11].XIC[8].icell.Ien 0.00338f
C1061 XThR.XTB6.A XThR.XTB7.A 0.44014f
C1062 XThC.Tn[10] Iout 0.83837f
C1063 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C1064 XThC.Tn[10] XThR.Tn[9] 0.28739f
C1065 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.SM 0.00168f
C1066 XA.XIR[4].XIC[1].icell.SM VPWR 0.00158f
C1067 XA.XIR[15].XIC[2].icell.PDM VPWR 0.0114f
C1068 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.15202f
C1069 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00214f
C1070 XA.XIR[6].XIC[11].icell.PDM VPWR 0.00799f
C1071 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PUM 0.00465f
C1072 XThC.Tn[6] XThR.Tn[12] 0.28739f
C1073 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02762f
C1074 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.15202f
C1075 XThR.XTB5.A XThR.Tn[8] 0.00204f
C1076 XA.XIR[14].XIC[8].icell.PDM VPWR 0.00799f
C1077 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C1078 XThR.XTB5.Y a_n997_1803# 0.06458f
C1079 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PDM 0.0059f
C1080 XA.XIR[11].XIC[4].icell.PDM Vbias 0.04261f
C1081 XA.XIR[15].XIC[12].icell.SM Iout 0.00388f
C1082 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Iout 0.00347f
C1083 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C1084 XA.XIR[5].XIC[6].icell.PDM Iout 0.00117f
C1085 XThR.Tn[11] XA.XIR[12].XIC[9].icell.SM 0.00121f
C1086 XThC.XTBN.Y XThC.Tn[4] 0.61061f
C1087 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00584f
C1088 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.15202f
C1089 XA.XIR[10].XIC[8].icell.PDM Vbias 0.04261f
C1090 XThC.Tn[1] XThR.Tn[4] 0.28739f
C1091 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00584f
C1092 XA.XIR[9].XIC[0].icell.PDM VPWR 0.00799f
C1093 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00214f
C1094 XA.XIR[13].XIC[0].icell.PDM Iout 0.00117f
C1095 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.SM 0.00168f
C1096 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PUM 0.00465f
C1097 XThR.Tn[1] XA.XIR[2].XIC[0].icell.Ien 0.00338f
C1098 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.SM 0.0039f
C1099 XA.XIR[6].XIC[5].icell.Ien Vbias 0.21098f
C1100 XA.XIR[9].XIC[4].icell.SM VPWR 0.00158f
C1101 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1102 XA.XIR[12].XIC[5].icell.PDM Iout 0.00117f
C1103 XA.XIR[12].XIC[12].icell.Ien Iout 0.06417f
C1104 XThC.XTB4.Y a_7651_9569# 0.00497f
C1105 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02762f
C1106 XA.XIR[11].XIC[12].icell.PDM VPWR 0.00799f
C1107 XThC.Tn[5] XThR.Tn[10] 0.28739f
C1108 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.03425f
C1109 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.03425f
C1110 XA.XIR[15].XIC[6].icell.SM Vbias 0.00701f
C1111 XA.XIR[5].XIC[8].icell.PUM Vbias 0.0031f
C1112 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00214f
C1113 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C1114 XThC.Tn[0] XA.XIR[4].XIC_dummy_left.icell.Iout 0.00109f
C1115 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00584f
C1116 XA.XIR[4].XIC[9].icell.SM Vbias 0.00701f
C1117 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.SM 0.0039f
C1118 XA.XIR[1].XIC[5].icell.PDM VPWR 0.00799f
C1119 XA.XIR[3].XIC[7].icell.Ien VPWR 0.1903f
C1120 XThR.Tn[8] XA.XIR[9].XIC[1].icell.Ien 0.00338f
C1121 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C1122 XA.XIR[8].XIC[1].icell.Ien Iout 0.06417f
C1123 XA.XIR[0].XIC[0].icell.SM Vbias 0.00691f
C1124 XA.XIR[6].XIC[12].icell.PUM VPWR 0.00937f
C1125 XA.XIR[14].XIC[13].icell.PDM VPWR 0.00799f
C1126 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00584f
C1127 XA.XIR[3].XIC[3].icell.Ien Iout 0.06417f
C1128 XA.XIR[2].XIC[0].icell.PDM Vbias 0.04207f
C1129 a_4861_9615# XThC.Tn[4] 0.00198f
C1130 XA.XIR[8].XIC[3].icell.SM Vbias 0.00701f
C1131 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[4].icell.Ien 0.00214f
C1132 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.SM 0.0039f
C1133 XA.XIR[4].XIC[5].icell.PDM VPWR 0.00799f
C1134 XA.XIR[5].XIC[13].icell.SM VPWR 0.00158f
C1135 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7] 0.00341f
C1136 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04031f
C1137 XA.XIR[10].XIC[13].icell.PDM Vbias 0.04261f
C1138 XThR.XTB5.Y XThR.Tn[13] 0.00145f
C1139 XA.XIR[15].XIC[9].icell.Ien Iout 0.06807f
C1140 XA.XIR[12].XIC[3].icell.PUM Vbias 0.0031f
C1141 XThC.XTBN.Y XA.XIR[0].XIC[11].icell.PDM 0.00104f
C1142 XA.XIR[1].XIC[2].icell.Ien VPWR 0.1903f
C1143 XA.XIR[5].XIC[9].icell.SM Iout 0.00388f
C1144 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07214f
C1145 XA.XIR[3].XIC[13].icell.PDM VPWR 0.00799f
C1146 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13] 0.00341f
C1147 XThC.XTB7.A data[2] 0.00198f
C1148 XA.XIR[14].XIC[6].icell.PUM VPWR 0.00937f
C1149 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.03426f
C1150 XA.XIR[11].XIC[4].icell.Ien Vbias 0.21098f
C1151 XA.XIR[4].XIC[12].icell.Ien Iout 0.06417f
C1152 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PUM 0.00465f
C1153 XA.XIR[8].XIC[3].icell.PDM Iout 0.00117f
C1154 XA.XIR[3].XIC[1].icell.PDM Iout 0.00117f
C1155 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04031f
C1156 XA.XIR[13].XIC[14].icell.PDM Vbias 0.04261f
C1157 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.SM 0.0039f
C1158 XA.XIR[9].XIC[12].icell.SM Vbias 0.00701f
C1159 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04031f
C1160 XA.XIR[13].XIC[8].icell.PUM VPWR 0.00937f
C1161 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C1162 XA.XIR[8].XIC[10].icell.Ien VPWR 0.1903f
C1163 XA.XIR[10].XIC[6].icell.Ien Vbias 0.21098f
C1164 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PUM 0.00444f
C1165 XThR.Tn[6] XA.XIR[7].XIC[8].icell.SM 0.00121f
C1166 XA.XIR[2].XIC[7].icell.PDM Iout 0.00117f
C1167 XA.XIR[12].XIC[8].icell.SM VPWR 0.00158f
C1168 XA.XIR[8].XIC[6].icell.Ien Iout 0.06417f
C1169 XThR.Tn[8] XA.XIR[9].XIC[6].icell.Ien 0.00338f
C1170 XA.XIR[0].XIC[5].icell.SM Vbias 0.00716f
C1171 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14] 0.00341f
C1172 XA.XIR[12].XIC[4].icell.SM Iout 0.00388f
C1173 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.SM 0.00168f
C1174 XThR.Tn[0] XA.XIR[0].XIC[4].icell.PDM 0.00341f
C1175 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.SM 0.0039f
C1176 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1177 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00214f
C1178 XA.XIR[3].XIC_15.icell.Ien Vbias 0.21234f
C1179 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PUM 0.00465f
C1180 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1181 XThR.Tn[1] XA.XIR[1].XIC[2].icell.PDM 0.00341f
C1182 XThR.Tn[0] XA.XIR[1].XIC[1].icell.Ien 0.00338f
C1183 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C1184 XThR.Tn[11] XA.XIR[12].XIC[13].icell.Ien 0.00338f
C1185 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C1186 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04031f
C1187 XA.XIR[1].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1188 XThR.Tn[14] XA.XIR[15].XIC[8].icell.SM 0.00121f
C1189 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02762f
C1190 XThC.Tn[3] XThR.Tn[14] 0.28739f
C1191 XA.XIR[7].XIC[8].icell.SM Vbias 0.00701f
C1192 XA.XIR[2].XIC[8].icell.Ien Vbias 0.21098f
C1193 XA.XIR[9].XIC_15.icell.Ien Iout 0.0642f
C1194 XA.XIR[0].XIC[12].icell.Ien VPWR 0.19211f
C1195 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C1196 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00214f
C1197 XThC.XTB5.Y a_6243_9615# 0.00907f
C1198 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.SM 0.00168f
C1199 XA.XIR[15].XIC[10].icell.SM Iout 0.00388f
C1200 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.SM 0.00168f
C1201 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5] 0.00341f
C1202 XA.XIR[8].XIC_dummy_left.icell.SM VPWR 0.00269f
C1203 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.03425f
C1204 XA.XIR[4].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1205 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Ien 0.00584f
C1206 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.SM 0.0039f
C1207 XA.XIR[1].XIC[10].icell.Ien Vbias 0.21104f
C1208 XThC.XTB7.A a_5155_9615# 0.02287f
C1209 XA.XIR[0].XIC[8].icell.Ien Iout 0.06389f
C1210 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C1211 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C1212 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00214f
C1213 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PUM 0.00465f
C1214 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.SM 0.0039f
C1215 XThR.Tn[13] XA.XIR[14].XIC[3].icell.Ien 0.00338f
C1216 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04035f
C1217 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01577f
C1218 XA.XIR[7].XIC_15.icell.Ien VPWR 0.25566f
C1219 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.SM 0.00168f
C1220 XA.XIR[12].XIC[10].icell.Ien Iout 0.06417f
C1221 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.15202f
C1222 XThC.XTB2.Y a_7651_9569# 0.00191f
C1223 XA.XIR[5].XIC[0].icell.Ien VPWR 0.1903f
C1224 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6] 0.00341f
C1225 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C1226 XA.XIR[7].XIC[11].icell.Ien Iout 0.06417f
C1227 XThR.Tn[0] XA.XIR[1].XIC[6].icell.Ien 0.00338f
C1228 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C1229 XThR.XTB7.B XThR.XTB6.A 1.47641f
C1230 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C1231 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PUM 0.00465f
C1232 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PUM 0.00465f
C1233 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00214f
C1234 XA.XIR[14].XIC[1].icell.PUM VPWR 0.00937f
C1235 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C1236 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.1106f
C1237 XThC.Tn[14] VPWR 6.85545f
C1238 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.SM 0.00168f
C1239 XThR.Tn[11] XA.XIR[12].XIC[14].icell.SM 0.00121f
C1240 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PUM 0.00465f
C1241 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.SM 0.00168f
C1242 XThR.Tn[7] XA.XIR[8].XIC[12].icell.Ien 0.00338f
C1243 XA.XIR[10].XIC[0].icell.SM Vbias 0.00675f
C1244 XA.XIR[7].XIC[0].icell.PDM Vbias 0.04207f
C1245 XThC.XTBN.Y a_6243_9615# 0.07731f
C1246 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02762f
C1247 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C1248 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C1249 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C1250 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PUM 0.00465f
C1251 XA.XIR[3].XIC[0].icell.Ien Iout 0.06411f
C1252 XThR.Tn[5] XA.XIR[6].XIC[8].icell.Ien 0.00338f
C1253 XThR.Tn[8] Iout 1.16233f
C1254 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PUM 0.00465f
C1255 XThR.Tn[8] XThR.Tn[9] 0.05786f
C1256 XA.XIR[6].XIC[7].icell.PDM Vbias 0.04261f
C1257 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C1258 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1259 XThR.Tn[2] XA.XIR[3].XIC[14].icell.SM 0.00121f
C1260 XA.XIR[6].XIC[2].icell.Ien VPWR 0.1903f
C1261 XA.XIR[14].XIC[4].icell.PDM Vbias 0.04261f
C1262 XA.XIR[5].XIC[14].icell.PDM Vbias 0.04261f
C1263 XA.XIR[15].XIC[3].icell.SM VPWR 0.00158f
C1264 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01734f
C1265 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00584f
C1266 XA.XIR[5].XIC[5].icell.PUM VPWR 0.00937f
C1267 XA.XIR[11].XIC[1].icell.Ien Iout 0.06417f
C1268 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C1269 XA.XIR[2].XIC_15.icell.SM Iout 0.0047f
C1270 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.SM 0.0039f
C1271 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1272 XA.XIR[13].XIC[8].icell.PDM Vbias 0.04261f
C1273 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01432f
C1274 XA.XIR[7].XIC[7].icell.PDM Iout 0.00117f
C1275 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01785f
C1276 XA.XIR[11].XIC[11].icell.PDM VPWR 0.00799f
C1277 XA.XIR[4].XIC[6].icell.SM VPWR 0.00158f
C1278 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00584f
C1279 XA.XIR[9].XIC[0].icell.SM Iout 0.00388f
C1280 XA.XIR[15].XIC[5].icell.PDM Iout 0.00117f
C1281 XA.XIR[6].XIC[14].icell.PDM Iout 0.00117f
C1282 XA.XIR[4].XIC[2].icell.SM Iout 0.00388f
C1283 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.15202f
C1284 XThR.XTB2.Y data[5] 0.017f
C1285 XA.XIR[9].XIC[4].icell.PUM Vbias 0.0031f
C1286 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C1287 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00214f
C1288 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PUM 0.00465f
C1289 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.SM 0.0039f
C1290 XA.XIR[14].XIC[12].icell.PDM VPWR 0.00799f
C1291 XThC.Tn[5] XThR.Tn[13] 0.28739f
C1292 XA.XIR[15].XIC[14].icell.Ien Iout 0.06807f
C1293 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07214f
C1294 XA.XIR[11].XIC[12].icell.SM Vbias 0.00701f
C1295 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PUM 0.00465f
C1296 XThR.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.00338f
C1297 XA.XIR[0].XIC[7].icell.PDM VPWR 0.00773f
C1298 XA.XIR[7].XIC[0].icell.SM VPWR 0.00158f
C1299 XA.XIR[10].XIC[12].icell.PDM Vbias 0.04261f
C1300 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.SM 0.00168f
C1301 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.SM 0.0039f
C1302 XA.XIR[9].XIC[3].icell.PDM Iout 0.00117f
C1303 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9] 0.00341f
C1304 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C1305 XA.XIR[3].XIC[5].icell.SM Vbias 0.00701f
C1306 XThR.Tn[0] XThR.Tn[2] 0.00536f
C1307 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C1308 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PUM 0.00465f
C1309 XA.XIR[1].XIC[1].icell.PDM Vbias 0.04261f
C1310 XA.XIR[9].XIC[9].icell.SM VPWR 0.00158f
C1311 XThR.Tn[12] XA.XIR[13].XIC[1].icell.Ien 0.00338f
C1312 XA.XIR[6].XIC[10].icell.Ien Vbias 0.21098f
C1313 XThC.Tn[4] XThR.Tn[8] 0.28739f
C1314 XA.XIR[10].XIC[3].icell.Ien VPWR 0.1903f
C1315 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.SM 0.00168f
C1316 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C1317 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C1318 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C1319 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00214f
C1320 XA.XIR[12].XIC[13].icell.SM VPWR 0.00158f
C1321 XA.XIR[4].XIC[1].icell.PDM Vbias 0.04261f
C1322 XA.XIR[5].XIC[13].icell.PUM Vbias 0.0031f
C1323 XA.XIR[13].XIC[13].icell.PDM Vbias 0.04261f
C1324 XA.XIR[9].XIC[5].icell.SM Iout 0.00388f
C1325 XA.XIR[0].XIC[2].icell.SM VPWR 0.00158f
C1326 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04031f
C1327 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.SM 0.0039f
C1328 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.SM 0.00168f
C1329 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04031f
C1330 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00214f
C1331 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04052f
C1332 XA.XIR[3].XIC[9].icell.PDM Vbias 0.04261f
C1333 XA.XIR[3].XIC[12].icell.Ien VPWR 0.1903f
C1334 XA.XIR[4].XIC[14].icell.SM Vbias 0.00701f
C1335 XA.XIR[8].XIC[11].icell.PDM Vbias 0.04261f
C1336 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C1337 XA.XIR[14].XIC[4].icell.Ien Vbias 0.21098f
C1338 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10] 0.00341f
C1339 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C1340 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14] 0.00341f
C1341 XA.XIR[2].XIC_15.icell.PDM Vbias 0.04401f
C1342 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C1343 XA.XIR[3].XIC[8].icell.Ien Iout 0.06417f
C1344 XA.XIR[13].XIC[6].icell.Ien Vbias 0.21098f
C1345 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C1346 XA.XIR[1].XIC[8].icell.PDM Iout 0.00117f
C1347 XThR.Tn[14] XA.XIR[15].XIC[13].icell.SM 0.00121f
C1348 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Iout 0.00347f
C1349 XA.XIR[8].XIC[8].icell.SM Vbias 0.00701f
C1350 XA.XIR[2].XIC[5].icell.Ien VPWR 0.1903f
C1351 XA.XIR[7].XIC[5].icell.SM VPWR 0.00158f
C1352 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00214f
C1353 XA.XIR[9].XIC[0].icell.PUM VPWR 0.00937f
C1354 XA.XIR[11].XIC_15.icell.PUM Vbias 0.0031f
C1355 XA.XIR[12].XIC[8].icell.PUM Vbias 0.0031f
C1356 a_6243_10571# VPWR 0.00653f
C1357 XA.XIR[1].XIC[7].icell.Ien VPWR 0.1903f
C1358 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.SM 0.0039f
C1359 XA.XIR[5].XIC[14].icell.SM Iout 0.00388f
C1360 XA.XIR[7].XIC[1].icell.SM Iout 0.00388f
C1361 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C1362 XA.XIR[4].XIC[8].icell.PDM Iout 0.00117f
C1363 XThC.Tn[5] XA.XIR[0].XIC[6].icell.PDM 0.00343f
C1364 XThC.XTB6.Y a_5949_9615# 0.26831f
C1365 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00214f
C1366 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.15202f
C1367 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C1368 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.03511f
C1369 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.04494f
C1370 XThC.Tn[1] XThC.Tn[2] 0.72045f
C1371 XA.XIR[11].XIC[9].icell.Ien Vbias 0.21098f
C1372 XThC.Tn[0] XThC.Tn[3] 0.12427f
C1373 XA.XIR[1].XIC[3].icell.Ien Iout 0.06417f
C1374 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02762f
C1375 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C1376 XThR.Tn[7] XA.XIR[8].XIC[2].icell.SM 0.00121f
C1377 XA.XIR[8].XIC_15.icell.Ien VPWR 0.25566f
C1378 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.15202f
C1379 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02762f
C1380 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02762f
C1381 XThR.Tn[6] XA.XIR[7].XIC[13].icell.SM 0.00121f
C1382 XA.XIR[12].XIC_15.icell.Ien Iout 0.0642f
C1383 XThR.XTB7.A a_n1049_5317# 0.02018f
C1384 XA.XIR[8].XIC[11].icell.Ien Iout 0.06417f
C1385 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.SM 0.00168f
C1386 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.SM 0.0039f
C1387 XThR.Tn[8] XA.XIR[9].XIC[11].icell.Ien 0.00338f
C1388 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C1389 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.PDM 0.00578f
C1390 XA.XIR[0].XIC[10].icell.SM Vbias 0.00716f
C1391 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00584f
C1392 XThC.XTB5.A XThC.XTB6.Y 0.00193f
C1393 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.SM 0.0039f
C1394 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.SM 0.0039f
C1395 XThR.Tn[4] XA.XIR[4].XIC[1].icell.PDM 0.00341f
C1396 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C1397 XA.XIR[5].XIC_dummy_left.icell.SM VPWR 0.00269f
C1398 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C1399 XThR.Tn[3] XA.XIR[3].XIC[2].icell.PDM 0.00341f
C1400 XThR.Tn[10] XA.XIR[11].XIC[3].icell.SM 0.00121f
C1401 XA.XIR[7].XIC[13].icell.SM Vbias 0.00701f
C1402 a_4067_9615# VPWR 0.70648f
C1403 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PUM 0.00465f
C1404 XA.XIR[2].XIC[13].icell.Ien Vbias 0.21098f
C1405 XThR.Tn[1] XA.XIR[2].XIC[4].icell.Ien 0.00338f
C1406 a_n997_3755# XThR.Tn[9] 0.19352f
C1407 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.SM 0.0039f
C1408 XThR.XTB2.Y XThR.Tn[9] 0.292f
C1409 XA.XIR[1].XIC[1].icell.PUM Vbias 0.0031f
C1410 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04031f
C1411 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00214f
C1412 XA.XIR[11].XIC[10].icell.SM Vbias 0.00701f
C1413 XA.XIR[15].XIC[12].icell.Ien Iout 0.06807f
C1414 XA.XIR[1].XIC_15.icell.Ien Vbias 0.2124f
C1415 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.SM 0.0039f
C1416 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.15202f
C1417 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C1418 XA.XIR[0].XIC[13].icell.Ien Iout 0.06389f
C1419 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.15202f
C1420 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.03425f
C1421 XA.XIR[5].XIC[5].icell.PDM VPWR 0.00799f
C1422 XA.XIR[4].XIC[1].icell.PUM Vbias 0.0031f
C1423 XThR.XTB5.Y a_n997_3979# 0.00418f
C1424 XThR.Tn[2] XA.XIR[2].XIC[14].icell.PDM 0.00341f
C1425 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C1426 XThC.XTB4.Y a_5949_9615# 0.00465f
C1427 XThR.Tn[13] XA.XIR[14].XIC[8].icell.Ien 0.00338f
C1428 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1429 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PDM 0.00172f
C1430 XA.XIR[0].XIC_dummy_right.icell.Ien Vbias 0.00307f
C1431 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02762f
C1432 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C1433 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PUM 0.00465f
C1434 XA.XIR[13].XIC[0].icell.SM Vbias 0.00675f
C1435 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.SM 0.00168f
C1436 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00584f
C1437 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C1438 XThC.XTB5.Y a_8963_9569# 0.00427f
C1439 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C1440 XA.XIR[12].XIC[4].icell.PDM VPWR 0.00799f
C1441 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00584f
C1442 XA.XIR[12].XIC[11].icell.SM VPWR 0.00158f
C1443 XA.XIR[7].XIC_dummy_right.icell.SM VPWR 0.00123f
C1444 XThR.Tn[0] XA.XIR[1].XIC[11].icell.Ien 0.00338f
C1445 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C1446 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C1447 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.03425f
C1448 XA.XIR[11].XIC[10].icell.PDM VPWR 0.00799f
C1449 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Iout 0.00347f
C1450 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C1451 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C1452 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C1453 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C1454 XA.XIR[14].XIC[1].icell.Ien Iout 0.06417f
C1455 XA.XIR[15].XIC[3].icell.PUM Vbias 0.0031f
C1456 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.SM 0.0039f
C1457 XA.XIR[5].XIC[3].icell.Ien Vbias 0.21098f
C1458 XA.XIR[7].XIC_15.icell.PDM Vbias 0.04401f
C1459 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PUM 0.00465f
C1460 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00584f
C1461 XA.XIR[8].XIC[0].icell.SM VPWR 0.00158f
C1462 XA.XIR[14].XIC[11].icell.PDM VPWR 0.00799f
C1463 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00214f
C1464 XThR.Tn[14] XA.XIR[15].XIC[11].icell.SM 0.00121f
C1465 XA.XIR[10].XIC[2].icell.PDM Iout 0.00117f
C1466 XThR.Tn[5] XA.XIR[6].XIC[13].icell.Ien 0.00338f
C1467 XThR.XTB7.B XThR.Tn[12] 0.00772f
C1468 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04031f
C1469 XA.XIR[3].XIC[2].icell.SM VPWR 0.00158f
C1470 XA.XIR[4].XIC[6].icell.PUM Vbias 0.0031f
C1471 XA.XIR[11].XIC[13].icell.PUM Vbias 0.0031f
C1472 XThC.XTB1.Y XThC.Tn[1] 0.01447f
C1473 XA.XIR[6].XIC[7].icell.Ien VPWR 0.1903f
C1474 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.SM 0.00168f
C1475 XA.XIR[10].XIC[11].icell.PDM Vbias 0.04261f
C1476 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C1477 XThR.XTB7.A a_n1049_6405# 0.02287f
C1478 XThR.Tn[6] XThR.XTBN.A 0.00131f
C1479 XThC.Tn[3] VPWR 5.90764f
C1480 XA.XIR[6].XIC[3].icell.Ien Iout 0.06417f
C1481 XA.XIR[15].XIC[8].icell.SM VPWR 0.00158f
C1482 XA.XIR[5].XIC[10].icell.PUM VPWR 0.00937f
C1483 XThC.XTBN.Y a_8963_9569# 0.22784f
C1484 XA.XIR[14].XIC[12].icell.SM Vbias 0.00701f
C1485 XA.XIR[15].XIC[4].icell.SM Iout 0.00388f
C1486 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02762f
C1487 XA.XIR[9].XIC[11].icell.PDM Vbias 0.04261f
C1488 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C1489 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00214f
C1490 XA.XIR[3].XIC[0].icell.PDM VPWR 0.00799f
C1491 XA.XIR[4].XIC[11].icell.SM VPWR 0.00158f
C1492 XA.XIR[8].XIC[2].icell.PDM VPWR 0.00799f
C1493 XA.XIR[12].XIC[14].icell.PUM VPWR 0.00937f
C1494 XA.XIR[0].XIC[3].icell.PDM Vbias 0.04278f
C1495 XA.XIR[13].XIC[12].icell.PDM Vbias 0.04261f
C1496 XThR.XTB5.A XThR.XTB7.Y 0.00179f
C1497 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C1498 XThR.XTB5.A data[4] 0.14415f
C1499 XThC.Tn[9] XThR.Tn[0] 0.28777f
C1500 XThC.Tn[11] XThR.Tn[5] 0.28739f
C1501 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C1502 XA.XIR[4].XIC[7].icell.SM Iout 0.00388f
C1503 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C1504 XA.XIR[2].XIC[6].icell.PDM VPWR 0.00799f
C1505 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.03425f
C1506 XA.XIR[1].XIC[0].icell.SM Vbias 0.00679f
C1507 XA.XIR[13].XIC[3].icell.Ien VPWR 0.1903f
C1508 XThR.XTB5.Y XThR.Tn[7] 0.00912f
C1509 XThR.Tn[1] XThR.Tn[2] 0.10497f
C1510 XA.XIR[9].XIC[9].icell.PUM Vbias 0.0031f
C1511 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.SM 0.0039f
C1512 XThR.XTB5.Y a_n997_2891# 0.00424f
C1513 XA.XIR[8].XIC[5].icell.SM VPWR 0.00158f
C1514 XA.XIR[10].XIC[1].icell.SM Vbias 0.00701f
C1515 XThR.XTB1.Y a_n997_3979# 0.06353f
C1516 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C1517 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.03425f
C1518 XA.XIR[12].XIC[5].icell.PUM VPWR 0.00937f
C1519 XA.XIR[8].XIC[1].icell.SM Iout 0.00388f
C1520 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12] 0.00341f
C1521 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00584f
C1522 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00584f
C1523 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.SM 0.00168f
C1524 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PUM 0.00465f
C1525 XThR.Tn[8] XA.XIR[9].XIC[1].icell.SM 0.00121f
C1526 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C1527 XA.XIR[11].XIC[6].icell.Ien VPWR 0.1903f
C1528 XA.XIR[11].XIC[14].icell.Ien Vbias 0.21098f
C1529 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38912f
C1530 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04031f
C1531 XThR.Tn[6] Vbias 3.74624f
C1532 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.SM 0.0039f
C1533 XThR.Tn[4] XA.XIR[5].XIC[3].icell.Ien 0.00338f
C1534 XA.XIR[3].XIC[10].icell.SM Vbias 0.00701f
C1535 XA.XIR[2].XIC[1].icell.Ien Iout 0.06417f
C1536 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.0353f
C1537 XA.XIR[9].XIC[14].icell.SM VPWR 0.00207f
C1538 XA.XIR[6].XIC_15.icell.Ien Vbias 0.21234f
C1539 XA.XIR[10].XIC[8].icell.Ien VPWR 0.1903f
C1540 XA.XIR[11].XIC[2].icell.Ien Iout 0.06417f
C1541 XA.XIR[15].XIC[10].icell.Ien Iout 0.06807f
C1542 XThR.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.00338f
C1543 XA.XIR[9].XIC[10].icell.SM Iout 0.00388f
C1544 XA.XIR[7].XIC[5].icell.PUM Vbias 0.0031f
C1545 XA.XIR[10].XIC[4].icell.Ien Iout 0.06417f
C1546 XA.XIR[2].XIC[3].icell.SM Vbias 0.00701f
C1547 XA.XIR[14].XIC_15.icell.PUM Vbias 0.0031f
C1548 XThC.XTB2.Y a_5949_9615# 0.00844f
C1549 XThC.XTB7.B a_6243_10571# 0.00108f
C1550 XA.XIR[0].XIC[7].icell.SM VPWR 0.00158f
C1551 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.SM 0.00168f
C1552 XThR.Tn[9] XA.XIR[10].XIC[4].icell.Ien 0.00338f
C1553 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PUM 0.00471f
C1554 XA.XIR[1].XIC[5].icell.SM Vbias 0.00704f
C1555 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00584f
C1556 XThR.XTB7.B a_n1049_5317# 0.01743f
C1557 XA.XIR[14].XIC[9].icell.Ien Vbias 0.21098f
C1558 XA.XIR[0].XIC[3].icell.SM Iout 0.00367f
C1559 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Iout 0.00347f
C1560 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04031f
C1561 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C1562 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02762f
C1563 XThR.Tn[1] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00122f
C1564 data[5] data[4] 0.64735f
C1565 XA.XIR[12].XIC[9].icell.SM VPWR 0.00158f
C1566 XA.XIR[3].XIC[13].icell.Ien Iout 0.06417f
C1567 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00584f
C1568 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C1569 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04031f
C1570 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8] 0.00341f
C1571 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[9].icell.Ien 0.00214f
C1572 XA.XIR[2].XIC[10].icell.Ien VPWR 0.1903f
C1573 XA.XIR[8].XIC[13].icell.SM Vbias 0.00701f
C1574 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.15202f
C1575 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.0404f
C1576 VPWR data[6] 0.21221f
C1577 XA.XIR[7].XIC[10].icell.SM VPWR 0.00158f
C1578 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C1579 XA.XIR[2].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1580 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C1581 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00214f
C1582 XA.XIR[3].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1583 XThC.Tn[8] XThR.Tn[2] 0.28739f
C1584 XA.XIR[7].XIC[6].icell.SM Iout 0.00388f
C1585 XA.XIR[1].XIC[12].icell.Ien VPWR 0.1903f
C1586 XA.XIR[2].XIC[6].icell.Ien Iout 0.06417f
C1587 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04031f
C1588 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C1589 XThR.Tn[0] XA.XIR[1].XIC[1].icell.SM 0.00121f
C1590 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.15202f
C1591 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00214f
C1592 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PUM 0.00465f
C1593 XThR.Tn[12] XA.XIR[13].XIC[2].icell.Ien 0.00338f
C1594 XThR.Tn[14] XA.XIR[15].XIC[9].icell.SM 0.00121f
C1595 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C1596 XA.XIR[1].XIC[8].icell.Ien Iout 0.06417f
C1597 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02762f
C1598 XA.XIR[11].XIC[11].icell.PUM Vbias 0.0031f
C1599 XThR.XTBN.Y XA.XIR[6].XIC_dummy_left.icell.Ien 0.00159f
C1600 XThR.Tn[7] XA.XIR[8].XIC[7].icell.SM 0.00121f
C1601 XThR.XTB1.Y XThR.Tn[7] 0.00426f
C1602 a_n1335_4229# VPWR 0.00633f
C1603 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PUM 0.00465f
C1604 XA.XIR[8].XIC_dummy_right.icell.SM VPWR 0.00123f
C1605 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C1606 XThR.Tn[5] XA.XIR[6].XIC[3].icell.SM 0.00121f
C1607 XThR.Tn[11] XA.XIR[12].XIC[5].icell.Ien 0.00338f
C1608 XThC.XTB6.A XThC.Tn[9] 0.00838f
C1609 XThC.XTB6.Y a_8739_9569# 0.00466f
C1610 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02762f
C1611 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.03425f
C1612 XThC.XTB7.A XThC.Tn[4] 0.0274f
C1613 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C1614 XA.XIR[14].XIC[10].icell.SM Vbias 0.00701f
C1615 XA.XIR[11].XIC[0].icell.SM VPWR 0.00158f
C1616 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.SM 0.00168f
C1617 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00214f
C1618 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.15202f
C1619 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04031f
C1620 XA.XIR[12].XIC[12].icell.PUM VPWR 0.00937f
C1621 XA.XIR[5].XIC[1].icell.PDM Vbias 0.04261f
C1622 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1623 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.SM 0.00168f
C1624 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C1625 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PUM 0.00465f
C1626 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C1627 XA.XIR[7].XIC[6].icell.PDM VPWR 0.00799f
C1628 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C1629 XThR.Tn[10] XA.XIR[11].XIC[8].icell.SM 0.00121f
C1630 XA.XIR[6].XIC[0].icell.SM Vbias 0.00675f
C1631 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.SM 0.0039f
C1632 XA.XIR[4].XIC[3].icell.PUM VPWR 0.00937f
C1633 XThR.Tn[4] Vbias 3.74761f
C1634 XThR.Tn[1] XA.XIR[2].XIC[9].icell.Ien 0.00338f
C1635 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C1636 XA.XIR[15].XIC[4].icell.PDM VPWR 0.0114f
C1637 XA.XIR[6].XIC[13].icell.PDM VPWR 0.00799f
C1638 XThR.XTB6.Y XThR.Tn[6] 0.00639f
C1639 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C1640 XA.XIR[12].XIC[0].icell.PDM Vbias 0.04207f
C1641 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PUM 0.00465f
C1642 XThC.Tn[13] XThR.Tn[6] 0.2874f
C1643 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.03425f
C1644 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C1645 XA.XIR[14].XIC[10].icell.PDM VPWR 0.00799f
C1646 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.15202f
C1647 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C1648 XA.XIR[6].XIC[1].icell.PDM Iout 0.00117f
C1649 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C1650 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02762f
C1651 XA.XIR[15].XIC[13].icell.SM VPWR 0.00158f
C1652 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00584f
C1653 XA.XIR[11].XIC[6].icell.PDM Vbias 0.04261f
C1654 XA.XIR[11].XIC[12].icell.Ien Vbias 0.21098f
C1655 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.SM 0.0039f
C1656 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C1657 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.SM 0.0039f
C1658 XA.XIR[5].XIC[8].icell.PDM Iout 0.00117f
C1659 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C1660 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PUM 0.00465f
C1661 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01432f
C1662 XA.XIR[10].XIC[10].icell.PDM Vbias 0.04261f
C1663 XThR.XTB7.B a_n1049_6405# 0.00268f
C1664 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00584f
C1665 XA.XIR[9].XIC[2].icell.PDM VPWR 0.00799f
C1666 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[1].icell.SM 0.0039f
C1667 XA.XIR[13].XIC[2].icell.PDM Iout 0.00117f
C1668 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C1669 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PUM 0.00465f
C1670 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00214f
C1671 XA.XIR[14].XIC[13].icell.PUM Vbias 0.0031f
C1672 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Iout 0.00347f
C1673 XThC.Tn[5] XThR.Tn[7] 0.28739f
C1674 XThR.Tn[3] Iout 1.16236f
C1675 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PUM 0.00465f
C1676 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.03425f
C1677 XThC.Tn[13] Vbias 2.40092f
C1678 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C1679 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1680 XA.XIR[6].XIC[5].icell.SM Vbias 0.00701f
C1681 XA.XIR[9].XIC[6].icell.PUM VPWR 0.00937f
C1682 XA.XIR[12].XIC[13].icell.Ien VPWR 0.1903f
C1683 XA.XIR[13].XIC[11].icell.PDM Vbias 0.04261f
C1684 XA.XIR[12].XIC[7].icell.PDM Iout 0.00117f
C1685 XThC.XTB7.B XThC.Tn[3] 0.00532f
C1686 XThC.XTB4.Y a_8739_9569# 0.00813f
C1687 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02762f
C1688 XThC.XTB7.Y XThC.Tn[7] 0.0835f
C1689 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00214f
C1690 XA.XIR[15].XIC[8].icell.PUM Vbias 0.0031f
C1691 XA.XIR[5].XIC[8].icell.Ien Vbias 0.21098f
C1692 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.SM 0.00168f
C1693 XThR.XTB4.Y XThR.Tn[12] 0.00209f
C1694 XThC.XTB6.Y XThC.Tn[11] 0.02513f
C1695 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04031f
C1696 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.SM 0.0039f
C1697 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C1698 XA.XIR[3].XIC[7].icell.SM VPWR 0.00158f
C1699 XA.XIR[4].XIC[11].icell.PUM Vbias 0.0031f
C1700 XA.XIR[1].XIC[7].icell.PDM VPWR 0.00799f
C1701 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00584f
C1702 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.0353f
C1703 XThR.Tn[14] XA.XIR[15].XIC[13].icell.Ien 0.00338f
C1704 XA.XIR[0].XIC[2].icell.PUM Vbias 0.0031f
C1705 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C1706 XA.XIR[6].XIC[12].icell.Ien VPWR 0.1903f
C1707 XThC.Tn[9] XThR.Tn[1] 0.28739f
C1708 XA.XIR[10].XIC[12].icell.SM Iout 0.00388f
C1709 XThR.XTB5.Y a_n997_1579# 0.00133f
C1710 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.SM 0.00168f
C1711 XA.XIR[2].XIC[2].icell.PDM Vbias 0.04261f
C1712 XThR.Tn[10] XThR.Tn[12] 0.00142f
C1713 XA.XIR[3].XIC[3].icell.SM Iout 0.00388f
C1714 XThR.Tn[9] XA.XIR[10].XIC[12].icell.SM 0.00121f
C1715 XA.XIR[15].XIC_15.icell.Ien Iout 0.0681f
C1716 XA.XIR[13].XIC[1].icell.SM Vbias 0.00701f
C1717 XA.XIR[6].XIC[8].icell.Ien Iout 0.06417f
C1718 XA.XIR[8].XIC[5].icell.PUM Vbias 0.0031f
C1719 XA.XIR[4].XIC[7].icell.PDM VPWR 0.00799f
C1720 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C1721 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7] 0.00341f
C1722 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01577f
C1723 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.SM 0.00168f
C1724 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.SM 0.0039f
C1725 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04031f
C1726 XA.XIR[12].XIC[3].icell.Ien Vbias 0.21098f
C1727 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.SM 0.0039f
C1728 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07214f
C1729 XThC.Tn[9] XThR.Tn[12] 0.28739f
C1730 XA.XIR[1].XIC[2].icell.SM VPWR 0.00158f
C1731 XA.XIR[14].XIC[6].icell.Ien VPWR 0.19084f
C1732 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13] 0.00341f
C1733 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00584f
C1734 XA.XIR[14].XIC[14].icell.Ien Vbias 0.21098f
C1735 XA.XIR[11].XIC[4].icell.SM Vbias 0.00701f
C1736 XA.XIR[12].XIC[14].icell.SM VPWR 0.00207f
C1737 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.03425f
C1738 XA.XIR[8].XIC[5].icell.PDM Iout 0.00117f
C1739 XThR.XTBN.Y a_n1049_5317# 0.07731f
C1740 XA.XIR[3].XIC[3].icell.PDM Iout 0.00117f
C1741 XA.XIR[4].XIC[12].icell.SM Iout 0.00388f
C1742 XA.XIR[14].XIC[2].icell.Ien Iout 0.06417f
C1743 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00584f
C1744 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04031f
C1745 XA.XIR[13].XIC[8].icell.Ien VPWR 0.1903f
C1746 XThC.Tn[4] XThR.Tn[3] 0.28739f
C1747 XA.XIR[9].XIC[14].icell.PUM Vbias 0.0031f
C1748 XA.XIR[10].XIC[6].icell.SM Vbias 0.00701f
C1749 XA.XIR[8].XIC[10].icell.SM VPWR 0.00158f
C1750 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.03546f
C1751 XThR.Tn[4] XThR.XTB6.Y 0.00264f
C1752 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C1753 XA.XIR[2].XIC[9].icell.PDM Iout 0.00117f
C1754 XA.XIR[12].XIC[10].icell.PUM VPWR 0.00937f
C1755 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00584f
C1756 XA.XIR[13].XIC[4].icell.Ien Iout 0.06417f
C1757 XA.XIR[4].XIC_15.icell.SM Vbias 0.00701f
C1758 XThC.Tn[13] XThR.Tn[4] 0.2874f
C1759 XA.XIR[8].XIC[6].icell.SM Iout 0.00388f
C1760 XA.XIR[0].XIC[7].icell.PUM Vbias 0.0031f
C1761 XThR.Tn[8] XA.XIR[9].XIC[6].icell.SM 0.00121f
C1762 XThR.XTB3.Y XThR.Tn[5] 0.00381f
C1763 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.03023f
C1764 XThR.Tn[0] XA.XIR[0].XIC[6].icell.PDM 0.00341f
C1765 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C1766 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C1767 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.03425f
C1768 XThR.Tn[14] XA.XIR[15].XIC[14].icell.SM 0.00121f
C1769 XThR.Tn[4] XA.XIR[5].XIC[8].icell.Ien 0.00338f
C1770 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.SM 0.00168f
C1771 XThC.XTB4.Y XThC.Tn[11] 0.30582f
C1772 XThC.Tn[8] XThR.Tn[10] 0.28739f
C1773 XA.XIR[11].XIC[7].icell.Ien Iout 0.06417f
C1774 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C1775 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PUM 0.00186f
C1776 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C1777 XThR.Tn[1] XA.XIR[1].XIC[4].icell.PDM 0.00341f
C1778 XThC.Tn[0] XThR.Tn[5] 0.28743f
C1779 XA.XIR[9].XIC[1].icell.PUM VPWR 0.00937f
C1780 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C1781 XThR.Tn[3] XA.XIR[4].XIC[8].icell.Ien 0.00338f
C1782 XThC.Tn[7] XThR.Tn[0] 0.2882f
C1783 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04031f
C1784 XA.XIR[5].XIC_15.icell.SM Iout 0.0047f
C1785 XA.XIR[2].XIC[8].icell.SM Vbias 0.00701f
C1786 XA.XIR[15].XIC[11].icell.SM VPWR 0.00158f
C1787 XA.XIR[7].XIC[10].icell.PUM Vbias 0.0031f
C1788 XA.XIR[10].XIC[9].icell.Ien Iout 0.06417f
C1789 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C1790 XThC.Tn[8] XThC.Tn[9] 0.05322f
C1791 XA.XIR[0].XIC[12].icell.SM VPWR 0.00158f
C1792 XA.XIR[11].XIC[10].icell.Ien Vbias 0.21098f
C1793 XThR.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.00338f
C1794 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00584f
C1795 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C1796 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5] 0.00341f
C1797 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00214f
C1798 XThR.XTB4.Y a_n1049_5317# 0.00463f
C1799 XA.XIR[3].XIC[0].icell.PUM VPWR 0.00937f
C1800 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.SM 0.0039f
C1801 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PUM 0.00465f
C1802 XA.XIR[1].XIC[10].icell.SM Vbias 0.00704f
C1803 XThC.Tn[12] XThC.Tn[14] 0.03994f
C1804 XA.XIR[0].XIC[8].icell.SM Iout 0.00367f
C1805 XThC.XTB7.A a_6243_9615# 0.02018f
C1806 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1807 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.03425f
C1808 XThR.Tn[2] XA.XIR[2].XIC[1].icell.PDM 0.00341f
C1809 XThC.XTB7.A data[1] 0.06544f
C1810 XA.XIR[14].XIC[11].icell.PUM Vbias 0.0031f
C1811 XThR.Tn[13] XA.XIR[14].XIC[3].icell.SM 0.00121f
C1812 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04031f
C1813 XThR.Tn[10] XA.XIR[11].XIC[13].icell.SM 0.00121f
C1814 XThC.XTBN.A Vbias 0.01661f
C1815 XA.XIR[2].XIC_15.icell.Ien VPWR 0.25566f
C1816 XA.XIR[12].XIC[11].icell.Ien VPWR 0.1903f
C1817 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C1818 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Iout 0.00347f
C1819 a_n1319_5611# VPWR 0.00674f
C1820 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.SM 0.0039f
C1821 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6] 0.00341f
C1822 XA.XIR[2].XIC[1].icell.PUM Vbias 0.0031f
C1823 XA.XIR[2].XIC[11].icell.Ien Iout 0.06417f
C1824 XA.XIR[7].XIC[11].icell.SM Iout 0.00388f
C1825 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.15202f
C1826 XThR.Tn[0] XA.XIR[1].XIC[6].icell.SM 0.00121f
C1827 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02762f
C1828 XA.XIR[14].XIC[0].icell.SM VPWR 0.00158f
C1829 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.03425f
C1830 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.SM 0.00168f
C1831 XThR.Tn[12] XA.XIR[13].XIC[7].icell.Ien 0.00338f
C1832 XA.XIR[11].XIC[0].icell.Ien Vbias 0.20951f
C1833 XA.XIR[1].XIC[13].icell.Ien Iout 0.06417f
C1834 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C1835 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PDM 0.00172f
C1836 XThR.Tn[7] XA.XIR[8].XIC[12].icell.SM 0.00121f
C1837 XThR.Tn[14] XA.XIR[15].XIC[11].icell.Ien 0.00338f
C1838 XA.XIR[10].XIC[1].icell.PDM VPWR 0.00799f
C1839 XA.XIR[10].XIC[2].icell.PUM Vbias 0.0031f
C1840 XA.XIR[7].XIC[2].icell.PDM Vbias 0.04261f
C1841 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.SM 0.0039f
C1842 XA.XIR[1].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1843 XA.XIR[10].XIC[10].icell.SM Iout 0.00388f
C1844 XA.XIR[15].XIC[14].icell.PUM VPWR 0.00937f
C1845 XThR.Tn[9] XA.XIR[10].XIC[10].icell.SM 0.00121f
C1846 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.SM 0.0039f
C1847 XThR.Tn[5] XA.XIR[6].XIC[8].icell.SM 0.00121f
C1848 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.03425f
C1849 XA.XIR[3].XIC[0].icell.SM Iout 0.00388f
C1850 XThR.Tn[12] a_n997_1803# 0.18719f
C1851 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.PUM 0.00121f
C1852 XA.XIR[15].XIC[0].icell.PDM Vbias 0.04207f
C1853 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.SM 0.00168f
C1854 XThR.XTBN.Y a_n1049_6405# 0.07602f
C1855 XA.XIR[6].XIC[9].icell.PDM Vbias 0.04261f
C1856 XA.XIR[6].XIC[2].icell.SM VPWR 0.00158f
C1857 XA.XIR[12].XIC[0].icell.Ien Iout 0.06411f
C1858 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.SM 0.0039f
C1859 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.15202f
C1860 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00214f
C1861 XA.XIR[14].XIC[6].icell.PDM Vbias 0.04261f
C1862 XThC.Tn[6] XThR.Tn[2] 0.28739f
C1863 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02762f
C1864 a_n1049_6699# XThR.XTB5.Y 0.0021f
C1865 XA.XIR[14].XIC[12].icell.Ien Vbias 0.21098f
C1866 XA.XIR[15].XIC[5].icell.PUM VPWR 0.00937f
C1867 XA.XIR[5].XIC[5].icell.Ien VPWR 0.1903f
C1868 XThR.Tn[11] Iout 1.16235f
C1869 XThR.Tn[9] XThR.Tn[11] 0.00252f
C1870 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1871 XA.XIR[13].XIC[10].icell.PDM Vbias 0.04261f
C1872 XA.XIR[7].XIC[9].icell.PDM Iout 0.00117f
C1873 XA.XIR[4].XIC[8].icell.PUM VPWR 0.00937f
C1874 XThR.Tn[1] XA.XIR[2].XIC[14].icell.Ien 0.00338f
C1875 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.SM 0.0039f
C1876 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00214f
C1877 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C1878 XA.XIR[15].XIC[7].icell.PDM Iout 0.00117f
C1879 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PUM 0.00102f
C1880 XA.XIR[9].XIC[4].icell.Ien Vbias 0.21098f
C1881 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.03425f
C1882 XThR.XTB4.Y a_n1049_6405# 0.01546f
C1883 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00584f
C1884 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02762f
C1885 XThR.Tn[5] VPWR 6.61445f
C1886 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00584f
C1887 XA.XIR[2].XIC[0].icell.SM VPWR 0.00158f
C1888 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.03425f
C1889 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00584f
C1890 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.15235f
C1891 XA.XIR[7].XIC[2].icell.PUM VPWR 0.00937f
C1892 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01093f
C1893 XA.XIR[11].XIC[1].icell.SM VPWR 0.00158f
C1894 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C1895 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C1896 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C1897 XA.XIR[15].XIC[9].icell.SM VPWR 0.00158f
C1898 XA.XIR[3].XIC[7].icell.PUM Vbias 0.0031f
C1899 XA.XIR[9].XIC[5].icell.PDM Iout 0.00117f
C1900 XThR.XTBN.Y XA.XIR[7].XIC_dummy_left.icell.Ien 0.00158f
C1901 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9] 0.00341f
C1902 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.03425f
C1903 XA.XIR[1].XIC[3].icell.PDM Vbias 0.04261f
C1904 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02762f
C1905 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.SM 0.00168f
C1906 XThC.Tn[2] XThR.Tn[6] 0.28739f
C1907 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.SM 0.0039f
C1908 XThR.Tn[12] XThR.Tn[13] 0.06297f
C1909 XA.XIR[6].XIC[10].icell.SM Vbias 0.00701f
C1910 XA.XIR[9].XIC[11].icell.PUM VPWR 0.00937f
C1911 XA.XIR[13].XIC[12].icell.SM Iout 0.00388f
C1912 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C1913 XA.XIR[10].XIC[3].icell.SM VPWR 0.00158f
C1914 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00214f
C1915 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.SM 0.0039f
C1916 XA.XIR[4].XIC[3].icell.PDM Vbias 0.04261f
C1917 XThC.XTB5.A data[1] 0.11102f
C1918 XA.XIR[5].XIC[13].icell.Ien Vbias 0.21098f
C1919 XThC.XTB6.A a_5949_10571# 0.00467f
C1920 XA.XIR[0].XIC[4].icell.PUM VPWR 0.00882f
C1921 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04031f
C1922 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C1923 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00214f
C1924 XThR.Tn[10] XA.XIR[11].XIC[11].icell.SM 0.00121f
C1925 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.SM 0.0039f
C1926 XThC.Tn[4] XThR.Tn[11] 0.28739f
C1927 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04031f
C1928 XA.XIR[3].XIC[11].icell.PDM Vbias 0.04261f
C1929 XThC.XTB3.Y Vbias 0.01225f
C1930 XA.XIR[3].XIC[12].icell.SM VPWR 0.00158f
C1931 XA.XIR[8].XIC[13].icell.PDM Vbias 0.04261f
C1932 XA.XIR[4].XIC_dummy_right.icell.PUM Vbias 0.00223f
C1933 XA.XIR[14].XIC[4].icell.SM Vbias 0.00701f
C1934 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10] 0.00341f
C1935 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00214f
C1936 XThC.Tn[2] Vbias 2.61718f
C1937 XA.XIR[1].XIC[10].icell.PDM Iout 0.00117f
C1938 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.SM 0.00168f
C1939 XA.XIR[13].XIC[6].icell.SM Vbias 0.00701f
C1940 XA.XIR[3].XIC[8].icell.SM Iout 0.00388f
C1941 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[6].icell.SM 0.0039f
C1942 XA.XIR[6].XIC[13].icell.Ien Iout 0.06417f
C1943 XA.XIR[2].XIC[5].icell.SM VPWR 0.00158f
C1944 XA.XIR[8].XIC[10].icell.PUM Vbias 0.0031f
C1945 XA.XIR[11].XIC_15.icell.PDM Vbias 0.04401f
C1946 XA.XIR[10].XIC[14].icell.Ien Iout 0.06417f
C1947 XA.XIR[7].XIC[7].icell.PUM VPWR 0.00937f
C1948 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02762f
C1949 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PUM 0.00465f
C1950 VPWR data[2] 0.21031f
C1951 XThR.Tn[9] XA.XIR[10].XIC[14].icell.Ien 0.00338f
C1952 XA.XIR[11].XIC_15.icell.Ien Vbias 0.21234f
C1953 XA.XIR[12].XIC[8].icell.Ien Vbias 0.21098f
C1954 XA.XIR[1].XIC[7].icell.SM VPWR 0.00158f
C1955 XA.XIR[4].XIC[10].icell.PDM Iout 0.00117f
C1956 XA.XIR[2].XIC[1].icell.SM Iout 0.00388f
C1957 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00214f
C1958 XA.XIR[9].XIC_15.icell.SM VPWR 0.00275f
C1959 XA.XIR[6].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1960 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.SM 0.0039f
C1961 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.SM 0.00168f
C1962 XA.XIR[15].XIC[12].icell.PUM VPWR 0.00937f
C1963 XThC.XTB5.Y XThC.Tn[5] 0.01095f
C1964 XThC.Tn[0] XA.XIR[11].XIC_dummy_left.icell.Iout 0.00109f
C1965 a_10915_9569# XThC.Tn[14] 0.20278f
C1966 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38996f
C1967 XA.XIR[1].XIC[3].icell.SM Iout 0.00388f
C1968 XThC.Tn[8] XThR.Tn[13] 0.28739f
C1969 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.SM 0.00168f
C1970 XA.XIR[14].XIC[7].icell.Ien Iout 0.06417f
C1971 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.SM 0.0039f
C1972 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00584f
C1973 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0404f
C1974 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.04498f
C1975 XThC.XTB2.Y data[0] 0.00267f
C1976 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00214f
C1977 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PUM 0.00186f
C1978 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.15202f
C1979 XThC.Tn[7] XThR.Tn[1] 0.2877f
C1980 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C1981 XA.XIR[13].XIC[9].icell.Ien Iout 0.06417f
C1982 XA.XIR[14].XIC[10].icell.Ien Vbias 0.21098f
C1983 XA.XIR[8].XIC[11].icell.SM Iout 0.00388f
C1984 XA.XIR[0].XIC[12].icell.PUM Vbias 0.0031f
C1985 XThR.Tn[8] XA.XIR[9].XIC[11].icell.SM 0.00121f
C1986 XThC.Tn[11] Iout 0.84142f
C1987 XThC.Tn[11] XThR.Tn[9] 0.28739f
C1988 XThR.Tn[2] XA.XIR[3].XIC[6].icell.Ien 0.00338f
C1989 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C1990 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Iout 0.00347f
C1991 XThR.Tn[4] XA.XIR[4].XIC[3].icell.PDM 0.00341f
C1992 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.SM 0.0039f
C1993 XThR.Tn[4] XA.XIR[5].XIC[13].icell.Ien 0.00338f
C1994 XThC.Tn[7] XThR.Tn[12] 0.28739f
C1995 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02762f
C1996 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02762f
C1997 XThR.Tn[3] XA.XIR[4].XIC[13].icell.Ien 0.00338f
C1998 XThR.Tn[3] XA.XIR[3].XIC[4].icell.PDM 0.00341f
C1999 XA.XIR[2].XIC[13].icell.SM Vbias 0.00701f
C2000 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04052f
C2001 XA.XIR[7].XIC_15.icell.PUM Vbias 0.0031f
C2002 a_5155_9615# VPWR 0.7051f
C2003 XThR.Tn[1] XA.XIR[2].XIC[4].icell.SM 0.00121f
C2004 XA.XIR[6].XIC[0].icell.PDM VPWR 0.00799f
C2005 XThC.Tn[2] XThR.Tn[4] 0.28739f
C2006 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02762f
C2007 XThC.XTBN.Y XThC.Tn[5] 0.60785f
C2008 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04031f
C2009 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.SM 0.00168f
C2010 XA.XIR[15].XIC[13].icell.Ien VPWR 0.32895f
C2011 XA.XIR[0].XIC[13].icell.SM Iout 0.00367f
C2012 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00584f
C2013 XA.XIR[5].XIC[7].icell.PDM VPWR 0.00799f
C2014 XA.XIR[4].XIC[1].icell.Ien Vbias 0.21098f
C2015 XThR.Tn[13] XA.XIR[14].XIC[8].icell.SM 0.00121f
C2016 XA.XIR[13].XIC[2].icell.PUM Vbias 0.0031f
C2017 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.SM 0.0039f
C2018 XA.XIR[13].XIC[1].icell.PDM VPWR 0.00799f
C2019 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C2020 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.03425f
C2021 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.SM 0.0039f
C2022 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[14].icell.Ien 0.00214f
C2023 XA.XIR[13].XIC[10].icell.SM Iout 0.00388f
C2024 a_8963_9569# XA.XIR[0].XIC[10].icell.PDM 0.0029f
C2025 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C2026 XThR.XTB7.B XThR.XTB7.A 0.35833f
C2027 XThC.Tn[6] XThR.Tn[10] 0.28739f
C2028 XThC.XTB5.Y a_10051_9569# 0.00133f
C2029 XA.XIR[12].XIC[6].icell.PDM VPWR 0.00799f
C2030 XA.XIR[2].XIC_dummy_right.icell.SM VPWR 0.00123f
C2031 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02762f
C2032 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PUM 0.00465f
C2033 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00214f
C2034 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.SM 0.00168f
C2035 XThR.Tn[0] XA.XIR[1].XIC[11].icell.SM 0.00121f
C2036 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.SM 0.00168f
C2037 XA.XIR[5].XIC[1].icell.Ien Iout 0.06417f
C2038 XThR.Tn[10] XA.XIR[11].XIC[9].icell.SM 0.00121f
C2039 XThC.Tn[7] XThC.Tn[8] 0.07597f
C2040 XThC.XTB1.Y Vbias 0.01234f
C2041 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00214f
C2042 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.SM 0.00168f
C2043 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00584f
C2044 XThR.Tn[14] Iout 1.16234f
C2045 XA.XIR[11].XIC[0].icell.PDM Iout 0.00117f
C2046 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PUM 0.00465f
C2047 XA.XIR[15].XIC[3].icell.Ien Vbias 0.17899f
C2048 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.03425f
C2049 XA.XIR[5].XIC[3].icell.SM Vbias 0.00701f
C2050 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C2051 a_4861_9615# XThC.Tn[5] 0.00208f
C2052 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Ien 0.00549f
C2053 XA.XIR[8].XIC[2].icell.PUM VPWR 0.00937f
C2054 XThR.Tn[5] XA.XIR[6].XIC[13].icell.SM 0.00121f
C2055 XThR.Tn[6] XA.XIR[7].XIC[0].icell.Ien 0.00338f
C2056 XA.XIR[10].XIC[4].icell.PDM Iout 0.00117f
C2057 XA.XIR[10].XIC[12].icell.Ien Iout 0.06417f
C2058 XA.XIR[15].XIC[14].icell.SM VPWR 0.00207f
C2059 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04031f
C2060 XA.XIR[3].XIC[4].icell.PUM VPWR 0.00937f
C2061 XA.XIR[4].XIC[6].icell.Ien Vbias 0.21098f
C2062 XThR.Tn[9] XA.XIR[10].XIC[12].icell.Ien 0.00338f
C2063 XA.XIR[6].XIC[7].icell.SM VPWR 0.00158f
C2064 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PUM 0.00429f
C2065 XThC.XTB6.Y VPWR 1.03148f
C2066 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00584f
C2067 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C2068 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C2069 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.SM 0.00168f
C2070 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.1106f
C2071 XA.XIR[15].XIC[10].icell.PUM VPWR 0.00937f
C2072 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02762f
C2073 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00214f
C2074 XA.XIR[5].XIC[10].icell.Ien VPWR 0.1903f
C2075 XA.XIR[6].XIC[3].icell.SM Iout 0.00388f
C2076 XThC.XTBN.Y a_10051_9569# 0.23006f
C2077 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C2078 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C2079 XThR.XTB7.A XThR.Tn[2] 0.12549f
C2080 XA.XIR[3].XIC[2].icell.PDM VPWR 0.00799f
C2081 XA.XIR[9].XIC[13].icell.PDM Vbias 0.04261f
C2082 XA.XIR[4].XIC[13].icell.PUM VPWR 0.00937f
C2083 XA.XIR[5].XIC[6].icell.Ien Iout 0.06417f
C2084 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02762f
C2085 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.15202f
C2086 XThR.Tn[14] XA.XIR[15].XIC[0].icell.Ien 0.00377f
C2087 XA.XIR[8].XIC[4].icell.PDM VPWR 0.00799f
C2088 XA.XIR[14].XIC[1].icell.SM VPWR 0.00158f
C2089 XA.XIR[0].XIC[5].icell.PDM Vbias 0.04275f
C2090 XA.XIR[7].XIC[0].icell.Ien Vbias 0.20951f
C2091 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.15202f
C2092 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02762f
C2093 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.15202f
C2094 XA.XIR[2].XIC[8].icell.PDM VPWR 0.00799f
C2095 XA.XIR[13].XIC[3].icell.SM VPWR 0.00158f
C2096 XA.XIR[1].XIC[2].icell.PUM Vbias 0.0031f
C2097 XA.XIR[9].XIC[9].icell.Ien Vbias 0.21098f
C2098 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00214f
C2099 XA.XIR[8].XIC[7].icell.PUM VPWR 0.00937f
C2100 XA.XIR[10].XIC[3].icell.PUM Vbias 0.0031f
C2101 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00214f
C2102 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.02762f
C2103 XThR.Tn[6] XA.XIR[7].XIC[5].icell.Ien 0.00338f
C2104 XA.XIR[12].XIC[5].icell.Ien VPWR 0.1903f
C2105 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C2106 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12] 0.00341f
C2107 XA.XIR[0].XIC[2].icell.Ien Vbias 0.2113f
C2108 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.03425f
C2109 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00584f
C2110 XThC.Tn[4] XThR.Tn[14] 0.28739f
C2111 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C2112 XA.XIR[11].XIC[14].icell.PDM Vbias 0.04261f
C2113 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.SM 0.00168f
C2114 XA.XIR[11].XIC[6].icell.SM VPWR 0.00158f
C2115 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04031f
C2116 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.SM 0.00168f
C2117 XA.XIR[3].XIC[12].icell.PUM Vbias 0.0031f
C2118 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.0353f
C2119 XThR.Tn[4] XA.XIR[5].XIC[3].icell.SM 0.00121f
C2120 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02762f
C2121 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Iout 0.00347f
C2122 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2123 XA.XIR[11].XIC[2].icell.SM Iout 0.00388f
C2124 XA.XIR[10].XIC[8].icell.SM VPWR 0.00158f
C2125 XA.XIR[15].XIC[11].icell.Ien VPWR 0.32895f
C2126 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00584f
C2127 XThR.Tn[3] XA.XIR[4].XIC[3].icell.SM 0.00121f
C2128 XA.XIR[14].XIC_15.icell.PDM Vbias 0.04401f
C2129 XThC.XTB7.B data[2] 0.07481f
C2130 XThR.Tn[14] XA.XIR[15].XIC[5].icell.Ien 0.00338f
C2131 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02762f
C2132 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.15202f
C2133 XA.XIR[13].XIC[14].icell.Ien Iout 0.06417f
C2134 XA.XIR[2].XIC[5].icell.PUM Vbias 0.0031f
C2135 XA.XIR[14].XIC_15.icell.Ien Vbias 0.21234f
C2136 XThC.XTB4.Y VPWR 0.91479f
C2137 XA.XIR[10].XIC[4].icell.SM Iout 0.00388f
C2138 XA.XIR[7].XIC[5].icell.Ien Vbias 0.21098f
C2139 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.03431f
C2140 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C2141 XThC.XTB2.Y XThC.Tn[0] 0.00125f
C2142 XThR.Tn[9] XA.XIR[10].XIC[4].icell.SM 0.00121f
C2143 XA.XIR[0].XIC[9].icell.PUM VPWR 0.00877f
C2144 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00214f
C2145 XA.XIR[12].XIC_15.icell.SM VPWR 0.00275f
C2146 XA.XIR[1].XIC[7].icell.PUM Vbias 0.0031f
C2147 XThC.Tn[0] XA.XIR[14].XIC_dummy_left.icell.Iout 0.00109f
C2148 XThR.Tn[10] XA.XIR[11].XIC[13].icell.Ien 0.00338f
C2149 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04031f
C2150 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C2151 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C2152 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00214f
C2153 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.SM 0.0039f
C2154 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C2155 XA.XIR[3].XIC[13].icell.SM Iout 0.00388f
C2156 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04031f
C2157 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.04591f
C2158 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8] 0.00341f
C2159 XA.XIR[2].XIC[10].icell.SM VPWR 0.00158f
C2160 XA.XIR[7].XIC[12].icell.PUM VPWR 0.00937f
C2161 XA.XIR[8].XIC_15.icell.PUM Vbias 0.0031f
C2162 XThR.XTB5.A VPWR 0.83112f
C2163 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00214f
C2164 XA.XIR[2].XIC[6].icell.SM Iout 0.00388f
C2165 XA.XIR[1].XIC[12].icell.SM VPWR 0.00158f
C2166 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.SM 0.00168f
C2167 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04031f
C2168 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.04036f
C2169 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C2170 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PUM 0.00465f
C2171 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PUM 0.00465f
C2172 XThR.Tn[12] XA.XIR[13].XIC[2].icell.SM 0.00121f
C2173 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2174 XA.XIR[1].XIC[8].icell.SM Iout 0.00388f
C2175 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C2176 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.SM 0.00168f
C2177 XA.XIR[10].XIC[10].icell.Ien Iout 0.06417f
C2178 XThR.Tn[13] XA.XIR[14].XIC[13].icell.SM 0.00121f
C2179 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00584f
C2180 XThR.Tn[9] XA.XIR[10].XIC[10].icell.Ien 0.00338f
C2181 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02762f
C2182 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.15202f
C2183 XA.XIR[3].XIC[1].icell.PUM VPWR 0.00937f
C2184 XThC.XTB7.B a_5155_9615# 0.00268f
C2185 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Ien 0.00584f
C2186 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.15202f
C2187 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PUM 0.00465f
C2188 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00584f
C2189 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02762f
C2190 XThR.Tn[11] XA.XIR[12].XIC[5].icell.SM 0.00121f
C2191 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02762f
C2192 a_2979_9615# Vbias 0.00736f
C2193 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C2194 XThC.XTB6.Y a_9827_9569# 0.00871f
C2195 XThR.Tn[10] XA.XIR[11].XIC[14].icell.SM 0.00121f
C2196 XThR.Tn[2] XA.XIR[3].XIC[11].icell.Ien 0.00338f
C2197 XA.XIR[11].XIC[2].icell.PUM VPWR 0.00937f
C2198 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C2199 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.SM 0.00168f
C2200 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PDM 0.00172f
C2201 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2202 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04031f
C2203 XA.XIR[5].XIC[3].icell.PDM Vbias 0.04261f
C2204 XA.XIR[7].XIC[8].icell.PDM VPWR 0.00799f
C2205 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.03425f
C2206 XThR.XTB3.Y XThR.Tn[9] 0.00285f
C2207 XA.XIR[9].XIC[1].icell.Ien VPWR 0.1903f
C2208 XA.XIR[6].XIC[2].icell.PUM Vbias 0.0031f
C2209 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.15202f
C2210 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.SM 0.0039f
C2211 XThC.Tn[6] XThR.Tn[13] 0.28739f
C2212 a_4067_9615# XThC.Tn[1] 0.00584f
C2213 XA.XIR[4].XIC[3].icell.Ien VPWR 0.1903f
C2214 XThR.Tn[1] XA.XIR[2].XIC[9].icell.SM 0.00121f
C2215 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07214f
C2216 VPWR data[5] 0.4402f
C2217 XA.XIR[15].XIC[6].icell.PDM VPWR 0.0114f
C2218 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.SM 0.00168f
C2219 XA.XIR[12].XIC[2].icell.PDM Vbias 0.04261f
C2220 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PUM 0.00179f
C2221 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.03023f
C2222 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C2223 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.SM 0.0039f
C2224 XThC.Tn[0] Iout 0.82523f
C2225 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C2226 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C2227 XThC.Tn[0] XThR.Tn[9] 0.28741f
C2228 XA.XIR[6].XIC[3].icell.PDM Iout 0.00117f
C2229 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00214f
C2230 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.SM 0.00168f
C2231 XA.XIR[11].XIC[8].icell.PDM Vbias 0.04261f
C2232 XA.XIR[14].XIC[0].icell.PDM Iout 0.00117f
C2233 XA.XIR[5].XIC[10].icell.PDM Iout 0.00117f
C2234 XThR.XTB5.Y a_n997_3755# 0.00418f
C2235 XThC.Tn[5] XThR.Tn[8] 0.28739f
C2236 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C2237 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C2238 XA.XIR[9].XIC[4].icell.PDM VPWR 0.00799f
C2239 a_7875_9569# VPWR 0.00639f
C2240 XA.XIR[13].XIC[4].icell.PDM Iout 0.00117f
C2241 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PUM 0.00465f
C2242 XA.XIR[13].XIC[12].icell.Ien Iout 0.06417f
C2243 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.SM 0.00168f
C2244 XThC.XTB2.Y VPWR 0.97668f
C2245 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.03425f
C2246 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PUM 0.00102f
C2247 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00214f
C2248 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.03425f
C2249 XA.XIR[3].XIC[2].icell.Ien Vbias 0.21098f
C2250 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C2251 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C2252 XThR.XTB7.A XThR.Tn[10] 0.00404f
C2253 XA.XIR[12].XIC[9].icell.PDM Iout 0.00117f
C2254 XA.XIR[6].XIC[7].icell.PUM Vbias 0.0031f
C2255 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.1106f
C2256 XA.XIR[9].XIC[6].icell.Ien VPWR 0.1903f
C2257 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.03023f
C2258 XThR.Tn[10] XA.XIR[11].XIC[11].icell.Ien 0.00338f
C2259 XA.XIR[15].XIC[8].icell.Ien Vbias 0.17899f
C2260 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PUM 0.00429f
C2261 XA.XIR[9].XIC[2].icell.Ien Iout 0.06417f
C2262 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.15202f
C2263 XA.XIR[5].XIC[8].icell.SM Vbias 0.00701f
C2264 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C2265 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00214f
C2266 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C2267 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02762f
C2268 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PUM 0.00465f
C2269 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04031f
C2270 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00584f
C2271 XA.XIR[4].XIC[11].icell.Ien Vbias 0.21098f
C2272 XA.XIR[3].XIC[9].icell.PUM VPWR 0.00937f
C2273 XThR.XTB5.Y a_n1049_5611# 0.0093f
C2274 XA.XIR[8].XIC[0].icell.PDM Vbias 0.04207f
C2275 XThC.XTB3.Y XThC.Tn[2] 0.1864f
C2276 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Ien 0.00584f
C2277 XA.XIR[1].XIC[9].icell.PDM VPWR 0.00799f
C2278 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02852f
C2279 XA.XIR[6].XIC[12].icell.SM VPWR 0.00158f
C2280 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.SM 0.0039f
C2281 XA.XIR[10].XIC[13].icell.SM VPWR 0.00158f
C2282 XA.XIR[11].XIC[13].icell.PDM Vbias 0.04261f
C2283 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C2284 XA.XIR[2].XIC[4].icell.PDM Vbias 0.04261f
C2285 XA.XIR[13].XIC[3].icell.PUM Vbias 0.0031f
C2286 XThC.Tn[1] XThC.Tn[3] 0.10977f
C2287 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00214f
C2288 XA.XIR[6].XIC[8].icell.SM Iout 0.00388f
C2289 XA.XIR[7].XIC[2].icell.Ien VPWR 0.1903f
C2290 XA.XIR[8].XIC[5].icell.Ien Vbias 0.21098f
C2291 XA.XIR[4].XIC[9].icell.PDM VPWR 0.00799f
C2292 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02762f
C2293 XA.XIR[5].XIC_15.icell.Ien VPWR 0.25566f
C2294 data[1] data[0] 0.64735f
C2295 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7] 0.00341f
C2296 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04031f
C2297 XThC.Tn[6] XThC.Tn[7] 0.1602f
C2298 XThR.Tn[13] XA.XIR[14].XIC[11].icell.SM 0.00121f
C2299 XA.XIR[12].XIC[3].icell.SM Vbias 0.00701f
C2300 XA.XIR[1].XIC[4].icell.PUM VPWR 0.00937f
C2301 XA.XIR[5].XIC[11].icell.Ien Iout 0.06417f
C2302 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.SM 0.0039f
C2303 XA.XIR[14].XIC[14].icell.PDM Vbias 0.04261f
C2304 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C2305 XA.XIR[14].XIC[6].icell.SM VPWR 0.00158f
C2306 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13] 0.00341f
C2307 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00214f
C2308 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C2309 XA.XIR[11].XIC[6].icell.PUM Vbias 0.0031f
C2310 Vbias bias[2] 0.05684f
C2311 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07214f
C2312 XA.XIR[3].XIC[5].icell.PDM Iout 0.00117f
C2313 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PUM 0.00465f
C2314 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2315 XA.XIR[14].XIC[2].icell.SM Iout 0.00388f
C2316 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02762f
C2317 XA.XIR[8].XIC[7].icell.PDM Iout 0.00117f
C2318 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C2319 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04031f
C2320 XA.XIR[13].XIC[8].icell.SM VPWR 0.00158f
C2321 XA.XIR[8].XIC[12].icell.PUM VPWR 0.00937f
C2322 XA.XIR[9].XIC[14].icell.Ien Vbias 0.21098f
C2323 XA.XIR[10].XIC[8].icell.PUM Vbias 0.0031f
C2324 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C2325 XA.XIR[2].XIC[11].icell.PDM Iout 0.00117f
C2326 XA.XIR[13].XIC[4].icell.SM Iout 0.00388f
C2327 XThR.Tn[6] XA.XIR[7].XIC[10].icell.Ien 0.00338f
C2328 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00584f
C2329 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00214f
C2330 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.SM 0.0039f
C2331 XA.XIR[0].XIC[7].icell.Ien Vbias 0.21134f
C2332 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C2333 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PUM 0.00465f
C2334 XThC.Tn[8] XThR.Tn[7] 0.28739f
C2335 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.SM 0.00168f
C2336 XA.XIR[12].XIC[6].icell.Ien Iout 0.06417f
C2337 XThR.Tn[0] XA.XIR[0].XIC[8].icell.PDM 0.00341f
C2338 XThR.Tn[2] XA.XIR[3].XIC[1].icell.SM 0.00121f
C2339 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00214f
C2340 XThR.Tn[4] XA.XIR[5].XIC[8].icell.SM 0.00121f
C2341 XThR.Tn[1] XA.XIR[1].XIC[6].icell.PDM 0.00341f
C2342 XA.XIR[10].XIC_15.icell.Ien Iout 0.0642f
C2343 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.SM 0.0039f
C2344 VPWR Iout 54.1536f
C2345 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04031f
C2346 XThC.XTB7.Y XThC.Tn[10] 0.07406f
C2347 XA.XIR[11].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2348 XA.XIR[11].XIC[7].icell.SM Iout 0.00388f
C2349 XThR.Tn[9] XA.XIR[10].XIC_15.icell.Ien 0.00117f
C2350 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.SM 0.00168f
C2351 XThR.Tn[9] VPWR 7.55029f
C2352 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04031f
C2353 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2354 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C2355 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.15202f
C2356 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C2357 XThR.Tn[3] XA.XIR[4].XIC[8].icell.SM 0.00121f
C2358 XA.XIR[2].XIC[10].icell.PUM Vbias 0.0031f
C2359 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00214f
C2360 XA.XIR[7].XIC[10].icell.Ien Vbias 0.21098f
C2361 XA.XIR[0].XIC[14].icell.PUM VPWR 0.00877f
C2362 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.15202f
C2363 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00214f
C2364 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.SM 0.00168f
C2365 XA.XIR[14].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2366 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.15202f
C2367 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5] 0.00341f
C2368 XA.XIR[1].XIC[12].icell.PUM Vbias 0.0031f
C2369 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Ien 0.0016f
C2370 XA.XIR[12].XIC[0].icell.PUM VPWR 0.00937f
C2371 XThR.Tn[2] XA.XIR[2].XIC[3].icell.PDM 0.00341f
C2372 XA.XIR[13].XIC[10].icell.Ien Iout 0.06417f
C2373 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C2374 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04031f
C2375 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[11].icell.SM 0.0039f
C2376 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04052f
C2377 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PUM 0.00465f
C2378 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00584f
C2379 XA.XIR[8].XIC[0].icell.Ien Vbias 0.20951f
C2380 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.15202f
C2381 XA.XIR[15].XIC[0].icell.Ien VPWR 0.32895f
C2382 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6] 0.00341f
C2383 XA.XIR[5].XIC[0].icell.SM VPWR 0.00158f
C2384 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C2385 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.03425f
C2386 XA.XIR[2].XIC[11].icell.SM Iout 0.00388f
C2387 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C2388 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.SM 0.0039f
C2389 XA.XIR[14].XIC[2].icell.PUM VPWR 0.00937f
C2390 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C2391 XThR.Tn[12] XA.XIR[13].XIC[7].icell.SM 0.00121f
C2392 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C2393 XA.XIR[1].XIC[13].icell.SM Iout 0.00388f
C2394 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.SM 0.00168f
C2395 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02762f
C2396 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.15202f
C2397 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00214f
C2398 XA.XIR[7].XIC[4].icell.PDM Vbias 0.04261f
C2399 XA.XIR[10].XIC[3].icell.PDM VPWR 0.00799f
C2400 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C2401 XThC.Tn[4] VPWR 5.88871f
C2402 XA.XIR[10].XIC[11].icell.SM VPWR 0.00158f
C2403 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PUM 0.00465f
C2404 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.15202f
C2405 XA.XIR[4].XIC[1].icell.SM Vbias 0.00701f
C2406 XA.XIR[15].XIC[2].icell.PDM Vbias 0.04261f
C2407 XA.XIR[6].XIC[11].icell.PDM Vbias 0.04261f
C2408 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C2409 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C2410 XThR.Tn[13] XA.XIR[14].XIC[9].icell.SM 0.00121f
C2411 XA.XIR[12].XIC[0].icell.SM Iout 0.00388f
C2412 XA.XIR[6].XIC[4].icell.PUM VPWR 0.00937f
C2413 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PUM 0.00465f
C2414 XA.XIR[14].XIC[8].icell.PDM Vbias 0.04261f
C2415 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C2416 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.SM 0.0039f
C2417 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Ien 0.00309f
C2418 XThC.Tn[10] XThR.Tn[0] 0.28747f
C2419 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Iout 0.00347f
C2420 XA.XIR[15].XIC[5].icell.Ien VPWR 0.32895f
C2421 XThC.Tn[12] XThR.Tn[5] 0.28739f
C2422 XA.XIR[5].XIC[5].icell.SM VPWR 0.00158f
C2423 XThR.XTB7.B XThR.Tn[10] 0.06102f
C2424 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.15202f
C2425 XThC.XTB7.B a_7875_9569# 0.01174f
C2426 XThR.Tn[1] XA.XIR[2].XIC[14].icell.SM 0.00121f
C2427 XA.XIR[7].XIC[11].icell.PDM Iout 0.00117f
C2428 XA.XIR[4].XIC[8].icell.Ien VPWR 0.1903f
C2429 XA.XIR[9].XIC[0].icell.PDM Vbias 0.04207f
C2430 XA.XIR[5].XIC[1].icell.SM Iout 0.00388f
C2431 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C2432 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.SM 0.00168f
C2433 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C2434 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.SM 0.0039f
C2435 XA.XIR[15].XIC[9].icell.PDM Iout 0.00117f
C2436 XA.XIR[4].XIC[4].icell.Ien Iout 0.06417f
C2437 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.SM 0.0039f
C2438 a_8963_9569# XThC.Tn[11] 0.19413f
C2439 XA.XIR[9].XIC[4].icell.SM Vbias 0.00701f
C2440 XA.XIR[8].XIC[2].icell.Ien VPWR 0.1903f
C2441 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PUM 0.00465f
C2442 XA.XIR[10].XIC[14].icell.PUM VPWR 0.00937f
C2443 XA.XIR[11].XIC[12].icell.PDM Vbias 0.04261f
C2444 XA.XIR[15].XIC_15.icell.SM VPWR 0.00275f
C2445 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C2446 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PUM 0.00465f
C2447 XThR.Tn[2] XThR.XTB4.Y 0.0021f
C2448 XA.XIR[2].XIC[2].icell.PUM VPWR 0.00937f
C2449 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.15202f
C2450 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.SM 0.00168f
C2451 XA.XIR[0].XIC[11].icell.PDM VPWR 0.00774f
C2452 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.03591f
C2453 XA.XIR[11].XIC[3].icell.PUM VPWR 0.00937f
C2454 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00214f
C2455 XA.XIR[3].XIC[7].icell.Ien Vbias 0.21098f
C2456 XA.XIR[9].XIC[7].icell.PDM Iout 0.00117f
C2457 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00214f
C2458 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9] 0.00341f
C2459 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C2460 XA.XIR[1].XIC[5].icell.PDM Vbias 0.04261f
C2461 XA.XIR[13].XIC[13].icell.SM VPWR 0.00158f
C2462 XA.XIR[14].XIC[13].icell.PDM Vbias 0.04261f
C2463 XA.XIR[6].XIC[12].icell.PUM Vbias 0.0031f
C2464 XThR.XTBN.Y XA.XIR[0].XIC_dummy_left.icell.Iout 0.00137f
C2465 XA.XIR[9].XIC[11].icell.Ien VPWR 0.1903f
C2466 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00584f
C2467 XA.XIR[10].XIC[5].icell.PUM VPWR 0.00937f
C2468 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11] 0.00341f
C2469 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C2470 XA.XIR[12].XIC[14].icell.PDM VPWR 0.00809f
C2471 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C2472 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02762f
C2473 XA.XIR[4].XIC[5].icell.PDM Vbias 0.04261f
C2474 XA.XIR[5].XIC[13].icell.SM Vbias 0.00701f
C2475 XA.XIR[9].XIC[7].icell.Ien Iout 0.06417f
C2476 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PUM 0.00465f
C2477 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.15202f
C2478 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18982f
C2479 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04031f
C2480 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C2481 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.SM 0.00168f
C2482 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PUM 0.00465f
C2483 XA.XIR[1].XIC[2].icell.Ien Vbias 0.21104f
C2484 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04031f
C2485 XA.XIR[3].XIC[13].icell.PDM Vbias 0.04261f
C2486 XA.XIR[14].XIC[6].icell.PUM Vbias 0.0031f
C2487 XA.XIR[8].XIC_15.icell.PDM Vbias 0.04401f
C2488 XA.XIR[3].XIC[14].icell.PUM VPWR 0.00937f
C2489 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02762f
C2490 XThC.Tn[9] XThR.Tn[2] 0.28739f
C2491 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C2492 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07555f
C2493 XA.XIR[1].XIC[12].icell.PDM Iout 0.00117f
C2494 XA.XIR[13].XIC[8].icell.PUM Vbias 0.0031f
C2495 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C2496 XA.XIR[8].XIC[10].icell.Ien Vbias 0.21098f
C2497 XA.XIR[7].XIC[7].icell.Ien VPWR 0.1903f
C2498 XA.XIR[6].XIC[13].icell.SM Iout 0.00388f
C2499 XA.XIR[2].XIC[7].icell.PUM VPWR 0.00937f
C2500 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.03425f
C2501 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04031f
C2502 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C2503 XA.XIR[12].XIC[8].icell.SM Vbias 0.00701f
C2504 XA.XIR[4].XIC[12].icell.PDM Iout 0.00117f
C2505 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01444f
C2506 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C2507 XA.XIR[5].XIC_dummy_right.icell.SM VPWR 0.00123f
C2508 XA.XIR[1].XIC[9].icell.PUM VPWR 0.00937f
C2509 XA.XIR[7].XIC[3].icell.Ien Iout 0.06417f
C2510 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C2511 XA.XIR[10].XIC[9].icell.SM VPWR 0.00158f
C2512 XThR.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.00338f
C2513 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02762f
C2514 XA.XIR[13].XIC_15.icell.Ien Iout 0.0642f
C2515 XThC.XTB7.B Iout 0.00967f
C2516 XA.XIR[14].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2517 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C2518 XA.XIR[14].XIC[7].icell.SM Iout 0.00388f
C2519 XThC.XTB7.A XThC.Tn[5] 0.02758f
C2520 XThR.Tn[7] XA.XIR[8].XIC[4].icell.Ien 0.00338f
C2521 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PUM 0.00465f
C2522 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38919f
C2523 XThR.Tn[6] XA.XIR[7].XIC_15.icell.Ien 0.00117f
C2524 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.SM 0.00168f
C2525 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00256f
C2526 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C2527 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C2528 XA.XIR[0].XIC[12].icell.Ien Vbias 0.2113f
C2529 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.04036f
C2530 XA.XIR[15].XIC_dummy_left.icell.SM VPWR 0.00269f
C2531 XThR.Tn[2] XA.XIR[3].XIC[6].icell.SM 0.00121f
C2532 XThR.XTB7.B a_n997_1803# 0.00228f
C2533 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.15202f
C2534 XThR.Tn[4] XA.XIR[4].XIC[5].icell.PDM 0.00341f
C2535 XThR.Tn[4] XA.XIR[5].XIC[13].icell.SM 0.00121f
C2536 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.03425f
C2537 XThC.Tn[14] XThR.Tn[6] 0.28745f
C2538 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.15202f
C2539 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PUM 0.00465f
C2540 XThR.Tn[10] XA.XIR[11].XIC[5].icell.Ien 0.00338f
C2541 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00584f
C2542 XThR.Tn[3] XA.XIR[3].XIC[6].icell.PDM 0.00341f
C2543 XThR.Tn[3] XA.XIR[4].XIC[13].icell.SM 0.00121f
C2544 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PUM 0.00465f
C2545 a_6243_9615# VPWR 0.70553f
C2546 XA.XIR[2].XIC_15.icell.PUM Vbias 0.0031f
C2547 XA.XIR[7].XIC_15.icell.Ien Vbias 0.21234f
C2548 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.15202f
C2549 XA.XIR[6].XIC[2].icell.PDM VPWR 0.00799f
C2550 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.03425f
C2551 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.15202f
C2552 VPWR data[1] 0.44103f
C2553 XA.XIR[5].XIC[0].icell.Ien Vbias 0.20951f
C2554 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04031f
C2555 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C2556 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C2557 XThR.Tn[13] XA.XIR[14].XIC[14].icell.SM 0.00121f
C2558 XA.XIR[10].XIC[12].icell.PUM VPWR 0.00937f
C2559 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C2560 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02762f
C2561 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.15202f
C2562 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.SM 0.00168f
C2563 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C2564 XA.XIR[5].XIC[9].icell.PDM VPWR 0.00799f
C2565 XA.XIR[14].XIC[1].icell.PUM Vbias 0.0031f
C2566 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02762f
C2567 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C2568 XThC.Tn[6] XThR.Tn[7] 0.28739f
C2569 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00214f
C2570 XThC.Tn[14] Vbias 2.45788f
C2571 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00214f
C2572 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Iout 0.00347f
C2573 XA.XIR[13].XIC[3].icell.PDM VPWR 0.00799f
C2574 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.SM 0.00168f
C2575 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.15202f
C2576 XA.XIR[13].XIC[11].icell.SM VPWR 0.00158f
C2577 XThC.XTB7.B XThC.Tn[4] 0.00356f
C2578 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PUM 0.00268f
C2579 a_9827_9569# XA.XIR[0].XIC[11].icell.PDM 0.00136f
C2580 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.0284f
C2581 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C2582 XThC.XTB5.Y XThC.Tn[8] 0.01728f
C2583 XThC.XTB7.Y a_7651_9569# 0.00477f
C2584 XThR.XTB1.Y data[4] 0.06453f
C2585 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02762f
C2586 XA.XIR[12].XIC[8].icell.PDM VPWR 0.00799f
C2587 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C2588 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C2589 XThR.XTB5.Y a_n997_2667# 0.00427f
C2590 XThC.XTB6.A a_5155_10571# 0.00306f
C2591 XA.XIR[15].XIC[1].icell.Ien Iout 0.06807f
C2592 XThC.XTB6.Y XThC.Tn[12] 0.02863f
C2593 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C2594 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C2595 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.0353f
C2596 XA.XIR[6].XIC[2].icell.Ien Vbias 0.21098f
C2597 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.03425f
C2598 XA.XIR[9].XIC[1].icell.SM VPWR 0.00158f
C2599 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00214f
C2600 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C2601 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00584f
C2602 XThR.XTB7.B XThR.Tn[13] 0.00276f
C2603 XThC.Tn[10] XThR.Tn[1] 0.28739f
C2604 XA.XIR[15].XIC[3].icell.SM Vbias 0.00701f
C2605 XA.XIR[11].XIC[2].icell.PDM Iout 0.00117f
C2606 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02762f
C2607 XA.XIR[5].XIC[5].icell.PUM Vbias 0.0031f
C2608 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.03425f
C2609 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.SM 0.0039f
C2610 a_5949_9615# XThC.Tn[5] 0.27124f
C2611 XThR.Tn[6] XA.XIR[7].XIC[0].icell.SM 0.00121f
C2612 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PUM 0.00186f
C2613 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00214f
C2614 XA.XIR[4].XIC[6].icell.SM Vbias 0.00701f
C2615 XA.XIR[10].XIC[6].icell.PDM Iout 0.00117f
C2616 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04031f
C2617 XA.XIR[3].XIC[4].icell.Ien VPWR 0.1903f
C2618 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2619 XA.XIR[10].XIC[13].icell.Ien VPWR 0.1903f
C2620 XA.XIR[11].XIC[11].icell.PDM Vbias 0.04261f
C2621 XThC.Tn[10] XThR.Tn[12] 0.28739f
C2622 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C2623 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02762f
C2624 XA.XIR[6].XIC[9].icell.PUM VPWR 0.00937f
C2625 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C2626 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C2627 XThR.Tn[13] XA.XIR[14].XIC[11].icell.Ien 0.00338f
C2628 XA.XIR[5].XIC[10].icell.SM VPWR 0.00158f
C2629 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7] 0.00341f
C2630 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00214f
C2631 XThR.Tn[4] XA.XIR[5].XIC[0].icell.Ien 0.00338f
C2632 XA.XIR[13].XIC[14].icell.PUM VPWR 0.00937f
C2633 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.15202f
C2634 XA.XIR[14].XIC[12].icell.PDM Vbias 0.04261f
C2635 XThC.XTBN.Y XThC.Tn[8] 0.50311f
C2636 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00214f
C2637 XThC.Tn[5] XThR.Tn[3] 0.28739f
C2638 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PUM 0.00465f
C2639 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C2640 XA.XIR[15].XIC[6].icell.Ien Iout 0.06807f
C2641 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C2642 XA.XIR[5].XIC[6].icell.SM Iout 0.00388f
C2643 XA.XIR[8].XIC[6].icell.PDM VPWR 0.00799f
C2644 XA.XIR[12].XIC[13].icell.PDM VPWR 0.00799f
C2645 XThR.Tn[14] XA.XIR[15].XIC[0].icell.SM 0.00128f
C2646 XA.XIR[4].XIC[13].icell.Ien VPWR 0.1903f
C2647 XA.XIR[3].XIC[4].icell.PDM VPWR 0.00799f
C2648 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.04563f
C2649 XA.XIR[9].XIC_15.icell.PDM Vbias 0.04401f
C2650 XThC.XTB1.Y a_2979_9615# 0.21263f
C2651 XThC.Tn[14] XThR.Tn[4] 0.28745f
C2652 XA.XIR[7].XIC[0].icell.SM Vbias 0.00675f
C2653 XA.XIR[14].XIC[3].icell.PUM VPWR 0.00937f
C2654 XA.XIR[0].XIC[7].icell.PDM Vbias 0.04278f
C2655 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.SM 0.0039f
C2656 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.SM 0.0039f
C2657 XA.XIR[4].XIC[9].icell.Ien Iout 0.06417f
C2658 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.SM 0.00168f
C2659 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C2660 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.04498f
C2661 XA.XIR[2].XIC[10].icell.PDM VPWR 0.00799f
C2662 XThC.Tn[0] XA.XIR[9].XIC_dummy_left.icell.Iout 0.00109f
C2663 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02762f
C2664 XA.XIR[13].XIC[5].icell.PUM VPWR 0.00937f
C2665 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04037f
C2666 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C2667 XA.XIR[9].XIC[9].icell.SM Vbias 0.00701f
C2668 XA.XIR[0].XIC[0].icell.Ien Iout 0.06382f
C2669 XA.XIR[8].XIC[7].icell.Ien VPWR 0.1903f
C2670 XA.XIR[10].XIC[3].icell.Ien Vbias 0.21098f
C2671 XThC.XTB4.Y XThC.Tn[12] 0.00209f
C2672 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01149f
C2673 XThR.Tn[6] XA.XIR[7].XIC[5].icell.SM 0.00121f
C2674 XThC.Tn[9] XThR.Tn[10] 0.28739f
C2675 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C2676 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.SM 0.0039f
C2677 XThC.Tn[1] XThR.Tn[5] 0.28739f
C2678 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.SM 0.00168f
C2679 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12] 0.00341f
C2680 XA.XIR[12].XIC[5].icell.SM VPWR 0.00158f
C2681 XA.XIR[12].XIC[13].icell.SM Vbias 0.00701f
C2682 XA.XIR[8].XIC[3].icell.Ien Iout 0.06417f
C2683 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.15202f
C2684 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02762f
C2685 XA.XIR[0].XIC[2].icell.SM Vbias 0.00716f
C2686 XThR.Tn[8] XA.XIR[9].XIC[3].icell.Ien 0.00338f
C2687 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C2688 XA.XIR[12].XIC[1].icell.SM Iout 0.00388f
C2689 XA.XIR[10].XIC[14].icell.SM VPWR 0.00207f
C2690 XA.XIR[11].XIC[8].icell.PUM VPWR 0.00937f
C2691 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C2692 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00214f
C2693 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02762f
C2694 XThC.Tn[8] XThC.Tn[10] 0.00465f
C2695 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04031f
C2696 XA.XIR[3].XIC[12].icell.Ien Vbias 0.21098f
C2697 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.SM 0.0039f
C2698 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2699 XThC.Tn[13] XThC.Tn[14] 0.38789f
C2700 XA.XIR[10].XIC[10].icell.PUM VPWR 0.00937f
C2701 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PUM 0.00465f
C2702 XThR.Tn[14] XA.XIR[15].XIC[5].icell.SM 0.00121f
C2703 XA.XIR[2].XIC[5].icell.Ien Vbias 0.21098f
C2704 XA.XIR[9].XIC[12].icell.Ien Iout 0.06417f
C2705 XA.XIR[7].XIC[5].icell.SM Vbias 0.00701f
C2706 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.SM 0.00168f
C2707 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.15202f
C2708 XA.XIR[0].XIC[9].icell.Ien VPWR 0.19115f
C2709 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.SM 0.0039f
C2710 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00214f
C2711 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2712 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02762f
C2713 XA.XIR[13].XIC[9].icell.SM VPWR 0.00158f
C2714 XA.XIR[1].XIC[7].icell.Ien Vbias 0.21104f
C2715 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C2716 XA.XIR[0].XIC[5].icell.Ien Iout 0.06389f
C2717 XThR.Tn[5] XA.XIR[6].XIC[0].icell.Ien 0.00338f
C2718 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04031f
C2719 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04031f
C2720 XThR.XTBN.Y a_n997_1803# 0.22873f
C2721 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04031f
C2722 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8] 0.00341f
C2723 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00214f
C2724 XA.XIR[8].XIC_15.icell.Ien Vbias 0.21234f
C2725 XA.XIR[7].XIC[12].icell.Ien VPWR 0.1903f
C2726 XA.XIR[2].XIC[12].icell.PUM VPWR 0.00937f
C2727 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C2728 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00584f
C2729 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.15202f
C2730 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00214f
C2731 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PUM 0.00465f
C2732 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00584f
C2733 XA.XIR[1].XIC[14].icell.PUM VPWR 0.00937f
C2734 XThR.Tn[0] XA.XIR[1].XIC[3].icell.Ien 0.00338f
C2735 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.SM 0.0039f
C2736 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04031f
C2737 XA.XIR[7].XIC[8].icell.Ien Iout 0.06417f
C2738 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.03425f
C2739 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C2740 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.03425f
C2741 XThR.XTB6.A a_n997_3755# 0.00149f
C2742 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C2743 XA.XIR[10].XIC[11].icell.Ien VPWR 0.1903f
C2744 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C2745 XThR.Tn[7] XA.XIR[8].XIC[9].icell.Ien 0.00338f
C2746 XA.XIR[3].XIC[1].icell.Ien VPWR 0.1903f
C2747 XThC.XTB7.B a_6243_9615# 0.01743f
C2748 XThC.Tn[7] XThR.Tn[2] 0.28746f
C2749 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.SM 0.0039f
C2750 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PUM 0.00465f
C2751 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00256f
C2752 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PUM 0.00465f
C2753 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02762f
C2754 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00214f
C2755 a_4067_9615# Vbias 0.00573f
C2756 XThC.XTB7.B data[1] 0.00593f
C2757 XA.XIR[12].XIC[1].icell.PUM VPWR 0.00937f
C2758 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C2759 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C2760 XThR.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.00338f
C2761 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PUM 0.00465f
C2762 XA.XIR[13].XIC[12].icell.PUM VPWR 0.00937f
C2763 XThR.Tn[2] XA.XIR[3].XIC[11].icell.SM 0.00121f
C2764 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02762f
C2765 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.SM 0.00168f
C2766 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.15202f
C2767 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00214f
C2768 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.04036f
C2769 XA.XIR[5].XIC[5].icell.PDM Vbias 0.04261f
C2770 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02799f
C2771 XA.XIR[7].XIC[10].icell.PDM VPWR 0.00799f
C2772 XThR.Tn[0] XThR.XTB2.Y 0.00125f
C2773 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C2774 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.1106f
C2775 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02762f
C2776 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C2777 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PUM 0.00465f
C2778 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C2779 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C2780 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.15202f
C2781 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C2782 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00214f
C2783 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00214f
C2784 XA.XIR[4].XIC[3].icell.SM VPWR 0.00158f
C2785 XA.XIR[15].XIC[8].icell.PDM VPWR 0.0114f
C2786 XA.XIR[10].XIC[0].icell.Ien Iout 0.06411f
C2787 XThR.Tn[9] XA.XIR[10].XIC[0].icell.Ien 0.0037f
C2788 XA.XIR[12].XIC[4].icell.PDM Vbias 0.04261f
C2789 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C2790 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.SM 0.00168f
C2791 XA.XIR[12].XIC[11].icell.SM Vbias 0.00701f
C2792 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.15202f
C2793 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.15202f
C2794 XA.XIR[6].XIC[5].icell.PDM Iout 0.00117f
C2795 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C2796 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C2797 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C2798 XA.XIR[11].XIC[10].icell.PDM Vbias 0.04261f
C2799 XThC.Tn[3] XThR.Tn[6] 0.28739f
C2800 XA.XIR[5].XIC[12].icell.PDM Iout 0.00117f
C2801 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02762f
C2802 XA.XIR[14].XIC[2].icell.PDM Iout 0.00117f
C2803 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C2804 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00584f
C2805 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.15202f
C2806 XA.XIR[9].XIC[6].icell.PDM VPWR 0.00799f
C2807 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00584f
C2808 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00584f
C2809 a_8963_9569# VPWR 0.0033f
C2810 XA.XIR[8].XIC[0].icell.SM Vbias 0.00675f
C2811 XThR.XTB7.A XThR.Tn[7] 0.00182f
C2812 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.SM 0.00168f
C2813 XA.XIR[13].XIC[6].icell.PDM Iout 0.00117f
C2814 XThR.XTB7.A a_n997_2891# 0.00342f
C2815 XA.XIR[13].XIC[13].icell.Ien VPWR 0.1903f
C2816 XA.XIR[14].XIC[11].icell.PDM Vbias 0.04261f
C2817 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C2818 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02762f
C2819 XA.XIR[3].XIC[2].icell.SM Vbias 0.00701f
C2820 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.SM 0.0039f
C2821 XThC.Tn[5] XThR.Tn[11] 0.28739f
C2822 XA.XIR[12].XIC[12].icell.PDM VPWR 0.00799f
C2823 XA.XIR[6].XIC[7].icell.Ien Vbias 0.21098f
C2824 XA.XIR[9].XIC[6].icell.SM VPWR 0.00158f
C2825 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C2826 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C2827 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.03579f
C2828 XA.XIR[15].XIC[8].icell.SM Vbias 0.00701f
C2829 XThC.Tn[3] Vbias 2.45762f
C2830 XA.XIR[9].XIC[2].icell.SM Iout 0.00388f
C2831 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00214f
C2832 XA.XIR[5].XIC[10].icell.PUM Vbias 0.0031f
C2833 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00214f
C2834 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.SM 0.00168f
C2835 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PDM 0.00587f
C2836 XA.XIR[15].XIC[13].icell.PDM VPWR 0.0114f
C2837 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.03425f
C2838 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04031f
C2839 XA.XIR[3].XIC[0].icell.PDM Vbias 0.04207f
C2840 XA.XIR[8].XIC[2].icell.PDM Vbias 0.04261f
C2841 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00584f
C2842 XThR.Tn[11] XA.XIR[12].XIC[1].icell.Ien 0.00338f
C2843 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00214f
C2844 XA.XIR[4].XIC[11].icell.SM Vbias 0.00701f
C2845 XA.XIR[3].XIC[9].icell.Ien VPWR 0.1903f
C2846 XA.XIR[12].XIC[14].icell.PUM Vbias 0.0031f
C2847 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.SM 0.0039f
C2848 XA.XIR[1].XIC[11].icell.PDM VPWR 0.00799f
C2849 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.03433f
C2850 XA.XIR[6].XIC[14].icell.PUM VPWR 0.00937f
C2851 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PUM 0.00465f
C2852 XThC.XTB5.Y XThC.Tn[6] 0.00352f
C2853 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00584f
C2854 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14] 0.00341f
C2855 XA.XIR[3].XIC[5].icell.Ien Iout 0.06417f
C2856 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.0353f
C2857 XA.XIR[2].XIC[6].icell.PDM Vbias 0.04261f
C2858 XA.XIR[13].XIC[3].icell.Ien Vbias 0.21098f
C2859 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[5].icell.Ien 0.00214f
C2860 XThC.Tn[9] XThR.Tn[13] 0.28739f
C2861 XA.XIR[8].XIC[5].icell.SM Vbias 0.00701f
C2862 XA.XIR[4].XIC[11].icell.PDM VPWR 0.00799f
C2863 XA.XIR[2].XIC[2].icell.Ien VPWR 0.1903f
C2864 XA.XIR[7].XIC[2].icell.SM VPWR 0.00158f
C2865 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C2866 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C2867 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04031f
C2868 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02762f
C2869 XA.XIR[12].XIC[5].icell.PUM Vbias 0.0031f
C2870 XA.XIR[5].XIC[11].icell.SM Iout 0.00388f
C2871 XA.XIR[13].XIC[14].icell.SM VPWR 0.00207f
C2872 XA.XIR[1].XIC[4].icell.Ien VPWR 0.1903f
C2873 XA.XIR[14].XIC[8].icell.PUM VPWR 0.00937f
C2874 XA.XIR[11].XIC[6].icell.Ien Vbias 0.21098f
C2875 XThC.Tn[12] Iout 0.84307f
C2876 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.03425f
C2877 XThC.Tn[12] XThR.Tn[9] 0.28739f
C2878 XA.XIR[4].XIC[14].icell.Ien Iout 0.06417f
C2879 XA.XIR[3].XIC[7].icell.PDM Iout 0.00117f
C2880 XA.XIR[9].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2881 XA.XIR[8].XIC[9].icell.PDM Iout 0.00117f
C2882 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.SM 0.0039f
C2883 XA.XIR[13].XIC[10].icell.PUM VPWR 0.00937f
C2884 XThC.Tn[8] XThR.Tn[8] 0.28739f
C2885 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04031f
C2886 XA.XIR[9].XIC[14].icell.SM Vbias 0.00701f
C2887 XA.XIR[8].XIC[12].icell.Ien VPWR 0.1903f
C2888 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00584f
C2889 XA.XIR[10].XIC[8].icell.Ien Vbias 0.21098f
C2890 XThR.Tn[6] XA.XIR[7].XIC[10].icell.SM 0.00121f
C2891 XA.XIR[2].XIC[13].icell.PDM Iout 0.00117f
C2892 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04031f
C2893 XA.XIR[8].XIC[8].icell.Ien Iout 0.06417f
C2894 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PUM 0.00465f
C2895 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.03425f
C2896 XA.XIR[0].XIC[7].icell.SM Vbias 0.00716f
C2897 XThR.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.00338f
C2898 XA.XIR[12].XIC[6].icell.SM Iout 0.00388f
C2899 XThR.Tn[0] XA.XIR[0].XIC[10].icell.PDM 0.00341f
C2900 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C2901 XThC.XTBN.Y XThC.Tn[6] 0.61358f
C2902 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C2903 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00214f
C2904 XThR.XTB7.B a_n997_3979# 0.01152f
C2905 XThC.Tn[3] XThR.Tn[4] 0.28739f
C2906 XA.XIR[10].XIC_15.icell.PDM Iout 0.00133f
C2907 XThR.Tn[1] XA.XIR[1].XIC[8].icell.PDM 0.00341f
C2908 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PDM 0.00172f
C2909 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C2910 XA.XIR[12].XIC[9].icell.SM Vbias 0.00701f
C2911 XThR.XTBN.Y XA.XIR[8].XIC_dummy_left.icell.Ien 0.00243f
C2912 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04031f
C2913 XA.XIR[2].XIC[10].icell.Ien Vbias 0.21098f
C2914 XA.XIR[7].XIC[10].icell.SM Vbias 0.00701f
C2915 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18971f
C2916 XThC.XTB7.Y a_5949_9615# 0.00153f
C2917 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C2918 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C2919 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5] 0.00341f
C2920 XThC.Tn[7] XThR.Tn[10] 0.28739f
C2921 XA.XIR[1].XIC[12].icell.Ien Vbias 0.21104f
C2922 XA.XIR[0].XIC[10].icell.Ien Iout 0.06389f
C2923 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.15202f
C2924 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Ien 0.00584f
C2925 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.15202f
C2926 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C2927 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.SM 0.0039f
C2928 XThR.Tn[2] XA.XIR[2].XIC[5].icell.PDM 0.00341f
C2929 XA.XIR[13].XIC[11].icell.Ien VPWR 0.1903f
C2930 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.SM 0.0039f
C2931 XThR.Tn[13] XA.XIR[14].XIC[5].icell.Ien 0.00338f
C2932 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04031f
C2933 a_7651_9569# XThC.Tn[8] 0.1927f
C2934 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PUM 0.00465f
C2935 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02762f
C2936 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.15202f
C2937 XThC.XTB5.A XThC.XTB7.Y 0.00179f
C2938 XA.XIR[15].XIC[0].icell.SM VPWR 0.00158f
C2939 XA.XIR[5].XIC[2].icell.PUM VPWR 0.00937f
C2940 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6] 0.00341f
C2941 XA.XIR[7].XIC[13].icell.Ien Iout 0.06417f
C2942 XThR.Tn[0] XA.XIR[1].XIC[8].icell.Ien 0.00338f
C2943 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C2944 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.SM 0.00168f
C2945 XA.XIR[11].XIC[1].icell.PDM VPWR 0.00799f
C2946 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00214f
C2947 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C2948 XA.XIR[11].XIC[0].icell.SM Vbias 0.00675f
C2949 XA.XIR[7].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2950 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.03425f
C2951 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02762f
C2952 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Iout 0.00347f
C2953 XA.XIR[12].XIC[12].icell.PUM Vbias 0.0031f
C2954 XThR.Tn[7] XA.XIR[8].XIC[14].icell.Ien 0.00338f
C2955 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PUM 0.00465f
C2956 XA.XIR[10].XIC[5].icell.PDM VPWR 0.00799f
C2957 XThR.Tn[13] a_n997_1803# 0.0021f
C2958 XA.XIR[7].XIC[6].icell.PDM Vbias 0.04261f
C2959 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C2960 XA.XIR[13].XIC[0].icell.Ien Iout 0.06411f
C2961 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.03425f
C2962 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02771f
C2963 XThR.Tn[5] XA.XIR[6].XIC[10].icell.Ien 0.00338f
C2964 XA.XIR[15].XIC[4].icell.PDM Vbias 0.04261f
C2965 XA.XIR[4].XIC[3].icell.PUM Vbias 0.0031f
C2966 XA.XIR[6].XIC[13].icell.PDM Vbias 0.04261f
C2967 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.SM 0.00168f
C2968 XThR.XTB7.B XThR.Tn[7] 0.07415f
C2969 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.03425f
C2970 XA.XIR[6].XIC[4].icell.Ien VPWR 0.1903f
C2971 XThR.XTB7.B a_n997_2891# 0.0168f
C2972 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02762f
C2973 XA.XIR[14].XIC[10].icell.PDM Vbias 0.04261f
C2974 XA.XIR[15].XIC[5].icell.SM VPWR 0.00158f
C2975 XA.XIR[15].XIC[13].icell.SM Vbias 0.00701f
C2976 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.03425f
C2977 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00256f
C2978 XA.XIR[12].XIC[11].icell.PDM VPWR 0.00799f
C2979 XA.XIR[5].XIC[7].icell.PUM VPWR 0.00937f
C2980 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.SM 0.0039f
C2981 XThC.XTB7.B a_8963_9569# 0.02071f
C2982 XThC.Tn[12] XA.XIR[0].XIC[11].icell.PDM 0.00106f
C2983 XA.XIR[15].XIC[1].icell.SM Iout 0.00388f
C2984 XA.XIR[9].XIC[2].icell.PDM Vbias 0.04261f
C2985 XA.XIR[7].XIC[13].icell.PDM Iout 0.00117f
C2986 XA.XIR[4].XIC[8].icell.SM VPWR 0.00158f
C2987 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00584f
C2988 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C2989 XThC.Tn[5] XThR.Tn[14] 0.28739f
C2990 XA.XIR[15].XIC[12].icell.PDM VPWR 0.0114f
C2991 XThC.XTB6.A XThC.XTB7.A 0.44014f
C2992 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.15202f
C2993 XA.XIR[4].XIC[4].icell.SM Iout 0.00388f
C2994 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C2995 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00214f
C2996 XA.XIR[9].XIC[6].icell.PUM Vbias 0.0031f
C2997 XA.XIR[12].XIC[13].icell.Ien Vbias 0.21098f
C2998 XThR.XTB6.A data[4] 0.48493f
C2999 XA.XIR[8].XIC[2].icell.SM VPWR 0.00158f
C3000 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C3001 XThR.Tn[13] XA.XIR[14].XIC[0].icell.Ien 0.0037f
C3002 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00584f
C3003 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C3004 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.03425f
C3005 XA.XIR[0].XIC[13].icell.PDM VPWR 0.00774f
C3006 XThC.XTB2.Y XThC.Tn[1] 0.17879f
C3007 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C3008 XA.XIR[11].XIC[3].icell.Ien VPWR 0.1903f
C3009 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C3010 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.SM 0.0039f
C3011 XA.XIR[9].XIC[9].icell.PDM Iout 0.00117f
C3012 XA.XIR[3].XIC[7].icell.SM Vbias 0.00701f
C3013 XThC.XTB5.Y data[3] 0.00931f
C3014 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.SM 0.00168f
C3015 XA.XIR[1].XIC[7].icell.PDM Vbias 0.04261f
C3016 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9] 0.00341f
C3017 XA.XIR[9].XIC[11].icell.SM VPWR 0.00158f
C3018 XA.XIR[6].XIC[12].icell.Ien Vbias 0.21098f
C3019 XA.XIR[10].XIC[5].icell.Ien VPWR 0.1903f
C3020 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00214f
C3021 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11] 0.00341f
C3022 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C3023 XA.XIR[5].XIC_15.icell.PUM Vbias 0.0031f
C3024 XA.XIR[9].XIC[7].icell.SM Iout 0.00388f
C3025 XA.XIR[4].XIC[7].icell.PDM Vbias 0.04261f
C3026 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.03425f
C3027 XA.XIR[0].XIC[4].icell.SM VPWR 0.00158f
C3028 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.SM 0.0039f
C3029 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04031f
C3030 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C3031 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04031f
C3032 XA.XIR[1].XIC[2].icell.SM Vbias 0.00704f
C3033 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00214f
C3034 XA.XIR[3].XIC_15.icell.PDM Vbias 0.04401f
C3035 XA.XIR[14].XIC[6].icell.Ien Vbias 0.21098f
C3036 XA.XIR[3].XIC[14].icell.Ien VPWR 0.19036f
C3037 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02762f
C3038 XA.XIR[3].XIC[10].icell.Ien Iout 0.06417f
C3039 XThR.XTB2.Y a_n1049_5317# 0.00844f
C3040 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.SM 0.00168f
C3041 XThR.XTBN.Y a_n997_3979# 0.23021f
C3042 XA.XIR[12].XIC[14].icell.SM Vbias 0.00701f
C3043 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C3044 XA.XIR[13].XIC[8].icell.Ien Vbias 0.21098f
C3045 XA.XIR[1].XIC[14].icell.PDM Iout 0.00117f
C3046 XA.XIR[8].XIC[10].icell.SM Vbias 0.00701f
C3047 XA.XIR[7].XIC[7].icell.SM VPWR 0.00158f
C3048 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.SM 0.0039f
C3049 XA.XIR[10].XIC_15.icell.SM VPWR 0.00275f
C3050 XA.XIR[2].XIC[7].icell.Ien VPWR 0.1903f
C3051 XA.XIR[10].XIC[14].icell.PDM Iout 0.00117f
C3052 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04052f
C3053 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00214f
C3054 XA.XIR[12].XIC[10].icell.PUM Vbias 0.0031f
C3055 XA.XIR[7].XIC[3].icell.SM Iout 0.00388f
C3056 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02762f
C3057 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.SM 0.0039f
C3058 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C3059 XA.XIR[1].XIC[9].icell.Ien VPWR 0.1903f
C3060 XA.XIR[4].XIC[14].icell.PDM Iout 0.00117f
C3061 XA.XIR[2].XIC[3].icell.Ien Iout 0.06417f
C3062 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.15202f
C3063 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.SM 0.00168f
C3064 XThR.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.00338f
C3065 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C3066 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02762f
C3067 XA.XIR[13].XIC_15.icell.PDM Iout 0.00133f
C3068 XA.XIR[1].XIC[5].icell.Ien Iout 0.06417f
C3069 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.SM 0.00168f
C3070 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C3071 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C3072 XA.XIR[9].XIC[1].icell.PUM Vbias 0.0031f
C3073 XThR.Tn[7] XA.XIR[8].XIC[4].icell.SM 0.00121f
C3074 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PUM 0.00465f
C3075 XThC.XTB3.Y a_4067_9615# 0.23056f
C3076 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.03425f
C3077 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C3078 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.SM 0.0039f
C3079 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PUM 0.00429f
C3080 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C3081 XA.XIR[8].XIC[13].icell.Ien Iout 0.06417f
C3082 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PUM 0.00465f
C3083 XThR.Tn[11] XA.XIR[12].XIC[2].icell.Ien 0.00338f
C3084 XThR.Tn[8] XA.XIR[9].XIC[13].icell.Ien 0.00338f
C3085 XA.XIR[15].XIC[11].icell.SM Vbias 0.00701f
C3086 a_4067_9615# XThC.Tn[2] 0.27699f
C3087 XA.XIR[0].XIC[12].icell.SM Vbias 0.00716f
C3088 XThC.Tn[7] XThR.Tn[13] 0.28739f
C3089 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.SM 0.00168f
C3090 XThR.XTB4.Y a_n997_3979# 0.00497f
C3091 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.SM 0.0039f
C3092 XA.XIR[8].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3093 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.15202f
C3094 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02762f
C3095 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.04036f
C3096 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PUM 0.00186f
C3097 XThC.Tn[1] Iout 0.84229f
C3098 XThR.Tn[4] XA.XIR[4].XIC[7].icell.PDM 0.00341f
C3099 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PUM 0.00465f
C3100 XThC.Tn[1] XThR.Tn[9] 0.28739f
C3101 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.03425f
C3102 XThC.XTB5.A XThC.XTB6.A 1.80461f
C3103 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PUM 0.00186f
C3104 XThR.Tn[10] XA.XIR[11].XIC[5].icell.SM 0.00121f
C3105 XThR.Tn[3] XA.XIR[3].XIC[8].icell.PDM 0.00341f
C3106 XA.XIR[2].XIC_15.icell.Ien Vbias 0.21234f
C3107 XThR.Tn[1] XA.XIR[2].XIC[6].icell.Ien 0.00338f
C3108 XA.XIR[12].XIC[11].icell.Ien Vbias 0.21098f
C3109 XThC.Tn[6] XThR.Tn[8] 0.28739f
C3110 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C3111 XA.XIR[6].XIC[4].icell.PDM VPWR 0.00799f
C3112 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.SM 0.0039f
C3113 XThR.XTB7.A a_n1049_6699# 0.02294f
C3114 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04052f
C3115 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00214f
C3116 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.15202f
C3117 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.15202f
C3118 XA.XIR[0].XIC_15.icell.Ien Iout 0.06388f
C3119 XA.XIR[14].XIC[0].icell.SM Vbias 0.00675f
C3120 XThR.XTB5.Y VPWR 1.0269f
C3121 XA.XIR[14].XIC[1].icell.PDM VPWR 0.00799f
C3122 XA.XIR[5].XIC[11].icell.PDM VPWR 0.00799f
C3123 XThR.XTBN.Y XThR.Tn[7] 0.8998f
C3124 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PUM 0.00465f
C3125 XThR.XTBN.Y a_n997_2891# 0.22804f
C3126 XA.XIR[13].XIC[5].icell.PDM VPWR 0.00799f
C3127 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02762f
C3128 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C3129 XA.XIR[10].XIC[1].icell.PDM Vbias 0.04261f
C3130 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00584f
C3131 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.SM 0.0039f
C3132 XA.XIR[15].XIC[14].icell.PUM Vbias 0.0031f
C3133 XThC.XTB7.Y a_8739_9569# 0.00474f
C3134 XA.XIR[6].XIC[0].icell.Ien Iout 0.06411f
C3135 XA.XIR[12].XIC[10].icell.PDM VPWR 0.00799f
C3136 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00584f
C3137 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.SM 0.00168f
C3138 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02762f
C3139 XThR.Tn[0] XA.XIR[1].XIC[13].icell.Ien 0.00338f
C3140 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.SM 0.00168f
C3141 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.SM 0.00168f
C3142 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.0353f
C3143 XThR.XTB2.Y a_n1049_6405# 0.00847f
C3144 XThR.XTB7.B a_n997_1579# 0.00209f
C3145 XA.XIR[6].XIC[2].icell.SM Vbias 0.00701f
C3146 XA.XIR[9].XIC[3].icell.PUM VPWR 0.00937f
C3147 XThC.XTB3.Y XThC.Tn[3] 0.01287f
C3148 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00584f
C3149 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.SM 0.00168f
C3150 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PUM 0.00465f
C3151 XA.XIR[15].XIC[11].icell.PDM VPWR 0.0114f
C3152 XA.XIR[15].XIC[5].icell.PUM Vbias 0.0031f
C3153 XA.XIR[11].XIC[4].icell.PDM Iout 0.00117f
C3154 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.SM 0.0039f
C3155 XA.XIR[5].XIC[5].icell.Ien Vbias 0.21098f
C3156 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00584f
C3157 XThR.Tn[5] XThR.Tn[6] 0.06649f
C3158 XThC.Tn[2] XThC.Tn[3] 0.33669f
C3159 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00214f
C3160 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.SM 0.00168f
C3161 XThR.Tn[5] XA.XIR[6].XIC_15.icell.Ien 0.00117f
C3162 XA.XIR[4].XIC[8].icell.PUM Vbias 0.0031f
C3163 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C3164 XA.XIR[10].XIC[8].icell.PDM Iout 0.00117f
C3165 XThR.XTB4.Y a_n997_2891# 0.00813f
C3166 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04031f
C3167 XA.XIR[3].XIC[4].icell.SM VPWR 0.00158f
C3168 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02762f
C3169 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C3170 XA.XIR[6].XIC[9].icell.Ien VPWR 0.1903f
C3171 XThC.Tn[0] XA.XIR[3].XIC_dummy_left.icell.Iout 0.00109f
C3172 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.SM 0.0039f
C3173 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.SM 0.00168f
C3174 XA.XIR[6].XIC[5].icell.Ien Iout 0.06417f
C3175 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[2].icell.SM 0.0039f
C3176 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7] 0.00341f
C3177 XA.XIR[5].XIC[12].icell.PUM VPWR 0.00937f
C3178 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00584f
C3179 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.03425f
C3180 XThR.Tn[10] a_n997_2891# 0.1927f
C3181 XThR.Tn[5] Vbias 3.74761f
C3182 XA.XIR[15].XIC[6].icell.SM Iout 0.00388f
C3183 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00214f
C3184 XThR.Tn[3] XA.XIR[4].XIC[0].icell.Ien 0.00338f
C3185 XA.XIR[3].XIC[6].icell.PDM VPWR 0.00799f
C3186 XA.XIR[4].XIC[13].icell.SM VPWR 0.00158f
C3187 XA.XIR[8].XIC[8].icell.PDM VPWR 0.00799f
C3188 XA.XIR[2].XIC[0].icell.SM Vbias 0.00675f
C3189 XA.XIR[7].XIC[2].icell.PUM Vbias 0.0031f
C3190 XA.XIR[14].XIC[3].icell.Ien VPWR 0.19084f
C3191 XA.XIR[0].XIC[9].icell.PDM Vbias 0.04282f
C3192 XThC.Tn[9] XThR.Tn[7] 0.28739f
C3193 XA.XIR[11].XIC[1].icell.SM Vbias 0.00701f
C3194 XA.XIR[2].XIC[12].icell.PDM VPWR 0.00799f
C3195 XA.XIR[4].XIC[9].icell.SM Iout 0.00388f
C3196 XA.XIR[15].XIC[9].icell.SM Vbias 0.00701f
C3197 XA.XIR[13].XIC[5].icell.Ien VPWR 0.1903f
C3198 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C3199 XA.XIR[9].XIC[11].icell.PUM Vbias 0.0031f
C3200 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04031f
C3201 XA.XIR[8].XIC[7].icell.SM VPWR 0.00158f
C3202 XA.XIR[10].XIC[3].icell.SM Vbias 0.00701f
C3203 XThR.XTB1.Y VPWR 1.12978f
C3204 XA.XIR[0].XIC[0].icell.SM Iout 0.00367f
C3205 XThC.XTB2.Y a_3523_10575# 0.01006f
C3206 XA.XIR[2].XIC[0].icell.PDM Iout 0.00117f
C3207 XThC.XTB7.Y XThC.Tn[11] 0.07471f
C3208 XA.XIR[12].XIC[7].icell.PUM VPWR 0.00937f
C3209 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00584f
C3210 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00584f
C3211 XThR.XTB6.Y a_n1319_5611# 0.01283f
C3212 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12] 0.00341f
C3213 XA.XIR[8].XIC[3].icell.SM Iout 0.00388f
C3214 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C3215 XThR.Tn[8] XA.XIR[9].XIC[3].icell.SM 0.00121f
C3216 XA.XIR[0].XIC[4].icell.PUM Vbias 0.0031f
C3217 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C3218 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3219 XA.XIR[10].XIC[13].icell.PDM Iout 0.00117f
C3220 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.04036f
C3221 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02762f
C3222 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PUM 0.00465f
C3223 XA.XIR[11].XIC[8].icell.Ien VPWR 0.1903f
C3224 XA.XIR[3].XIC[12].icell.SM Vbias 0.00701f
C3225 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.SM 0.0039f
C3226 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02762f
C3227 XThR.Tn[4] XA.XIR[5].XIC[5].icell.Ien 0.00338f
C3228 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C3229 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.03425f
C3230 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PUM 0.00465f
C3231 XA.XIR[11].XIC[4].icell.Ien Iout 0.06417f
C3232 XThR.Tn[3] XA.XIR[4].XIC[5].icell.Ien 0.00338f
C3233 XA.XIR[13].XIC[14].icell.PDM Iout 0.00117f
C3234 XA.XIR[13].XIC_15.icell.SM VPWR 0.00275f
C3235 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02803f
C3236 XA.XIR[7].XIC[7].icell.PUM Vbias 0.0031f
C3237 XA.XIR[9].XIC[12].icell.SM Iout 0.00388f
C3238 XA.XIR[2].XIC[5].icell.SM Vbias 0.00701f
C3239 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C3240 XA.XIR[10].XIC[6].icell.Ien Iout 0.06417f
C3241 XA.XIR[0].XIC[9].icell.SM VPWR 0.00158f
C3242 XThR.Tn[9] XA.XIR[10].XIC[6].icell.Ien 0.00338f
C3243 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02762f
C3244 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5] 0.00341f
C3245 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02762f
C3246 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00584f
C3247 XA.XIR[1].XIC[7].icell.SM Vbias 0.00704f
C3248 XA.XIR[9].XIC_15.icell.SM Vbias 0.00701f
C3249 XA.XIR[0].XIC[5].icell.SM Iout 0.00367f
C3250 XA.XIR[15].XIC[12].icell.PUM Vbias 0.0031f
C3251 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04031f
C3252 XThR.Tn[5] XA.XIR[6].XIC[0].icell.SM 0.00121f
C3253 XA.XIR[3].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3254 XThR.Tn[4] XThR.Tn[5] 0.07388f
C3255 XA.XIR[3].XIC_15.icell.Ien Iout 0.0642f
C3256 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00584f
C3257 XThC.XTB5.A XThC.Tn[8] 0.00205f
C3258 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04031f
C3259 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8] 0.00341f
C3260 XThC.Tn[8] XThR.Tn[3] 0.28739f
C3261 XA.XIR[2].XIC[12].icell.Ien VPWR 0.1903f
C3262 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.PDM 0.00591f
C3263 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[10].icell.Ien 0.00214f
C3264 XA.XIR[7].XIC[12].icell.SM VPWR 0.00158f
C3265 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Ien 0.00584f
C3266 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PUM 0.00465f
C3267 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6] 0.00341f
C3268 XA.XIR[10].XIC[0].icell.PUM VPWR 0.00937f
C3269 XA.XIR[1].XIC[14].icell.Ien VPWR 0.19036f
C3270 XA.XIR[7].XIC[8].icell.SM Iout 0.00388f
C3271 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.03023f
C3272 XA.XIR[2].XIC[8].icell.Ien Iout 0.06417f
C3273 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04052f
C3274 XThC.Tn[5] VPWR 5.90052f
C3275 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.15202f
C3276 XThR.Tn[0] XA.XIR[1].XIC[3].icell.SM 0.00121f
C3277 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.SM 0.00168f
C3278 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.SM 0.00168f
C3279 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00214f
C3280 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.SM 0.0039f
C3281 XThR.Tn[12] XA.XIR[13].XIC[4].icell.Ien 0.00338f
C3282 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02762f
C3283 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PUM 0.00465f
C3284 XA.XIR[1].XIC[10].icell.Ien Iout 0.06417f
C3285 XThR.XTB7.B a_n1049_6699# 0.0036f
C3286 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00584f
C3287 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.SM 0.00168f
C3288 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C3289 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11336f
C3290 XThR.Tn[7] XA.XIR[8].XIC[9].icell.SM 0.00121f
C3291 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C3292 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.03425f
C3293 XThC.Tn[11] XThR.Tn[0] 0.28749f
C3294 XThC.Tn[13] XThR.Tn[5] 0.2874f
C3295 a_5155_9615# Vbias 0.00695f
C3296 XA.XIR[12].XIC[1].icell.Ien VPWR 0.1903f
C3297 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.03425f
C3298 XThR.Tn[5] XA.XIR[6].XIC[5].icell.SM 0.00121f
C3299 XThR.Tn[11] XA.XIR[12].XIC[7].icell.Ien 0.00338f
C3300 XA.XIR[6].XIC[0].icell.PDM Vbias 0.04207f
C3301 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.03425f
C3302 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00584f
C3303 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C3304 XA.XIR[15].XIC[13].icell.Ien Vbias 0.17899f
C3305 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PDM 0.00172f
C3306 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00214f
C3307 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.15202f
C3308 XA.XIR[5].XIC[7].icell.PDM Vbias 0.04261f
C3309 XThR.XTBN.Y a_n997_1579# 0.23006f
C3310 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C3311 XA.XIR[5].XIC[2].icell.Ien VPWR 0.1903f
C3312 XA.XIR[7].XIC[12].icell.PDM VPWR 0.00799f
C3313 XThR.XTB7.Y a_n1049_5317# 0.27822f
C3314 XA.XIR[13].XIC[1].icell.PDM Vbias 0.04261f
C3315 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C3316 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.03425f
C3317 XA.XIR[7].XIC[0].icell.PDM Iout 0.00117f
C3318 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PUM 0.00465f
C3319 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C3320 XThR.Tn[1] XA.XIR[2].XIC[11].icell.Ien 0.00338f
C3321 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.SM 0.00168f
C3322 XA.XIR[4].XIC[5].icell.PUM VPWR 0.00937f
C3323 XA.XIR[10].XIC[0].icell.SM Iout 0.00388f
C3324 XA.XIR[15].XIC[10].icell.PDM VPWR 0.0114f
C3325 XThR.Tn[9] XA.XIR[10].XIC[0].icell.SM 0.00127f
C3326 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02762f
C3327 XA.XIR[12].XIC[6].icell.PDM Vbias 0.04261f
C3328 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02762f
C3329 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C3330 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.15202f
C3331 XA.XIR[6].XIC[7].icell.PDM Iout 0.00117f
C3332 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.SM 0.0039f
C3333 XA.XIR[14].XIC[4].icell.PDM Iout 0.00117f
C3334 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PUM 0.00465f
C3335 XA.XIR[5].XIC[14].icell.PDM Iout 0.00117f
C3336 a_10051_9569# VPWR 0.00319f
C3337 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00584f
C3338 XA.XIR[9].XIC[8].icell.PDM VPWR 0.00799f
C3339 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PUM 0.00465f
C3340 XA.XIR[8].XIC[2].icell.PUM Vbias 0.0031f
C3341 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C3342 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.SM 0.00168f
C3343 XA.XIR[0].XIC[0].icell.PDM VPWR 0.00774f
C3344 XA.XIR[13].XIC[8].icell.PDM Iout 0.00117f
C3345 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Iout 0.00347f
C3346 XA.XIR[3].XIC[4].icell.PUM Vbias 0.0031f
C3347 XA.XIR[15].XIC[14].icell.SM Vbias 0.00701f
C3348 XA.XIR[9].XIC[8].icell.PUM VPWR 0.00937f
C3349 XA.XIR[6].XIC[7].icell.SM Vbias 0.00701f
C3350 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.SM 0.00168f
C3351 XThC.Tn[10] XThR.Tn[2] 0.28739f
C3352 XThC.XTB6.Y Vbias 0.01503f
C3353 XA.XIR[15].XIC[10].icell.PUM Vbias 0.0031f
C3354 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.15202f
C3355 XA.XIR[5].XIC[10].icell.Ien Vbias 0.21098f
C3356 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C3357 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04031f
C3358 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.SM 0.0039f
C3359 XThR.Tn[11] XThR.Tn[12] 0.11452f
C3360 XA.XIR[4].XIC[13].icell.PUM Vbias 0.0031f
C3361 XA.XIR[11].XIC[12].icell.SM Iout 0.00388f
C3362 XA.XIR[3].XIC[9].icell.SM VPWR 0.00158f
C3363 XA.XIR[3].XIC[2].icell.PDM Vbias 0.04261f
C3364 XA.XIR[8].XIC[4].icell.PDM Vbias 0.04261f
C3365 XA.XIR[14].XIC[1].icell.SM Vbias 0.00701f
C3366 XA.XIR[1].XIC[13].icell.PDM VPWR 0.00799f
C3367 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10] 0.00341f
C3368 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.SM 0.00168f
C3369 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.SM 0.00168f
C3370 XA.XIR[6].XIC[14].icell.Ien VPWR 0.19036f
C3371 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.03425f
C3372 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04031f
C3373 XA.XIR[10].XIC[12].icell.PDM Iout 0.00117f
C3374 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14] 0.00341f
C3375 XA.XIR[3].XIC[5].icell.SM Iout 0.00388f
C3376 XThR.Tn[3] a_n1049_6405# 0.00542f
C3377 XA.XIR[2].XIC[8].icell.PDM Vbias 0.04261f
C3378 XA.XIR[1].XIC[1].icell.PDM Iout 0.00117f
C3379 XA.XIR[13].XIC[3].icell.SM Vbias 0.00701f
C3380 XA.XIR[8].XIC[7].icell.PUM Vbias 0.0031f
C3381 XA.XIR[2].XIC[2].icell.SM VPWR 0.00158f
C3382 XA.XIR[6].XIC[10].icell.Ien Iout 0.06417f
C3383 XA.XIR[7].XIC[4].icell.PUM VPWR 0.00937f
C3384 XThC.XTB7.A XThC.Tn[6] 0.10589f
C3385 XA.XIR[4].XIC[13].icell.PDM VPWR 0.00799f
C3386 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.SM 0.0039f
C3387 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04031f
C3388 XA.XIR[12].XIC[5].icell.Ien Vbias 0.21098f
C3389 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3390 XA.XIR[4].XIC[1].icell.PDM Iout 0.00117f
C3391 XA.XIR[1].XIC[4].icell.SM VPWR 0.00158f
C3392 XA.XIR[13].XIC[13].icell.PDM Iout 0.00117f
C3393 XA.XIR[14].XIC[8].icell.Ien VPWR 0.19084f
C3394 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02762f
C3395 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00584f
C3396 XThR.XTB5.A XThR.XTBN.A 0.06303f
C3397 XA.XIR[11].XIC[6].icell.SM Vbias 0.00701f
C3398 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.03023f
C3399 XA.XIR[3].XIC[9].icell.PDM Iout 0.00117f
C3400 XA.XIR[4].XIC[14].icell.SM Iout 0.00388f
C3401 XA.XIR[8].XIC[11].icell.PDM Iout 0.00117f
C3402 XA.XIR[14].XIC[4].icell.Ien Iout 0.06417f
C3403 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04031f
C3404 XA.XIR[9].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3405 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00584f
C3406 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C3407 XA.XIR[8].XIC[12].icell.SM VPWR 0.00158f
C3408 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.SM 0.0039f
C3409 XA.XIR[10].XIC[8].icell.SM Vbias 0.00701f
C3410 XA.XIR[15].XIC[11].icell.Ien Vbias 0.17899f
C3411 XA.XIR[2].XIC_15.icell.PDM Iout 0.00133f
C3412 XA.XIR[13].XIC[6].icell.Ien Iout 0.06417f
C3413 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02762f
C3414 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00584f
C3415 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C3416 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00214f
C3417 XA.XIR[8].XIC[8].icell.SM Iout 0.00388f
C3418 XThC.XTB4.Y Vbias 0.01548f
C3419 XThR.Tn[12] XA.XIR[13].XIC[12].icell.SM 0.00121f
C3420 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.03425f
C3421 XA.XIR[0].XIC[9].icell.PUM Vbias 0.0031f
C3422 XThR.Tn[8] XA.XIR[9].XIC[8].icell.SM 0.00121f
C3423 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PUM 0.00465f
C3424 XThC.Tn[8] XThR.Tn[11] 0.28739f
C3425 XThR.Tn[2] XA.XIR[3].XIC[3].icell.Ien 0.00338f
C3426 XThR.Tn[0] XA.XIR[0].XIC[12].icell.PDM 0.00341f
C3427 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.SM 0.00168f
C3428 XA.XIR[12].XIC_15.icell.SM Vbias 0.00701f
C3429 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39003f
C3430 XThR.Tn[4] XA.XIR[5].XIC[10].icell.Ien 0.00338f
C3431 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PUM 0.00444f
C3432 XThR.Tn[1] XA.XIR[1].XIC[10].icell.PDM 0.00341f
C3433 XA.XIR[11].XIC[9].icell.Ien Iout 0.06417f
C3434 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C3435 XThR.XTBN.Y a_n1049_6699# 0.07601f
C3436 XThC.Tn[7] XThR.Tn[7] 0.28739f
C3437 XThR.Tn[3] XA.XIR[4].XIC[10].icell.Ien 0.00338f
C3438 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C3439 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04031f
C3440 XA.XIR[7].XIC[12].icell.PUM Vbias 0.0031f
C3441 XA.XIR[2].XIC[10].icell.SM Vbias 0.00701f
C3442 XA.XIR[0].XIC[14].icell.SM VPWR 0.00207f
C3443 XThR.Tn[1] XA.XIR[2].XIC[1].icell.SM 0.00121f
C3444 XA.XIR[13].XIC[0].icell.PUM VPWR 0.00937f
C3445 XThC.XTB7.B XThC.Tn[5] 0.00714f
C3446 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.SM 0.00168f
C3447 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04031f
C3448 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PUM 0.00465f
C3449 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.SM 0.0039f
C3450 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C3451 XA.XIR[1].XIC[12].icell.SM Vbias 0.00704f
C3452 XA.XIR[0].XIC[10].icell.SM Iout 0.00367f
C3453 XThC.XTB6.Y XThC.Tn[13] 0.32552f
C3454 XThR.XTBN.A data[5] 0.0148f
C3455 XThR.Tn[2] XA.XIR[2].XIC[7].icell.PDM 0.00341f
C3456 XThC.XTB6.A data[0] 0.48493f
C3457 XThR.Tn[13] XA.XIR[14].XIC[5].icell.SM 0.00121f
C3458 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04031f
C3459 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.SM 0.00168f
C3460 XA.XIR[3].XIC[1].icell.PUM Vbias 0.0031f
C3461 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PUM 0.00186f
C3462 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.03425f
C3463 XThC.Tn[11] XThR.Tn[1] 0.28739f
C3464 XA.XIR[15].XIC[2].icell.PUM VPWR 0.00937f
C3465 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.SM 0.00168f
C3466 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6] 0.00341f
C3467 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C3468 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PUM 0.00465f
C3469 a_5949_9615# XThC.Tn[6] 0.0018f
C3470 XA.XIR[2].XIC[13].icell.Ien Iout 0.06417f
C3471 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.SM 0.0039f
C3472 XA.XIR[7].XIC[13].icell.SM Iout 0.00388f
C3473 XThR.Tn[0] XA.XIR[1].XIC[8].icell.SM 0.00121f
C3474 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.15202f
C3475 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C3476 XThR.XTB4.Y a_n1049_6699# 0.23756f
C3477 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C3478 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C3479 XThR.Tn[12] XA.XIR[13].XIC[9].icell.Ien 0.00338f
C3480 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C3481 XA.XIR[11].XIC[2].icell.PUM Vbias 0.0031f
C3482 XA.XIR[11].XIC[3].icell.PDM VPWR 0.00799f
C3483 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.SM 0.00168f
C3484 XA.XIR[1].XIC_15.icell.Ien Iout 0.0642f
C3485 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Ien 0.00232f
C3486 XThC.Tn[11] XThR.Tn[12] 0.28739f
C3487 XA.XIR[2].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3488 XA.XIR[11].XIC[10].icell.SM Iout 0.00388f
C3489 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.03425f
C3490 XThR.Tn[7] XA.XIR[8].XIC[14].icell.SM 0.00121f
C3491 XThR.XTB7.B XThR.Tn[8] 0.05091f
C3492 XA.XIR[10].XIC[7].icell.PDM VPWR 0.00799f
C3493 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C3494 XA.XIR[7].XIC[8].icell.PDM Vbias 0.04261f
C3495 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C3496 XA.XIR[9].XIC[1].icell.Ien Vbias 0.21098f
C3497 XThR.XTB1.Y a_n1335_8331# 0.0097f
C3498 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PUM 0.00465f
C3499 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.SM 0.0039f
C3500 XA.XIR[13].XIC[0].icell.SM Iout 0.00388f
C3501 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PUM 0.00465f
C3502 XThR.Tn[5] XA.XIR[6].XIC[10].icell.SM 0.00121f
C3503 XThC.XTBN.Y XThC.Tn[9] 0.49745f
C3504 XA.XIR[6].XIC_15.icell.PDM Vbias 0.04401f
C3505 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02762f
C3506 XThC.Tn[6] XThR.Tn[3] 0.28739f
C3507 XA.XIR[15].XIC[6].icell.PDM Vbias 0.04261f
C3508 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00584f
C3509 XA.XIR[4].XIC[3].icell.Ien Vbias 0.21098f
C3510 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C3511 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.SM 0.0039f
C3512 XA.XIR[6].XIC[4].icell.SM VPWR 0.00158f
C3513 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.15202f
C3514 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08441f
C3515 XA.XIR[15].XIC[7].icell.PUM VPWR 0.00937f
C3516 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PUM 0.00465f
C3517 XA.XIR[5].XIC[7].icell.Ien VPWR 0.1903f
C3518 XThR.XTB7.A a_n1049_5611# 0.01824f
C3519 XThC.XTB7.B a_10051_9569# 0.00209f
C3520 XThC.Tn[10] XThR.Tn[10] 0.28739f
C3521 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.SM 0.00168f
C3522 XThC.Tn[0] XThR.Tn[0] 0.28807f
C3523 XA.XIR[5].XIC[3].icell.Ien Iout 0.06417f
C3524 XA.XIR[7].XIC_15.icell.PDM Iout 0.00133f
C3525 XA.XIR[9].XIC[4].icell.PDM Vbias 0.04261f
C3526 a_7875_9569# Vbias 0.00315f
C3527 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.SM 0.0039f
C3528 XA.XIR[4].XIC[10].icell.PUM VPWR 0.00937f
C3529 XThC.Tn[2] XThR.Tn[5] 0.28739f
C3530 XA.XIR[0].XIC[1].icell.PUM VPWR 0.00877f
C3531 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00214f
C3532 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02762f
C3533 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PUM 0.00465f
C3534 XThR.Tn[12] XA.XIR[13].XIC[10].icell.SM 0.00121f
C3535 XThC.XTB2.Y Vbias 0.0123f
C3536 XThC.Tn[9] XThC.Tn[10] 0.07959f
C3537 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C3538 XA.XIR[9].XIC[6].icell.Ien Vbias 0.21098f
C3539 XA.XIR[8].XIC[4].icell.PUM VPWR 0.00937f
C3540 XThR.XTB5.A XThR.XTB6.Y 0.00193f
C3541 XThR.Tn[6] XA.XIR[7].XIC[2].icell.Ien 0.00338f
C3542 XThR.Tn[2] XA.XIR[3].XIC[0].icell.Ien 0.00338f
C3543 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00584f
C3544 XThR.Tn[13] a_n997_1579# 0.19413f
C3545 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00584f
C3546 XA.XIR[10].XIC[11].icell.PDM Iout 0.00117f
C3547 XA.XIR[12].XIC[2].icell.Ien VPWR 0.1903f
C3548 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04031f
C3549 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00256f
C3550 XA.XIR[14].XIC[12].icell.SM Iout 0.00388f
C3551 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07079f
C3552 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00584f
C3553 XA.XIR[11].XIC[3].icell.SM VPWR 0.00158f
C3554 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.SM 0.00168f
C3555 XThC.XTB7.Y VPWR 1.07717f
C3556 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00214f
C3557 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C3558 XA.XIR[9].XIC[11].icell.PDM Iout 0.00117f
C3559 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9] 0.00341f
C3560 XA.XIR[3].XIC[9].icell.PUM Vbias 0.0031f
C3561 XA.XIR[1].XIC[9].icell.PDM Vbias 0.04261f
C3562 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PUM 0.00465f
C3563 XA.XIR[13].XIC[12].icell.PDM Iout 0.00117f
C3564 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.SM 0.0039f
C3565 XA.XIR[6].XIC[12].icell.SM Vbias 0.00701f
C3566 XA.XIR[9].XIC[13].icell.PUM VPWR 0.00937f
C3567 XA.XIR[10].XIC[5].icell.SM VPWR 0.00158f
C3568 XA.XIR[10].XIC[13].icell.SM Vbias 0.00701f
C3569 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C3570 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11] 0.00341f
C3571 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C3572 XThR.Tn[14] XA.XIR[15].XIC[2].icell.Ien 0.00338f
C3573 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.15202f
C3574 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.SM 0.0039f
C3575 XA.XIR[1].XIC[0].icell.SM Iout 0.00388f
C3576 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PUM 0.00465f
C3577 XA.XIR[7].XIC[2].icell.Ien Vbias 0.21098f
C3578 XA.XIR[4].XIC[9].icell.PDM Vbias 0.04261f
C3579 XA.XIR[10].XIC[1].icell.SM Iout 0.00388f
C3580 XA.XIR[5].XIC_15.icell.Ien Vbias 0.21234f
C3581 XThR.Tn[9] XA.XIR[10].XIC[1].icell.SM 0.00121f
C3582 XA.XIR[0].XIC[6].icell.PUM VPWR 0.00877f
C3583 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C3584 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.SM 0.00168f
C3585 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00214f
C3586 XThR.XTBN.A XThR.Tn[9] 0.12398f
C3587 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PUM 0.00465f
C3588 XA.XIR[1].XIC[4].icell.PUM Vbias 0.0031f
C3589 XA.XIR[3].XIC[14].icell.SM VPWR 0.00207f
C3590 XA.XIR[14].XIC[6].icell.SM Vbias 0.00701f
C3591 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C3592 XA.XIR[12].XIC_15.icell.PDM Vbias 0.04401f
C3593 XThR.Tn[6] Iout 1.1623f
C3594 XA.XIR[11].XIC[14].icell.Ien Iout 0.06417f
C3595 XA.XIR[3].XIC[10].icell.SM Iout 0.00388f
C3596 XA.XIR[12].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3597 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C3598 XA.XIR[13].XIC[8].icell.SM Vbias 0.00701f
C3599 XA.XIR[2].XIC[7].icell.SM VPWR 0.00158f
C3600 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.SM 0.00168f
C3601 XA.XIR[6].XIC_15.icell.Ien Iout 0.0642f
C3602 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3603 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[7].icell.SM 0.0039f
C3604 XA.XIR[8].XIC[12].icell.PUM Vbias 0.0031f
C3605 XA.XIR[7].XIC[9].icell.PUM VPWR 0.00937f
C3606 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02764f
C3607 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.SM 0.00168f
C3608 XA.XIR[1].XIC[9].icell.SM VPWR 0.00158f
C3609 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C3610 XA.XIR[2].XIC[3].icell.SM Iout 0.00388f
C3611 XThC.Tn[8] XThR.Tn[14] 0.28739f
C3612 XThR.XTB6.A VPWR 0.68638f
C3613 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00214f
C3614 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04031f
C3615 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C3616 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.SM 0.0039f
C3617 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39f
C3618 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C3619 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C3620 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02762f
C3621 XA.XIR[1].XIC[5].icell.SM Iout 0.00388f
C3622 XA.XIR[14].XIC[9].icell.Ien Iout 0.06417f
C3623 XThC.Tn[8] data[0] 0.01643f
C3624 Vbias Iout 83.1596f
C3625 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00214f
C3626 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.SM 0.0039f
C3627 XThR.Tn[9] Vbias 3.74874f
C3628 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.03023f
C3629 XThR.XTB1.Y a_n1049_8581# 0.21263f
C3630 XThC.XTB3.Y a_5155_9615# 0.00913f
C3631 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.0352f
C3632 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.15202f
C3633 XA.XIR[8].XIC[13].icell.SM Iout 0.00388f
C3634 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.SM 0.00168f
C3635 XA.XIR[0].XIC[14].icell.PUM Vbias 0.0031f
C3636 XThR.Tn[8] XA.XIR[9].XIC[13].icell.SM 0.00121f
C3637 XThR.Tn[11] XA.XIR[12].XIC[2].icell.SM 0.00121f
C3638 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C3639 XA.XIR[6].XIC[0].icell.PUM VPWR 0.00937f
C3640 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C3641 XThR.Tn[0] VPWR 6.66912f
C3642 XThR.Tn[12] XA.XIR[13].XIC[14].icell.Ien 0.00338f
C3643 XThR.Tn[2] XA.XIR[3].XIC[8].icell.Ien 0.00338f
C3644 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C3645 XThR.Tn[4] XA.XIR[4].XIC[9].icell.PDM 0.00341f
C3646 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.SM 0.0039f
C3647 XThR.Tn[4] XA.XIR[5].XIC_15.icell.Ien 0.00117f
C3648 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04031f
C3649 XThR.XTB7.B a_n997_3755# 0.01174f
C3650 XA.XIR[10].XIC[1].icell.PUM VPWR 0.00937f
C3651 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C3652 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C3653 XThR.Tn[3] XA.XIR[3].XIC[10].icell.PDM 0.00341f
C3654 XThR.Tn[3] XA.XIR[4].XIC_15.icell.Ien 0.00117f
C3655 XThC.Tn[4] XThR.Tn[6] 0.28739f
C3656 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C3657 XThR.Tn[1] XA.XIR[2].XIC[6].icell.SM 0.00121f
C3658 XThR.XTBN.Y XThR.Tn[8] 0.47811f
C3659 XA.XIR[15].XIC[0].icell.Ien Vbias 0.17752f
C3660 XA.XIR[6].XIC[6].icell.PDM VPWR 0.00799f
C3661 XA.XIR[5].XIC[0].icell.SM Vbias 0.00675f
C3662 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C3663 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00256f
C3664 XA.XIR[5].XIC[13].icell.PDM VPWR 0.00799f
C3665 XA.XIR[14].XIC[3].icell.PDM VPWR 0.00799f
C3666 XA.XIR[14].XIC[2].icell.PUM Vbias 0.0031f
C3667 XA.XIR[14].XIC[10].icell.SM Iout 0.00388f
C3668 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.03425f
C3669 XThC.Tn[6] XThR.Tn[11] 0.28739f
C3670 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PUM 0.00465f
C3671 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.SM 0.00168f
C3672 XA.XIR[13].XIC[7].icell.PDM VPWR 0.00799f
C3673 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C3674 XA.XIR[5].XIC[1].icell.PDM Iout 0.00117f
C3675 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.SM 0.00168f
C3676 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC_15.icell.Ien 0.00214f
C3677 XA.XIR[10].XIC[3].icell.PDM Vbias 0.04261f
C3678 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C3679 XA.XIR[10].XIC[11].icell.SM Vbias 0.00701f
C3680 XThC.Tn[4] Vbias 2.48532f
C3681 XThC.XTB7.Y a_9827_9569# 0.00571f
C3682 XA.XIR[6].XIC[0].icell.SM Iout 0.00388f
C3683 XThR.XTB7.B a_n1049_5611# 0.00927f
C3684 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PUM 0.00465f
C3685 XThR.Tn[4] Iout 1.16233f
C3686 XThR.Tn[0] XA.XIR[1].XIC[13].icell.SM 0.00121f
C3687 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C3688 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C3689 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00584f
C3690 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C3691 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00214f
C3692 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02762f
C3693 XA.XIR[12].XIC[0].icell.PDM Iout 0.00117f
C3694 XA.XIR[6].XIC[4].icell.PUM Vbias 0.0031f
C3695 XA.XIR[9].XIC[3].icell.Ien VPWR 0.1903f
C3696 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PUM 0.00465f
C3697 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C3698 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00584f
C3699 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00584f
C3700 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C3701 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.03425f
C3702 XThR.XTB2.Y XThR.Tn[2] 0.00271f
C3703 XThC.XTB5.Y XThC.Tn[7] 0.00912f
C3704 XA.XIR[11].XIC[6].icell.PDM Iout 0.00117f
C3705 XA.XIR[15].XIC[5].icell.Ien Vbias 0.17899f
C3706 XA.XIR[5].XIC[5].icell.SM Vbias 0.00701f
C3707 XA.XIR[11].XIC[12].icell.Ien Iout 0.06417f
C3708 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.SM 0.00168f
C3709 XThC.Tn[10] XThR.Tn[13] 0.28739f
C3710 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02762f
C3711 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.03425f
C3712 XA.XIR[10].XIC[10].icell.PDM Iout 0.00117f
C3713 XThC.Tn[0] XThR.Tn[1] 0.28748f
C3714 XA.XIR[3].XIC[6].icell.PUM VPWR 0.00937f
C3715 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04031f
C3716 XA.XIR[4].XIC[8].icell.Ien Vbias 0.21098f
C3717 XThR.Tn[8] XThR.Tn[10] 0.00255f
C3718 XA.XIR[1].XIC[0].icell.PDM VPWR 0.00799f
C3719 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02762f
C3720 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C3721 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02762f
C3722 XA.XIR[6].XIC[9].icell.SM VPWR 0.00158f
C3723 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C3724 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C3725 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PUM 0.00465f
C3726 XThC.Tn[13] Iout 0.84238f
C3727 XThR.XTB7.A XThR.Tn[3] 0.0306f
C3728 XThC.Tn[13] XThR.Tn[9] 0.2874f
C3729 XThR.Tn[4] XA.XIR[5].XIC[0].icell.SM 0.00121f
C3730 XThC.Tn[0] XThR.Tn[12] 0.28741f
C3731 XA.XIR[4].XIC[0].icell.PDM VPWR 0.00799f
C3732 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C3733 XA.XIR[8].XIC[2].icell.Ien Vbias 0.21098f
C3734 XA.XIR[5].XIC[12].icell.Ien VPWR 0.1903f
C3735 XA.XIR[6].XIC[5].icell.SM Iout 0.00388f
C3736 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7] 0.00341f
C3737 XThC.Tn[9] XThR.Tn[8] 0.28739f
C3738 XA.XIR[13].XIC[11].icell.PDM Iout 0.00117f
C3739 XThR.Tn[10] XA.XIR[11].XIC[1].icell.Ien 0.00338f
C3740 XA.XIR[10].XIC[14].icell.PUM Vbias 0.0031f
C3741 XA.XIR[15].XIC_15.icell.SM Vbias 0.00701f
C3742 XThR.Tn[3] XA.XIR[4].XIC[0].icell.SM 0.00121f
C3743 XThC.XTB6.A VPWR 0.68179f
C3744 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C3745 XA.XIR[3].XIC[8].icell.PDM VPWR 0.00799f
C3746 XA.XIR[5].XIC[8].icell.Ien Iout 0.06417f
C3747 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01577f
C3748 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00584f
C3749 XA.XIR[8].XIC[10].icell.PDM VPWR 0.00799f
C3750 XA.XIR[2].XIC[2].icell.PUM Vbias 0.0031f
C3751 XA.XIR[14].XIC[3].icell.SM VPWR 0.00158f
C3752 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C3753 XA.XIR[0].XIC[11].icell.PDM Vbias 0.04282f
C3754 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13] 0.00341f
C3755 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.0353f
C3756 XA.XIR[11].XIC[3].icell.PUM Vbias 0.0031f
C3757 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C3758 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.SM 0.00168f
C3759 XThC.XTBN.A a_7875_9569# 0.01939f
C3760 XA.XIR[2].XIC[14].icell.PDM VPWR 0.00809f
C3761 XThR.XTB7.A data[4] 0.8689f
C3762 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C3763 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C3764 XA.XIR[13].XIC[5].icell.SM VPWR 0.00158f
C3765 XA.XIR[13].XIC[13].icell.SM Vbias 0.00701f
C3766 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00214f
C3767 XThC.XTBN.Y XThC.Tn[7] 0.91493f
C3768 XA.XIR[9].XIC[11].icell.Ien Vbias 0.21098f
C3769 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04031f
C3770 XThC.Tn[4] XThR.Tn[4] 0.28739f
C3771 XThR.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.00338f
C3772 XA.XIR[8].XIC[9].icell.PUM VPWR 0.00937f
C3773 XA.XIR[10].XIC[5].icell.PUM Vbias 0.0031f
C3774 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C3775 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C3776 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C3777 XA.XIR[12].XIC[14].icell.PDM Vbias 0.04261f
C3778 XA.XIR[2].XIC[2].icell.PDM Iout 0.00117f
C3779 XThR.Tn[6] XA.XIR[7].XIC[7].icell.Ien 0.00338f
C3780 XA.XIR[13].XIC[1].icell.SM Iout 0.00388f
C3781 XA.XIR[12].XIC[7].icell.Ien VPWR 0.1903f
C3782 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.SM 0.00168f
C3783 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12] 0.00341f
C3784 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00584f
C3785 XA.XIR[0].XIC[4].icell.Ien Vbias 0.21127f
C3786 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3787 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Iout 0.00347f
C3788 XThC.XTB4.Y XThC.Tn[2] 0.0021f
C3789 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.03425f
C3790 XA.XIR[11].XIC[8].icell.SM VPWR 0.00158f
C3791 XA.XIR[12].XIC[3].icell.Ien Iout 0.06417f
C3792 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C3793 XThR.Tn[4] XA.XIR[5].XIC[5].icell.SM 0.00121f
C3794 XA.XIR[3].XIC[14].icell.PUM Vbias 0.0031f
C3795 XA.XIR[14].XIC[14].icell.Ien Iout 0.06417f
C3796 XA.XIR[15].XIC_15.icell.PDM Vbias 0.04401f
C3797 XA.XIR[11].XIC[4].icell.SM Iout 0.00388f
C3798 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.03425f
C3799 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C3800 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00584f
C3801 XThR.Tn[3] XA.XIR[4].XIC[5].icell.SM 0.00121f
C3802 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Iout 0.00347f
C3803 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.15202f
C3804 XThR.Tn[14] XA.XIR[15].XIC[7].icell.Ien 0.00338f
C3805 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PUM 0.00465f
C3806 XA.XIR[2].XIC[7].icell.PUM Vbias 0.0031f
C3807 XA.XIR[10].XIC[6].icell.SM Iout 0.00388f
C3808 XA.XIR[7].XIC[7].icell.Ien Vbias 0.21098f
C3809 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.SM 0.00168f
C3810 XA.XIR[0].XIC[11].icell.PUM VPWR 0.00878f
C3811 XThR.Tn[9] XA.XIR[10].XIC[6].icell.SM 0.00121f
C3812 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.15202f
C3813 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5] 0.00341f
C3814 XA.XIR[4].XIC_15.icell.SM Iout 0.0047f
C3815 XA.XIR[1].XIC[9].icell.PUM Vbias 0.0031f
C3816 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C3817 XThC.XTB7.A a_8739_10571# 0.00995f
C3818 XA.XIR[10].XIC[9].icell.SM Vbias 0.00701f
C3819 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04031f
C3820 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38993f
C3821 XThR.XTB3.Y a_n1049_5317# 0.00899f
C3822 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PUM 0.00465f
C3823 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PUM 0.00465f
C3824 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00214f
C3825 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04031f
C3826 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PUM 0.00471f
C3827 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C3828 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8] 0.00341f
C3829 XA.XIR[12].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3830 XA.XIR[2].XIC[12].icell.SM VPWR 0.00158f
C3831 XThR.XTBN.Y a_n997_3755# 0.229f
C3832 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C3833 XA.XIR[7].XIC[14].icell.PUM VPWR 0.00937f
C3834 XA.XIR[1].XIC[0].icell.Ien VPWR 0.1903f
C3835 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C3836 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6] 0.00341f
C3837 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.15202f
C3838 XA.XIR[1].XIC[14].icell.SM VPWR 0.00207f
C3839 XA.XIR[2].XIC[8].icell.SM Iout 0.00388f
C3840 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C3841 XA.XIR[11].XIC[10].icell.Ien Iout 0.06417f
C3842 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C3843 XThR.Tn[12] XA.XIR[13].XIC[4].icell.SM 0.00121f
C3844 XA.XIR[4].XIC[0].icell.Ien VPWR 0.1903f
C3845 XThR.Tn[1] VPWR 6.67344f
C3846 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02762f
C3847 XA.XIR[1].XIC[10].icell.SM Iout 0.00388f
C3848 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00584f
C3849 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PUM 0.00465f
C3850 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C3851 XA.XIR[13].XIC[1].icell.PUM VPWR 0.00937f
C3852 XA.XIR[0].XIC_15.icell.SM VPWR 0.00257f
C3853 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.15202f
C3854 XThC.XTBN.Y a_3773_9615# 0.08456f
C3855 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00584f
C3856 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.15202f
C3857 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C3858 XThR.Tn[12] VPWR 7.57625f
C3859 a_6243_9615# Vbias 0.01019f
C3860 XThR.XTB3.Y a_n1335_7243# 0.00941f
C3861 XThR.Tn[11] XA.XIR[12].XIC[7].icell.SM 0.00121f
C3862 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C3863 XA.XIR[6].XIC[2].icell.PDM Vbias 0.04261f
C3864 Vbias data[1] 0.00255f
C3865 XThR.XTBN.Y a_n1049_5611# 0.0768f
C3866 XThR.Tn[2] XA.XIR[3].XIC[13].icell.Ien 0.00338f
C3867 XA.XIR[10].XIC[12].icell.PUM Vbias 0.0031f
C3868 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C3869 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.SM 0.00168f
C3870 XThR.XTB4.Y a_n997_3755# 0.00497f
C3871 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C3872 XA.XIR[5].XIC[9].icell.PDM Vbias 0.04261f
C3873 XA.XIR[15].XIC[2].icell.Ien VPWR 0.32895f
C3874 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PUM 0.00465f
C3875 XThC.Tn[6] XThR.Tn[14] 0.28739f
C3876 XA.XIR[5].XIC[2].icell.SM VPWR 0.00158f
C3877 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C3878 XA.XIR[11].XIC[0].icell.Ien Iout 0.06411f
C3879 XA.XIR[7].XIC[14].icell.PDM VPWR 0.00809f
C3880 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C3881 a_10051_9569# XThC.Tn[12] 0.00623f
C3882 XA.XIR[13].XIC[3].icell.PDM Vbias 0.04261f
C3883 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.15202f
C3884 XThC.XTB3.Y a_7875_9569# 0.0061f
C3885 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00214f
C3886 XA.XIR[13].XIC[11].icell.SM Vbias 0.00701f
C3887 XA.XIR[7].XIC[2].icell.PDM Iout 0.00117f
C3888 XA.XIR[4].XIC[5].icell.Ien VPWR 0.1903f
C3889 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C3890 XThR.Tn[12] XA.XIR[13].XIC[10].icell.Ien 0.00338f
C3891 XThR.Tn[1] XA.XIR[2].XIC[11].icell.SM 0.00121f
C3892 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.03425f
C3893 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C3894 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C3895 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C3896 XThR.XTB2.Y XThR.Tn[10] 0.00106f
C3897 XA.XIR[12].XIC[8].icell.PDM Vbias 0.04261f
C3898 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.SM 0.0039f
C3899 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02762f
C3900 XA.XIR[15].XIC[0].icell.PDM Iout 0.00117f
C3901 XA.XIR[6].XIC[9].icell.PDM Iout 0.00117f
C3902 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C3903 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PUM 0.00465f
C3904 XThC.XTB2.Y XThC.Tn[2] 0.01113f
C3905 XA.XIR[9].XIC[1].icell.SM Vbias 0.00701f
C3906 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3907 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C3908 XA.XIR[14].XIC[6].icell.PDM Iout 0.00117f
C3909 XA.XIR[14].XIC[12].icell.Ien Iout 0.06417f
C3910 XThR.XTB4.Y a_n1049_5611# 0.00465f
C3911 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02762f
C3912 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PUM 0.00465f
C3913 XThR.XTB7.B XThR.Tn[3] 0.00532f
C3914 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.03425f
C3915 XThC.Tn[8] VPWR 6.8418f
C3916 XA.XIR[9].XIC[10].icell.PDM VPWR 0.00799f
C3917 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3918 XThR.XTB3.Y a_n1049_6405# 0.00913f
C3919 XA.XIR[13].XIC[10].icell.PDM Iout 0.00117f
C3920 XA.XIR[0].XIC[2].icell.PDM VPWR 0.00774f
C3921 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00214f
C3922 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02762f
C3923 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C3924 XA.XIR[3].XIC[4].icell.Ien Vbias 0.21098f
C3925 XA.XIR[10].XIC[13].icell.Ien Vbias 0.21098f
C3926 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00214f
C3927 XA.XIR[15].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3928 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.15202f
C3929 XA.XIR[9].XIC[8].icell.Ien VPWR 0.1903f
C3930 XA.XIR[6].XIC[9].icell.PUM Vbias 0.0031f
C3931 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C3932 XA.XIR[7].XIC[0].icell.PUM VPWR 0.00937f
C3933 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PUM 0.00465f
C3934 XThR.XTB7.B data[4] 0.01382f
C3935 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C3936 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C3937 XA.XIR[9].XIC[4].icell.Ien Iout 0.06417f
C3938 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.15202f
C3939 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.SM 0.00168f
C3940 XA.XIR[5].XIC[10].icell.SM Vbias 0.00701f
C3941 XA.XIR[13].XIC[14].icell.PUM Vbias 0.0031f
C3942 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PUM 0.00465f
C3943 XThC.XTB6.A XThC.XTB7.B 1.47641f
C3944 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00214f
C3945 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.03425f
C3946 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.SM 0.0039f
C3947 XThR.XTB5.Y a_n1319_6405# 0.01188f
C3948 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04031f
C3949 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C3950 XA.XIR[3].XIC[4].icell.PDM Vbias 0.04261f
C3951 a_n1049_5317# VPWR 0.72036f
C3952 XA.XIR[11].XIC[13].icell.SM VPWR 0.00158f
C3953 XA.XIR[12].XIC[13].icell.PDM Vbias 0.04261f
C3954 XA.XIR[3].XIC[11].icell.PUM VPWR 0.00937f
C3955 XA.XIR[4].XIC[13].icell.Ien Vbias 0.21098f
C3956 XA.XIR[14].XIC[3].icell.PUM Vbias 0.0031f
C3957 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.0353f
C3958 XA.XIR[8].XIC[6].icell.PDM Vbias 0.04261f
C3959 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10] 0.00341f
C3960 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07214f
C3961 XA.XIR[6].XIC[14].icell.SM VPWR 0.00207f
C3962 XA.XIR[2].XIC[10].icell.PDM Vbias 0.04261f
C3963 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14] 0.00341f
C3964 XA.XIR[1].XIC[3].icell.PDM Iout 0.00117f
C3965 XA.XIR[13].XIC[5].icell.PUM Vbias 0.0031f
C3966 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07214f
C3967 XA.XIR[2].XIC[4].icell.PUM VPWR 0.00937f
C3968 XA.XIR[8].XIC[7].icell.Ien Vbias 0.21098f
C3969 XA.XIR[6].XIC[10].icell.SM Iout 0.00388f
C3970 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C3971 XA.XIR[7].XIC[4].icell.Ien VPWR 0.1903f
C3972 XA.XIR[15].XIC[14].icell.PDM Vbias 0.04261f
C3973 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C3974 XA.XIR[12].XIC[5].icell.SM Vbias 0.00701f
C3975 XThR.Tn[2] XThR.Tn[3] 0.10553f
C3976 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C3977 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3978 XA.XIR[4].XIC[3].icell.PDM Iout 0.00117f
C3979 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C3980 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.SM 0.0039f
C3981 XA.XIR[1].XIC[6].icell.PUM VPWR 0.00937f
C3982 XA.XIR[5].XIC[13].icell.Ien Iout 0.06417f
C3983 XA.XIR[14].XIC[8].icell.SM VPWR 0.00158f
C3984 XA.XIR[10].XIC[14].icell.SM Vbias 0.00701f
C3985 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.15235f
C3986 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00214f
C3987 XA.XIR[11].XIC[8].icell.PUM Vbias 0.0031f
C3988 XA.XIR[8].XIC[13].icell.PDM Iout 0.00117f
C3989 XA.XIR[3].XIC[11].icell.PDM Iout 0.00117f
C3990 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04052f
C3991 XA.XIR[5].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3992 XA.XIR[14].XIC[4].icell.SM Iout 0.00388f
C3993 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.SM 0.00168f
C3994 XA.XIR[8].XIC[14].icell.PUM VPWR 0.00937f
C3995 XA.XIR[10].XIC[10].icell.PUM Vbias 0.0031f
C3996 XThC.Tn[2] Iout 0.84806f
C3997 XThR.Tn[6] XA.XIR[7].XIC[12].icell.Ien 0.00338f
C3998 XThC.Tn[2] XThR.Tn[9] 0.28739f
C3999 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00584f
C4000 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00214f
C4001 XA.XIR[3].XIC_15.icell.SM VPWR 0.00275f
C4002 XA.XIR[13].XIC[6].icell.SM Iout 0.00388f
C4003 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.SM 0.00168f
C4004 XA.XIR[0].XIC[9].icell.Ien Vbias 0.2113f
C4005 XA.XIR[11].XIC_15.icell.PDM Iout 0.00133f
C4006 XThR.XTBN.Y a_n997_715# 0.21503f
C4007 XA.XIR[11].XIC_15.icell.Ien Iout 0.0642f
C4008 XThR.Tn[0] XA.XIR[0].XIC[14].icell.PDM 0.00341f
C4009 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.15202f
C4010 XA.XIR[12].XIC[8].icell.Ien Iout 0.06417f
C4011 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.03425f
C4012 XThR.Tn[2] XA.XIR[3].XIC[3].icell.SM 0.00121f
C4013 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C4014 XThC.Tn[7] XThR.Tn[8] 0.28739f
C4015 VPWR data[7] 0.212f
C4016 XA.XIR[1].XIC_dummy_left.icell.SM VPWR 0.00269f
C4017 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C4018 XA.XIR[13].XIC[9].icell.SM Vbias 0.00701f
C4019 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.SM 0.00168f
C4020 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00214f
C4021 XThR.Tn[4] XA.XIR[5].XIC[10].icell.SM 0.00121f
C4022 XThR.Tn[1] XA.XIR[1].XIC[12].icell.PDM 0.00341f
C4023 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C4024 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.03547f
C4025 XThR.Tn[10] XA.XIR[11].XIC[2].icell.Ien 0.00338f
C4026 XA.XIR[4].XIC_dummy_left.icell.SM VPWR 0.00269f
C4027 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04031f
C4028 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.15202f
C4029 XThR.Tn[3] XA.XIR[4].XIC[10].icell.SM 0.00121f
C4030 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.SM 0.00168f
C4031 XA.XIR[2].XIC[12].icell.PUM Vbias 0.0031f
C4032 XA.XIR[7].XIC[12].icell.Ien Vbias 0.21098f
C4033 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.15202f
C4034 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C4035 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.03425f
C4036 XThR.XTB7.B a_n997_2667# 0.02071f
C4037 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C4038 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00214f
C4039 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.15202f
C4040 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04031f
C4041 XA.XIR[1].XIC[14].icell.PUM Vbias 0.0031f
C4042 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02762f
C4043 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.03425f
C4044 XA.XIR[14].XIC[10].icell.Ien Iout 0.06417f
C4045 XA.XIR[5].XIC[0].icell.PDM VPWR 0.00799f
C4046 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C4047 XThR.Tn[2] XA.XIR[2].XIC[9].icell.PDM 0.00341f
C4048 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PUM 0.00465f
C4049 XA.XIR[6].XIC[1].icell.PUM VPWR 0.00937f
C4050 XA.XIR[10].XIC[11].icell.Ien Vbias 0.21098f
C4051 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04031f
C4052 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.03425f
C4053 XThC.XTB3.Y XThC.Tn[4] 0.00382f
C4054 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[12].icell.SM 0.0039f
C4055 XA.XIR[3].XIC[1].icell.Ien Vbias 0.21098f
C4056 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C4057 a_n1049_6405# VPWR 0.72095f
C4058 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.15202f
C4059 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00584f
C4060 XThR.Tn[12] XA.XIR[13].XIC_15.icell.Ien 0.00117f
C4061 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.01438f
C4062 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C4063 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02762f
C4064 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C4065 XA.XIR[12].XIC[1].icell.PUM Vbias 0.0031f
C4066 XThC.Tn[2] XThC.Tn[4] 0.02725f
C4067 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.03425f
C4068 XA.XIR[2].XIC[13].icell.SM Iout 0.00388f
C4069 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.SM 0.0039f
C4070 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.SM 0.0039f
C4071 XA.XIR[13].XIC[12].icell.PUM Vbias 0.0031f
C4072 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C4073 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C4074 XA.XIR[11].XIC[5].icell.PDM VPWR 0.00799f
C4075 XA.XIR[11].XIC[11].icell.SM VPWR 0.00158f
C4076 XA.XIR[4].XIC[1].icell.Ien Iout 0.06417f
C4077 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00214f
C4078 XA.XIR[10].XIC[9].icell.PDM VPWR 0.00799f
C4079 XA.XIR[7].XIC[10].icell.PDM Vbias 0.04261f
C4080 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.03425f
C4081 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C4082 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.03425f
C4083 XA.XIR[15].XIC[8].icell.PDM Vbias 0.04261f
C4084 XA.XIR[4].XIC[3].icell.SM Vbias 0.00701f
C4085 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.SM 0.0039f
C4086 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01432f
C4087 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C4088 XThR.XTBN.Y XThR.Tn[3] 0.62502f
C4089 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.SM 0.00168f
C4090 a_n1049_8581# XThR.Tn[0] 0.2685f
C4091 XA.XIR[6].XIC[6].icell.PUM VPWR 0.00937f
C4092 XThR.XTB7.B XThR.Tn[11] 0.03888f
C4093 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00584f
C4094 XThC.Tn[10] XThR.Tn[7] 0.28739f
C4095 XThC.XTBN.A data[1] 0.01444f
C4096 XA.XIR[15].XIC[7].icell.Ien VPWR 0.32895f
C4097 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C4098 XA.XIR[5].XIC[7].icell.SM VPWR 0.00158f
C4099 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.03425f
C4100 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.03425f
C4101 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.15202f
C4102 XThC.XTB7.B XThC.Tn[8] 0.09736f
C4103 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.389f
C4104 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C4105 XA.XIR[15].XIC[3].icell.Ien Iout 0.06807f
C4106 XA.XIR[9].XIC[6].icell.PDM Vbias 0.04261f
C4107 a_8963_9569# Vbias 0.00243f
C4108 XA.XIR[4].XIC[10].icell.Ien VPWR 0.1903f
C4109 XA.XIR[5].XIC[3].icell.SM Iout 0.00388f
C4110 XThC.XTB7.Y XThC.Tn[12] 0.07222f
C4111 XA.XIR[13].XIC[13].icell.Ien Vbias 0.21098f
C4112 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PUM 0.00465f
C4113 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18966f
C4114 XA.XIR[2].XIC[1].icell.PDM VPWR 0.00799f
C4115 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Iout 0.00347f
C4116 XA.XIR[4].XIC[6].icell.Ien Iout 0.06417f
C4117 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00214f
C4118 XA.XIR[12].XIC[12].icell.PDM Vbias 0.04261f
C4119 XA.XIR[11].XIC[14].icell.PUM VPWR 0.00937f
C4120 XA.XIR[9].XIC[6].icell.SM Vbias 0.00701f
C4121 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.SM 0.0039f
C4122 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C4123 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PUM 0.00465f
C4124 XA.XIR[8].XIC[4].icell.Ien VPWR 0.1903f
C4125 XThR.Tn[13] XA.XIR[14].XIC[1].icell.Ien 0.00338f
C4126 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C4127 XThR.Tn[6] XA.XIR[7].XIC[2].icell.SM 0.00121f
C4128 XThR.Tn[2] XA.XIR[3].XIC[0].icell.SM 0.00121f
C4129 XA.XIR[12].XIC[2].icell.SM VPWR 0.00158f
C4130 XA.XIR[15].XIC[13].icell.PDM Vbias 0.04261f
C4131 XA.XIR[14].XIC[13].icell.SM VPWR 0.00158f
C4132 XThC.Tn[2] XA.XIR[0].XIC[4].icell.Ien 0.00191f
C4133 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C4134 XA.XIR[11].XIC[5].icell.PUM VPWR 0.00937f
C4135 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PUM 0.00465f
C4136 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04031f
C4137 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C4138 XA.XIR[9].XIC[13].icell.PDM Iout 0.00117f
C4139 XA.XIR[3].XIC[9].icell.Ien Vbias 0.21098f
C4140 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00214f
C4141 XA.XIR[1].XIC[11].icell.PDM Vbias 0.04261f
C4142 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9] 0.00341f
C4143 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.03425f
C4144 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00214f
C4145 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.SM 0.0039f
C4146 XA.XIR[7].XIC[0].icell.Ien Iout 0.06411f
C4147 XA.XIR[9].XIC[13].icell.Ien VPWR 0.1903f
C4148 XA.XIR[6].XIC[14].icell.PUM Vbias 0.0031f
C4149 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00584f
C4150 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C4151 XA.XIR[10].XIC[7].icell.PUM VPWR 0.00937f
C4152 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11] 0.00341f
C4153 XThR.Tn[14] XA.XIR[15].XIC[2].icell.SM 0.00121f
C4154 XA.XIR[9].XIC[9].icell.Ien Iout 0.06417f
C4155 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.03425f
C4156 XA.XIR[2].XIC[2].icell.Ien Vbias 0.21098f
C4157 XA.XIR[4].XIC[11].icell.PDM Vbias 0.04261f
C4158 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.15202f
C4159 XThC.Tn[9] XThR.Tn[3] 0.28739f
C4160 XA.XIR[7].XIC[2].icell.SM Vbias 0.00701f
C4161 XA.XIR[0].XIC[6].icell.Ien VPWR 0.18973f
C4162 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00584f
C4163 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C4164 XThR.Tn[7] XA.XIR[8].XIC[1].icell.Ien 0.00338f
C4165 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.03425f
C4166 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C4167 XA.XIR[13].XIC[14].icell.SM Vbias 0.00701f
C4168 XA.XIR[1].XIC[4].icell.Ien Vbias 0.21104f
C4169 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C4170 XA.XIR[14].XIC[8].icell.PUM Vbias 0.0031f
C4171 XA.XIR[0].XIC[2].icell.Ien Iout 0.06389f
C4172 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4173 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Iout 0.00347f
C4174 XA.XIR[11].XIC[14].icell.PDM Iout 0.00117f
C4175 XThC.Tn[6] VPWR 5.90436f
C4176 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.SM 0.0039f
C4177 XA.XIR[13].XIC[10].icell.PUM Vbias 0.0031f
C4178 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C4179 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8] 0.00341f
C4180 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.15222f
C4181 XA.XIR[7].XIC[9].icell.Ien VPWR 0.1903f
C4182 XA.XIR[2].XIC[9].icell.PUM VPWR 0.00937f
C4183 XA.XIR[8].XIC[12].icell.Ien Vbias 0.21098f
C4184 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.15202f
C4185 XA.XIR[11].XIC[9].icell.SM VPWR 0.00158f
C4186 XThC.Tn[12] XThR.Tn[0] 0.28786f
C4187 XA.XIR[14].XIC_15.icell.PDM Iout 0.00133f
C4188 XA.XIR[14].XIC_15.icell.Ien Iout 0.0642f
C4189 XA.XIR[7].XIC[5].icell.Ien Iout 0.06417f
C4190 XA.XIR[1].XIC[11].icell.PUM VPWR 0.00937f
C4191 XThC.Tn[14] XThR.Tn[5] 0.28745f
C4192 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.SM 0.00168f
C4193 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04031f
C4194 XThR.XTBN.Y a_n997_2667# 0.22784f
C4195 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.SM 0.00168f
C4196 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PUM 0.00465f
C4197 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C4198 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.SM 0.0039f
C4199 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C4200 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C4201 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C4202 XThR.Tn[7] XA.XIR[8].XIC[6].icell.Ien 0.00338f
C4203 XThC.XTB3.Y a_6243_9615# 0.00899f
C4204 XThR.Tn[8] a_n997_3979# 0.1927f
C4205 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C4206 XThR.Tn[5] XA.XIR[6].XIC[2].icell.Ien 0.00338f
C4207 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PUM 0.00186f
C4208 XA.XIR[2].XIC[0].icell.Ien VPWR 0.1903f
C4209 XA.XIR[0].XIC[14].icell.Ien Vbias 0.2113f
C4210 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.03425f
C4211 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.SM 0.00168f
C4212 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02762f
C4213 XThR.Tn[2] XA.XIR[3].XIC[8].icell.SM 0.00121f
C4214 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.15202f
C4215 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02762f
C4216 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04031f
C4217 XThR.Tn[4] XA.XIR[4].XIC[11].icell.PDM 0.00341f
C4218 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01746f
C4219 XA.XIR[13].XIC[11].icell.Ien Vbias 0.21098f
C4220 XA.XIR[7].XIC[1].icell.PDM VPWR 0.00799f
C4221 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00584f
C4222 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.03425f
C4223 XThR.Tn[10] XA.XIR[11].XIC[7].icell.Ien 0.00338f
C4224 XA.XIR[10].XIC[1].icell.Ien VPWR 0.1903f
C4225 XA.XIR[1].XIC_15.icell.SM VPWR 0.00275f
C4226 XThR.Tn[3] XA.XIR[3].XIC[12].icell.PDM 0.00341f
C4227 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00214f
C4228 XA.XIR[11].XIC[12].icell.PUM VPWR 0.00937f
C4229 XThR.XTB4.Y a_n997_2667# 0.07199f
C4230 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.15202f
C4231 XA.XIR[15].XIC[0].icell.SM Vbias 0.00675f
C4232 XA.XIR[6].XIC[8].icell.PDM VPWR 0.00799f
C4233 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.15202f
C4234 XA.XIR[5].XIC[2].icell.PUM Vbias 0.0031f
C4235 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02762f
C4236 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C4237 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.SM 0.00168f
C4238 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.15202f
C4239 XA.XIR[14].XIC[5].icell.PDM VPWR 0.00799f
C4240 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07214f
C4241 XA.XIR[14].XIC[11].icell.SM VPWR 0.00158f
C4242 XA.XIR[11].XIC[1].icell.PDM Vbias 0.04261f
C4243 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00214f
C4244 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.03425f
C4245 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C4246 XThR.XTBN.Y XThR.Tn[11] 0.52266f
C4247 XA.XIR[13].XIC[9].icell.PDM VPWR 0.00799f
C4248 XA.XIR[5].XIC[3].icell.PDM Iout 0.00117f
C4249 XThC.Tn[11] XThR.Tn[2] 0.28739f
C4250 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00214f
C4251 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C4252 XA.XIR[10].XIC[5].icell.PDM Vbias 0.04261f
C4253 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.15202f
C4254 XThC.XTB7.Y a_10915_9569# 0.06874f
C4255 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C4256 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PUM 0.00186f
C4257 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.SM 0.00168f
C4258 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.SM 0.00168f
C4259 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C4260 XA.XIR[12].XIC[2].icell.PDM Iout 0.00117f
C4261 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PUM 0.00465f
C4262 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.SM 0.00168f
C4263 XA.XIR[6].XIC[4].icell.Ien Vbias 0.21098f
C4264 XA.XIR[9].XIC[3].icell.SM VPWR 0.00158f
C4265 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.03425f
C4266 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.SM 0.00168f
C4267 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00584f
C4268 XA.XIR[15].XIC[5].icell.SM Vbias 0.00701f
C4269 XA.XIR[5].XIC[7].icell.PUM Vbias 0.0031f
C4270 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C4271 XA.XIR[11].XIC[8].icell.PDM Iout 0.00117f
C4272 XA.XIR[11].XIC[13].icell.Ien VPWR 0.1903f
C4273 XA.XIR[12].XIC[11].icell.PDM Vbias 0.04261f
C4274 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C4275 XThR.Tn[7] XThR.Tn[8] 0.07425f
C4276 XThR.XTB7.Y a_n997_1803# 0.00571f
C4277 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.SM 0.0039f
C4278 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C4279 XThC.XTB7.A XThC.Tn[7] 0.00184f
C4280 XA.XIR[4].XIC[8].icell.SM Vbias 0.00701f
C4281 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00214f
C4282 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C4283 XA.XIR[3].XIC[6].icell.Ien VPWR 0.1903f
C4284 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.15202f
C4285 XA.XIR[1].XIC[2].icell.PDM VPWR 0.00799f
C4286 XA.XIR[6].XIC[11].icell.PUM VPWR 0.00937f
C4287 XA.XIR[14].XIC[14].icell.PUM VPWR 0.00937f
C4288 XA.XIR[15].XIC[12].icell.PDM Vbias 0.04261f
C4289 XA.XIR[3].XIC[2].icell.Ien Iout 0.06417f
C4290 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PUM 0.00465f
C4291 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00584f
C4292 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.03425f
C4293 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.SM 0.00168f
C4294 XA.XIR[8].XIC[2].icell.SM Vbias 0.00701f
C4295 XA.XIR[4].XIC[2].icell.PDM VPWR 0.00799f
C4296 XA.XIR[5].XIC[12].icell.SM VPWR 0.00158f
C4297 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7] 0.00341f
C4298 XThR.Tn[10] XThR.Tn[11] 0.05908f
C4299 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00214f
C4300 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.SM 0.0039f
C4301 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.SM 0.00168f
C4302 XA.XIR[15].XIC[8].icell.Ien Iout 0.06807f
C4303 XA.XIR[8].XIC[12].icell.PDM VPWR 0.00799f
C4304 XA.XIR[5].XIC[8].icell.SM Iout 0.00388f
C4305 XA.XIR[3].XIC[10].icell.PDM VPWR 0.00799f
C4306 XA.XIR[4].XIC_15.icell.Ien VPWR 0.25566f
C4307 XA.XIR[14].XIC[5].icell.PUM VPWR 0.00937f
C4308 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.SM 0.00168f
C4309 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C4310 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PUM 0.00429f
C4311 XA.XIR[0].XIC[13].icell.PDM Vbias 0.04282f
C4312 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13] 0.00341f
C4313 XA.XIR[11].XIC[3].icell.Ien Vbias 0.21098f
C4314 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C4315 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.SM 0.0039f
C4316 XThC.Tn[9] XThR.Tn[11] 0.28739f
C4317 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C4318 XThC.XTBN.A a_8963_9569# 0.01679f
C4319 XA.XIR[8].XIC[0].icell.PDM Iout 0.00117f
C4320 XA.XIR[4].XIC[11].icell.Ien Iout 0.06417f
C4321 XA.XIR[13].XIC[7].icell.PUM VPWR 0.00937f
C4322 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04031f
C4323 XA.XIR[8].XIC[9].icell.Ien VPWR 0.1903f
C4324 XA.XIR[9].XIC[11].icell.SM Vbias 0.00701f
C4325 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04031f
C4326 XA.XIR[10].XIC[5].icell.Ien Vbias 0.21098f
C4327 XThR.Tn[6] XA.XIR[7].XIC[7].icell.SM 0.00121f
C4328 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02762f
C4329 XA.XIR[2].XIC[4].icell.PDM Iout 0.00117f
C4330 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C4331 XA.XIR[11].XIC[13].icell.PDM Iout 0.00117f
C4332 XA.XIR[11].XIC[14].icell.SM VPWR 0.00207f
C4333 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C4334 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C4335 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.SM 0.0039f
C4336 XA.XIR[12].XIC[7].icell.SM VPWR 0.00158f
C4337 XA.XIR[8].XIC[5].icell.Ien Iout 0.06417f
C4338 XA.XIR[6].XIC_15.icell.SM VPWR 0.00275f
C4339 XA.XIR[0].XIC[4].icell.SM Vbias 0.00716f
C4340 XThR.Tn[8] XA.XIR[9].XIC[5].icell.Ien 0.00338f
C4341 XThR.XTB6.A a_n1319_5317# 0.00295f
C4342 XA.XIR[12].XIC[3].icell.SM Iout 0.00388f
C4343 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C4344 XThR.Tn[0] XA.XIR[0].XIC[1].icell.PDM 0.00341f
C4345 XA.XIR[11].XIC[10].icell.PUM VPWR 0.00937f
C4346 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00214f
C4347 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00584f
C4348 XA.XIR[3].XIC[14].icell.Ien Vbias 0.21098f
C4349 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.SM 0.0039f
C4350 XThC.XTB7.B XThC.Tn[6] 0.05039f
C4351 XA.XIR[14].XIC[14].icell.PDM Iout 0.00117f
C4352 VPWR data[3] 0.20846f
C4353 XThC.XTB5.Y XThC.Tn[10] 0.01742f
C4354 XThR.XTB2.Y a_n997_3979# 0.00191f
C4355 XThR.Tn[14] XA.XIR[15].XIC[7].icell.SM 0.00121f
C4356 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.03425f
C4357 XThC.XTB6.Y XThC.Tn[14] 0.00128f
C4358 XA.XIR[14].XIC[9].icell.SM VPWR 0.00158f
C4359 XA.XIR[9].XIC[14].icell.Ien Iout 0.06417f
C4360 XA.XIR[2].XIC[7].icell.Ien Vbias 0.21098f
C4361 XA.XIR[7].XIC[7].icell.SM Vbias 0.00701f
C4362 XA.XIR[10].XIC_15.icell.SM Vbias 0.00701f
C4363 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C4364 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.15202f
C4365 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.0404f
C4366 XA.XIR[0].XIC[11].icell.Ien VPWR 0.19072f
C4367 XThC.XTB5.Y a_4861_9615# 0.0021f
C4368 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.SM 0.0039f
C4369 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C4370 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5] 0.00341f
C4371 XA.XIR[1].XIC[9].icell.Ien Vbias 0.21104f
C4372 XThC.Tn[12] XThR.Tn[1] 0.28739f
C4373 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00214f
C4374 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.SM 0.00168f
C4375 XA.XIR[0].XIC[7].icell.Ien Iout 0.06389f
C4376 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04052f
C4377 XA.XIR[2].XIC_dummy_left.icell.SM VPWR 0.00269f
C4378 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C4379 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.03431f
C4380 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.04036f
C4381 XThR.Tn[13] XA.XIR[14].XIC[2].icell.Ien 0.00338f
C4382 XA.XIR[11].XIC[0].icell.PUM VPWR 0.00937f
C4383 XA.XIR[2].XIC[14].icell.PUM VPWR 0.00937f
C4384 XThC.Tn[12] XThR.Tn[12] 0.28739f
C4385 XA.XIR[7].XIC[14].icell.Ien VPWR 0.19036f
C4386 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C4387 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00584f
C4388 XThR.XTB7.A VPWR 0.88595f
C4389 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.15202f
C4390 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6] 0.00341f
C4391 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.15202f
C4392 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00214f
C4393 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00584f
C4394 XA.XIR[7].XIC[10].icell.Ien Iout 0.06417f
C4395 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.04497f
C4396 XThR.Tn[0] XA.XIR[1].XIC[5].icell.Ien 0.00338f
C4397 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02762f
C4398 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4399 XA.XIR[11].XIC[11].icell.Ien VPWR 0.1903f
C4400 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.SM 0.00168f
C4401 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.SM 0.00168f
C4402 XA.XIR[4].XIC[0].icell.SM VPWR 0.00158f
C4403 XThC.Tn[7] XThR.Tn[3] 0.28739f
C4404 XThR.XTB5.Y XThR.Tn[6] 0.00349f
C4405 XThC.XTBN.Y XThC.Tn[10] 0.51405f
C4406 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C4407 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02762f
C4408 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.SM 0.00168f
C4409 XA.XIR[13].XIC[1].icell.Ien VPWR 0.1903f
C4410 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.SM 0.0039f
C4411 XThR.Tn[7] XA.XIR[8].XIC[11].icell.Ien 0.00338f
C4412 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00584f
C4413 XA.XIR[14].XIC[12].icell.PUM VPWR 0.00937f
C4414 XThC.XTBN.Y a_4861_9615# 0.07601f
C4415 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00584f
C4416 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00214f
C4417 XThR.Tn[5] XA.XIR[6].XIC[7].icell.Ien 0.00338f
C4418 XA.XIR[8].XIC[0].icell.Ien Iout 0.06411f
C4419 XA.XIR[6].XIC[4].icell.PDM Vbias 0.04261f
C4420 XThR.Tn[8] XA.XIR[9].XIC[0].icell.Ien 0.00338f
C4421 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.SM 0.0039f
C4422 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.02762f
C4423 XThC.Tn[1] XThR.Tn[0] 0.28784f
C4424 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.SM 0.0039f
C4425 XThC.Tn[11] XThR.Tn[10] 0.28739f
C4426 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[1].icell.Ien 0.00214f
C4427 XThC.Tn[3] XThR.Tn[5] 0.28739f
C4428 XThR.Tn[2] XA.XIR[3].XIC[13].icell.SM 0.00121f
C4429 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C4430 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00214f
C4431 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C4432 XA.XIR[5].XIC[11].icell.PDM Vbias 0.04261f
C4433 XA.XIR[14].XIC[1].icell.PDM Vbias 0.04261f
C4434 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C4435 XThC.XTB5.Y a_5155_10571# 0.01188f
C4436 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.SM 0.00168f
C4437 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.03425f
C4438 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C4439 XA.XIR[15].XIC[2].icell.SM VPWR 0.00158f
C4440 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PUM 0.00465f
C4441 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C4442 XA.XIR[5].XIC[4].icell.PUM VPWR 0.00937f
C4443 XThC.Tn[9] XThC.Tn[11] 0.00252f
C4444 XA.XIR[13].XIC[5].icell.PDM Vbias 0.04261f
C4445 XThC.XTB3.Y a_8963_9569# 0.002f
C4446 XThR.XTB6.A a_n1319_6405# 0.00306f
C4447 XA.XIR[4].XIC[5].icell.SM VPWR 0.00158f
C4448 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C4449 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02762f
C4450 XA.XIR[7].XIC[4].icell.PDM Iout 0.00117f
C4451 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00214f
C4452 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.SM 0.0039f
C4453 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00214f
C4454 XA.XIR[12].XIC[10].icell.PDM Vbias 0.04261f
C4455 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.SM 0.0039f
C4456 XA.XIR[4].XIC[1].icell.SM Iout 0.00388f
C4457 XA.XIR[15].XIC[2].icell.PDM Iout 0.00117f
C4458 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.15202f
C4459 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.03425f
C4460 XA.XIR[6].XIC[11].icell.PDM Iout 0.00117f
C4461 XA.XIR[9].XIC[3].icell.PUM Vbias 0.0031f
C4462 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00584f
C4463 XA.XIR[14].XIC[8].icell.PDM Iout 0.00117f
C4464 XA.XIR[14].XIC[13].icell.Ien VPWR 0.19084f
C4465 XA.XIR[15].XIC[11].icell.PDM Vbias 0.04261f
C4466 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C4467 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00584f
C4468 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.03023f
C4469 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00584f
C4470 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00584f
C4471 XA.XIR[9].XIC[12].icell.PDM VPWR 0.00799f
C4472 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C4473 XA.XIR[0].XIC[4].icell.PDM VPWR 0.00777f
C4474 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.SM 0.00168f
C4475 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C4476 XA.XIR[3].XIC[4].icell.SM Vbias 0.00701f
C4477 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.SM 0.0039f
C4478 XA.XIR[9].XIC[0].icell.PDM Iout 0.00117f
C4479 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9] 0.00341f
C4480 XA.XIR[1].XIC[1].icell.Ien VPWR 0.1903f
C4481 XA.XIR[9].XIC[8].icell.SM VPWR 0.00158f
C4482 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C4483 XThR.Tn[12] XA.XIR[13].XIC[0].icell.Ien 0.00368f
C4484 XA.XIR[6].XIC[9].icell.Ien Vbias 0.21098f
C4485 XA.XIR[10].XIC[2].icell.Ien VPWR 0.1903f
C4486 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.03425f
C4487 XThR.Tn[11] XThR.Tn[13] 0.00153f
C4488 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00214f
C4489 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.SM 0.00168f
C4490 XA.XIR[5].XIC[12].icell.PUM Vbias 0.0031f
C4491 XA.XIR[9].XIC[4].icell.SM Iout 0.00388f
C4492 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C4493 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.03425f
C4494 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04031f
C4495 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.03425f
C4496 XA.XIR[0].XIC[1].icell.SM VPWR 0.00158f
C4497 XThC.Tn[0] XThR.Tn[2] 0.28748f
C4498 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C4499 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04031f
C4500 XA.XIR[11].XIC[12].icell.PDM Iout 0.00117f
C4501 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04031f
C4502 XA.XIR[4].XIC[13].icell.SM Vbias 0.00701f
C4503 XA.XIR[3].XIC[6].icell.PDM Vbias 0.04261f
C4504 XA.XIR[14].XIC[3].icell.Ien Vbias 0.21098f
C4505 XA.XIR[3].XIC[11].icell.Ien VPWR 0.1903f
C4506 XA.XIR[8].XIC[8].icell.PDM Vbias 0.04261f
C4507 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00584f
C4508 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10] 0.00341f
C4509 XThC.Tn[9] XThR.Tn[14] 0.28739f
C4510 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4511 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.15202f
C4512 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02762f
C4513 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00584f
C4514 XA.XIR[2].XIC[12].icell.PDM Vbias 0.04261f
C4515 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14] 0.00341f
C4516 XA.XIR[3].XIC[7].icell.Ien Iout 0.06417f
C4517 XA.XIR[1].XIC[5].icell.PDM Iout 0.00117f
C4518 XA.XIR[13].XIC[5].icell.Ien Vbias 0.21098f
C4519 XA.XIR[14].XIC[13].icell.PDM Iout 0.00117f
C4520 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[6].icell.Ien 0.00214f
C4521 XA.XIR[8].XIC[7].icell.SM Vbias 0.00701f
C4522 XA.XIR[2].XIC[4].icell.Ien VPWR 0.1903f
C4523 XA.XIR[14].XIC[14].icell.SM VPWR 0.00207f
C4524 XA.XIR[7].XIC[4].icell.SM VPWR 0.00158f
C4525 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PUM 0.00465f
C4526 XThR.Tn[1] a_n1049_7787# 0.26879f
C4527 XA.XIR[12].XIC[7].icell.PUM Vbias 0.0031f
C4528 XA.XIR[4].XIC[5].icell.PDM Iout 0.00117f
C4529 XThC.XTB6.A XThC.Tn[1] 0.00411f
C4530 XA.XIR[1].XIC[6].icell.Ien VPWR 0.1903f
C4531 XA.XIR[5].XIC[13].icell.SM Iout 0.00388f
C4532 XA.XIR[14].XIC[10].icell.PUM VPWR 0.00937f
C4533 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00214f
C4534 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C4535 XA.XIR[10].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4536 XA.XIR[11].XIC[8].icell.Ien Vbias 0.21098f
C4537 a_5155_9615# XThC.Tn[3] 0.00508f
C4538 XA.XIR[3].XIC[13].icell.PDM Iout 0.00117f
C4539 XA.XIR[4].XIC_dummy_right.icell.SM VPWR 0.00123f
C4540 XA.XIR[1].XIC[2].icell.Ien Iout 0.06417f
C4541 XA.XIR[8].XIC_15.icell.PDM Iout 0.00133f
C4542 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C4543 XA.XIR[8].XIC[14].icell.Ien VPWR 0.19036f
C4544 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C4545 XThR.Tn[7] XA.XIR[8].XIC[1].icell.SM 0.00121f
C4546 XThR.Tn[6] XA.XIR[7].XIC[12].icell.SM 0.00121f
C4547 XA.XIR[13].XIC_15.icell.SM Vbias 0.00701f
C4548 XThC.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00109f
C4549 XA.XIR[8].XIC[10].icell.Ien Iout 0.06417f
C4550 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38912f
C4551 XThR.Tn[8] XA.XIR[9].XIC[10].icell.Ien 0.00338f
C4552 XA.XIR[0].XIC[9].icell.SM Vbias 0.00716f
C4553 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PUM 0.00465f
C4554 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04675f
C4555 XThC.Tn[5] XThR.Tn[6] 0.28739f
C4556 XA.XIR[12].XIC[8].icell.SM Iout 0.00388f
C4557 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.SM 0.00168f
C4558 XThR.XTB7.B VPWR 1.67379f
C4559 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00214f
C4560 XThR.Tn[1] XA.XIR[1].XIC[14].icell.PDM 0.00341f
C4561 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C4562 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C4563 XThR.Tn[10] XA.XIR[11].XIC[2].icell.SM 0.00121f
C4564 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.04036f
C4565 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PUM 0.00465f
C4566 XA.XIR[2].XIC[12].icell.Ien Vbias 0.21098f
C4567 XThC.Tn[7] XThR.Tn[11] 0.28739f
C4568 XA.XIR[7].XIC[12].icell.SM Vbias 0.00701f
C4569 XThR.Tn[1] XA.XIR[2].XIC[3].icell.Ien 0.00338f
C4570 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.SM 0.00168f
C4571 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04031f
C4572 XA.XIR[14].XIC[11].icell.Ien VPWR 0.19084f
C4573 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PUM 0.00465f
C4574 XA.XIR[1].XIC[14].icell.Ien Vbias 0.21104f
C4575 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.15202f
C4576 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.15202f
C4577 XA.XIR[0].XIC[12].icell.Ien Iout 0.06389f
C4578 XThC.Tn[5] Vbias 2.31635f
C4579 XA.XIR[5].XIC[2].icell.PDM VPWR 0.00799f
C4580 XThR.Tn[2] XA.XIR[2].XIC[11].icell.PDM 0.00341f
C4581 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.SM 0.0039f
C4582 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02762f
C4583 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Ien 0.00232f
C4584 XA.XIR[6].XIC[1].icell.Ien VPWR 0.1903f
C4585 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04031f
C4586 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C4587 XThR.Tn[13] XA.XIR[14].XIC[7].icell.Ien 0.00338f
C4588 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PDM 0.00172f
C4589 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.03425f
C4590 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00584f
C4591 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.15202f
C4592 XThC.XTB5.Y a_7651_9569# 0.00418f
C4593 XA.XIR[12].XIC[1].icell.PDM VPWR 0.00799f
C4594 XA.XIR[12].XIC[1].icell.Ien Vbias 0.21098f
C4595 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C4596 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.SM 0.00168f
C4597 XA.XIR[7].XIC_15.icell.Ien Iout 0.0642f
C4598 XThC.Tn[11] XThR.Tn[13] 0.28739f
C4599 XThR.Tn[0] XA.XIR[1].XIC[10].icell.Ien 0.00338f
C4600 XThR.Tn[2] VPWR 6.62952f
C4601 XA.XIR[5].XIC[0].icell.Ien Iout 0.06411f
C4602 XThC.Tn[1] XThR.Tn[1] 0.28739f
C4603 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C4604 XThR.Tn[13] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00107f
C4605 XA.XIR[11].XIC[7].icell.PDM VPWR 0.00799f
C4606 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C4607 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.SM 0.00168f
C4608 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PUM 0.00465f
C4609 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.0353f
C4610 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.15202f
C4611 XThR.XTB7.Y a_n997_3979# 0.00477f
C4612 XA.XIR[7].XIC[12].icell.PDM Vbias 0.04261f
C4613 XA.XIR[5].XIC[2].icell.Ien Vbias 0.21098f
C4614 XThC.Tn[14] Iout 0.84284f
C4615 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C4616 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00214f
C4617 XThC.Tn[14] XThR.Tn[9] 0.28745f
C4618 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PUM 0.00465f
C4619 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02762f
C4620 XThC.Tn[1] XThR.Tn[12] 0.28739f
C4621 XThC.Tn[10] XThR.Tn[8] 0.28739f
C4622 XThR.Tn[5] XA.XIR[6].XIC[12].icell.Ien 0.00338f
C4623 XA.XIR[4].XIC[5].icell.PUM Vbias 0.0031f
C4624 XA.XIR[15].XIC[10].icell.PDM Vbias 0.04261f
C4625 XA.XIR[3].XIC[1].icell.SM VPWR 0.00158f
C4626 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PUM 0.00442f
C4627 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C4628 XA.XIR[6].XIC[6].icell.Ien VPWR 0.1903f
C4629 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_15.icell.SM 0.0039f
C4630 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.SM 0.0039f
C4631 XA.XIR[15].XIC[7].icell.SM VPWR 0.00158f
C4632 XA.XIR[5].XIC[9].icell.PUM VPWR 0.00937f
C4633 XA.XIR[6].XIC[2].icell.Ien Iout 0.06417f
C4634 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C4635 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.SM 0.0039f
C4636 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.SM 0.0039f
C4637 XThC.XTBN.Y a_7651_9569# 0.23021f
C4638 XThC.Tn[5] XThR.Tn[4] 0.28739f
C4639 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C4640 XA.XIR[15].XIC[3].icell.SM Iout 0.00388f
C4641 XA.XIR[4].XIC[10].icell.SM VPWR 0.00158f
C4642 XA.XIR[9].XIC[8].icell.PDM Vbias 0.04261f
C4643 a_10051_9569# Vbias 0.00678f
C4644 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C4645 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00584f
C4646 XA.XIR[0].XIC[0].icell.PDM Vbias 0.04227f
C4647 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00214f
C4648 XThC.XTB4.Y XThC.Tn[3] 0.18952f
C4649 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PDM 0.00555f
C4650 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.11857f
C4651 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.15202f
C4652 XA.XIR[4].XIC[6].icell.SM Iout 0.00388f
C4653 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.15202f
C4654 XA.XIR[11].XIC[11].icell.PDM Iout 0.00117f
C4655 XA.XIR[2].XIC[3].icell.PDM VPWR 0.00799f
C4656 XThC.Tn[0] XThR.Tn[10] 0.28736f
C4657 XA.XIR[13].XIC[2].icell.Ien VPWR 0.1903f
C4658 XA.XIR[8].XIC[4].icell.SM VPWR 0.00158f
C4659 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00214f
C4660 XA.XIR[9].XIC[8].icell.PUM Vbias 0.0031f
C4661 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C4662 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.03425f
C4663 XThR.Tn[13] XThR.Tn[14] 0.1554f
C4664 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00584f
C4665 XA.XIR[12].XIC[4].icell.PUM VPWR 0.00937f
C4666 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00214f
C4667 XA.XIR[14].XIC[12].icell.PDM Iout 0.00117f
C4668 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.SM 0.00168f
C4669 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.SM 0.0039f
C4670 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04031f
C4671 XA.XIR[11].XIC[5].icell.Ien VPWR 0.1903f
C4672 XA.XIR[3].XIC[9].icell.SM Vbias 0.00701f
C4673 XA.XIR[9].XIC_15.icell.PDM Iout 0.00133f
C4674 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9] 0.00341f
C4675 XA.XIR[1].XIC[13].icell.PDM Vbias 0.04261f
C4676 XThR.Tn[4] XA.XIR[5].XIC[2].icell.Ien 0.00338f
C4677 XA.XIR[9].XIC[13].icell.SM VPWR 0.00158f
C4678 XA.XIR[7].XIC[0].icell.SM Iout 0.00388f
C4679 XA.XIR[6].XIC[14].icell.Ien Vbias 0.21098f
C4680 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.15202f
C4681 XA.XIR[10].XIC[7].icell.Ien VPWR 0.1903f
C4682 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.SM 0.00168f
C4683 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.SM 0.0039f
C4684 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11] 0.00341f
C4685 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C4686 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C4687 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C4688 XThR.Tn[3] XA.XIR[4].XIC[2].icell.Ien 0.00338f
C4689 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C4690 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00214f
C4691 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PUM 0.00465f
C4692 XA.XIR[4].XIC[13].icell.PDM Vbias 0.04261f
C4693 XA.XIR[2].XIC[2].icell.SM Vbias 0.00701f
C4694 XA.XIR[9].XIC[9].icell.SM Iout 0.00388f
C4695 XA.XIR[7].XIC[4].icell.PUM Vbias 0.0031f
C4696 XA.XIR[10].XIC[3].icell.Ien Iout 0.06417f
C4697 XThR.XTB7.Y a_n997_2891# 0.00474f
C4698 XThC.XTB2.Y a_4067_9615# 0.02133f
C4699 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.SM 0.0039f
C4700 XThR.Tn[9] XA.XIR[10].XIC[3].icell.Ien 0.00338f
C4701 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C4702 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.SM 0.00168f
C4703 XA.XIR[0].XIC[6].icell.SM VPWR 0.00158f
C4704 XA.XIR[12].XIC[13].icell.SM Iout 0.00388f
C4705 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C4706 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02762f
C4707 XA.XIR[1].XIC[4].icell.SM Vbias 0.00704f
C4708 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00214f
C4709 XA.XIR[13].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4710 XA.XIR[0].XIC[2].icell.SM Iout 0.00367f
C4711 XA.XIR[14].XIC[8].icell.Ien Vbias 0.21098f
C4712 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04031f
C4713 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C4714 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C4715 XThR.XTBN.Y VPWR 4.54127f
C4716 XA.XIR[11].XIC_15.icell.SM VPWR 0.00275f
C4717 XA.XIR[3].XIC[12].icell.Ien Iout 0.06417f
C4718 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PUM 0.00465f
C4719 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.04036f
C4720 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8] 0.00341f
C4721 XA.XIR[2].XIC[9].icell.Ien VPWR 0.1903f
C4722 XA.XIR[7].XIC[9].icell.SM VPWR 0.00158f
C4723 XA.XIR[8].XIC[12].icell.SM Vbias 0.00701f
C4724 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.SM 0.0039f
C4725 XA.XIR[2].XIC[5].icell.Ien Iout 0.06417f
C4726 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C4727 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04031f
C4728 XA.XIR[7].XIC[5].icell.SM Iout 0.00388f
C4729 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PUM 0.00465f
C4730 XA.XIR[1].XIC[11].icell.Ien VPWR 0.1903f
C4731 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C4732 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.15202f
C4733 XA.XIR[1].XIC[7].icell.Ien Iout 0.06417f
C4734 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.03425f
C4735 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C4736 XA.XIR[10].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4737 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02762f
C4738 XThR.Tn[7] XA.XIR[8].XIC[6].icell.SM 0.00121f
C4739 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PUM 0.00465f
C4740 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C4741 XThC.Tn[7] XThR.Tn[14] 0.28739f
C4742 XThR.XTB2.Y a_n1049_6699# 0.00851f
C4743 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.SM 0.0039f
C4744 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.SM 0.00168f
C4745 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.15202f
C4746 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02762f
C4747 XThR.Tn[11] XA.XIR[12].XIC[4].icell.Ien 0.00338f
C4748 a_10051_9569# XThC.Tn[13] 0.19413f
C4749 XThR.Tn[5] XA.XIR[6].XIC[2].icell.SM 0.00121f
C4750 XA.XIR[8].XIC_15.icell.Ien Iout 0.0642f
C4751 XThR.Tn[8] XA.XIR[9].XIC_15.icell.Ien 0.00117f
C4752 XThR.XTB4.Y VPWR 0.92827f
C4753 XA.XIR[0].XIC[14].icell.SM Vbias 0.00716f
C4754 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C4755 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04052f
C4756 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C4757 XA.XIR[11].XIC[1].icell.PUM VPWR 0.00937f
C4758 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00214f
C4759 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.SM 0.0039f
C4760 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.15202f
C4761 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04031f
C4762 XThR.Tn[4] XA.XIR[4].XIC[13].icell.PDM 0.00341f
C4763 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PUM 0.00465f
C4764 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PUM 0.00465f
C4765 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C4766 XThR.Tn[10] VPWR 7.53208f
C4767 XA.XIR[7].XIC[3].icell.PDM VPWR 0.00799f
C4768 XThR.Tn[3] XA.XIR[3].XIC[14].icell.PDM 0.00341f
C4769 XThR.Tn[10] XA.XIR[11].XIC[7].icell.SM 0.00121f
C4770 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01745f
C4771 XThR.Tn[1] XA.XIR[2].XIC[8].icell.Ien 0.00338f
C4772 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.SM 0.0039f
C4773 XA.XIR[6].XIC[10].icell.PDM VPWR 0.00799f
C4774 XA.XIR[15].XIC[2].icell.PUM Vbias 0.0031f
C4775 XA.XIR[15].XIC[1].icell.PDM VPWR 0.0114f
C4776 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.SM 0.0039f
C4777 XThC.Tn[9] VPWR 6.83084f
C4778 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C4779 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00214f
C4780 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00214f
C4781 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02762f
C4782 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.15202f
C4783 XThR.XTB5.A a_n1335_4229# 0.01243f
C4784 XA.XIR[14].XIC[7].icell.PDM VPWR 0.00799f
C4785 XA.XIR[11].XIC[3].icell.PDM Vbias 0.04261f
C4786 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PUM 0.00465f
C4787 XA.XIR[5].XIC[5].icell.PDM Iout 0.00117f
C4788 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PUM 0.00465f
C4789 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02762f
C4790 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.SM 0.00168f
C4791 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00584f
C4792 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00584f
C4793 XA.XIR[10].XIC[7].icell.PDM Vbias 0.04261f
C4794 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C4795 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.SM 0.0039f
C4796 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00584f
C4797 XThR.Tn[0] XA.XIR[1].XIC_15.icell.Ien 0.00117f
C4798 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C4799 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C4800 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C4801 XA.XIR[9].XIC[5].icell.PUM VPWR 0.00937f
C4802 XA.XIR[12].XIC[4].icell.PDM Iout 0.00117f
C4803 XA.XIR[6].XIC[4].icell.SM Vbias 0.00701f
C4804 XA.XIR[12].XIC[11].icell.SM Iout 0.00388f
C4805 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C4806 data[5] data[6] 0.01513f
C4807 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C4808 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C4809 XA.XIR[15].XIC[7].icell.PUM Vbias 0.0031f
C4810 XA.XIR[11].XIC[10].icell.PDM Iout 0.00117f
C4811 XA.XIR[5].XIC[7].icell.Ien Vbias 0.21098f
C4812 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.SM 0.0039f
C4813 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00584f
C4814 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.SM 0.00168f
C4815 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02762f
C4816 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C4817 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.03425f
C4818 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00214f
C4819 XA.XIR[4].XIC[10].icell.PUM Vbias 0.0031f
C4820 XA.XIR[3].XIC[6].icell.SM VPWR 0.00158f
C4821 XA.XIR[1].XIC[4].icell.PDM VPWR 0.00799f
C4822 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C4823 XA.XIR[8].XIC[0].icell.SM Iout 0.00388f
C4824 XA.XIR[0].XIC[1].icell.PUM Vbias 0.0031f
C4825 XThR.Tn[8] XA.XIR[9].XIC[0].icell.SM 0.00121f
C4826 XA.XIR[14].XIC[11].icell.PDM Iout 0.00117f
C4827 XA.XIR[6].XIC[11].icell.Ien VPWR 0.1903f
C4828 XThC.Tn[0] XThR.Tn[13] 0.28746f
C4829 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C4830 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C4831 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.03425f
C4832 XA.XIR[3].XIC[2].icell.SM Iout 0.00388f
C4833 a_4067_9615# XThC.Tn[4] 0.00141f
C4834 XA.XIR[6].XIC[7].icell.Ien Iout 0.06417f
C4835 XA.XIR[8].XIC[4].icell.PUM Vbias 0.0031f
C4836 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[3].icell.SM 0.0039f
C4837 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7] 0.00341f
C4838 XA.XIR[4].XIC[4].icell.PDM VPWR 0.00799f
C4839 XA.XIR[5].XIC[14].icell.PUM VPWR 0.00937f
C4840 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04037f
C4841 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C4842 XA.XIR[15].XIC[8].icell.SM Iout 0.00388f
C4843 XA.XIR[12].XIC[2].icell.Ien Vbias 0.21098f
C4844 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C4845 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C4846 XThC.Tn[3] Iout 0.8384f
C4847 XA.XIR[1].XIC[1].icell.SM VPWR 0.00158f
C4848 XThC.Tn[3] XThR.Tn[9] 0.28739f
C4849 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C4850 XA.XIR[3].XIC[12].icell.PDM VPWR 0.00799f
C4851 XA.XIR[8].XIC[14].icell.PDM VPWR 0.00809f
C4852 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00214f
C4853 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13] 0.00341f
C4854 XThC.Tn[12] data[3] 0.00161f
C4855 XA.XIR[14].XIC[5].icell.Ien VPWR 0.19084f
C4856 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C4857 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.03589f
C4858 XA.XIR[0].XIC_15.icell.PDM Vbias 0.04422f
C4859 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.15202f
C4860 XThC.XTB7.Y Vbias 0.01727f
C4861 XA.XIR[11].XIC[3].icell.SM Vbias 0.00701f
C4862 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C4863 XA.XIR[4].XIC[11].icell.SM Iout 0.00388f
C4864 XThC.XTBN.A a_10051_9569# 0.00199f
C4865 XA.XIR[3].XIC[0].icell.PDM Iout 0.00117f
C4866 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02762f
C4867 XA.XIR[8].XIC[2].icell.PDM Iout 0.00117f
C4868 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04031f
C4869 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04031f
C4870 XA.XIR[13].XIC[7].icell.Ien VPWR 0.1903f
C4871 XA.XIR[9].XIC[13].icell.PUM Vbias 0.0031f
C4872 XThR.XTB6.A XThR.XTBN.A 0.0512f
C4873 XA.XIR[8].XIC[9].icell.SM VPWR 0.00158f
C4874 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C4875 XA.XIR[10].XIC[5].icell.SM Vbias 0.00701f
C4876 XA.XIR[2].XIC[6].icell.PDM Iout 0.00117f
C4877 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4878 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C4879 XA.XIR[13].XIC[3].icell.Ien Iout 0.06417f
C4880 XThR.XTB7.Y a_n997_1579# 0.013f
C4881 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02762f
C4882 XA.XIR[12].XIC[9].icell.PUM VPWR 0.00937f
C4883 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.SM 0.00168f
C4884 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00584f
C4885 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00584f
C4886 XA.XIR[8].XIC[5].icell.SM Iout 0.00388f
C4887 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.PDM 0.00591f
C4888 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02762f
C4889 XThR.Tn[8] XA.XIR[9].XIC[5].icell.SM 0.00121f
C4890 XA.XIR[0].XIC[6].icell.PUM Vbias 0.0031f
C4891 XThR.Tn[0] XA.XIR[0].XIC[3].icell.PDM 0.00341f
C4892 a_n997_1803# VPWR 0.01991f
C4893 XA.XIR[3].XIC[14].icell.SM Vbias 0.00701f
C4894 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.SM 0.0039f
C4895 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02762f
C4896 XThR.Tn[4] XA.XIR[5].XIC[7].icell.Ien 0.00338f
C4897 XA.XIR[14].XIC_15.icell.SM VPWR 0.00275f
C4898 XThR.Tn[0] XA.XIR[1].XIC[0].icell.SM 0.00121f
C4899 XThR.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.00341f
C4900 XA.XIR[11].XIC[6].icell.Ien Iout 0.06417f
C4901 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.03023f
C4902 XThR.Tn[11] XA.XIR[12].XIC[12].icell.SM 0.00121f
C4903 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Iout 0.00347f
C4904 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01432f
C4905 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.04036f
C4906 XThR.Tn[3] XA.XIR[4].XIC[7].icell.Ien 0.00338f
C4907 XThC.XTB7.A XThC.Tn[10] 0.00406f
C4908 XA.XIR[9].XIC[14].icell.SM Iout 0.00388f
C4909 XA.XIR[7].XIC[9].icell.PUM Vbias 0.0031f
C4910 XA.XIR[2].XIC[7].icell.SM Vbias 0.00701f
C4911 XA.XIR[0].XIC[11].icell.SM VPWR 0.00158f
C4912 XA.XIR[10].XIC[8].icell.Ien Iout 0.06417f
C4913 XThC.XTB5.Y a_5949_9615# 0.0093f
C4914 XThR.Tn[9] XA.XIR[10].XIC[8].icell.Ien 0.00338f
C4915 XThC.XTB3.Y XThC.Tn[5] 0.00384f
C4916 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.SM 0.0039f
C4917 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PUM 0.00465f
C4918 XA.XIR[8].XIC[0].icell.PUM VPWR 0.00937f
C4919 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5] 0.00341f
C4920 XThC.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.00109f
C4921 XThC.XTB7.A a_4861_9615# 0.02294f
C4922 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00584f
C4923 XA.XIR[1].XIC[9].icell.SM Vbias 0.00704f
C4924 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02762f
C4925 XA.XIR[0].XIC[7].icell.SM Iout 0.00367f
C4926 XThC.Tn[3] XThC.Tn[4] 0.49877f
C4927 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PUM 0.00465f
C4928 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.SM 0.0039f
C4929 XA.XIR[13].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4930 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.04036f
C4931 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02762f
C4932 XThR.Tn[13] XA.XIR[14].XIC[2].icell.SM 0.00121f
C4933 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PUM 0.00465f
C4934 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.SM 0.0039f
C4935 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PDM 0.00172f
C4936 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[11].icell.Ien 0.00214f
C4937 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.SM 0.00168f
C4938 XA.XIR[7].XIC[14].icell.SM VPWR 0.00207f
C4939 XA.XIR[2].XIC[14].icell.Ien VPWR 0.19036f
C4940 XA.XIR[12].XIC[9].icell.SM Iout 0.00388f
C4941 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C4942 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C4943 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02762f
C4944 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6] 0.00341f
C4945 XA.XIR[2].XIC[10].icell.Ien Iout 0.06417f
C4946 XA.XIR[7].XIC[10].icell.SM Iout 0.00388f
C4947 XThR.Tn[0] XA.XIR[1].XIC[5].icell.SM 0.00121f
C4948 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.15202f
C4949 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00214f
C4950 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C4951 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C4952 XA.XIR[14].XIC[0].icell.Ien VPWR 0.19084f
C4953 XThR.Tn[12] XA.XIR[13].XIC[6].icell.Ien 0.00338f
C4954 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.SM 0.0039f
C4955 XA.XIR[4].XIC[2].icell.PUM VPWR 0.00937f
C4956 XThR.Tn[0] Vbias 3.75791f
C4957 XA.XIR[1].XIC[12].icell.Ien Iout 0.06417f
C4958 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.SM 0.0039f
C4959 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00584f
C4960 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C4961 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PUM 0.00186f
C4962 XThR.Tn[7] XA.XIR[8].XIC[11].icell.SM 0.00121f
C4963 XThR.Tn[13] VPWR 7.61336f
C4964 XThC.XTBN.Y a_5949_9615# 0.0768f
C4965 XThC.Tn[11] XThR.Tn[7] 0.28739f
C4966 XA.XIR[10].XIC[1].icell.PUM Vbias 0.0031f
C4967 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.03425f
C4968 XThR.Tn[11] XA.XIR[12].XIC[9].icell.Ien 0.00338f
C4969 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C4970 XThC.XTB7.B XThC.Tn[9] 0.09571f
C4971 XThR.Tn[5] XA.XIR[6].XIC[7].icell.SM 0.00121f
C4972 XA.XIR[6].XIC[6].icell.PDM Vbias 0.04261f
C4973 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Iout 0.00347f
C4974 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C4975 XThR.XTB2.Y XThR.Tn[8] 0.00167f
C4976 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PUM 0.00186f
C4977 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C4978 XThC.XTB7.Y XThC.Tn[13] 0.11626f
C4979 XA.XIR[6].XIC[1].icell.SM VPWR 0.00158f
C4980 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.SM 0.00168f
C4981 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00214f
C4982 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.15202f
C4983 XA.XIR[14].XIC[3].icell.PDM Vbias 0.04261f
C4984 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.SM 0.00168f
C4985 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C4986 XA.XIR[5].XIC[13].icell.PDM Vbias 0.04261f
C4987 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PUM 0.00465f
C4988 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.15202f
C4989 XA.XIR[15].XIC[4].icell.PUM VPWR 0.00937f
C4990 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02762f
C4991 XA.XIR[11].XIC[0].icell.SM Iout 0.00388f
C4992 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C4993 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PUM 0.00465f
C4994 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.03425f
C4995 XA.XIR[5].XIC[4].icell.Ien VPWR 0.1903f
C4996 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02762f
C4997 XThC.XTB5.A XThC.XTBN.Y 0.00282f
C4998 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00214f
C4999 XA.XIR[13].XIC[7].icell.PDM Vbias 0.04261f
C5000 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C5001 XA.XIR[7].XIC[6].icell.PDM Iout 0.00117f
C5002 XThR.Tn[1] XA.XIR[2].XIC[13].icell.Ien 0.00338f
C5003 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PUM 0.00465f
C5004 XThR.Tn[3] a_n1049_6699# 0.27008f
C5005 XA.XIR[4].XIC[7].icell.PUM VPWR 0.00937f
C5006 XA.XIR[15].XIC[4].icell.PDM Iout 0.00117f
C5007 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C5008 XA.XIR[6].XIC[13].icell.PDM Iout 0.00117f
C5009 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C5010 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PUM 0.00471f
C5011 XA.XIR[9].XIC[3].icell.Ien Vbias 0.21098f
C5012 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00214f
C5013 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02762f
C5014 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.SM 0.0039f
C5015 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.SM 0.00168f
C5016 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PUM 0.00465f
C5017 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C5018 XA.XIR[14].XIC[10].icell.PDM Iout 0.00117f
C5019 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C5020 XA.XIR[15].XIC[13].icell.SM Iout 0.00388f
C5021 XA.XIR[9].XIC[14].icell.PDM VPWR 0.00809f
C5022 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00584f
C5023 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C5024 XThR.Tn[11] XA.XIR[12].XIC[10].icell.SM 0.00121f
C5025 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00214f
C5026 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00214f
C5027 XA.XIR[7].XIC[1].icell.PUM VPWR 0.00937f
C5028 XA.XIR[0].XIC[6].icell.PDM VPWR 0.0078f
C5029 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C5030 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C5031 XThC.Tn[10] XThR.Tn[3] 0.28739f
C5032 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PDM 0.0059f
C5033 XA.XIR[3].XIC[6].icell.PUM Vbias 0.0031f
C5034 XA.XIR[9].XIC[2].icell.PDM Iout 0.00117f
C5035 XA.XIR[1].XIC[0].icell.PDM Vbias 0.04207f
C5036 XThC.Tn[0] XA.XIR[6].XIC_dummy_left.icell.Iout 0.00109f
C5037 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9] 0.00341f
C5038 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11154f
C5039 XA.XIR[6].XIC[9].icell.SM Vbias 0.00701f
C5040 XA.XIR[9].XIC[10].icell.PUM VPWR 0.00937f
C5041 XThR.Tn[12] XA.XIR[13].XIC[0].icell.SM 0.00127f
C5042 XA.XIR[10].XIC[2].icell.SM VPWR 0.00158f
C5043 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00584f
C5044 XThC.Tn[7] VPWR 6.29093f
C5045 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.SM 0.0039f
C5046 XA.XIR[4].XIC[0].icell.PDM Vbias 0.04207f
C5047 XA.XIR[12].XIC[13].icell.Ien Iout 0.06417f
C5048 XA.XIR[5].XIC[12].icell.Ien Vbias 0.21098f
C5049 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C5050 XA.XIR[0].XIC[3].icell.PUM VPWR 0.00877f
C5051 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.SM 0.00168f
C5052 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04031f
C5053 XThC.XTB6.A Vbias 0.00648f
C5054 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.04036f
C5055 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.SM 0.0039f
C5056 XA.XIR[3].XIC[8].icell.PDM Vbias 0.04261f
C5057 XA.XIR[4].XIC_15.icell.PUM Vbias 0.0031f
C5058 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04031f
C5059 XA.XIR[8].XIC[10].icell.PDM Vbias 0.04261f
C5060 XA.XIR[14].XIC[3].icell.SM Vbias 0.00701f
C5061 XA.XIR[3].XIC[11].icell.SM VPWR 0.00158f
C5062 XThC.Tn[13] XThR.Tn[0] 0.28789f
C5063 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10] 0.00341f
C5064 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C5065 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C5066 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14] 0.00341f
C5067 XA.XIR[3].XIC[7].icell.SM Iout 0.00388f
C5068 XA.XIR[2].XIC[14].icell.PDM Vbias 0.04261f
C5069 XA.XIR[1].XIC[7].icell.PDM Iout 0.00117f
C5070 XA.XIR[13].XIC[5].icell.SM Vbias 0.00701f
C5071 XA.XIR[8].XIC[9].icell.PUM Vbias 0.0031f
C5072 XA.XIR[6].XIC[12].icell.Ien Iout 0.06417f
C5073 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5074 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5075 XA.XIR[7].XIC[6].icell.PUM VPWR 0.00937f
C5076 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02762f
C5077 XA.XIR[2].XIC[4].icell.SM VPWR 0.00158f
C5078 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C5079 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.03425f
C5080 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.SM 0.0039f
C5081 XA.XIR[12].XIC[7].icell.Ien Vbias 0.21098f
C5082 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C5083 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.PDM 0.00591f
C5084 XA.XIR[1].XIC[6].icell.SM VPWR 0.00158f
C5085 a_5949_10571# VPWR 0.00653f
C5086 XA.XIR[4].XIC[7].icell.PDM Iout 0.00117f
C5087 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.SM 0.0039f
C5088 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02827f
C5089 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00584f
C5090 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PUM 0.00465f
C5091 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C5092 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01451f
C5093 XA.XIR[11].XIC[8].icell.SM Vbias 0.00701f
C5094 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02762f
C5095 XA.XIR[1].XIC[2].icell.SM Iout 0.00388f
C5096 XA.XIR[3].XIC_15.icell.PDM Iout 0.00133f
C5097 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38997f
C5098 XThC.XTB4.Y data[2] 0.0086f
C5099 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00214f
C5100 XA.XIR[14].XIC[6].icell.Ien Iout 0.06417f
C5101 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00584f
C5102 XA.XIR[8].XIC[14].icell.SM VPWR 0.00207f
C5103 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C5104 XThC.XTB6.A a_7331_10587# 0.00304f
C5105 XA.XIR[12].XIC[14].icell.SM Iout 0.00388f
C5106 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04031f
C5107 XA.XIR[13].XIC[8].icell.Ien Iout 0.06417f
C5108 XThR.XTB7.A a_n1319_5317# 0.0017f
C5109 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00584f
C5110 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.15202f
C5111 XA.XIR[8].XIC[10].icell.SM Iout 0.00388f
C5112 XThR.Tn[8] XA.XIR[9].XIC[10].icell.SM 0.00121f
C5113 XA.XIR[0].XIC[11].icell.PUM Vbias 0.0031f
C5114 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.03425f
C5115 XThR.Tn[2] XA.XIR[3].XIC[5].icell.Ien 0.00338f
C5116 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02762f
C5117 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C5118 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C5119 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00214f
C5120 XA.XIR[5].XIC[0].icell.PUM VPWR 0.00937f
C5121 XThR.Tn[4] XA.XIR[4].XIC[0].icell.PDM 0.00346f
C5122 XA.XIR[6].XIC_dummy_left.icell.Ien Vbias 0.00329f
C5123 XThR.Tn[4] XA.XIR[5].XIC[12].icell.Ien 0.00338f
C5124 XThR.XTB3.Y a_n997_3979# 0.00604f
C5125 XThR.XTBN.A XThR.Tn[12] 0.22096f
C5126 XA.XIR[14].XIC_dummy_left.icell.SM VPWR 0.00269f
C5127 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C5128 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PUM 0.00465f
C5129 XThR.Tn[3] XA.XIR[4].XIC[12].icell.Ien 0.00338f
C5130 XThR.Tn[3] XA.XIR[3].XIC[1].icell.PDM 0.00341f
C5131 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PDM 0.00172f
C5132 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.03425f
C5133 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PUM 0.00465f
C5134 XA.XIR[7].XIC[14].icell.PUM Vbias 0.0031f
C5135 XA.XIR[2].XIC[12].icell.SM Vbias 0.00701f
C5136 a_3773_9615# VPWR 0.70508f
C5137 XThR.Tn[1] XA.XIR[2].XIC[3].icell.SM 0.00121f
C5138 XThR.Tn[11] XA.XIR[12].XIC[14].icell.Ien 0.00338f
C5139 XThR.XTB2.Y a_n997_3755# 0.06476f
C5140 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C5141 XA.XIR[1].XIC[0].icell.Ien Vbias 0.20957f
C5142 XThC.Tn[12] XThR.Tn[2] 0.28739f
C5143 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04031f
C5144 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PUM 0.00465f
C5145 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.SM 0.0039f
C5146 XA.XIR[15].XIC[11].icell.SM Iout 0.00388f
C5147 XA.XIR[1].XIC[14].icell.SM Vbias 0.00704f
C5148 XA.XIR[0].XIC[12].icell.SM Iout 0.00367f
C5149 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C5150 XA.XIR[5].XIC[4].icell.PDM VPWR 0.00799f
C5151 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C5152 XA.XIR[4].XIC[0].icell.Ien Vbias 0.20951f
C5153 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C5154 XThR.Tn[2] XA.XIR[2].XIC[13].icell.PDM 0.00341f
C5155 XThR.XTBN.Y a_n1049_8581# 0.0607f
C5156 XThR.Tn[1] Vbias 3.74871f
C5157 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C5158 XThC.XTB4.Y a_5155_9615# 0.01546f
C5159 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C5160 XThR.Tn[13] XA.XIR[14].XIC[7].icell.SM 0.00121f
C5161 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Iout 0.00347f
C5162 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04052f
C5163 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11115f
C5164 XA.XIR[0].XIC_15.icell.SM Vbias 0.00716f
C5165 XA.XIR[13].XIC[1].icell.PUM Vbias 0.0031f
C5166 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Ien 0.00232f
C5167 XThC.XTB5.Y a_8739_9569# 0.00424f
C5168 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C5169 XA.XIR[12].XIC[3].icell.PDM VPWR 0.00799f
C5170 XThR.Tn[12] Vbias 3.74784f
C5171 XA.XIR[2].XIC_15.icell.Ien Iout 0.0642f
C5172 XA.XIR[12].XIC[11].icell.Ien Iout 0.06417f
C5173 XThR.Tn[0] XA.XIR[1].XIC[10].icell.SM 0.00121f
C5174 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C5175 XThR.XTB2.Y a_n1049_5611# 0.00844f
C5176 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.PUM 0.00121f
C5177 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02762f
C5178 XA.XIR[11].XIC[9].icell.PDM VPWR 0.00799f
C5179 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C5180 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.03425f
C5181 XA.XIR[14].XIC[0].icell.SM Iout 0.00388f
C5182 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PUM 0.00465f
C5183 XA.XIR[15].XIC[2].icell.Ien Vbias 0.17899f
C5184 XA.XIR[7].XIC[14].icell.PDM Vbias 0.04261f
C5185 XA.XIR[5].XIC[2].icell.SM Vbias 0.00701f
C5186 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.SM 0.00168f
C5187 XThC.Tn[8] XThR.Tn[6] 0.28739f
C5188 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.03425f
C5189 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.SM 0.0039f
C5190 XThR.Tn[5] XA.XIR[6].XIC[12].icell.SM 0.00121f
C5191 XA.XIR[4].XIC[5].icell.Ien Vbias 0.21098f
C5192 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.SM 0.00168f
C5193 XA.XIR[10].XIC[1].icell.PDM Iout 0.00117f
C5194 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04031f
C5195 XA.XIR[3].XIC[3].icell.PUM VPWR 0.00937f
C5196 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.0355f
C5197 XA.XIR[6].XIC[6].icell.SM VPWR 0.00158f
C5198 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C5199 XThR.XTB3.Y XThR.Tn[7] 0.00819f
C5200 XThR.XTB3.Y a_n997_2891# 0.07285f
C5201 XThC.Tn[10] XThR.Tn[11] 0.28739f
C5202 XA.XIR[15].XIC[9].icell.PUM VPWR 0.00937f
C5203 XA.XIR[6].XIC[2].icell.SM Iout 0.00388f
C5204 XA.XIR[5].XIC[9].icell.Ien VPWR 0.1903f
C5205 XThC.XTBN.Y a_8739_9569# 0.22804f
C5206 XThC.Tn[0] XThR.Tn[7] 0.2874f
C5207 XThC.Tn[8] Vbias 2.30271f
C5208 XA.XIR[9].XIC[10].icell.PDM Vbias 0.04261f
C5209 XA.XIR[5].XIC[5].icell.Ien Iout 0.06417f
C5210 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.SM 0.0039f
C5211 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.15222f
C5212 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C5213 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C5214 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C5215 XA.XIR[4].XIC[12].icell.PUM VPWR 0.00937f
C5216 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.03425f
C5217 XA.XIR[8].XIC[1].icell.PDM VPWR 0.00799f
C5218 a_n1049_5317# XThR.Tn[6] 0.26047f
C5219 XA.XIR[0].XIC[2].icell.PDM Vbias 0.04282f
C5220 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.15202f
C5221 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00214f
C5222 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.15235f
C5223 XA.XIR[2].XIC[5].icell.PDM VPWR 0.00799f
C5224 XThR.Tn[1] a_n1049_7493# 0.00444f
C5225 XA.XIR[13].XIC[2].icell.SM VPWR 0.00158f
C5226 XA.XIR[9].XIC[8].icell.Ien Vbias 0.21098f
C5227 XThC.XTB7.B XThC.Tn[7] 0.08407f
C5228 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C5229 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C5230 XA.XIR[8].XIC[6].icell.PUM VPWR 0.00937f
C5231 XThR.XTB1.Y bias[2] 0.00266f
C5232 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00584f
C5233 XThC.XTB5.Y XThC.Tn[11] 0.02206f
C5234 XThR.Tn[6] XA.XIR[7].XIC[4].icell.Ien 0.00338f
C5235 XA.XIR[12].XIC[4].icell.Ien VPWR 0.1903f
C5236 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12] 0.00341f
C5237 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C5238 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.SM 0.00168f
C5239 XThR.Tn[5] Iout 1.16233f
C5240 a_8739_9569# XThC.Tn[10] 0.19671f
C5241 XA.XIR[11].XIC[5].icell.SM VPWR 0.00158f
C5242 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00256f
C5243 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C5244 a_n997_3979# VPWR 0.01662f
C5245 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00214f
C5246 XA.XIR[11].XIC[13].icell.SM Vbias 0.00701f
C5247 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C5248 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04031f
C5249 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C5250 XThR.Tn[8] data[4] 0.01643f
C5251 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.SM 0.0039f
C5252 XThR.Tn[11] XA.XIR[12].XIC[12].icell.Ien 0.00338f
C5253 XA.XIR[3].XIC[11].icell.PUM Vbias 0.0031f
C5254 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.03425f
C5255 XA.XIR[1].XIC_15.icell.PDM Vbias 0.04401f
C5256 XThR.Tn[4] XA.XIR[5].XIC[2].icell.SM 0.00121f
C5257 XA.XIR[2].XIC[0].icell.SM Iout 0.00388f
C5258 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01577f
C5259 XThC.Tn[13] XThR.Tn[1] 0.2874f
C5260 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.04617f
C5261 XA.XIR[6].XIC[14].icell.SM Vbias 0.00701f
C5262 XA.XIR[11].XIC[1].icell.SM Iout 0.00388f
C5263 XA.XIR[10].XIC[7].icell.SM VPWR 0.00158f
C5264 XA.XIR[15].XIC[9].icell.SM Iout 0.00388f
C5265 XThR.Tn[14] XA.XIR[15].XIC[4].icell.Ien 0.00338f
C5266 XThR.Tn[3] XA.XIR[4].XIC[2].icell.SM 0.00121f
C5267 XThR.XTBN.A data[7] 0.07741f
C5268 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5269 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.15202f
C5270 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.03425f
C5271 XA.XIR[2].XIC[4].icell.PUM Vbias 0.0031f
C5272 XA.XIR[7].XIC[4].icell.Ien Vbias 0.21098f
C5273 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C5274 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C5275 XA.XIR[4].XIC_15.icell.PDM Vbias 0.04401f
C5276 XA.XIR[0].XIC[8].icell.PUM VPWR 0.00881f
C5277 XA.XIR[10].XIC[3].icell.SM Iout 0.00388f
C5278 XThC.XTB2.Y a_5155_9615# 0.00847f
C5279 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C5280 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00214f
C5281 XThR.Tn[9] XA.XIR[10].XIC[3].icell.SM 0.00121f
C5282 XThC.Tn[13] XThR.Tn[12] 0.2874f
C5283 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04031f
C5284 XA.XIR[1].XIC[6].icell.PUM Vbias 0.0031f
C5285 XThR.XTB7.B a_n1319_5317# 0.00108f
C5286 XA.XIR[14].XIC[8].icell.SM Vbias 0.00701f
C5287 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04031f
C5288 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C5289 XThC.XTB6.A XThC.XTBN.A 0.0513f
C5290 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.03425f
C5291 XThC.XTBN.Y XThC.Tn[11] 0.53369f
C5292 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02762f
C5293 XA.XIR[3].XIC[12].icell.SM Iout 0.00388f
C5294 XThC.Tn[8] XThR.Tn[4] 0.28739f
C5295 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04031f
C5296 a_n1049_7787# XThR.Tn[2] 0.00158f
C5297 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8] 0.00341f
C5298 XA.XIR[8].XIC[14].icell.PUM Vbias 0.0031f
C5299 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38936f
C5300 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[8].icell.SM 0.0039f
C5301 XA.XIR[2].XIC[9].icell.SM VPWR 0.00158f
C5302 XA.XIR[7].XIC[11].icell.PUM VPWR 0.00937f
C5303 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.SM 0.0039f
C5304 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02762f
C5305 XA.XIR[3].XIC_15.icell.SM Vbias 0.00701f
C5306 XA.XIR[2].XIC[5].icell.SM Iout 0.00388f
C5307 XA.XIR[1].XIC[11].icell.SM VPWR 0.00158f
C5308 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00214f
C5309 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04031f
C5310 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.SM 0.0039f
C5311 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.SM 0.00168f
C5312 XThR.Tn[12] XA.XIR[13].XIC[1].icell.SM 0.00121f
C5313 XA.XIR[1].XIC[7].icell.SM Iout 0.00388f
C5314 XThC.Tn[2] XThR.Tn[0] 0.28882f
C5315 XThC.Tn[12] XThR.Tn[10] 0.28739f
C5316 XA.XIR[9].XIC_15.icell.SM Iout 0.0047f
C5317 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.SM 0.00168f
C5318 XThC.Tn[4] XThR.Tn[5] 0.28739f
C5319 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00214f
C5320 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.15202f
C5321 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00214f
C5322 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PUM 0.00465f
C5323 XA.XIR[8].XIC[1].icell.PUM VPWR 0.00937f
C5324 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.SM 0.0039f
C5325 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.15202f
C5326 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C5327 XThC.Tn[10] XThC.Tn[11] 0.09949f
C5328 XThR.Tn[11] XA.XIR[12].XIC[4].icell.SM 0.00121f
C5329 XA.XIR[0].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5330 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02762f
C5331 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.SM 0.00168f
C5332 XThC.XTB6.Y a_7875_9569# 0.0046f
C5333 XThR.Tn[7] VPWR 6.97893f
C5334 XThR.Tn[2] XA.XIR[3].XIC[10].icell.Ien 0.00338f
C5335 a_n997_2891# VPWR 0.01347f
C5336 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04031f
C5337 XThR.Tn[4] XA.XIR[4].XIC_15.icell.PDM 0.00341f
C5338 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.SM 0.0039f
C5339 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PUM 0.00465f
C5340 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C5341 XA.XIR[5].XIC[0].icell.PDM Vbias 0.04207f
C5342 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.03425f
C5343 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C5344 XA.XIR[7].XIC_15.icell.SM VPWR 0.00275f
C5345 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.03425f
C5346 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10] 0.00341f
C5347 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PUM 0.00429f
C5348 XA.XIR[7].XIC[5].icell.PDM VPWR 0.00799f
C5349 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.15202f
C5350 XA.XIR[6].XIC[1].icell.PUM Vbias 0.0031f
C5351 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C5352 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Iout 0.00347f
C5353 XThR.Tn[1] XA.XIR[2].XIC[8].icell.SM 0.00121f
C5354 XA.XIR[4].XIC[2].icell.Ien VPWR 0.1903f
C5355 XThR.XTB6.Y a_n1049_5317# 0.01199f
C5356 XA.XIR[6].XIC[12].icell.PDM VPWR 0.00799f
C5357 XA.XIR[15].XIC[3].icell.PDM VPWR 0.0114f
C5358 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C5359 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PUM 0.00465f
C5360 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.03425f
C5361 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C5362 XA.XIR[14].XIC[9].icell.PDM VPWR 0.00799f
C5363 XA.XIR[6].XIC[0].icell.PDM Iout 0.00117f
C5364 XA.XIR[11].XIC[5].icell.PDM Vbias 0.04261f
C5365 XA.XIR[15].XIC[13].icell.Ien Iout 0.06807f
C5366 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.03425f
C5367 XA.XIR[11].XIC[11].icell.SM Vbias 0.00701f
C5368 XA.XIR[5].XIC[7].icell.PDM Iout 0.00117f
C5369 XThR.Tn[11] XA.XIR[12].XIC[10].icell.Ien 0.00338f
C5370 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C5371 XA.XIR[10].XIC[9].icell.PDM Vbias 0.04261f
C5372 XA.XIR[9].XIC[1].icell.PDM VPWR 0.00799f
C5373 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Ien 0.00232f
C5374 XA.XIR[13].XIC[1].icell.PDM Iout 0.00117f
C5375 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02762f
C5376 XThC.Tn[1] XThR.Tn[2] 0.28739f
C5377 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.SM 0.0039f
C5378 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.SM 0.00168f
C5379 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.SM 0.00168f
C5380 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PUM 0.00465f
C5381 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00214f
C5382 XA.XIR[12].XIC[6].icell.PDM Iout 0.00117f
C5383 XA.XIR[6].XIC[6].icell.PUM Vbias 0.0031f
C5384 XA.XIR[12].XIC[12].icell.SM VPWR 0.00158f
C5385 XA.XIR[9].XIC[5].icell.Ien VPWR 0.1903f
C5386 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.SM 0.00168f
C5387 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00584f
C5388 XThR.XTB5.A data[5] 0.11096f
C5389 XThC.Tn[10] XThR.Tn[14] 0.28739f
C5390 XThC.XTB4.Y a_7875_9569# 0.00497f
C5391 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00584f
C5392 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.SM 0.0039f
C5393 XA.XIR[15].XIC[7].icell.Ien Vbias 0.17899f
C5394 XA.XIR[5].XIC[7].icell.SM Vbias 0.00701f
C5395 XThC.XTB1.Y a_3299_10575# 0.0097f
C5396 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02762f
C5397 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C5398 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C5399 XThR.XTBN.Y a_n1049_7787# 0.08456f
C5400 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C5401 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.04036f
C5402 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00584f
C5403 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C5404 XThR.XTB2.Y data[4] 0.00267f
C5405 XThR.XTB7.Y a_n997_3755# 0.00476f
C5406 XA.XIR[7].XIC_dummy_left.icell.Ien Vbias 0.00329f
C5407 XA.XIR[4].XIC[10].icell.Ien Vbias 0.21098f
C5408 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00214f
C5409 XA.XIR[3].XIC[8].icell.PUM VPWR 0.00937f
C5410 XA.XIR[1].XIC[6].icell.PDM VPWR 0.00799f
C5411 XThC.XTB6.A XThC.Tn[2] 0.00108f
C5412 XThR.Tn[14] XA.XIR[15].XIC[12].icell.SM 0.00121f
C5413 XA.XIR[0].XIC[1].icell.Ien Vbias 0.2113f
C5414 XA.XIR[6].XIC[11].icell.SM VPWR 0.00158f
C5415 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02762f
C5416 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C5417 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.15202f
C5418 XA.XIR[15].XIC[14].icell.SM Iout 0.00388f
C5419 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.SM 0.00168f
C5420 a_n1049_6405# XThR.Tn[4] 0.26564f
C5421 XA.XIR[2].XIC[1].icell.PDM Vbias 0.04261f
C5422 a_5155_9615# XThC.Tn[4] 0.26653f
C5423 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5424 XA.XIR[11].XIC[14].icell.PUM Vbias 0.0031f
C5425 XA.XIR[8].XIC[4].icell.Ien Vbias 0.21098f
C5426 XA.XIR[6].XIC[7].icell.SM Iout 0.00388f
C5427 XA.XIR[4].XIC[6].icell.PDM VPWR 0.00799f
C5428 XA.XIR[5].XIC[14].icell.Ien VPWR 0.19036f
C5429 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7] 0.00341f
C5430 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04031f
C5431 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.0353f
C5432 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.SM 0.00168f
C5433 XA.XIR[12].XIC[2].icell.SM Vbias 0.00701f
C5434 XA.XIR[3].XIC[14].icell.PDM VPWR 0.00809f
C5435 XA.XIR[5].XIC[10].icell.Ien Iout 0.06417f
C5436 XA.XIR[1].XIC[3].icell.PUM VPWR 0.00937f
C5437 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5438 XA.XIR[14].XIC[5].icell.SM VPWR 0.00158f
C5439 XA.XIR[14].XIC[13].icell.SM Vbias 0.00701f
C5440 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13] 0.00341f
C5441 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.SM 0.00168f
C5442 XA.XIR[11].XIC[5].icell.PUM Vbias 0.0031f
C5443 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.SM 0.00168f
C5444 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C5445 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.SM 0.00168f
C5446 XA.XIR[8].XIC[4].icell.PDM Iout 0.00117f
C5447 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01577f
C5448 XA.XIR[3].XIC[2].icell.PDM Iout 0.00117f
C5449 XThC.Tn[6] XThR.Tn[6] 0.28739f
C5450 XThC.XTBN.A XThC.Tn[8] 0.1369f
C5451 XA.XIR[13].XIC[7].icell.SM VPWR 0.00158f
C5452 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04031f
C5453 XA.XIR[14].XIC[1].icell.SM Iout 0.00388f
C5454 XA.XIR[9].XIC[13].icell.Ien Vbias 0.21098f
C5455 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00584f
C5456 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00214f
C5457 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04031f
C5458 a_n1049_5611# XThR.XTB7.Y 0.00153f
C5459 XA.XIR[10].XIC[7].icell.PUM Vbias 0.0031f
C5460 XA.XIR[8].XIC[11].icell.PUM VPWR 0.00937f
C5461 XA.XIR[2].XIC[8].icell.PDM Iout 0.00117f
C5462 XThR.Tn[6] XA.XIR[7].XIC[9].icell.Ien 0.00338f
C5463 XA.XIR[12].XIC[9].icell.Ien VPWR 0.1903f
C5464 XA.XIR[13].XIC[3].icell.SM Iout 0.00388f
C5465 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C5466 XA.XIR[0].XIC[6].icell.Ien Vbias 0.21134f
C5467 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00584f
C5468 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5469 XThR.Tn[0] XA.XIR[0].XIC[5].icell.PDM 0.00341f
C5470 XA.XIR[12].XIC[5].icell.Ien Iout 0.06417f
C5471 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.SM 0.00168f
C5472 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02762f
C5473 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PUM 0.00186f
C5474 XA.XIR[3].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5475 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00214f
C5476 XThR.Tn[4] XA.XIR[5].XIC[7].icell.SM 0.00121f
C5477 XThC.Tn[6] Vbias 2.22871f
C5478 XThR.Tn[1] XA.XIR[1].XIC[3].icell.PDM 0.00341f
C5479 XA.XIR[9].XIC[0].icell.Ien VPWR 0.1903f
C5480 XA.XIR[11].XIC[6].icell.SM Iout 0.00388f
C5481 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C5482 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00584f
C5483 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.15202f
C5484 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04031f
C5485 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.SM 0.00168f
C5486 XThR.Tn[3] XA.XIR[4].XIC[7].icell.SM 0.00121f
C5487 XThR.Tn[14] XA.XIR[15].XIC[9].icell.Ien 0.00338f
C5488 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02762f
C5489 XA.XIR[2].XIC[9].icell.PUM Vbias 0.0031f
C5490 XA.XIR[7].XIC[9].icell.Ien Vbias 0.21098f
C5491 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PUM 0.00465f
C5492 XA.XIR[15].XIC[11].icell.Ien Iout 0.06807f
C5493 XThR.Tn[9] XA.XIR[10].XIC[8].icell.SM 0.00121f
C5494 XA.XIR[0].XIC[13].icell.PUM VPWR 0.00877f
C5495 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02762f
C5496 XA.XIR[11].XIC[9].icell.SM Vbias 0.00701f
C5497 XA.XIR[10].XIC[8].icell.SM Iout 0.00388f
C5498 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.15202f
C5499 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5] 0.00341f
C5500 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.SM 0.0039f
C5501 XThC.XTB6.Y XThC.Tn[4] 0.00264f
C5502 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00214f
C5503 XThC.XTB7.A a_5949_9615# 0.01824f
C5504 XA.XIR[1].XIC[11].icell.PUM Vbias 0.0031f
C5505 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PUM 0.00465f
C5506 XA.XIR[8].XIC_15.icell.SM VPWR 0.00275f
C5507 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.03425f
C5508 XA.XIR[12].XIC_15.icell.SM Iout 0.0047f
C5509 XThC.Tn[12] XThR.Tn[13] 0.28739f
C5510 XThR.Tn[2] XA.XIR[2].XIC[0].icell.PDM 0.00347f
C5511 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00214f
C5512 XThC.Tn[2] XThR.Tn[1] 0.28742f
C5513 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04031f
C5514 XA.XIR[2].XIC[14].icell.SM VPWR 0.00207f
C5515 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C5516 XA.XIR[12].XIC[10].icell.SM VPWR 0.00158f
C5517 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.15202f
C5518 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5519 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02762f
C5520 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10] 0.00341f
C5521 XThC.XTB2.Y a_7875_9569# 0.06476f
C5522 XA.XIR[5].XIC[1].icell.PUM VPWR 0.00937f
C5523 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6] 0.00341f
C5524 XA.XIR[2].XIC[10].icell.SM Iout 0.00388f
C5525 XThC.Tn[2] XThR.Tn[12] 0.28739f
C5526 XA.XIR[2].XIC[0].icell.Ien Vbias 0.20951f
C5527 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.SM 0.00168f
C5528 a_n997_1579# VPWR 0.02417f
C5529 XThC.XTB5.A XThC.XTB7.A 0.07824f
C5530 XThC.Tn[11] XThR.Tn[8] 0.28739f
C5531 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.SM 0.00168f
C5532 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C5533 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.SM 0.00168f
C5534 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C5535 XThR.Tn[12] XA.XIR[13].XIC[6].icell.SM 0.00121f
C5536 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00584f
C5537 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.03425f
C5538 XA.XIR[1].XIC[12].icell.SM Iout 0.00388f
C5539 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.SM 0.00168f
C5540 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00214f
C5541 XThR.XTB3.Y a_n1049_6699# 0.0093f
C5542 XThR.Tn[11] XA.XIR[12].XIC_15.icell.Ien 0.00117f
C5543 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C5544 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00584f
C5545 XThR.Tn[14] XA.XIR[15].XIC[10].icell.SM 0.00121f
C5546 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.15202f
C5547 data[1] data[2] 0.01393f
C5548 XA.XIR[10].XIC[1].icell.Ien Vbias 0.21098f
C5549 XA.XIR[10].XIC[0].icell.PDM VPWR 0.00799f
C5550 XA.XIR[7].XIC[1].icell.PDM Vbias 0.04261f
C5551 XThC.XTBN.Y XThC.Tn[0] 0.53577f
C5552 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C5553 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.03023f
C5554 XA.XIR[11].XIC[12].icell.PUM Vbias 0.0031f
C5555 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00584f
C5556 XA.XIR[1].XIC_15.icell.SM Vbias 0.00704f
C5557 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.15202f
C5558 XThC.Tn[6] XThR.Tn[4] 0.28739f
C5559 XA.XIR[6].XIC[8].icell.PDM Vbias 0.04261f
C5560 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PUM 0.00465f
C5561 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PUM 0.00465f
C5562 XThR.Tn[2] XA.XIR[3].XIC_15.icell.Ien 0.00117f
C5563 XA.XIR[6].XIC[3].icell.PUM VPWR 0.00937f
C5564 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C5565 XA.XIR[14].XIC[5].icell.PDM Vbias 0.04261f
C5566 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.03425f
C5567 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C5568 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.SM 0.00168f
C5569 XA.XIR[5].XIC_15.icell.PDM Vbias 0.04401f
C5570 XA.XIR[14].XIC[11].icell.SM Vbias 0.00701f
C5571 XThC.XTB4.Y XThC.Tn[4] 0.00758f
C5572 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C5573 XA.XIR[15].XIC[4].icell.Ien VPWR 0.32895f
C5574 XThC.Tn[1] XThR.Tn[10] 0.28739f
C5575 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02762f
C5576 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.03425f
C5577 XA.XIR[5].XIC[4].icell.SM VPWR 0.00158f
C5578 XA.XIR[12].XIC[13].icell.PUM VPWR 0.00937f
C5579 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00214f
C5580 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.15202f
C5581 XThC.XTB3.Y XThC.Tn[8] 0.00178f
C5582 XA.XIR[13].XIC[9].icell.PDM Vbias 0.04261f
C5583 XA.XIR[7].XIC[8].icell.PDM Iout 0.00117f
C5584 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02762f
C5585 XA.XIR[4].XIC[7].icell.Ien VPWR 0.1903f
C5586 XThR.Tn[1] XA.XIR[2].XIC[13].icell.SM 0.00121f
C5587 XA.XIR[9].XIC[1].icell.Ien Iout 0.06417f
C5588 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.15202f
C5589 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.SM 0.0039f
C5590 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02823f
C5591 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.PDM 0.00591f
C5592 XA.XIR[6].XIC_15.icell.PDM Iout 0.00133f
C5593 XThR.XTB7.Y a_n997_715# 0.06874f
C5594 XA.XIR[15].XIC[6].icell.PDM Iout 0.00117f
C5595 XA.XIR[4].XIC[3].icell.Ien Iout 0.06417f
C5596 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.0343f
C5597 XA.XIR[9].XIC[3].icell.SM Vbias 0.00701f
C5598 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00214f
C5599 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02762f
C5600 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.03425f
C5601 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02762f
C5602 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00584f
C5603 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C5604 XA.XIR[11].XIC[13].icell.Ien Vbias 0.21098f
C5605 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5606 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.SM 0.00168f
C5607 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.15202f
C5608 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01093f
C5609 XA.XIR[7].XIC[1].icell.Ien VPWR 0.1903f
C5610 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00214f
C5611 XThC.XTB5.Y VPWR 1.01191f
C5612 XA.XIR[9].XIC[4].icell.PDM Iout 0.00117f
C5613 XA.XIR[1].XIC[2].icell.PDM Vbias 0.04261f
C5614 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9] 0.00341f
C5615 XA.XIR[3].XIC[6].icell.Ien Vbias 0.21098f
C5616 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02762f
C5617 XA.XIR[9].XIC[10].icell.Ien VPWR 0.1903f
C5618 XA.XIR[6].XIC[11].icell.PUM Vbias 0.0031f
C5619 XA.XIR[14].XIC[14].icell.PUM Vbias 0.0031f
C5620 XA.XIR[10].XIC[4].icell.PUM VPWR 0.00937f
C5621 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PUM 0.00465f
C5622 XA.XIR[9].XIC[6].icell.Ien Iout 0.06417f
C5623 XA.XIR[12].XIC[14].icell.Ien VPWR 0.19036f
C5624 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.SM 0.0039f
C5625 XA.XIR[5].XIC[12].icell.SM Vbias 0.00701f
C5626 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.15202f
C5627 XA.XIR[4].XIC[2].icell.PDM Vbias 0.04261f
C5628 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.0353f
C5629 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18966f
C5630 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C5631 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.SM 0.0039f
C5632 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00214f
C5633 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04031f
C5634 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PDM 0.00172f
C5635 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04031f
C5636 XA.XIR[8].XIC[12].icell.PDM Vbias 0.04261f
C5637 XA.XIR[3].XIC[13].icell.PUM VPWR 0.00937f
C5638 XA.XIR[4].XIC_15.icell.Ien Vbias 0.21234f
C5639 XA.XIR[3].XIC[10].icell.PDM Vbias 0.04261f
C5640 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.SM 0.0039f
C5641 XA.XIR[14].XIC[5].icell.PUM Vbias 0.0031f
C5642 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10] 0.00341f
C5643 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PUM 0.00465f
C5644 XA.XIR[1].XIC[9].icell.PDM Iout 0.00117f
C5645 XThR.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.00338f
C5646 XA.XIR[13].XIC[7].icell.PUM Vbias 0.0031f
C5647 XA.XIR[6].XIC[12].icell.SM Iout 0.00388f
C5648 XA.XIR[8].XIC[9].icell.Ien Vbias 0.21098f
C5649 XA.XIR[2].XIC[6].icell.PUM VPWR 0.00937f
C5650 XA.XIR[7].XIC[6].icell.Ien VPWR 0.1903f
C5651 XA.XIR[10].XIC[13].icell.SM Iout 0.00388f
C5652 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00584f
C5653 XA.XIR[11].XIC[14].icell.SM Vbias 0.00701f
C5654 XThR.Tn[9] XA.XIR[10].XIC[13].icell.SM 0.00121f
C5655 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00584f
C5656 XA.XIR[12].XIC[7].icell.SM Vbias 0.00701f
C5657 XA.XIR[9].XIC_dummy_left.icell.SM VPWR 0.00269f
C5658 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00214f
C5659 XA.XIR[4].XIC[9].icell.PDM Iout 0.00117f
C5660 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.SM 0.0039f
C5661 XA.XIR[5].XIC_15.icell.Ien Iout 0.0642f
C5662 XThC.XTBN.Y VPWR 4.08849f
C5663 XA.XIR[1].XIC[8].icell.PUM VPWR 0.00937f
C5664 XA.XIR[7].XIC[2].icell.Ien Iout 0.06417f
C5665 XA.XIR[6].XIC_15.icell.SM Vbias 0.00701f
C5666 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.03425f
C5667 XThC.XTB6.Y a_6243_9615# 0.01199f
C5668 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C5669 XA.XIR[11].XIC[10].icell.PUM Vbias 0.0031f
C5670 XThR.XTB7.A XThR.XTBN.A 0.19736f
C5671 a_n1049_6699# VPWR 0.72162f
C5672 XA.XIR[14].XIC[6].icell.SM Iout 0.00388f
C5673 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C5674 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02762f
C5675 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5676 XThR.Tn[7] XA.XIR[8].XIC[3].icell.Ien 0.00338f
C5677 XA.XIR[12].XIC_15.icell.PDM Iout 0.00133f
C5678 XThR.Tn[6] XA.XIR[7].XIC[14].icell.Ien 0.00338f
C5679 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.SM 0.0039f
C5680 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00584f
C5681 XThR.XTB7.A XThR.Tn[6] 0.1056f
C5682 XA.XIR[13].XIC[8].icell.SM Iout 0.00388f
C5683 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00214f
C5684 XA.XIR[14].XIC[9].icell.SM Vbias 0.00701f
C5685 XA.XIR[0].XIC[11].icell.Ien Vbias 0.2113f
C5686 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00214f
C5687 XThC.XTB1.Y XThC.Tn[8] 0.29191f
C5688 XA.XIR[12].XIC[11].icell.PUM VPWR 0.00937f
C5689 XThR.Tn[2] XA.XIR[3].XIC[5].icell.SM 0.00121f
C5690 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10] 0.00341f
C5691 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00214f
C5692 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.15202f
C5693 XThR.Tn[4] XA.XIR[5].XIC[12].icell.SM 0.00121f
C5694 XThR.Tn[4] XA.XIR[4].XIC[2].icell.PDM 0.00341f
C5695 XThC.Tn[10] VPWR 6.83631f
C5696 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.03425f
C5697 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.SM 0.0039f
C5698 XThR.Tn[10] XA.XIR[11].XIC[4].icell.Ien 0.00338f
C5699 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C5700 XThR.Tn[3] XA.XIR[4].XIC[12].icell.SM 0.00121f
C5701 XThR.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.00341f
C5702 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.03425f
C5703 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.03425f
C5704 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PUM 0.00465f
C5705 a_4861_9615# VPWR 0.70525f
C5706 XA.XIR[7].XIC[14].icell.Ien Vbias 0.21098f
C5707 XThR.Tn[9] Iout 1.16233f
C5708 XA.XIR[2].XIC[14].icell.PUM Vbias 0.0031f
C5709 XThC.XTBN.A XThC.Tn[6] 0.00131f
C5710 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.SM 0.0039f
C5711 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00214f
C5712 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.SM 0.00168f
C5713 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C5714 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.15202f
C5715 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.15202f
C5716 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5717 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Ien 0.00584f
C5718 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04031f
C5719 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PUM 0.0044f
C5720 XA.XIR[15].XIC[12].icell.SM VPWR 0.00158f
C5721 XA.XIR[1].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5722 XA.XIR[11].XIC[11].icell.Ien Vbias 0.21098f
C5723 XA.XIR[5].XIC[6].icell.PDM VPWR 0.00799f
C5724 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.03425f
C5725 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13] 0.00341f
C5726 XA.XIR[4].XIC[0].icell.SM Vbias 0.00675f
C5727 XThR.Tn[2] XA.XIR[2].XIC_15.icell.PDM 0.00341f
C5728 XThC.XTB4.Y a_6243_9615# 0.00463f
C5729 XA.XIR[13].XIC[1].icell.Ien Vbias 0.21098f
C5730 XA.XIR[13].XIC[0].icell.PDM VPWR 0.00799f
C5731 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PUM 0.00465f
C5732 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[13].icell.SM 0.0039f
C5733 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00584f
C5734 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.15202f
C5735 XA.XIR[14].XIC[12].icell.PUM Vbias 0.0031f
C5736 XThC.XTB5.Y a_9827_9569# 0.06458f
C5737 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.SM 0.00168f
C5738 XA.XIR[12].XIC[5].icell.PDM VPWR 0.00799f
C5739 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C5740 XA.XIR[12].XIC[12].icell.Ien VPWR 0.1903f
C5741 XThC.XTB7.A a_8739_9569# 0.00342f
C5742 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.SM 0.0039f
C5743 XA.XIR[15].XIC[0].icell.Ien Iout 0.06801f
C5744 XA.XIR[5].XIC[0].icell.SM Iout 0.00388f
C5745 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.SM 0.00168f
C5746 XThC.Tn[1] XThR.Tn[13] 0.28739f
C5747 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.SM 0.00168f
C5748 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02762f
C5749 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.03425f
C5750 XA.XIR[15].XIC[2].icell.SM Vbias 0.00701f
C5751 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00214f
C5752 XA.XIR[5].XIC[4].icell.PUM Vbias 0.0031f
C5753 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C5754 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PUM 0.00465f
C5755 XA.XIR[8].XIC[1].icell.Ien VPWR 0.1903f
C5756 XThR.XTB3.Y XThR.Tn[8] 0.00178f
C5757 XThR.Tn[14] XA.XIR[15].XIC[12].icell.Ien 0.00338f
C5758 XA.XIR[10].XIC[3].icell.PDM Iout 0.00117f
C5759 XA.XIR[4].XIC[5].icell.SM Vbias 0.00701f
C5760 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01577f
C5761 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00584f
C5762 XA.XIR[10].XIC[11].icell.SM Iout 0.00388f
C5763 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04031f
C5764 XA.XIR[3].XIC[3].icell.Ien VPWR 0.1903f
C5765 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00584f
C5766 XThC.Tn[4] Iout 0.83918f
C5767 XThR.Tn[9] XA.XIR[10].XIC[11].icell.SM 0.00121f
C5768 XThC.Tn[4] XThR.Tn[9] 0.28739f
C5769 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02762f
C5770 XA.XIR[6].XIC[8].icell.PUM VPWR 0.00937f
C5771 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.03425f
C5772 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00584f
C5773 XThC.Tn[0] XThR.Tn[8] 0.2874f
C5774 a_5155_10571# VPWR 0.00653f
C5775 XThR.XTB7.Y a_n997_2667# 0.00474f
C5776 XThR.XTB7.A XThR.Tn[4] 0.02736f
C5777 XA.XIR[15].XIC[9].icell.Ien VPWR 0.32895f
C5778 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.SM 0.0039f
C5779 XA.XIR[5].XIC[9].icell.SM VPWR 0.00158f
C5780 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.15202f
C5781 XThC.XTBN.Y a_9827_9569# 0.22873f
C5782 XA.XIR[14].XIC[13].icell.Ien Vbias 0.21098f
C5783 XThR.XTB7.A a_n1049_7493# 0.0127f
C5784 XA.XIR[15].XIC[5].icell.Ien Iout 0.06807f
C5785 XA.XIR[3].XIC[1].icell.PDM VPWR 0.00799f
C5786 XA.XIR[9].XIC[12].icell.PDM Vbias 0.04261f
C5787 XA.XIR[4].XIC[12].icell.Ien VPWR 0.1903f
C5788 XA.XIR[5].XIC[5].icell.SM Iout 0.00388f
C5789 XA.XIR[8].XIC[3].icell.PDM VPWR 0.00799f
C5790 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C5791 XA.XIR[0].XIC[4].icell.PDM Vbias 0.04271f
C5792 XA.XIR[2].XIC[7].icell.PDM VPWR 0.00799f
C5793 XA.XIR[4].XIC[8].icell.Ien Iout 0.06417f
C5794 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.15202f
C5795 XA.XIR[1].XIC[1].icell.Ien Vbias 0.21104f
C5796 XA.XIR[13].XIC[4].icell.PUM VPWR 0.00937f
C5797 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00214f
C5798 XA.XIR[9].XIC[8].icell.SM Vbias 0.00701f
C5799 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.SM 0.0039f
C5800 XA.XIR[10].XIC[2].icell.Ien Vbias 0.21098f
C5801 XA.XIR[8].XIC[6].icell.Ien VPWR 0.1903f
C5802 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.SM 0.0039f
C5803 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C5804 XThR.Tn[6] XA.XIR[7].XIC[4].icell.SM 0.00121f
C5805 XA.XIR[12].XIC[4].icell.SM VPWR 0.00158f
C5806 XA.XIR[8].XIC[2].icell.Ien Iout 0.06417f
C5807 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12] 0.00341f
C5808 XThR.Tn[8] XA.XIR[9].XIC[2].icell.Ien 0.00338f
C5809 XA.XIR[0].XIC[1].icell.SM Vbias 0.00716f
C5810 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PUM 0.00465f
C5811 XA.XIR[15].XIC_15.icell.SM Iout 0.0047f
C5812 XA.XIR[11].XIC[7].icell.PUM VPWR 0.00937f
C5813 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.SM 0.00168f
C5814 XThC.XTB3.Y XThC.Tn[6] 0.00301f
C5815 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04031f
C5816 XA.XIR[3].XIC[11].icell.Ien Vbias 0.21098f
C5817 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00214f
C5818 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C5819 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00256f
C5820 XA.XIR[9].XIC_15.icell.Ien VPWR 0.25566f
C5821 XA.XIR[6].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5822 XA.XIR[15].XIC[10].icell.SM VPWR 0.00158f
C5823 XA.XIR[10].XIC[9].icell.PUM VPWR 0.00937f
C5824 XThC.Tn[3] XThC.Tn[5] 0.00492f
C5825 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00584f
C5826 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C5827 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5828 XThR.Tn[14] XA.XIR[15].XIC[4].icell.SM 0.00121f
C5829 XThR.XTB7.B XThR.XTBN.A 0.35142f
C5830 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C5831 XA.XIR[2].XIC[4].icell.Ien Vbias 0.21098f
C5832 XA.XIR[9].XIC[11].icell.Ien Iout 0.06417f
C5833 XA.XIR[13].XIC[13].icell.SM Iout 0.00388f
C5834 XA.XIR[14].XIC[14].icell.SM Vbias 0.00701f
C5835 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C5836 XA.XIR[7].XIC[4].icell.SM Vbias 0.00701f
C5837 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.15202f
C5838 XThC.XTB2.Y a_6243_9615# 0.00844f
C5839 XA.XIR[0].XIC[8].icell.Ien VPWR 0.19149f
C5840 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.SM 0.00168f
C5841 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C5842 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.SM 0.0039f
C5843 XA.XIR[12].XIC[14].icell.PDM Iout 0.00117f
C5844 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.SM 0.00168f
C5845 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PUM 0.00465f
C5846 XThC.XTB2.Y data[1] 0.017f
C5847 XA.XIR[1].XIC[6].icell.Ien Vbias 0.21104f
C5848 XThR.XTB7.B XThR.Tn[6] 0.04822f
C5849 XA.XIR[0].XIC[4].icell.Ien Iout 0.06389f
C5850 XThR.Tn[10] XA.XIR[11].XIC[12].icell.SM 0.00121f
C5851 XA.XIR[14].XIC[10].icell.PUM Vbias 0.0031f
C5852 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C5853 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04031f
C5854 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PUM 0.00465f
C5855 XA.XIR[12].XIC[10].icell.Ien VPWR 0.1903f
C5856 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.SM 0.0039f
C5857 XThC.XTB3.Y a_4387_10575# 0.00941f
C5858 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10] 0.00341f
C5859 XA.XIR[15].XIC_15.icell.PDM Iout 0.00133f
C5860 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04031f
C5861 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8] 0.00341f
C5862 XA.XIR[2].XIC[11].icell.PUM VPWR 0.00937f
C5863 XA.XIR[8].XIC[14].icell.Ien Vbias 0.21098f
C5864 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PUM 0.00465f
C5865 XA.XIR[7].XIC[11].icell.Ien VPWR 0.1903f
C5866 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.SM 0.00168f
C5867 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.SM 0.0039f
C5868 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C5869 XThC.Tn[12] XThR.Tn[7] 0.28739f
C5870 XA.XIR[7].XIC[7].icell.Ien Iout 0.06417f
C5871 XA.XIR[1].XIC[13].icell.PUM VPWR 0.00937f
C5872 XA.XIR[11].XIC_dummy_left.icell.Ien Vbias 0.00329f
C5873 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02762f
C5874 XThR.Tn[0] XA.XIR[1].XIC[2].icell.Ien 0.00338f
C5875 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04031f
C5876 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C5877 XThC.XTB7.B XThC.Tn[10] 0.14845f
C5878 XThR.Tn[14] XA.XIR[15].XIC[10].icell.Ien 0.00338f
C5879 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C5880 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C5881 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.SM 0.00168f
C5882 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00584f
C5883 XA.XIR[15].XIC[13].icell.PUM VPWR 0.00937f
C5884 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C5885 XA.XIR[10].XIC[9].icell.SM Iout 0.00388f
C5886 XThR.Tn[9] XA.XIR[10].XIC[9].icell.SM 0.00121f
C5887 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Iout 0.00347f
C5888 XA.XIR[3].XIC[0].icell.Ien VPWR 0.1903f
C5889 XThR.Tn[7] XA.XIR[8].XIC[8].icell.Ien 0.00338f
C5890 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.15202f
C5891 XThR.Tn[8] VPWR 7.51456f
C5892 XThC.XTB7.B a_4861_9615# 0.0036f
C5893 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C5894 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.03425f
C5895 XThC.XTBN.A data[3] 0.07741f
C5896 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13] 0.00341f
C5897 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02762f
C5898 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.SM 0.00168f
C5899 XThR.Tn[5] XA.XIR[6].XIC[4].icell.Ien 0.00338f
C5900 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C5901 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C5902 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5903 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02762f
C5904 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C5905 XThC.XTB7.A data[0] 0.86893f
C5906 XThC.XTB6.Y a_8963_9569# 0.00468f
C5907 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PUM 0.00186f
C5908 XA.XIR[14].XIC[11].icell.Ien Vbias 0.21098f
C5909 XThR.Tn[2] XA.XIR[3].XIC[10].icell.SM 0.00121f
C5910 XA.XIR[11].XIC[1].icell.Ien VPWR 0.1903f
C5911 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04031f
C5912 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.03023f
C5913 XA.XIR[2].XIC_15.icell.SM VPWR 0.00275f
C5914 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.15202f
C5915 XA.XIR[5].XIC[2].icell.PDM Vbias 0.04261f
C5916 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.03529f
C5917 XA.XIR[7].XIC[7].icell.PDM VPWR 0.00799f
C5918 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00584f
C5919 XThR.Tn[10] XA.XIR[11].XIC[9].icell.Ien 0.00338f
C5920 XA.XIR[9].XIC[0].icell.SM VPWR 0.00158f
C5921 XThR.XTB3.Y a_n997_3755# 0.0061f
C5922 XA.XIR[6].XIC[1].icell.Ien Vbias 0.21098f
C5923 a_3773_9615# XThC.Tn[1] 0.27139f
C5924 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C5925 XThR.Tn[14] a_n997_715# 0.1927f
C5926 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00214f
C5927 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00214f
C5928 XA.XIR[4].XIC[2].icell.SM VPWR 0.00158f
C5929 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.15202f
C5930 XA.XIR[6].XIC[14].icell.PDM VPWR 0.00809f
C5931 XA.XIR[15].XIC[5].icell.PDM VPWR 0.0114f
C5932 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00584f
C5933 XA.XIR[12].XIC[1].icell.PDM Vbias 0.04261f
C5934 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.03425f
C5935 XThR.Tn[11] a_n997_2667# 0.19413f
C5936 XThR.Tn[2] Vbias 3.74868f
C5937 XA.XIR[6].XIC[2].icell.PDM Iout 0.00117f
C5938 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.15202f
C5939 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C5940 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.SM 0.0039f
C5941 XThC.Tn[11] XThR.Tn[3] 0.28739f
C5942 XA.XIR[11].XIC[7].icell.PDM Vbias 0.04261f
C5943 XA.XIR[15].XIC[14].icell.Ien VPWR 0.329f
C5944 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00214f
C5945 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00214f
C5946 XA.XIR[5].XIC[9].icell.PDM Iout 0.00117f
C5947 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01757f
C5948 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.15202f
C5949 XA.XIR[9].XIC[3].icell.PDM VPWR 0.00799f
C5950 a_7651_9569# VPWR 0.00385f
C5951 XThR.XTB7.B XThR.Tn[4] 0.00356f
C5952 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[2].icell.Ien 0.00214f
C5953 XA.XIR[13].XIC[3].icell.PDM Iout 0.00117f
C5954 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.SM 0.00168f
C5955 XA.XIR[13].XIC[11].icell.SM Iout 0.00388f
C5956 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C5957 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.SM 0.0039f
C5958 XThR.XTB3.Y a_n1049_5611# 0.009f
C5959 XA.XIR[3].XIC[1].icell.SM Vbias 0.00701f
C5960 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C5961 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.03425f
C5962 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PUM 0.00465f
C5963 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PUM 0.00102f
C5964 XA.XIR[12].XIC[8].icell.PDM Iout 0.00117f
C5965 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.SM 0.00168f
C5966 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02787f
C5967 XA.XIR[9].XIC[5].icell.SM VPWR 0.00158f
C5968 XA.XIR[6].XIC[6].icell.Ien Vbias 0.21098f
C5969 XThC.Tn[14] XThR.Tn[0] 0.28766f
C5970 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C5971 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00584f
C5972 XThC.XTB4.Y a_8963_9569# 0.07199f
C5973 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C5974 XThR.Tn[10] XA.XIR[11].XIC[10].icell.SM 0.00121f
C5975 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C5976 XA.XIR[9].XIC[1].icell.SM Iout 0.00388f
C5977 XA.XIR[15].XIC[7].icell.SM Vbias 0.00701f
C5978 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C5979 XA.XIR[5].XIC[9].icell.PUM Vbias 0.0031f
C5980 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.SM 0.0039f
C5981 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.SM 0.00168f
C5982 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02762f
C5983 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.SM 0.00168f
C5984 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04031f
C5985 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00214f
C5986 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C5987 XThR.Tn[11] XA.XIR[12].XIC[0].icell.Ien 0.0037f
C5988 XA.XIR[3].XIC[8].icell.Ien VPWR 0.1903f
C5989 XA.XIR[4].XIC[10].icell.SM Vbias 0.00701f
C5990 XA.XIR[1].XIC[8].icell.PDM VPWR 0.00799f
C5991 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PUM 0.00465f
C5992 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C5993 XA.XIR[6].XIC[13].icell.PUM VPWR 0.00937f
C5994 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C5995 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.SM 0.00168f
C5996 XA.XIR[2].XIC[3].icell.PDM Vbias 0.04261f
C5997 XA.XIR[10].XIC[13].icell.Ien Iout 0.06417f
C5998 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Iout 0.00347f
C5999 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C6000 XA.XIR[13].XIC[2].icell.Ien Vbias 0.21098f
C6001 XThR.Tn[9] XA.XIR[10].XIC[13].icell.Ien 0.00338f
C6002 XA.XIR[3].XIC[4].icell.Ien Iout 0.06417f
C6003 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.SM 0.0039f
C6004 XA.XIR[4].XIC[8].icell.PDM VPWR 0.00799f
C6005 XA.XIR[5].XIC[14].icell.SM VPWR 0.00207f
C6006 XA.XIR[8].XIC[4].icell.SM Vbias 0.00701f
C6007 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7] 0.00341f
C6008 XA.XIR[7].XIC[1].icell.SM VPWR 0.00158f
C6009 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00214f
C6010 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C6011 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04031f
C6012 XA.XIR[12].XIC[4].icell.PUM Vbias 0.0031f
C6013 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C6014 XA.XIR[15].XIC[11].icell.PUM VPWR 0.00937f
C6015 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00214f
C6016 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6017 XA.XIR[1].XIC[3].icell.Ien VPWR 0.1903f
C6018 XA.XIR[5].XIC[10].icell.SM Iout 0.00388f
C6019 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C6020 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02762f
C6021 XA.XIR[14].XIC[7].icell.PUM VPWR 0.00937f
C6022 XThC.XTB7.Y a_6243_10571# 0.01283f
C6023 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13] 0.00341f
C6024 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C6025 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C6026 a_n1049_7493# XThR.Tn[2] 0.26564f
C6027 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.SM 0.0039f
C6028 XA.XIR[11].XIC[5].icell.Ien Vbias 0.21098f
C6029 XA.XIR[12].XIC[13].icell.PDM Iout 0.00117f
C6030 XA.XIR[3].XIC[4].icell.PDM Iout 0.00117f
C6031 XA.XIR[12].XIC_15.icell.Ien VPWR 0.25566f
C6032 XThR.XTBN.Y XThR.Tn[6] 0.59882f
C6033 XA.XIR[8].XIC[6].icell.PDM Iout 0.00117f
C6034 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C6035 XA.XIR[4].XIC[13].icell.Ien Iout 0.06417f
C6036 XA.XIR[13].XIC[9].icell.PUM VPWR 0.00937f
C6037 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04031f
C6038 XThC.XTB5.A data[0] 0.14415f
C6039 XA.XIR[9].XIC[13].icell.SM Vbias 0.00701f
C6040 XA.XIR[10].XIC[7].icell.Ien Vbias 0.21098f
C6041 XA.XIR[8].XIC[11].icell.Ien VPWR 0.1903f
C6042 XA.XIR[2].XIC[10].icell.PDM Iout 0.00117f
C6043 XThR.Tn[6] XA.XIR[7].XIC[9].icell.SM 0.00121f
C6044 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C6045 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.SM 0.0039f
C6046 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.SM 0.00168f
C6047 XA.XIR[4].XIC_dummy_right.icell.Ien Vbias 0.00288f
C6048 XA.XIR[8].XIC[7].icell.Ien Iout 0.06417f
C6049 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10] 0.00341f
C6050 XA.XIR[15].XIC[14].icell.PDM Iout 0.00117f
C6051 XA.XIR[0].XIC[6].icell.SM Vbias 0.00716f
C6052 XThR.Tn[8] XA.XIR[9].XIC[7].icell.Ien 0.00338f
C6053 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C6054 XThR.Tn[0] XA.XIR[0].XIC[7].icell.PDM 0.00341f
C6055 XA.XIR[12].XIC[5].icell.SM Iout 0.00388f
C6056 XThC.Tn[13] XThR.Tn[2] 0.2874f
C6057 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C6058 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.SM 0.0039f
C6059 XThR.Tn[14] XA.XIR[15].XIC_15.icell.Ien 0.00117f
C6060 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Ien 0.00584f
C6061 XA.XIR[10].XIC[14].icell.SM Iout 0.00388f
C6062 XThR.Tn[1] XA.XIR[1].XIC[5].icell.PDM 0.00341f
C6063 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00584f
C6064 XA.XIR[11].XIC_15.icell.SM Vbias 0.00701f
C6065 XThR.XTBN.Y Vbias 0.00722f
C6066 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C6067 XThR.Tn[9] XA.XIR[10].XIC[14].icell.SM 0.00121f
C6068 a_n997_3755# VPWR 0.0133f
C6069 XThR.XTB2.Y VPWR 0.98816f
C6070 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04031f
C6071 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.SM 0.0039f
C6072 XA.XIR[9].XIC_dummy_right.icell.SM VPWR 0.00123f
C6073 XThC.Tn[0] XA.XIR[7].XIC_dummy_left.icell.Iout 0.00109f
C6074 XA.XIR[2].XIC[9].icell.Ien Vbias 0.21098f
C6075 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.03425f
C6076 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02762f
C6077 XA.XIR[7].XIC[9].icell.SM Vbias 0.00701f
C6078 XA.XIR[15].XIC[12].icell.Ien VPWR 0.32895f
C6079 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C6080 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18966f
C6081 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C6082 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00214f
C6083 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5] 0.00341f
C6084 XThR.XTB4.Y XThR.Tn[6] 0.00605f
C6085 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.SM 0.0039f
C6086 XA.XIR[3].XIC_dummy_left.icell.SM VPWR 0.00269f
C6087 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02762f
C6088 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13] 0.00341f
C6089 XA.XIR[1].XIC[11].icell.Ien Vbias 0.21104f
C6090 XThR.XTBN.A XThR.Tn[10] 0.12147f
C6091 XA.XIR[0].XIC[9].icell.Ien Iout 0.06389f
C6092 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.15202f
C6093 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.15202f
C6094 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.03425f
C6095 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6096 XThR.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.00341f
C6097 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PUM 0.00465f
C6098 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02762f
C6099 XA.XIR[13].XIC[9].icell.SM Iout 0.00388f
C6100 XThR.Tn[10] XA.XIR[11].XIC[14].icell.Ien 0.00338f
C6101 XThR.Tn[13] XA.XIR[14].XIC[4].icell.Ien 0.00338f
C6102 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04031f
C6103 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02762f
C6104 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02762f
C6105 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6106 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.SM 0.00168f
C6107 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00584f
C6108 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C6109 a_n1049_5611# VPWR 0.71817f
C6110 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6] 0.00341f
C6111 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.15202f
C6112 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00584f
C6113 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00214f
C6114 XA.XIR[7].XIC[12].icell.Ien Iout 0.06417f
C6115 XThR.Tn[0] XA.XIR[1].XIC[7].icell.Ien 0.00338f
C6116 XThC.Tn[9] XThR.Tn[6] 0.28739f
C6117 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C6118 XA.XIR[14].XIC[1].icell.Ien VPWR 0.19084f
C6119 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.SM 0.0039f
C6120 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C6121 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PUM 0.0047f
C6122 XA.XIR[11].XIC[1].icell.PUM Vbias 0.0031f
C6123 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C6124 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PUM 0.00465f
C6125 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.SM 0.0039f
C6126 XThR.Tn[7] XA.XIR[8].XIC[13].icell.Ien 0.00338f
C6127 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00584f
C6128 XA.XIR[10].XIC[2].icell.PDM VPWR 0.00799f
C6129 XA.XIR[7].XIC[3].icell.PDM Vbias 0.04261f
C6130 XThR.Tn[10] Vbias 3.7463f
C6131 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00214f
C6132 XA.XIR[10].XIC[11].icell.Ien Iout 0.06417f
C6133 XThC.Tn[11] XThR.Tn[11] 0.28739f
C6134 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00214f
C6135 XThR.Tn[9] XA.XIR[10].XIC[11].icell.Ien 0.00338f
C6136 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C6137 XThR.Tn[5] XA.XIR[6].XIC[9].icell.Ien 0.00338f
C6138 XA.XIR[15].XIC[1].icell.PDM Vbias 0.04261f
C6139 XA.XIR[3].XIC[1].icell.Ien Iout 0.06417f
C6140 XA.XIR[6].XIC[10].icell.PDM Vbias 0.04261f
C6141 XThR.XTBN.Y XThR.Tn[4] 0.60351f
C6142 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00214f
C6143 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.03425f
C6144 XThC.Tn[1] XThR.Tn[7] 0.28739f
C6145 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C6146 XA.XIR[6].XIC[3].icell.Ien VPWR 0.1903f
C6147 XThC.Tn[9] Vbias 2.3038f
C6148 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00214f
C6149 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.SM 0.00168f
C6150 XA.XIR[14].XIC[7].icell.PDM Vbias 0.04261f
C6151 XThR.XTBN.Y a_n1049_7493# 0.08456f
C6152 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C6153 XA.XIR[15].XIC[4].icell.SM VPWR 0.00158f
C6154 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C6155 XA.XIR[5].XIC[6].icell.PUM VPWR 0.00937f
C6156 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Ien 0.00618f
C6157 XThC.XTB7.B a_7651_9569# 0.01152f
C6158 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C6159 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PUM 0.00465f
C6160 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PUM 0.00186f
C6161 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00214f
C6162 XA.XIR[7].XIC[10].icell.PDM Iout 0.00117f
C6163 XA.XIR[4].XIC[7].icell.SM VPWR 0.00158f
C6164 XThC.XTB5.Y XThC.Tn[12] 0.32495f
C6165 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PUM 0.00465f
C6166 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.0353f
C6167 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.04041f
C6168 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00584f
C6169 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PUM 0.00465f
C6170 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.15202f
C6171 XThC.Tn[2] XA.XIR[0].XIC[4].icell.PDM 0.00353f
C6172 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C6173 XA.XIR[15].XIC[8].icell.PDM Iout 0.00117f
C6174 XA.XIR[4].XIC[3].icell.SM Iout 0.00388f
C6175 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C6176 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Iout 0.00347f
C6177 XA.XIR[9].XIC[5].icell.PUM Vbias 0.0031f
C6178 XA.XIR[8].XIC[1].icell.SM VPWR 0.00158f
C6179 XThC.Tn[14] XThR.Tn[1] 0.28745f
C6180 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.03425f
C6181 XThR.XTB4.Y XThR.Tn[4] 0.00757f
C6182 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C6183 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C6184 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00584f
C6185 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00584f
C6186 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02762f
C6187 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.1106f
C6188 XA.XIR[2].XIC[1].icell.Ien VPWR 0.1903f
C6189 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C6190 XThR.XTBN.Y XA.XIR[10].XIC_dummy_left.icell.Iout 0.00376f
C6191 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C6192 XA.XIR[0].XIC[10].icell.PDM VPWR 0.00774f
C6193 XA.XIR[11].XIC[2].icell.Ien VPWR 0.1903f
C6194 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.SM 0.0039f
C6195 XA.XIR[3].XIC[6].icell.SM Vbias 0.00701f
C6196 XThC.Tn[14] XThR.Tn[12] 0.28745f
C6197 XA.XIR[15].XIC[10].icell.Ien VPWR 0.32895f
C6198 XA.XIR[9].XIC[6].icell.PDM Iout 0.00117f
C6199 XA.XIR[1].XIC[4].icell.PDM Vbias 0.04261f
C6200 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9] 0.00341f
C6201 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.SM 0.0039f
C6202 XA.XIR[13].XIC[13].icell.Ien Iout 0.06417f
C6203 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00214f
C6204 XA.XIR[6].XIC[11].icell.Ien Vbias 0.21098f
C6205 XA.XIR[9].XIC[10].icell.SM VPWR 0.00158f
C6206 XThC.XTB7.A VPWR 0.87301f
C6207 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11] 0.00341f
C6208 XThC.Tn[0] XThR.Tn[3] 0.28747f
C6209 XA.XIR[10].XIC[4].icell.Ien VPWR 0.1903f
C6210 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.SM 0.00168f
C6211 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PUM 0.00465f
C6212 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.03425f
C6213 XA.XIR[12].XIC[12].icell.PDM Iout 0.00117f
C6214 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00214f
C6215 XA.XIR[4].XIC[4].icell.PDM Vbias 0.04261f
C6216 XA.XIR[9].XIC[6].icell.SM Iout 0.00388f
C6217 XThR.XTBN.A a_n997_1803# 0.09118f
C6218 XA.XIR[5].XIC[14].icell.PUM Vbias 0.0031f
C6219 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.SM 0.00168f
C6220 XThR.XTB3.Y data[4] 0.03253f
C6221 XThC.XTBN.Y XThC.Tn[12] 0.56523f
C6222 XThC.Tn[9] XThR.Tn[4] 0.28739f
C6223 XThC.XTB6.A a_6243_10571# 0.00295f
C6224 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04031f
C6225 XA.XIR[0].XIC[3].icell.SM VPWR 0.00158f
C6226 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C6227 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C6228 XThR.Tn[10] XA.XIR[11].XIC[12].icell.Ien 0.00338f
C6229 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02762f
C6230 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04031f
C6231 XA.XIR[3].XIC[12].icell.PDM Vbias 0.04261f
C6232 XA.XIR[1].XIC[1].icell.SM Vbias 0.00704f
C6233 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00584f
C6234 XA.XIR[8].XIC[14].icell.PDM Vbias 0.04261f
C6235 XA.XIR[14].XIC[5].icell.Ien Vbias 0.21098f
C6236 XA.XIR[3].XIC[13].icell.Ien VPWR 0.1903f
C6237 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10] 0.00341f
C6238 XA.XIR[15].XIC[13].icell.PDM Iout 0.00117f
C6239 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00256f
C6240 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PUM 0.00465f
C6241 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00584f
C6242 XA.XIR[1].XIC[11].icell.PDM Iout 0.00117f
C6243 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C6244 XA.XIR[13].XIC[7].icell.Ien Vbias 0.21098f
C6245 XA.XIR[3].XIC[9].icell.Ien Iout 0.06417f
C6246 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PUM 0.00465f
C6247 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[7].icell.Ien 0.00214f
C6248 XThC.Tn[0] XA.XIR[8].XIC_dummy_left.icell.Iout 0.00109f
C6249 XThC.Tn[13] XThR.Tn[10] 0.2874f
C6250 XA.XIR[8].XIC[9].icell.SM Vbias 0.00701f
C6251 XThC.Tn[3] XThR.Tn[0] 0.28743f
C6252 XA.XIR[7].XIC[6].icell.SM VPWR 0.00158f
C6253 XA.XIR[2].XIC[6].icell.Ien VPWR 0.1903f
C6254 a_n997_715# VPWR 0.02818f
C6255 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C6256 XA.XIR[11].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6257 XThC.Tn[5] XThR.Tn[5] 0.28739f
C6258 XA.XIR[12].XIC[9].icell.PUM Vbias 0.0031f
C6259 XA.XIR[2].XIC[2].icell.Ien Iout 0.06417f
C6260 XA.XIR[4].XIC[11].icell.PDM Iout 0.00117f
C6261 XA.XIR[7].XIC[2].icell.SM Iout 0.00388f
C6262 XA.XIR[1].XIC[8].icell.Ien VPWR 0.1903f
C6263 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.15202f
C6264 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6265 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00214f
C6266 XThC.Tn[6] XA.XIR[0].XIC[7].icell.Ien 0.002f
C6267 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.SM 0.0039f
C6268 XThC.Tn[10] XThC.Tn[12] 0.00453f
C6269 XThR.Tn[13] XA.XIR[14].XIC[12].icell.SM 0.00121f
C6270 XA.XIR[1].XIC[4].icell.Ien Iout 0.06417f
C6271 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.0404f
C6272 XA.XIR[13].XIC[14].icell.SM Iout 0.00388f
C6273 XA.XIR[14].XIC_15.icell.SM Vbias 0.00701f
C6274 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13] 0.00341f
C6275 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00214f
C6276 XThR.Tn[7] XA.XIR[8].XIC[3].icell.SM 0.00121f
C6277 XA.XIR[12].XIC_dummy_right.icell.SM VPWR 0.00123f
C6278 XThR.Tn[6] XA.XIR[7].XIC[14].icell.SM 0.00121f
C6279 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02762f
C6280 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00584f
C6281 XA.XIR[8].XIC[12].icell.Ien Iout 0.06417f
C6282 XThR.Tn[8] XA.XIR[9].XIC[12].icell.Ien 0.00338f
C6283 XA.XIR[0].XIC[11].icell.SM Vbias 0.00716f
C6284 XThR.XTBN.A XThR.Tn[13] 0.00106f
C6285 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C6286 XA.XIR[15].XIC[0].icell.PUM VPWR 0.00937f
C6287 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.SM 0.00168f
C6288 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.15202f
C6289 XThR.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.00341f
C6290 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PUM 0.00465f
C6291 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00214f
C6292 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02762f
C6293 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Ien 0.00584f
C6294 XThR.Tn[10] XA.XIR[11].XIC[4].icell.SM 0.00121f
C6295 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C6296 XThR.Tn[3] XA.XIR[3].XIC[5].icell.PDM 0.00341f
C6297 a_5949_9615# VPWR 0.7053f
C6298 XA.XIR[2].XIC[14].icell.Ien Vbias 0.21098f
C6299 XA.XIR[7].XIC[14].icell.SM Vbias 0.00701f
C6300 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.03425f
C6301 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.03425f
C6302 XThR.Tn[1] XA.XIR[2].XIC[5].icell.Ien 0.00338f
C6303 XA.XIR[6].XIC[1].icell.PDM VPWR 0.00799f
C6304 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C6305 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04031f
C6306 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.03554f
C6307 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PUM 0.00186f
C6308 XThR.XTB3.Y a_n997_2667# 0.002f
C6309 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C6310 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.15202f
C6311 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.15202f
C6312 XA.XIR[0].XIC[14].icell.Ien Iout 0.06389f
C6313 XA.XIR[14].XIC[0].icell.Ien Vbias 0.20951f
C6314 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C6315 XA.XIR[5].XIC[8].icell.PDM VPWR 0.00799f
C6316 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C6317 XA.XIR[4].XIC[2].icell.PUM Vbias 0.0031f
C6318 XThC.Tn[2] XThR.Tn[2] 0.28739f
C6319 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.SM 0.0039f
C6320 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.SM 0.0039f
C6321 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.SM 0.0039f
C6322 XThR.XTB6.A a_n1335_4229# 0.00304f
C6323 XThR.Tn[13] XA.XIR[14].XIC[9].icell.Ien 0.00338f
C6324 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C6325 XThR.Tn[13] Vbias 3.74874f
C6326 XA.XIR[13].XIC[2].icell.PDM VPWR 0.00799f
C6327 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00214f
C6328 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.03425f
C6329 XA.XIR[13].XIC[11].icell.Ien Iout 0.06417f
C6330 XThC.Tn[11] XThR.Tn[14] 0.28739f
C6331 XThR.Tn[3] VPWR 6.64542f
C6332 XThC.XTB5.A VPWR 0.82807f
C6333 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PUM 0.00465f
C6334 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C6335 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00584f
C6336 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C6337 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PUM 0.00465f
C6338 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C6339 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C6340 XA.XIR[12].XIC[7].icell.PDM VPWR 0.00799f
C6341 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00189f
C6342 XThR.Tn[0] XA.XIR[1].XIC[12].icell.Ien 0.00338f
C6343 XA.XIR[15].XIC[0].icell.SM Iout 0.00388f
C6344 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C6345 XThR.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.00338f
C6346 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.SM 0.0039f
C6347 XA.XIR[6].XIC[1].icell.SM Vbias 0.00701f
C6348 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C6349 XThR.XTB7.Y VPWR 1.14768f
C6350 XA.XIR[15].XIC[4].icell.PUM Vbias 0.0031f
C6351 VPWR data[4] 0.5303f
C6352 XA.XIR[5].XIC[4].icell.Ien Vbias 0.21098f
C6353 XA.XIR[11].XIC[1].icell.PDM Iout 0.00117f
C6354 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.SM 0.00168f
C6355 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Iout 0.00347f
C6356 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11107f
C6357 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.03425f
C6358 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C6359 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.SM 0.00168f
C6360 XThR.Tn[5] XA.XIR[6].XIC[14].icell.Ien 0.00338f
C6361 XA.XIR[4].XIC[7].icell.PUM Vbias 0.0031f
C6362 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.SM 0.0039f
C6363 XA.XIR[10].XIC[5].icell.PDM Iout 0.00117f
C6364 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C6365 XThR.XTB6.Y a_n997_1803# 0.00871f
C6366 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04031f
C6367 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C6368 XA.XIR[15].XIC_15.icell.Ien VPWR 0.36724f
C6369 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.SM 0.0039f
C6370 XA.XIR[10].XIC[12].icell.SM VPWR 0.00158f
C6371 XA.XIR[3].XIC[3].icell.SM VPWR 0.00158f
C6372 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.SM 0.00168f
C6373 XA.XIR[6].XIC[8].icell.Ien VPWR 0.1903f
C6374 XThR.Tn[13] XA.XIR[14].XIC[10].icell.SM 0.00121f
C6375 XA.XIR[6].XIC[4].icell.Ien Iout 0.06417f
C6376 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.03425f
C6377 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.SM 0.0039f
C6378 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.03425f
C6379 XA.XIR[5].XIC[11].icell.PUM VPWR 0.00937f
C6380 XThC.Tn[7] XThR.Tn[6] 0.28739f
C6381 XThC.XTBN.A XThC.Tn[9] 0.12399f
C6382 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7] 0.00341f
C6383 XThC.XTBN.Y a_10915_9569# 0.21503f
C6384 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.SM 0.0039f
C6385 XThR.Tn[10] XA.XIR[11].XIC[0].icell.Ien 0.00338f
C6386 XA.XIR[15].XIC[5].icell.SM Iout 0.00388f
C6387 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00584f
C6388 XA.XIR[4].XIC[12].icell.SM VPWR 0.00158f
C6389 XA.XIR[3].XIC[3].icell.PDM VPWR 0.00799f
C6390 XThR.XTBN.Y XA.XIR[13].XIC_dummy_left.icell.Iout 0.00446f
C6391 XThC.Tn[0] XThR.Tn[11] 0.28744f
C6392 XA.XIR[12].XIC[11].icell.PDM Iout 0.00117f
C6393 XA.XIR[9].XIC[14].icell.PDM Vbias 0.04261f
C6394 XA.XIR[8].XIC[5].icell.PDM VPWR 0.00799f
C6395 XA.XIR[14].XIC[2].icell.Ien VPWR 0.19084f
C6396 XA.XIR[7].XIC[1].icell.PUM Vbias 0.0031f
C6397 XA.XIR[0].XIC[6].icell.PDM Vbias 0.04282f
C6398 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00584f
C6399 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C6400 XA.XIR[4].XIC[8].icell.SM Iout 0.00388f
C6401 XThC.XTB7.A XThC.XTB7.B 0.35844f
C6402 XA.XIR[2].XIC[9].icell.PDM VPWR 0.00799f
C6403 XA.XIR[13].XIC[4].icell.Ien VPWR 0.1903f
C6404 XA.XIR[8].XIC[6].icell.SM VPWR 0.00158f
C6405 XA.XIR[9].XIC[10].icell.PUM Vbias 0.0031f
C6406 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C6407 XA.XIR[10].XIC[2].icell.SM Vbias 0.00701f
C6408 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.SM 0.00168f
C6409 XA.XIR[15].XIC[12].icell.PDM Iout 0.00117f
C6410 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00584f
C6411 XThC.Tn[7] Vbias 2.28836f
C6412 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12] 0.00341f
C6413 XA.XIR[12].XIC[6].icell.PUM VPWR 0.00937f
C6414 XA.XIR[8].XIC[2].icell.SM Iout 0.00388f
C6415 XA.XIR[0].XIC[3].icell.PUM Vbias 0.0031f
C6416 XThR.Tn[8] XA.XIR[9].XIC[2].icell.SM 0.00121f
C6417 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02762f
C6418 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.03425f
C6419 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C6420 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01577f
C6421 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C6422 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.SM 0.0039f
C6423 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04031f
C6424 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C6425 XA.XIR[11].XIC[7].icell.Ien VPWR 0.1903f
C6426 XA.XIR[3].XIC[11].icell.SM Vbias 0.00701f
C6427 XA.XIR[5].XIC_15.icell.SM VPWR 0.00275f
C6428 XThR.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.00338f
C6429 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PUM 0.00465f
C6430 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C6431 XThC.XTB6.Y XThC.Tn[5] 0.20189f
C6432 XA.XIR[11].XIC[3].icell.Ien Iout 0.06417f
C6433 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C6434 XA.XIR[10].XIC[9].icell.Ien VPWR 0.1903f
C6435 XThC.Tn[13] XThR.Tn[13] 0.2874f
C6436 XThR.Tn[3] XA.XIR[4].XIC[4].icell.Ien 0.00338f
C6437 XA.XIR[2].XIC[4].icell.SM Vbias 0.00701f
C6438 XA.XIR[9].XIC[11].icell.SM Iout 0.00388f
C6439 XA.XIR[14].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6440 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13] 0.00341f
C6441 XA.XIR[7].XIC[6].icell.PUM Vbias 0.0031f
C6442 XA.XIR[10].XIC[5].icell.Ien Iout 0.06417f
C6443 XThC.Tn[3] XThR.Tn[1] 0.28739f
C6444 XThR.Tn[9] XA.XIR[10].XIC[5].icell.Ien 0.00338f
C6445 XA.XIR[0].XIC[8].icell.SM VPWR 0.00158f
C6446 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.SM 0.00168f
C6447 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C6448 a_n997_2667# VPWR 0.01642f
C6449 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.SM 0.0039f
C6450 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.03425f
C6451 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6452 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C6453 XA.XIR[1].XIC[6].icell.SM Vbias 0.00704f
C6454 XA.XIR[0].XIC[4].icell.SM Iout 0.00367f
C6455 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04031f
C6456 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.SM 0.00168f
C6457 XThC.Tn[3] XThR.Tn[12] 0.28739f
C6458 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.03425f
C6459 XA.XIR[8].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6460 XThC.Tn[12] XThR.Tn[8] 0.28739f
C6461 XA.XIR[3].XIC[14].icell.Ien Iout 0.06417f
C6462 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38708f
C6463 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04031f
C6464 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8] 0.00341f
C6465 XA.XIR[2].XIC[11].icell.Ien VPWR 0.1903f
C6466 XA.XIR[8].XIC[14].icell.SM Vbias 0.00701f
C6467 XA.XIR[7].XIC[11].icell.SM VPWR 0.00158f
C6468 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PUM 0.00465f
C6469 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.SM 0.0039f
C6470 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.03425f
C6471 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.SM 0.0039f
C6472 XThC.XTBN.Y XThC.Tn[1] 0.7252f
C6473 XA.XIR[2].XIC[7].icell.Ien Iout 0.06417f
C6474 XA.XIR[10].XIC_15.icell.SM Iout 0.0047f
C6475 XThR.Tn[0] XA.XIR[1].XIC[2].icell.SM 0.00121f
C6476 XA.XIR[1].XIC[13].icell.Ien VPWR 0.1903f
C6477 XA.XIR[7].XIC[7].icell.SM Iout 0.00388f
C6478 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04031f
C6479 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.15202f
C6480 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.SM 0.00168f
C6481 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PUM 0.00465f
C6482 XThR.Tn[12] XA.XIR[13].XIC[3].icell.Ien 0.00338f
C6483 XThC.Tn[7] XThR.Tn[4] 0.28739f
C6484 a_n1049_7493# XA.XIR[1].XIC_dummy_left.icell.Iout 0.0013f
C6485 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C6486 XA.XIR[1].XIC[9].icell.Ien Iout 0.06417f
C6487 XThR.Tn[13] XA.XIR[14].XIC[14].icell.Ien 0.00338f
C6488 XA.XIR[10].XIC[10].icell.SM VPWR 0.00158f
C6489 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.04432f
C6490 XA.XIR[3].XIC[0].icell.SM VPWR 0.00158f
C6491 XThR.Tn[7] XA.XIR[8].XIC[8].icell.SM 0.00121f
C6492 XThC.XTB7.B a_5949_9615# 0.00927f
C6493 XThC.XTB4.Y XThC.Tn[5] 0.00814f
C6494 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C6495 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.SM 0.0039f
C6496 XThC.Tn[2] XThR.Tn[10] 0.28739f
C6497 XThR.Tn[11] XA.XIR[12].XIC[6].icell.Ien 0.00338f
C6498 a_3773_9615# Vbias 0.00846f
C6499 XThR.Tn[5] XA.XIR[6].XIC[4].icell.SM 0.00121f
C6500 XA.XIR[12].XIC[0].icell.Ien VPWR 0.1903f
C6501 XThC.XTB3.Y XThC.Tn[9] 0.00285f
C6502 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.SM 0.00168f
C6503 XThC.XTB6.Y a_10051_9569# 0.07626f
C6504 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PDM 0.00172f
C6505 XThR.Tn[10] XA.XIR[11].XIC_15.icell.Ien 0.00117f
C6506 XThR.Tn[11] VPWR 7.58404f
C6507 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.15202f
C6508 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.SM 0.0039f
C6509 XA.XIR[5].XIC[4].icell.PDM Vbias 0.04261f
C6510 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04031f
C6511 XA.XIR[7].XIC[9].icell.PDM VPWR 0.00799f
C6512 XA.XIR[9].XIC[2].icell.PUM VPWR 0.00937f
C6513 XThC.XTB5.A XThC.XTB7.B 0.30355f
C6514 XThR.XTB6.A a_n1319_5611# 0.00467f
C6515 XThR.Tn[1] XA.XIR[2].XIC[10].icell.Ien 0.00338f
C6516 XA.XIR[4].XIC[4].icell.PUM VPWR 0.00937f
C6517 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.SM 0.0039f
C6518 XA.XIR[15].XIC[7].icell.PDM VPWR 0.0114f
C6519 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6520 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.SM 0.0039f
C6521 XA.XIR[12].XIC[3].icell.PDM Vbias 0.04261f
C6522 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00214f
C6523 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.15202f
C6524 XA.XIR[6].XIC[4].icell.PDM Iout 0.00117f
C6525 XA.XIR[10].XIC[13].icell.PUM VPWR 0.00937f
C6526 XA.XIR[11].XIC[9].icell.PDM Vbias 0.04261f
C6527 XA.XIR[14].XIC[1].icell.PDM Iout 0.00117f
C6528 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00584f
C6529 XA.XIR[5].XIC[11].icell.PDM Iout 0.00117f
C6530 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C6531 a_8739_9569# VPWR 0.00583f
C6532 XA.XIR[9].XIC[5].icell.PDM VPWR 0.00799f
C6533 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00584f
C6534 XA.XIR[13].XIC[5].icell.PDM Iout 0.00117f
C6535 XThR.XTB7.A a_n1331_2891# 0.00995f
C6536 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C6537 XA.XIR[13].XIC[12].icell.SM VPWR 0.00158f
C6538 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00584f
C6539 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.SM 0.00168f
C6540 XA.XIR[3].XIC[3].icell.PUM Vbias 0.0031f
C6541 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.SM 0.00168f
C6542 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.03425f
C6543 XA.XIR[12].XIC[10].icell.PDM Iout 0.00117f
C6544 XA.XIR[6].XIC[6].icell.SM Vbias 0.00701f
C6545 XA.XIR[9].XIC[7].icell.PUM VPWR 0.00937f
C6546 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.SM 0.00168f
C6547 XA.XIR[15].XIC[9].icell.PUM Vbias 0.0031f
C6548 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.SM 0.0039f
C6549 XThR.XTBN.A a_n997_3979# 0.02087f
C6550 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.SM 0.0039f
C6551 XA.XIR[5].XIC[9].icell.Ien Vbias 0.21098f
C6552 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00584f
C6553 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.03425f
C6554 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C6555 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C6556 XA.XIR[15].XIC[11].icell.PDM Iout 0.00117f
C6557 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C6558 XThC.Tn[0] XThR.Tn[14] 0.28742f
C6559 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04031f
C6560 XA.XIR[4].XIC[12].icell.PUM Vbias 0.0031f
C6561 XThR.Tn[11] XA.XIR[12].XIC[0].icell.SM 0.00127f
C6562 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.SM 0.0039f
C6563 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02762f
C6564 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C6565 XA.XIR[3].XIC[8].icell.SM VPWR 0.00158f
C6566 XA.XIR[8].XIC[1].icell.PDM Vbias 0.04261f
C6567 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.SM 0.00168f
C6568 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.03425f
C6569 XA.XIR[1].XIC[10].icell.PDM VPWR 0.00799f
C6570 XA.XIR[6].XIC[13].icell.Ien VPWR 0.1903f
C6571 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PUM 0.00429f
C6572 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00214f
C6573 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14] 0.00341f
C6574 XA.XIR[2].XIC[5].icell.PDM Vbias 0.04261f
C6575 XA.XIR[10].XIC[14].icell.Ien VPWR 0.19036f
C6576 XA.XIR[3].XIC[4].icell.SM Iout 0.00388f
C6577 XA.XIR[15].XIC_dummy_right.icell.SM VPWR 0.00123f
C6578 XA.XIR[13].XIC[2].icell.SM Vbias 0.00701f
C6579 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.SM 0.00168f
C6580 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.SM 0.00168f
C6581 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[4].icell.SM 0.0039f
C6582 XA.XIR[4].XIC[10].icell.PDM VPWR 0.00799f
C6583 XA.XIR[2].XIC[1].icell.SM VPWR 0.00158f
C6584 XA.XIR[8].XIC[6].icell.PUM Vbias 0.0031f
C6585 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02762f
C6586 XA.XIR[6].XIC[9].icell.Ien Iout 0.06417f
C6587 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7] 0.00341f
C6588 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6589 XA.XIR[7].XIC[3].icell.PUM VPWR 0.00937f
C6590 XThR.XTB6.A XThR.Tn[5] 0.00361f
C6591 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04031f
C6592 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02762f
C6593 XThR.Tn[13] XA.XIR[14].XIC[12].icell.Ien 0.00338f
C6594 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.SM 0.00168f
C6595 XA.XIR[12].XIC[4].icell.Ien Vbias 0.21098f
C6596 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02762f
C6597 XA.XIR[1].XIC[3].icell.SM VPWR 0.00158f
C6598 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01577f
C6599 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00214f
C6600 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.SM 0.00168f
C6601 XA.XIR[14].XIC[7].icell.Ien VPWR 0.19084f
C6602 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13] 0.00341f
C6603 XA.XIR[11].XIC[5].icell.SM Vbias 0.00701f
C6604 XA.XIR[3].XIC[6].icell.PDM Iout 0.00117f
C6605 XA.XIR[4].XIC[13].icell.SM Iout 0.00388f
C6606 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6607 XA.XIR[14].XIC[3].icell.Ien Iout 0.06417f
C6608 XA.XIR[8].XIC[8].icell.PDM Iout 0.00117f
C6609 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.SM 0.00168f
C6610 XA.XIR[13].XIC[9].icell.Ien VPWR 0.1903f
C6611 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04031f
C6612 XA.XIR[8].XIC[11].icell.SM VPWR 0.00158f
C6613 XA.XIR[9].XIC_15.icell.PUM Vbias 0.0031f
C6614 XThC.Tn[11] VPWR 6.86576f
C6615 XA.XIR[10].XIC[7].icell.SM Vbias 0.00701f
C6616 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.03023f
C6617 XA.XIR[2].XIC[12].icell.PDM Iout 0.00117f
C6618 XA.XIR[13].XIC[5].icell.Ien Iout 0.06417f
C6619 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C6620 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00584f
C6621 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C6622 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00584f
C6623 XA.XIR[8].XIC[7].icell.SM Iout 0.00388f
C6624 XThR.Tn[8] XA.XIR[9].XIC[7].icell.SM 0.00121f
C6625 XA.XIR[0].XIC[8].icell.PUM Vbias 0.0031f
C6626 XThR.Tn[0] XA.XIR[0].XIC[9].icell.PDM 0.00341f
C6627 XThC.XTBN.A XThC.Tn[7] 0.01439f
C6628 XThR.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.00338f
C6629 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.15202f
C6630 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.SM 0.0039f
C6631 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.0404f
C6632 XThR.Tn[4] XA.XIR[5].XIC[9].icell.Ien 0.00338f
C6633 XThR.Tn[1] XA.XIR[1].XIC[7].icell.PDM 0.00341f
C6634 XA.XIR[11].XIC[8].icell.Ien Iout 0.06417f
C6635 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00214f
C6636 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04031f
C6637 XThR.XTBN.A XThR.Tn[7] 0.01439f
C6638 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PUM 0.00465f
C6639 XA.XIR[5].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6640 XThC.Tn[0] XA.XIR[2].XIC_dummy_left.icell.Iout 0.00109f
C6641 XThR.Tn[3] XA.XIR[4].XIC[9].icell.Ien 0.00338f
C6642 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00584f
C6643 XA.XIR[2].XIC[9].icell.SM Vbias 0.00701f
C6644 XThR.XTBN.A a_n997_2891# 0.01719f
C6645 XA.XIR[7].XIC[11].icell.PUM Vbias 0.0031f
C6646 XA.XIR[10].XIC[11].icell.PUM VPWR 0.00937f
C6647 XA.XIR[0].XIC[13].icell.SM VPWR 0.00158f
C6648 XA.XIR[13].XIC_15.icell.SM Iout 0.0047f
C6649 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5] 0.00341f
C6650 XA.XIR[1].XIC[11].icell.SM Vbias 0.00704f
C6651 XThR.Tn[6] XThR.Tn[7] 0.06617f
C6652 XA.XIR[0].XIC[9].icell.SM Iout 0.00367f
C6653 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00584f
C6654 XA.XIR[12].XIC_dummy_left.icell.SM VPWR 0.00269f
C6655 XThR.Tn[2] XA.XIR[2].XIC[4].icell.PDM 0.00341f
C6656 XA.XIR[13].XIC[10].icell.SM VPWR 0.00158f
C6657 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.03425f
C6658 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PUM 0.00465f
C6659 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04052f
C6660 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04031f
C6661 XThR.Tn[13] XA.XIR[14].XIC[4].icell.SM 0.00121f
C6662 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C6663 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[12].icell.Ien 0.00214f
C6664 data[6] data[7] 0.04128f
C6665 XA.XIR[8].XIC[1].icell.PUM Vbias 0.0031f
C6666 XThC.Tn[2] XThR.Tn[13] 0.28739f
C6667 XA.XIR[15].XIC[1].icell.PUM VPWR 0.00937f
C6668 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6] 0.00341f
C6669 XA.XIR[5].XIC[1].icell.Ien VPWR 0.1903f
C6670 XA.XIR[2].XIC[12].icell.Ien Iout 0.06417f
C6671 XA.XIR[7].XIC[12].icell.SM Iout 0.00388f
C6672 XThR.Tn[0] XA.XIR[1].XIC[7].icell.SM 0.00121f
C6673 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.SM 0.00168f
C6674 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.SM 0.00168f
C6675 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00214f
C6676 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.15202f
C6677 XThR.Tn[7] Vbias 3.74624f
C6678 XThR.Tn[14] VPWR 7.78627f
C6679 XThR.Tn[12] XA.XIR[13].XIC[8].icell.Ien 0.00338f
C6680 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.03425f
C6681 XA.XIR[11].XIC[0].icell.PDM VPWR 0.00799f
C6682 XA.XIR[1].XIC[14].icell.Ien Iout 0.06417f
C6683 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PUM 0.00102f
C6684 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.SM 0.0039f
C6685 XThC.Tn[5] Iout 0.83957f
C6686 XThC.Tn[5] XThR.Tn[9] 0.28739f
C6687 XA.XIR[7].XIC_15.icell.SM Vbias 0.00701f
C6688 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00584f
C6689 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.SM 0.00168f
C6690 VPWR data[0] 0.52929f
C6691 XThC.Tn[1] XThR.Tn[8] 0.28739f
C6692 XA.XIR[7].XIC[5].icell.PDM Vbias 0.04261f
C6693 XA.XIR[10].XIC[4].icell.PDM VPWR 0.00799f
C6694 XThR.Tn[7] XA.XIR[8].XIC[13].icell.SM 0.00121f
C6695 XThR.XTB2.Y a_n1335_8107# 0.01006f
C6696 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.SM 0.00168f
C6697 XA.XIR[10].XIC[12].icell.Ien VPWR 0.1903f
C6698 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C6699 XThR.Tn[5] XA.XIR[6].XIC[9].icell.SM 0.00121f
C6700 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.0353f
C6701 XA.XIR[4].XIC[2].icell.Ien Vbias 0.21098f
C6702 XA.XIR[6].XIC[12].icell.PDM Vbias 0.04261f
C6703 XA.XIR[15].XIC[3].icell.PDM Vbias 0.04261f
C6704 XThR.XTB6.Y a_n997_3979# 0.0046f
C6705 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02762f
C6706 XA.XIR[12].XIC[1].icell.Ien Iout 0.06417f
C6707 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.03425f
C6708 XA.XIR[6].XIC[3].icell.SM VPWR 0.00158f
C6709 XThR.Tn[13] XA.XIR[14].XIC[10].icell.Ien 0.00338f
C6710 VPWR bias[1] 1.23968f
C6711 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Ien 0.00232f
C6712 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00214f
C6713 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.15202f
C6714 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C6715 XA.XIR[14].XIC[9].icell.PDM Vbias 0.04261f
C6716 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C6717 XA.XIR[13].XIC[13].icell.PUM VPWR 0.00937f
C6718 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.SM 0.00168f
C6719 XA.XIR[15].XIC[6].icell.PUM VPWR 0.00937f
C6720 XA.XIR[5].XIC[6].icell.Ien VPWR 0.1903f
C6721 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PUM 0.00465f
C6722 XThC.XTB7.B a_8739_9569# 0.0168f
C6723 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.SM 0.00168f
C6724 XA.XIR[5].XIC[2].icell.Ien Iout 0.06417f
C6725 XThR.Tn[1] XA.XIR[2].XIC_15.icell.Ien 0.00117f
C6726 XA.XIR[7].XIC[12].icell.PDM Iout 0.00117f
C6727 XA.XIR[4].XIC[9].icell.PUM VPWR 0.00937f
C6728 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PUM 0.00465f
C6729 XA.XIR[9].XIC[1].icell.PDM Vbias 0.04261f
C6730 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.03425f
C6731 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.03425f
C6732 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00214f
C6733 XA.XIR[15].XIC[10].icell.PDM Iout 0.00117f
C6734 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00214f
C6735 XThC.XTB3.Y XThC.Tn[7] 0.00819f
C6736 XA.XIR[12].XIC[12].icell.SM Vbias 0.00701f
C6737 XA.XIR[9].XIC[5].icell.Ien Vbias 0.21098f
C6738 XA.XIR[8].XIC[3].icell.PUM VPWR 0.00937f
C6739 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.SM 0.0039f
C6740 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.15202f
C6741 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C6742 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00584f
C6743 XThC.Tn[4] XThC.Tn[5] 0.4169f
C6744 XThR.XTB2.Y a_n1049_7787# 0.2342f
C6745 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.1106f
C6746 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02762f
C6747 XA.XIR[0].XIC[12].icell.PDM VPWR 0.011f
C6748 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.SM 0.00168f
C6749 XA.XIR[11].XIC[2].icell.SM VPWR 0.00158f
C6750 XA.XIR[3].XIC[8].icell.PUM Vbias 0.0031f
C6751 XA.XIR[9].XIC[8].icell.PDM Iout 0.00117f
C6752 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9] 0.00341f
C6753 XA.XIR[1].XIC[6].icell.PDM Vbias 0.04261f
C6754 XA.XIR[6].XIC[11].icell.SM Vbias 0.00701f
C6755 XA.XIR[13].XIC[14].icell.Ien VPWR 0.19036f
C6756 XA.XIR[9].XIC[12].icell.PUM VPWR 0.00937f
C6757 XA.XIR[10].XIC[4].icell.SM VPWR 0.00158f
C6758 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.SM 0.0039f
C6759 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.03023f
C6760 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11] 0.00341f
C6761 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00584f
C6762 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02762f
C6763 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.15202f
C6764 XA.XIR[4].XIC[6].icell.PDM Vbias 0.04261f
C6765 XA.XIR[5].XIC[14].icell.Ien Vbias 0.21098f
C6766 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C6767 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C6768 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04031f
C6769 XA.XIR[0].XIC[5].icell.PUM VPWR 0.00877f
C6770 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Ien 0.00232f
C6771 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C6772 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C6773 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04031f
C6774 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.SM 0.0039f
C6775 XThR.XTB6.Y a_n997_2891# 0.00466f
C6776 XA.XIR[3].XIC[14].icell.PDM Vbias 0.04261f
C6777 XA.XIR[1].XIC[3].icell.PUM Vbias 0.0031f
C6778 XA.XIR[14].XIC[5].icell.SM Vbias 0.00701f
C6779 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C6780 XA.XIR[3].XIC[13].icell.SM VPWR 0.00158f
C6781 XThC.Tn[13] XThR.Tn[7] 0.2874f
C6782 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C6783 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.03425f
C6784 XA.XIR[12].XIC_15.icell.PUM Vbias 0.0031f
C6785 XA.XIR[3].XIC[9].icell.SM Iout 0.00388f
C6786 XA.XIR[1].XIC[13].icell.PDM Iout 0.00117f
C6787 XA.XIR[13].XIC[7].icell.SM Vbias 0.00701f
C6788 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.03425f
C6789 XThC.XTB7.B XThC.Tn[11] 0.03903f
C6790 XA.XIR[8].XIC[11].icell.PUM Vbias 0.0031f
C6791 XA.XIR[2].XIC[6].icell.SM VPWR 0.00158f
C6792 XA.XIR[6].XIC[14].icell.Ien Iout 0.06417f
C6793 XA.XIR[7].XIC[8].icell.PUM VPWR 0.00937f
C6794 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.SM 0.00168f
C6795 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.SM 0.00168f
C6796 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C6797 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.SM 0.0039f
C6798 XA.XIR[12].XIC[9].icell.Ien Vbias 0.21098f
C6799 XA.XIR[2].XIC[2].icell.SM Iout 0.00388f
C6800 XA.XIR[4].XIC[13].icell.PDM Iout 0.00117f
C6801 XA.XIR[1].XIC[8].icell.SM VPWR 0.00158f
C6802 XA.XIR[10].XIC[10].icell.Ien VPWR 0.1903f
C6803 XThR.Tn[1] XA.XIR[2].XIC[0].icell.SM 0.00121f
C6804 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.SM 0.00168f
C6805 XA.XIR[1].XIC[4].icell.SM Iout 0.00388f
C6806 XA.XIR[14].XIC[8].icell.Ien Iout 0.06417f
C6807 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C6808 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PUM 0.00465f
C6809 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00584f
C6810 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.SM 0.00168f
C6811 XThC.XTB3.Y a_3773_9615# 0.00124f
C6812 XA.XIR[9].XIC[0].icell.Ien Vbias 0.20951f
C6813 XThR.XTBN.A a_n997_1579# 0.00199f
C6814 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00584f
C6815 XA.XIR[13].XIC[11].icell.PUM VPWR 0.00937f
C6816 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.15202f
C6817 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.04036f
C6818 XA.XIR[8].XIC[12].icell.SM Iout 0.00388f
C6819 XThR.Tn[11] XA.XIR[12].XIC[1].icell.SM 0.00121f
C6820 a_3773_9615# XThC.Tn[2] 0.01175f
C6821 XThR.Tn[8] XA.XIR[9].XIC[12].icell.SM 0.00121f
C6822 XA.XIR[0].XIC[13].icell.PUM Vbias 0.0031f
C6823 XThR.Tn[2] XA.XIR[3].XIC[7].icell.Ien 0.00338f
C6824 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C6825 XThR.Tn[4] XA.XIR[5].XIC[14].icell.Ien 0.00338f
C6826 XThR.XTB3.Y VPWR 1.07975f
C6827 XA.XIR[8].XIC_15.icell.SM Vbias 0.00701f
C6828 XThR.Tn[4] XA.XIR[4].XIC[6].icell.PDM 0.00341f
C6829 XThC.Tn[12] XThR.Tn[3] 0.28739f
C6830 XThR.XTB5.A XThR.XTB6.A 1.80461f
C6831 XThR.Tn[3] XA.XIR[3].XIC[7].icell.PDM 0.00341f
C6832 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6833 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Ien 0.00728f
C6834 XThR.Tn[3] XA.XIR[4].XIC[14].icell.Ien 0.00338f
C6835 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PUM 0.00465f
C6836 XThC.Tn[0] VPWR 5.95931f
C6837 XA.XIR[7].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6838 XA.XIR[2].XIC[14].icell.SM Vbias 0.00701f
C6839 XThC.XTB1.Y XThC.Tn[7] 0.0045f
C6840 XThR.Tn[1] XA.XIR[2].XIC[5].icell.SM 0.00121f
C6841 XA.XIR[12].XIC[10].icell.SM Vbias 0.00701f
C6842 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.SM 0.00168f
C6843 XA.XIR[6].XIC[3].icell.PDM VPWR 0.00799f
C6844 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PDM 0.00172f
C6845 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.04036f
C6846 XA.XIR[5].XIC[1].icell.PUM Vbias 0.0031f
C6847 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.SM 0.0039f
C6848 XThR.Tn[13] XA.XIR[14].XIC_15.icell.Ien 0.00117f
C6849 XA.XIR[0].XIC[14].icell.SM Iout 0.00367f
C6850 XA.XIR[5].XIC[10].icell.PDM VPWR 0.00799f
C6851 XA.XIR[14].XIC[0].icell.PDM VPWR 0.00799f
C6852 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PUM 0.00465f
C6853 XThC.Tn[8] XThR.Tn[5] 0.28739f
C6854 XThC.XTB7.B data[0] 0.0138f
C6855 XA.XIR[13].XIC[4].icell.PDM VPWR 0.00799f
C6856 XA.XIR[13].XIC[12].icell.Ien VPWR 0.1903f
C6857 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02762f
C6858 XA.XIR[10].XIC[0].icell.PDM Vbias 0.04207f
C6859 XThC.XTB7.Y a_7875_9569# 0.00476f
C6860 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.03425f
C6861 XA.XIR[12].XIC[9].icell.PDM VPWR 0.00799f
C6862 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C6863 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.SM 0.00168f
C6864 XThR.Tn[0] XA.XIR[1].XIC[12].icell.SM 0.00121f
C6865 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C6866 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.03425f
C6867 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C6868 XA.XIR[9].XIC[2].icell.Ien VPWR 0.1903f
C6869 XA.XIR[6].XIC[3].icell.PUM Vbias 0.0031f
C6870 XA.XIR[15].XIC[4].icell.Ien Vbias 0.17899f
C6871 XA.XIR[11].XIC[3].icell.PDM Iout 0.00117f
C6872 XA.XIR[5].XIC[4].icell.SM Vbias 0.00701f
C6873 a_6243_9615# XThC.Tn[5] 0.00158f
C6874 XThR.Tn[5] a_n1049_5317# 0.00158f
C6875 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C6876 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00214f
C6877 XThR.XTB6.A data[5] 0.37233f
C6878 XA.XIR[12].XIC[13].icell.PUM Vbias 0.0031f
C6879 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.SM 0.0039f
C6880 XThR.Tn[5] XA.XIR[6].XIC[14].icell.SM 0.00121f
C6881 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PUM 0.00102f
C6882 XThR.Tn[6] XA.XIR[7].XIC[1].icell.Ien 0.00338f
C6883 XA.XIR[10].XIC[7].icell.PDM Iout 0.00117f
C6884 XA.XIR[4].XIC[7].icell.Ien Vbias 0.21098f
C6885 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04031f
C6886 XA.XIR[3].XIC[5].icell.PUM VPWR 0.00937f
C6887 XA.XIR[6].XIC[8].icell.SM VPWR 0.00158f
C6888 XA.XIR[6].XIC[4].icell.SM Iout 0.00388f
C6889 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PUM 0.00465f
C6890 XA.XIR[5].XIC[11].icell.Ien VPWR 0.1903f
C6891 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7] 0.00341f
C6892 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00584f
C6893 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PUM 0.00441f
C6894 XA.XIR[5].XIC[7].icell.Ien Iout 0.06417f
C6895 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.SM 0.0039f
C6896 XA.XIR[4].XIC[14].icell.PUM VPWR 0.00937f
C6897 XThR.Tn[14] XA.XIR[15].XIC[1].icell.Ien 0.00338f
C6898 XA.XIR[8].XIC[7].icell.PDM VPWR 0.00799f
C6899 XA.XIR[3].XIC[5].icell.PDM VPWR 0.00799f
C6900 XA.XIR[7].XIC[1].icell.Ien Vbias 0.21098f
C6901 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.SM 0.00168f
C6902 XA.XIR[14].XIC[2].icell.SM VPWR 0.00158f
C6903 XA.XIR[0].XIC[8].icell.PDM Vbias 0.04282f
C6904 XThC.XTB5.Y Vbias 0.01575f
C6905 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C6906 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00214f
C6907 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00214f
C6908 XA.XIR[2].XIC[11].icell.PDM VPWR 0.00799f
C6909 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04031f
C6910 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C6911 XA.XIR[13].XIC[4].icell.SM VPWR 0.00158f
C6912 XThC.Tn[14] XThR.Tn[2] 0.28745f
C6913 XA.XIR[9].XIC[10].icell.Ien Vbias 0.21098f
C6914 XA.XIR[8].XIC[8].icell.PUM VPWR 0.00937f
C6915 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PUM 0.00465f
C6916 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C6917 XA.XIR[10].XIC[4].icell.PUM Vbias 0.0031f
C6918 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00584f
C6919 XThR.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.00338f
C6920 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00214f
C6921 XA.XIR[12].XIC[6].icell.Ien VPWR 0.1903f
C6922 XA.XIR[12].XIC[14].icell.Ien Vbias 0.21098f
C6923 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12] 0.00341f
C6924 XA.XIR[0].XIC[3].icell.Ien Vbias 0.21128f
C6925 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.03425f
C6926 XA.XIR[10].XIC_15.icell.Ien VPWR 0.25566f
C6927 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.SM 0.00168f
C6928 XA.XIR[11].XIC[7].icell.SM VPWR 0.00158f
C6929 XThR.XTB6.Y a_n997_1579# 0.07626f
C6930 XA.XIR[12].XIC[2].icell.Ien Iout 0.06417f
C6931 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00214f
C6932 XA.XIR[3].XIC[13].icell.PUM Vbias 0.0031f
C6933 XThR.Tn[4] XA.XIR[5].XIC[4].icell.SM 0.00121f
C6934 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.03425f
C6935 XA.XIR[11].XIC[3].icell.SM Iout 0.00388f
C6936 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C6937 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.SM 0.00168f
C6938 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C6939 XThR.Tn[3] XA.XIR[4].XIC[4].icell.SM 0.00121f
C6940 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.15202f
C6941 XThR.Tn[14] XA.XIR[15].XIC[6].icell.Ien 0.00338f
C6942 XA.XIR[7].XIC[6].icell.Ien Vbias 0.21098f
C6943 XA.XIR[2].XIC[6].icell.PUM Vbias 0.0031f
C6944 XA.XIR[0].XIC[10].icell.PUM VPWR 0.00877f
C6945 XA.XIR[10].XIC[5].icell.SM Iout 0.00388f
C6946 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00214f
C6947 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C6948 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.SM 0.00168f
C6949 XThR.Tn[9] XA.XIR[10].XIC[5].icell.SM 0.00121f
C6950 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5] 0.00346f
C6951 XThC.XTBN.Y Vbias 0.16321f
C6952 XA.XIR[13].XIC[10].icell.Ien VPWR 0.1903f
C6953 XA.XIR[1].XIC[8].icell.PUM Vbias 0.0031f
C6954 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04031f
C6955 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04031f
C6956 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C6957 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C6958 XThC.Tn[10] XThR.Tn[6] 0.28739f
C6959 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PUM 0.00465f
C6960 XA.XIR[3].XIC[14].icell.SM Iout 0.00388f
C6961 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00584f
C6962 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04031f
C6963 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8] 0.00341f
C6964 XA.XIR[8].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6965 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[9].icell.SM 0.0039f
C6966 XA.XIR[7].XIC[13].icell.PUM VPWR 0.00937f
C6967 XA.XIR[2].XIC[11].icell.SM VPWR 0.00158f
C6968 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PUM 0.00465f
C6969 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C6970 XA.XIR[2].XIC[7].icell.SM Iout 0.00388f
C6971 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6972 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00214f
C6973 XThC.Tn[12] XThR.Tn[11] 0.28739f
C6974 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PUM 0.00179f
C6975 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.04036f
C6976 XA.XIR[1].XIC[13].icell.SM VPWR 0.00158f
C6977 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C6978 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.SM 0.0039f
C6979 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PUM 0.00465f
C6980 XA.XIR[12].XIC[11].icell.PUM Vbias 0.0031f
C6981 XThR.Tn[12] XA.XIR[13].XIC[3].icell.SM 0.00121f
C6982 XA.XIR[1].XIC[9].icell.SM Iout 0.00388f
C6983 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.SM 0.00168f
C6984 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04052f
C6985 XThC.Tn[2] XThR.Tn[7] 0.28739f
C6986 XThC.Tn[10] Vbias 2.36503f
C6987 XThR.XTB6.A XThR.Tn[9] 0.00838f
C6988 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.15202f
C6989 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.SM 0.00168f
C6990 XA.XIR[3].XIC[2].icell.PUM VPWR 0.00937f
C6991 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C6992 XThC.XTB7.B XThC.Tn[0] 0.00139f
C6993 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00214f
C6994 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C6995 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.15202f
C6996 XA.XIR[12].XIC[0].icell.SM VPWR 0.00158f
C6997 a_4861_9615# Vbias 0.00548f
C6998 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.SM 0.00168f
C6999 XThR.Tn[11] XA.XIR[12].XIC[6].icell.SM 0.00121f
C7000 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C7001 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00584f
C7002 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C7003 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00584f
C7004 XThC.XTB6.Y XThC.Tn[8] 0.02461f
C7005 XThC.XTB5.Y XThC.Tn[13] 0.00145f
C7006 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.03425f
C7007 XThR.Tn[2] XA.XIR[3].XIC[12].icell.Ien 0.00338f
C7008 XA.XIR[15].XIC[12].icell.SM Vbias 0.00701f
C7009 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04052f
C7010 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.SM 0.0039f
C7011 XThR.XTB7.A data[6] 0.00197f
C7012 XA.XIR[5].XIC[6].icell.PDM Vbias 0.04261f
C7013 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C7014 XThR.Tn[0] Iout 1.16239f
C7015 XA.XIR[5].XIC[1].icell.SM VPWR 0.00158f
C7016 XA.XIR[7].XIC[11].icell.PDM VPWR 0.00799f
C7017 XThR.XTB7.Y a_n1319_5317# 0.01283f
C7018 XThC.XTB6.A a_7875_9569# 0.00149f
C7019 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.15202f
C7020 XA.XIR[13].XIC[0].icell.PDM Vbias 0.04207f
C7021 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PUM 0.00465f
C7022 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02762f
C7023 XThR.Tn[1] XA.XIR[2].XIC[10].icell.SM 0.00121f
C7024 XA.XIR[4].XIC[4].icell.Ien VPWR 0.1903f
C7025 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C7026 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00214f
C7027 XA.XIR[15].XIC[9].icell.PDM VPWR 0.0114f
C7028 a_n1049_6699# XThR.Tn[4] 0.00158f
C7029 XA.XIR[12].XIC[5].icell.PDM Vbias 0.04261f
C7030 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02762f
C7031 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PUM 0.00465f
C7032 XA.XIR[12].XIC[12].icell.Ien Vbias 0.21098f
C7033 XA.XIR[6].XIC[6].icell.PDM Iout 0.00117f
C7034 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Ien 0.00553f
C7035 XA.XIR[5].XIC[13].icell.PDM Iout 0.00117f
C7036 XA.XIR[14].XIC[3].icell.PDM Iout 0.00117f
C7037 XThC.Tn[1] XThR.Tn[3] 0.28739f
C7038 a_9827_9569# VPWR 0.0017f
C7039 XA.XIR[9].XIC[7].icell.PDM VPWR 0.00799f
C7040 XA.XIR[8].XIC[1].icell.Ien Vbias 0.21098f
C7041 XThC.XTBN.Y XThC.Tn[13] 0.62331f
C7042 XA.XIR[13].XIC[7].icell.PDM Iout 0.00117f
C7043 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.SM 0.00168f
C7044 XThC.Tn[10] XThR.Tn[4] 0.28739f
C7045 XA.XIR[3].XIC[3].icell.Ien Vbias 0.21098f
C7046 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C7047 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00214f
C7048 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C7049 XA.XIR[15].XIC_15.icell.PUM Vbias 0.0031f
C7050 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00584f
C7051 XA.XIR[6].XIC[8].icell.PUM Vbias 0.0031f
C7052 XA.XIR[9].XIC[7].icell.Ien VPWR 0.1903f
C7053 XThC.XTB4.Y XThC.Tn[8] 0.01306f
C7054 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C7055 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00584f
C7056 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00584f
C7057 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C7058 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C7059 XA.XIR[15].XIC[9].icell.Ien Vbias 0.17899f
C7060 XThC.Tn[0] XA.XIR[5].XIC_dummy_left.icell.Iout 0.00109f
C7061 XA.XIR[9].XIC[3].icell.Ien Iout 0.06417f
C7062 XA.XIR[5].XIC[9].icell.SM Vbias 0.00701f
C7063 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.15202f
C7064 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C7065 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.SM 0.00168f
C7066 XThC.Tn[4] XThR.Tn[0] 0.28741f
C7067 XThC.Tn[14] XThR.Tn[10] 0.28745f
C7068 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02762f
C7069 XThC.Tn[6] XThR.Tn[5] 0.28739f
C7070 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04031f
C7071 XA.XIR[3].XIC[1].icell.PDM Vbias 0.04261f
C7072 XA.XIR[8].XIC[3].icell.PDM Vbias 0.04261f
C7073 XA.XIR[4].XIC[12].icell.Ien Vbias 0.21098f
C7074 XA.XIR[1].XIC[12].icell.PDM VPWR 0.008f
C7075 XA.XIR[3].XIC[10].icell.PUM VPWR 0.00937f
C7076 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00214f
C7077 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C7078 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C7079 XA.XIR[6].XIC[13].icell.SM VPWR 0.00158f
C7080 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.03504f
C7081 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14] 0.00341f
C7082 XA.XIR[2].XIC[7].icell.PDM Vbias 0.04261f
C7083 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C7084 XThC.Tn[11] XThC.Tn[12] 0.22144f
C7085 XA.XIR[13].XIC[4].icell.PUM Vbias 0.0031f
C7086 XA.XIR[1].XIC[0].icell.PDM Iout 0.00117f
C7087 XA.XIR[8].XIC[6].icell.Ien Vbias 0.21098f
C7088 XA.XIR[6].XIC[9].icell.SM Iout 0.00388f
C7089 XA.XIR[7].XIC[3].icell.Ien VPWR 0.1903f
C7090 XA.XIR[2].XIC[3].icell.PUM VPWR 0.00937f
C7091 XA.XIR[4].XIC[12].icell.PDM VPWR 0.00799f
C7092 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04031f
C7093 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C7094 XA.XIR[12].XIC[4].icell.SM Vbias 0.00701f
C7095 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C7096 XA.XIR[5].XIC[12].icell.Ien Iout 0.06417f
C7097 XThC.XTB7.B VPWR 1.32988f
C7098 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C7099 XA.XIR[1].XIC[5].icell.PUM VPWR 0.00937f
C7100 XA.XIR[4].XIC[0].icell.PDM Iout 0.00117f
C7101 XA.XIR[13].XIC_15.icell.Ien VPWR 0.25566f
C7102 XA.XIR[14].XIC[7].icell.SM VPWR 0.00158f
C7103 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C7104 XA.XIR[11].XIC[7].icell.PUM Vbias 0.0031f
C7105 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Iout 0.00347f
C7106 XA.XIR[3].XIC[8].icell.PDM Iout 0.00117f
C7107 bias[1] bias[0] 0.13857f
C7108 XA.XIR[8].XIC[10].icell.PDM Iout 0.00117f
C7109 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00584f
C7110 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04031f
C7111 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C7112 XA.XIR[14].XIC[3].icell.SM Iout 0.00388f
C7113 XA.XIR[9].XIC_15.icell.Ien Vbias 0.21234f
C7114 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00214f
C7115 XA.XIR[8].XIC[13].icell.PUM VPWR 0.00937f
C7116 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04031f
C7117 XA.XIR[10].XIC[9].icell.PUM Vbias 0.0031f
C7118 XA.XIR[15].XIC[10].icell.SM Vbias 0.00701f
C7119 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C7120 XThR.Tn[6] XA.XIR[7].XIC[11].icell.Ien 0.00338f
C7121 XA.XIR[2].XIC[14].icell.PDM Iout 0.00117f
C7122 XA.XIR[13].XIC[5].icell.SM Iout 0.00388f
C7123 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.SM 0.0039f
C7124 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.SM 0.00168f
C7125 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.03589f
C7126 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00584f
C7127 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C7128 XA.XIR[0].XIC[8].icell.Ien Vbias 0.2113f
C7129 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.15202f
C7130 XThR.XTBN.A XThR.Tn[8] 0.1369f
C7131 XThR.Tn[0] XA.XIR[0].XIC[11].icell.PDM 0.00341f
C7132 XA.XIR[12].XIC[7].icell.Ien Iout 0.06417f
C7133 XThR.Tn[2] XA.XIR[3].XIC[2].icell.SM 0.00121f
C7134 XA.XIR[10].XIC_dummy_right.icell.SM VPWR 0.00123f
C7135 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.SM 0.00168f
C7136 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02762f
C7137 XThR.Tn[4] XA.XIR[5].XIC[9].icell.SM 0.00121f
C7138 XThR.Tn[1] XA.XIR[1].XIC[9].icell.PDM 0.00341f
C7139 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.SM 0.00168f
C7140 XA.XIR[11].XIC[8].icell.SM Iout 0.00388f
C7141 XA.XIR[12].XIC[10].icell.Ien Vbias 0.21098f
C7142 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00584f
C7143 XThR.Tn[3] XA.XIR[4].XIC[9].icell.SM 0.00121f
C7144 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04031f
C7145 XThC.Tn[3] XThR.Tn[2] 0.28739f
C7146 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.15202f
C7147 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.04036f
C7148 XA.XIR[7].XIC[11].icell.Ien Vbias 0.21098f
C7149 XA.XIR[2].XIC[11].icell.PUM Vbias 0.0031f
C7150 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01499f
C7151 XThC.XTB7.Y a_6243_9615# 0.27822f
C7152 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PUM 0.00465f
C7153 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.15202f
C7154 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5] 0.00341f
C7155 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C7156 XThC.Tn[12] XThR.Tn[14] 0.28739f
C7157 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.04036f
C7158 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.15202f
C7159 XA.XIR[1].XIC[13].icell.PUM Vbias 0.0031f
C7160 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02762f
C7161 XThR.Tn[2] XA.XIR[2].XIC[6].icell.PDM 0.00341f
C7162 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C7163 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00214f
C7164 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.03425f
C7165 XA.XIR[15].XIC[13].icell.PUM Vbias 0.0031f
C7166 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04031f
C7167 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.SM 0.00168f
C7168 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Ien 0.00584f
C7169 XA.XIR[3].XIC[0].icell.Ien Vbias 0.20951f
C7170 XThR.XTB7.B data[6] 0.07481f
C7171 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.15202f
C7172 XThR.Tn[8] Vbias 3.74624f
C7173 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C7174 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00214f
C7175 XThC.XTB2.Y XThC.Tn[8] 0.00167f
C7176 XA.XIR[15].XIC[1].icell.Ien VPWR 0.32895f
C7177 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11117f
C7178 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6] 0.00341f
C7179 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PUM 0.00465f
C7180 XA.XIR[2].XIC[12].icell.SM Iout 0.00388f
C7181 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12] 0.00341f
C7182 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.03425f
C7183 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C7184 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C7185 XA.XIR[1].XIC[0].icell.Ien Iout 0.06411f
C7186 XThR.Tn[12] XA.XIR[13].XIC[8].icell.SM 0.00121f
C7187 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.SM 0.0039f
C7188 XA.XIR[11].XIC[2].icell.PDM VPWR 0.00799f
C7189 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Iout 0.00347f
C7190 XA.XIR[11].XIC[1].icell.Ien Vbias 0.21098f
C7191 XA.XIR[1].XIC[14].icell.SM Iout 0.00388f
C7192 XA.XIR[2].XIC_15.icell.SM Vbias 0.00701f
C7193 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C7194 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00584f
C7195 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PUM 0.00186f
C7196 XA.XIR[4].XIC[0].icell.Ien Iout 0.06411f
C7197 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PUM 0.00429f
C7198 XA.XIR[7].XIC[7].icell.PDM Vbias 0.04261f
C7199 XA.XIR[10].XIC[6].icell.PDM VPWR 0.00799f
C7200 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PUM 0.00179f
C7201 XThR.Tn[1] Iout 1.16236f
C7202 XA.XIR[9].XIC[0].icell.SM Vbias 0.00675f
C7203 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C7204 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00584f
C7205 XThC.XTBN.A XThC.Tn[10] 0.12148f
C7206 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02762f
C7207 XA.XIR[0].XIC_15.icell.SM Iout 0.00367f
C7208 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C7209 XA.XIR[15].XIC[5].icell.PDM Vbias 0.04261f
C7210 XA.XIR[6].XIC[14].icell.PDM Vbias 0.04261f
C7211 XA.XIR[4].XIC[2].icell.SM Vbias 0.00701f
C7212 XThC.Tn[1] XThR.Tn[11] 0.28739f
C7213 XThR.Tn[12] Iout 1.16233f
C7214 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02762f
C7215 XA.XIR[6].XIC[5].icell.PUM VPWR 0.00937f
C7216 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C7217 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C7218 XA.XIR[15].XIC[6].icell.Ien VPWR 0.32895f
C7219 XA.XIR[15].XIC[14].icell.Ien Vbias 0.17899f
C7220 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.03425f
C7221 XA.XIR[5].XIC[6].icell.SM VPWR 0.00158f
C7222 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Ien 0.00232f
C7223 XThC.XTB7.B a_9827_9569# 0.00228f
C7224 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.15202f
C7225 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00214f
C7226 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00584f
C7227 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.02762f
C7228 XA.XIR[15].XIC[2].icell.Ien Iout 0.06807f
C7229 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C7230 a_7651_9569# Vbias 0.00376f
C7231 XA.XIR[5].XIC[2].icell.SM Iout 0.00388f
C7232 XA.XIR[7].XIC[14].icell.PDM Iout 0.00117f
C7233 XA.XIR[9].XIC[3].icell.PDM Vbias 0.04261f
C7234 XA.XIR[4].XIC[9].icell.Ien VPWR 0.1903f
C7235 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C7236 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.03425f
C7237 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.SM 0.0039f
C7238 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18966f
C7239 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PUM 0.00465f
C7240 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C7241 XA.XIR[4].XIC[5].icell.Ien Iout 0.06417f
C7242 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.03425f
C7243 XA.XIR[9].XIC[5].icell.SM Vbias 0.00701f
C7244 XA.XIR[8].XIC[3].icell.Ien VPWR 0.1903f
C7245 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C7246 XThC.XTB6.Y XThC.Tn[6] 0.00689f
C7247 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C7248 XThR.Tn[6] XA.XIR[7].XIC[1].icell.SM 0.00121f
C7249 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02762f
C7250 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C7251 XA.XIR[12].XIC[1].icell.SM VPWR 0.00158f
C7252 XThC.Tn[14] XThR.Tn[13] 0.28745f
C7253 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02762f
C7254 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C7255 XA.XIR[0].XIC[14].icell.PDM VPWR 0.00783f
C7256 XThC.Tn[4] XThR.Tn[1] 0.2874f
C7257 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PUM 0.0047f
C7258 XA.XIR[11].XIC[4].icell.PUM VPWR 0.00937f
C7259 XThC.Tn[8] Iout 0.8379f
C7260 XA.XIR[9].XIC[10].icell.PDM Iout 0.00117f
C7261 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00214f
C7262 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.SM 0.0039f
C7263 XThC.Tn[8] XThR.Tn[9] 0.28739f
C7264 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9] 0.00341f
C7265 XA.XIR[3].XIC[8].icell.Ien Vbias 0.21098f
C7266 XA.XIR[1].XIC[8].icell.PDM Vbias 0.04261f
C7267 XA.XIR[9].XIC[12].icell.Ien VPWR 0.1903f
C7268 XA.XIR[6].XIC[13].icell.PUM Vbias 0.0031f
C7269 XA.XIR[10].XIC[6].icell.PUM VPWR 0.00937f
C7270 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C7271 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PUM 0.00465f
C7272 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11] 0.00341f
C7273 XThR.Tn[14] XA.XIR[15].XIC[1].icell.SM 0.00121f
C7274 XThC.Tn[13] XThR.Tn[8] 0.2874f
C7275 XThC.Tn[4] XThR.Tn[12] 0.28739f
C7276 XA.XIR[5].XIC[14].icell.SM Vbias 0.00701f
C7277 XA.XIR[7].XIC[1].icell.SM Vbias 0.00701f
C7278 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.15202f
C7279 XA.XIR[9].XIC[8].icell.Ien Iout 0.06417f
C7280 XA.XIR[4].XIC[8].icell.PDM Vbias 0.04261f
C7281 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.SM 0.00168f
C7282 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C7283 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18987f
C7284 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.SM 0.0039f
C7285 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00214f
C7286 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04031f
C7287 XThR.XTBN.A a_n997_3755# 0.01939f
C7288 XA.XIR[15].XIC[11].icell.PUM Vbias 0.0031f
C7289 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C7290 XA.XIR[1].XIC[3].icell.Ien Vbias 0.21104f
C7291 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01577f
C7292 XA.XIR[14].XIC[7].icell.PUM Vbias 0.0031f
C7293 XThC.XTBN.Y XThC.Tn[2] 0.64352f
C7294 XA.XIR[11].XIC[13].icell.SM Iout 0.00388f
C7295 XThR.XTB7.A XThR.Tn[5] 0.02751f
C7296 XA.XIR[12].XIC_15.icell.Ien Vbias 0.21234f
C7297 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Ien 0.00246f
C7298 XA.XIR[1].XIC_15.icell.PDM Iout 0.00133f
C7299 XA.XIR[13].XIC[9].icell.PUM Vbias 0.0031f
C7300 XA.XIR[2].XIC[8].icell.PUM VPWR 0.00937f
C7301 XA.XIR[6].XIC[14].icell.SM Iout 0.00388f
C7302 XA.XIR[8].XIC[11].icell.Ien Vbias 0.21098f
C7303 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00214f
C7304 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C7305 XA.XIR[7].XIC[8].icell.Ien VPWR 0.1903f
C7306 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C7307 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C7308 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00584f
C7309 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C7310 XThC.Tn[0] XA.XIR[12].XIC_dummy_left.icell.Iout 0.00109f
C7311 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00584f
C7312 data[2] data[3] 0.04128f
C7313 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.SM 0.0039f
C7314 XThC.XTB4.Y XThC.Tn[6] 0.00608f
C7315 XA.XIR[4].XIC_15.icell.PDM Iout 0.00133f
C7316 XA.XIR[0].XIC[0].icell.PUM VPWR 0.00877f
C7317 XA.XIR[7].XIC[4].icell.Ien Iout 0.06417f
C7318 XA.XIR[1].XIC[10].icell.PUM VPWR 0.00937f
C7319 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00214f
C7320 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04031f
C7321 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02762f
C7322 XThC.Tn[3] XThR.Tn[10] 0.28739f
C7323 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.04036f
C7324 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02762f
C7325 XThC.XTB3.Y XThC.Tn[10] 0.29462f
C7326 XA.XIR[13].XIC_dummy_right.icell.SM VPWR 0.00123f
C7327 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.PDM 0.00591f
C7328 XA.XIR[14].XIC[8].icell.SM Iout 0.00388f
C7329 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.03425f
C7330 XThR.Tn[7] XA.XIR[8].XIC[5].icell.Ien 0.00338f
C7331 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.SM 0.0039f
C7332 XThC.XTB3.Y a_4861_9615# 0.0093f
C7333 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00584f
C7334 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PUM 0.00465f
C7335 XThC.XTB6.A data[1] 0.37233f
C7336 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00214f
C7337 a_n1049_5611# XThR.Tn[6] 0.00158f
C7338 XA.XIR[15].XIC[12].icell.Ien Vbias 0.17899f
C7339 XA.XIR[0].XIC[13].icell.Ien Vbias 0.2113f
C7340 XThR.Tn[12] XA.XIR[13].XIC[13].icell.SM 0.00121f
C7341 XA.XIR[3].XIC_15.icell.SM Iout 0.0047f
C7342 a_n1049_8581# VPWR 0.71705f
C7343 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00584f
C7344 XThR.Tn[2] XA.XIR[3].XIC[7].icell.SM 0.00121f
C7345 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.SM 0.00168f
C7346 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.SM 0.0039f
C7347 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00214f
C7348 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C7349 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.15202f
C7350 XThR.Tn[4] XA.XIR[4].XIC[8].icell.PDM 0.00341f
C7351 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04031f
C7352 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C7353 XThR.Tn[4] XA.XIR[5].XIC[14].icell.SM 0.00121f
C7354 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12] 0.00341f
C7355 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.03425f
C7356 XA.XIR[10].XIC[0].icell.Ien VPWR 0.1903f
C7357 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C7358 XThR.Tn[3] XA.XIR[3].XIC[9].icell.PDM 0.00341f
C7359 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C7360 XThR.Tn[10] XA.XIR[11].XIC[6].icell.Ien 0.00338f
C7361 XThR.Tn[3] XA.XIR[4].XIC[14].icell.SM 0.00121f
C7362 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C7363 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.03425f
C7364 XA.XIR[2].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7365 XA.XIR[6].XIC[5].icell.PDM VPWR 0.00799f
C7366 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.15202f
C7367 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00214f
C7368 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C7369 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.15202f
C7370 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PDM 0.00172f
C7371 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.03425f
C7372 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.SM 0.00168f
C7373 VPWR bias[0] 1.93694f
C7374 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.SM 0.00168f
C7375 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C7376 XA.XIR[14].XIC[2].icell.PDM VPWR 0.00799f
C7377 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.15202f
C7378 XA.XIR[5].XIC[12].icell.PDM VPWR 0.00799f
C7379 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C7380 XA.XIR[14].XIC[1].icell.Ien Vbias 0.21098f
C7381 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PUM 0.00465f
C7382 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PUM 0.00465f
C7383 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.03425f
C7384 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00584f
C7385 XThR.XTB4.Y data[6] 0.0086f
C7386 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C7387 XA.XIR[13].XIC[6].icell.PDM VPWR 0.00799f
C7388 XA.XIR[5].XIC[0].icell.PDM Iout 0.00117f
C7389 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC[14].icell.SM 0.0039f
C7390 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.15202f
C7391 XA.XIR[10].XIC[2].icell.PDM Vbias 0.04261f
C7392 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00584f
C7393 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PUM 0.00465f
C7394 XThC.XTB7.Y a_8963_9569# 0.00474f
C7395 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.03425f
C7396 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00214f
C7397 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C7398 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C7399 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02762f
C7400 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.SM 0.0039f
C7401 XThC.Tn[1] XThR.Tn[14] 0.28739f
C7402 XA.XIR[9].XIC[2].icell.SM VPWR 0.00158f
C7403 XA.XIR[6].XIC[3].icell.Ien Vbias 0.21098f
C7404 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01432f
C7405 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C7406 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02893f
C7407 XA.XIR[0].XIC_dummy_left.icell.SM VPWR 0.00269f
C7408 XThR.XTB2.Y a_n1049_7493# 0.02133f
C7409 XA.XIR[15].XIC[4].icell.SM Vbias 0.00701f
C7410 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00214f
C7411 XThR.Tn[7] XA.XIR[8].XIC[0].icell.Ien 0.00338f
C7412 XA.XIR[11].XIC[5].icell.PDM Iout 0.00117f
C7413 XA.XIR[5].XIC[6].icell.PUM Vbias 0.0031f
C7414 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.SM 0.00168f
C7415 XA.XIR[11].XIC[11].icell.SM Iout 0.00388f
C7416 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C7417 XA.XIR[10].XIC[9].icell.PDM Iout 0.00117f
C7418 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C7419 XA.XIR[3].XIC[5].icell.Ien VPWR 0.1903f
C7420 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04031f
C7421 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.11103f
C7422 XA.XIR[4].XIC[7].icell.SM Vbias 0.00701f
C7423 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00584f
C7424 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.SM 0.00168f
C7425 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.03425f
C7426 XA.XIR[6].XIC[10].icell.PUM VPWR 0.00937f
C7427 XThR.XTB6.Y a_n997_3755# 0.0046f
C7428 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C7429 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00584f
C7430 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00214f
C7431 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.03425f
C7432 XA.XIR[8].XIC[1].icell.SM Vbias 0.00701f
C7433 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[3].icell.Ien 0.00214f
C7434 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02762f
C7435 XA.XIR[5].XIC[11].icell.SM VPWR 0.00158f
C7436 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7] 0.00341f
C7437 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C7438 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C7439 XThR.Tn[10] XA.XIR[11].XIC[0].icell.SM 0.00121f
C7440 XA.XIR[15].XIC[7].icell.Ien Iout 0.06807f
C7441 XThC.Tn[12] VPWR 6.85795f
C7442 XA.XIR[3].XIC[7].icell.PDM VPWR 0.00799f
C7443 XA.XIR[5].XIC[7].icell.SM Iout 0.00388f
C7444 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C7445 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.03549f
C7446 XA.XIR[4].XIC[14].icell.Ien VPWR 0.19036f
C7447 XA.XIR[8].XIC[9].icell.PDM VPWR 0.00799f
C7448 XA.XIR[14].XIC[4].icell.PUM VPWR 0.00937f
C7449 XA.XIR[2].XIC[1].icell.Ien Vbias 0.21098f
C7450 XA.XIR[0].XIC[10].icell.PDM Vbias 0.04282f
C7451 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C7452 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00584f
C7453 XA.XIR[11].XIC[2].icell.Ien Vbias 0.21098f
C7454 XA.XIR[4].XIC[10].icell.Ien Iout 0.06417f
C7455 XA.XIR[2].XIC[13].icell.PDM VPWR 0.00799f
C7456 XA.XIR[15].XIC[10].icell.Ien Vbias 0.17899f
C7457 XThC.XTBN.A a_7651_9569# 0.02087f
C7458 XA.XIR[13].XIC[6].icell.PUM VPWR 0.00937f
C7459 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04031f
C7460 XA.XIR[9].XIC[10].icell.SM Vbias 0.00701f
C7461 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.SM 0.0039f
C7462 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.03426f
C7463 XA.XIR[10].XIC[4].icell.Ien Vbias 0.21098f
C7464 XThC.XTB7.A Vbias 0.0149f
C7465 XA.XIR[8].XIC[8].icell.Ien VPWR 0.1903f
C7466 XA.XIR[0].XIC[1].icell.Ien Iout 0.06389f
C7467 XThR.Tn[12] XA.XIR[13].XIC[11].icell.SM 0.00121f
C7468 XThR.Tn[6] XA.XIR[7].XIC[6].icell.SM 0.00121f
C7469 XA.XIR[2].XIC[1].icell.PDM Iout 0.00117f
C7470 a_n1049_7787# XThR.XTB3.Y 0.00124f
C7471 XA.XIR[12].XIC[6].icell.SM VPWR 0.00158f
C7472 XA.XIR[8].XIC[4].icell.Ien Iout 0.06417f
C7473 XThR.XTB6.Y a_n1049_5611# 0.26831f
C7474 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12] 0.00341f
C7475 XThR.XTB7.B XThR.Tn[5] 0.00705f
C7476 XThR.Tn[8] XA.XIR[9].XIC[4].icell.Ien 0.00338f
C7477 XA.XIR[0].XIC[3].icell.SM Vbias 0.00716f
C7478 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C7479 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07214f
C7480 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C7481 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C7482 XA.XIR[11].XIC[9].icell.PUM VPWR 0.00937f
C7483 XA.XIR[12].XIC[2].icell.SM Iout 0.00388f
C7484 XA.XIR[3].XIC[13].icell.Ien Vbias 0.21098f
C7485 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00214f
C7486 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.38919f
C7487 XA.XIR[14].XIC[13].icell.SM Iout 0.00388f
C7488 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04031f
C7489 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.PDM 0.00586f
C7490 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00584f
C7491 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C7492 XThR.Tn[14] XA.XIR[15].XIC[6].icell.SM 0.00121f
C7493 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00584f
C7494 XA.XIR[9].XIC[13].icell.Ien Iout 0.06417f
C7495 XA.XIR[7].XIC[6].icell.SM Vbias 0.00701f
C7496 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.15202f
C7497 XA.XIR[2].XIC[6].icell.Ien Vbias 0.21098f
C7498 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18966f
C7499 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C7500 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5] 0.00341f
C7501 XThC.Tn[3] XThR.Tn[13] 0.28739f
C7502 XA.XIR[9].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7503 XA.XIR[1].XIC[8].icell.Ien Vbias 0.21104f
C7504 XA.XIR[0].XIC[6].icell.Ien Iout 0.06389f
C7505 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04031f
C7506 XThR.Tn[5] XA.XIR[6].XIC[1].icell.Ien 0.00338f
C7507 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.03425f
C7508 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.SM 0.0039f
C7509 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04031f
C7510 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8] 0.00341f
C7511 XA.XIR[2].XIC[13].icell.PUM VPWR 0.00937f
C7512 XThC.Tn[6] Iout 0.83892f
C7513 XThC.Tn[6] XThR.Tn[9] 0.28739f
C7514 XA.XIR[7].XIC[13].icell.Ien VPWR 0.1903f
C7515 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12] 0.00341f
C7516 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02762f
C7517 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.15202f
C7518 XThC.Tn[2] XThR.Tn[8] 0.28739f
C7519 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6] 0.00341f
C7520 XA.XIR[10].XIC_dummy_left.icell.SM VPWR 0.00269f
C7521 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01577f
C7522 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.SM 0.0039f
C7523 XA.XIR[7].XIC[9].icell.Ien Iout 0.06417f
C7524 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PDM 0.00172f
C7525 XThR.Tn[0] XA.XIR[1].XIC[4].icell.Ien 0.00338f
C7526 XA.XIR[11].XIC[9].icell.SM Iout 0.00388f
C7527 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.SM 0.00168f
C7528 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.03425f
C7529 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C7530 XA.XIR[13].XIC[0].icell.Ien VPWR 0.1903f
C7531 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C7532 XThR.Tn[7] XA.XIR[8].XIC[10].icell.Ien 0.00338f
C7533 XThC.XTBN.Y a_2979_9615# 0.0607f
C7534 XA.XIR[12].XIC[2].icell.PUM VPWR 0.00937f
C7535 a_5949_9615# Vbias 0.00634f
C7536 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C7537 XThR.Tn[5] XA.XIR[6].XIC[6].icell.Ien 0.00338f
C7538 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00584f
C7539 XA.XIR[6].XIC[1].icell.PDM Vbias 0.04261f
C7540 XThR.XTBN.A data[4] 0.02581f
C7541 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.SM 0.00168f
C7542 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C7543 XThR.Tn[2] XA.XIR[3].XIC[12].icell.SM 0.00121f
C7544 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Iout 0.00347f
C7545 XA.XIR[2].XIC[0].icell.Ien Iout 0.06411f
C7546 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.15202f
C7547 XThR.XTB5.A XThR.XTB7.A 0.07862f
C7548 XA.XIR[5].XIC[8].icell.PDM Vbias 0.04261f
C7549 XA.XIR[15].XIC[1].icell.SM VPWR 0.00158f
C7550 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00214f
C7551 XA.XIR[7].XIC[13].icell.PDM VPWR 0.00799f
C7552 XA.XIR[5].XIC[3].icell.PUM VPWR 0.00937f
C7553 a_9827_9569# XThC.Tn[12] 0.19481f
C7554 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C7555 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00584f
C7556 XThC.XTB3.Y a_7651_9569# 0.00604f
C7557 XThC.Tn[0] XThC.Tn[1] 1.15401f
C7558 XA.XIR[13].XIC[2].icell.PDM Vbias 0.04261f
C7559 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.03425f
C7560 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PUM 0.00465f
C7561 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.SM 0.00168f
C7562 XA.XIR[10].XIC[1].icell.Ien Iout 0.06417f
C7563 XA.XIR[7].XIC[1].icell.PDM Iout 0.00117f
C7564 XThC.XTB5.A Vbias 0.00557f
C7565 XA.XIR[4].XIC[4].icell.SM VPWR 0.00158f
C7566 XThR.Tn[12] XA.XIR[13].XIC[9].icell.SM 0.00121f
C7567 XThR.Tn[3] Vbias 3.74868f
C7568 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.15202f
C7569 XThR.Tn[9] XA.XIR[10].XIC[1].icell.Ien 0.00338f
C7570 XA.XIR[12].XIC[7].icell.PDM Vbias 0.04261f
C7571 XA.XIR[1].XIC_15.icell.SM Iout 0.0047f
C7572 XThC.Tn[4] XThC.Tn[6] 0.00202f
C7573 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.03425f
C7574 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.15202f
C7575 XA.XIR[6].XIC[8].icell.PDM Iout 0.00117f
C7576 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PUM 0.00429f
C7577 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PUM 0.00465f
C7578 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Ien 0.00232f
C7579 a_n1049_7787# VPWR 0.72173f
C7580 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00214f
C7581 XA.XIR[5].XIC_15.icell.PDM Iout 0.00133f
C7582 XA.XIR[14].XIC[5].icell.PDM Iout 0.00117f
C7583 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.SM 0.00168f
C7584 XA.XIR[14].XIC[11].icell.SM Iout 0.00388f
C7585 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C7586 a_10915_9569# VPWR 0.00307f
C7587 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PUM 0.00465f
C7588 XA.XIR[9].XIC[9].icell.PDM VPWR 0.00799f
C7589 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.SM 0.0039f
C7590 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02762f
C7591 XA.XIR[0].XIC[1].icell.PDM VPWR 0.00774f
C7592 XA.XIR[13].XIC[9].icell.PDM Iout 0.00117f
C7593 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C7594 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00584f
C7595 XA.XIR[10].XIC[12].icell.SM Vbias 0.00701f
C7596 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.SM 0.0039f
C7597 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.SM 0.00168f
C7598 XA.XIR[15].XIC_15.icell.Ien Vbias 0.17891f
C7599 XA.XIR[3].XIC[3].icell.SM Vbias 0.00701f
C7600 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C7601 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.SM 0.00168f
C7602 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.03425f
C7603 XA.XIR[6].XIC[8].icell.Ien Vbias 0.21098f
C7604 XA.XIR[9].XIC[7].icell.SM VPWR 0.00158f
C7605 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02762f
C7606 XThC.Tn[14] XThR.Tn[7] 0.28745f
C7607 XThC.XTB5.A a_7331_10587# 0.01243f
C7608 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.SM 0.00168f
C7609 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C7610 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00256f
C7611 XThC.Tn[0] XA.XIR[15].XIC_dummy_left.icell.Iout 0.00109f
C7612 XThR.XTB7.A data[5] 0.06538f
C7613 XA.XIR[9].XIC[3].icell.SM Iout 0.00388f
C7614 XA.XIR[5].XIC[11].icell.PUM Vbias 0.0031f
C7615 XThC.XTB7.B XThC.Tn[12] 0.00772f
C7616 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.SM 0.0039f
C7617 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C7618 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04031f
C7619 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PUM 0.00465f
C7620 XThR.XTBN.Y XThR.Tn[5] 0.59912f
C7621 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00214f
C7622 XA.XIR[4].XIC[12].icell.SM Vbias 0.00701f
C7623 XA.XIR[3].XIC[3].icell.PDM Vbias 0.04261f
C7624 a_n1319_5317# VPWR 0.00672f
C7625 XA.XIR[8].XIC[5].icell.PDM Vbias 0.04261f
C7626 XA.XIR[11].XIC[13].icell.Ien Iout 0.06417f
C7627 XA.XIR[3].XIC[10].icell.Ien VPWR 0.1903f
C7628 XA.XIR[14].XIC[2].icell.Ien Vbias 0.21098f
C7629 XA.XIR[1].XIC[14].icell.PDM VPWR 0.00809f
C7630 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10] 0.00341f
C7631 XA.XIR[10].XIC[14].icell.PDM VPWR 0.00809f
C7632 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C7633 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01577f
C7634 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14] 0.00341f
C7635 XThR.XTBN.A a_n997_2667# 0.01679f
C7636 XA.XIR[2].XIC[9].icell.PDM Vbias 0.04261f
C7637 XA.XIR[3].XIC[6].icell.Ien Iout 0.06417f
C7638 XThR.Tn[3] XThR.Tn[4] 0.06967f
C7639 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.SM 0.00168f
C7640 XA.XIR[1].XIC[2].icell.PDM Iout 0.00117f
C7641 XA.XIR[13].XIC[4].icell.Ien Vbias 0.21098f
C7642 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02762f
C7643 XA.XIR[2].XIC[3].icell.Ien VPWR 0.1903f
C7644 XA.XIR[4].XIC[14].icell.PDM VPWR 0.00809f
C7645 XA.XIR[8].XIC[6].icell.SM Vbias 0.00701f
C7646 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C7647 XA.XIR[7].XIC[3].icell.SM VPWR 0.00158f
C7648 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04031f
C7649 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00214f
C7650 XA.XIR[12].XIC[6].icell.PUM Vbias 0.0031f
C7651 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07214f
C7652 XA.XIR[1].XIC[5].icell.Ien VPWR 0.1903f
C7653 XA.XIR[5].XIC[12].icell.SM Iout 0.00388f
C7654 XA.XIR[4].XIC[2].icell.PDM Iout 0.00117f
C7655 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00256f
C7656 XA.XIR[14].XIC[9].icell.PUM VPWR 0.00937f
C7657 XA.XIR[10].XIC_15.icell.PUM Vbias 0.0031f
C7658 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.SM 0.00168f
C7659 XA.XIR[11].XIC[7].icell.Ien Vbias 0.21098f
C7660 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.SM 0.0039f
C7661 XA.XIR[4].XIC_15.icell.Ien Iout 0.0642f
C7662 XA.XIR[3].XIC[10].icell.PDM Iout 0.00117f
C7663 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.SM 0.00168f
C7664 XA.XIR[8].XIC[12].icell.PDM Iout 0.00117f
C7665 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Ien 0.00584f
C7666 XA.XIR[5].XIC_15.icell.SM Vbias 0.00701f
C7667 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.04036f
C7668 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00214f
C7669 XA.XIR[10].XIC[9].icell.Ien Vbias 0.21098f
C7670 XA.XIR[8].XIC[13].icell.Ien VPWR 0.1903f
C7671 XThR.XTB4.Y XThR.Tn[5] 0.00751f
C7672 XThR.Tn[6] XA.XIR[7].XIC[11].icell.SM 0.00121f
C7673 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C7674 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.SM 0.0039f
C7675 XThC.Tn[13] XThR.Tn[3] 0.2874f
C7676 XThR.Tn[12] XA.XIR[13].XIC[13].icell.Ien 0.00338f
C7677 XA.XIR[8].XIC[9].icell.Ien Iout 0.06417f
C7678 XA.XIR[0].XIC[8].icell.SM Vbias 0.00716f
C7679 XThC.XTB7.A XThC.XTBN.A 0.197f
C7680 XThR.Tn[8] XA.XIR[9].XIC[9].icell.Ien 0.00338f
C7681 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02762f
C7682 XThC.XTB1.Y a_7651_9569# 0.06353f
C7683 XThR.Tn[0] XA.XIR[0].XIC[13].icell.PDM 0.00341f
C7684 XA.XIR[12].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7685 XThC.Tn[1] VPWR 5.91915f
C7686 XA.XIR[11].XIC[14].icell.SM Iout 0.00388f
C7687 XA.XIR[12].XIC[7].icell.SM Iout 0.00388f
C7688 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12] 0.00341f
C7689 XA.XIR[1].XIC[0].icell.PUM VPWR 0.00937f
C7690 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.SM 0.00168f
C7691 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.SM 0.0039f
C7692 XA.XIR[6].XIC_15.icell.SM Iout 0.0047f
C7693 XThR.Tn[1] XA.XIR[1].XIC[11].icell.PDM 0.00341f
C7694 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02762f
C7695 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C7696 XA.XIR[4].XIC[0].icell.PUM VPWR 0.00937f
C7697 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04031f
C7698 XThR.Tn[10] XA.XIR[11].XIC[1].icell.SM 0.00121f
C7699 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C7700 XA.XIR[15].XIC_dummy_left.icell.Ien Vbias 0.00329f
C7701 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02762f
C7702 XThR.XTBN.A XThR.Tn[11] 0.11968f
C7703 XThC.Tn[9] XThR.Tn[5] 0.28739f
C7704 XA.XIR[7].XIC[11].icell.SM Vbias 0.00701f
C7705 XA.XIR[2].XIC[11].icell.Ien Vbias 0.21098f
C7706 XA.XIR[13].XIC_dummy_left.icell.SM VPWR 0.00269f
C7707 XA.XIR[0].XIC_15.icell.Ien VPWR 0.2554f
C7708 XThR.Tn[1] XA.XIR[2].XIC[2].icell.Ien 0.00338f
C7709 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.03425f
C7710 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.SM 0.0039f
C7711 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02834f
C7712 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04031f
C7713 XA.XIR[1].XIC[13].icell.Ien Vbias 0.21104f
C7714 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00214f
C7715 XA.XIR[14].XIC[9].icell.SM Iout 0.00388f
C7716 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.15202f
C7717 XA.XIR[0].XIC[11].icell.Ien Iout 0.06389f
C7718 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.15202f
C7719 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.15202f
C7720 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02762f
C7721 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C7722 XThR.Tn[2] XA.XIR[2].XIC[8].icell.PDM 0.00341f
C7723 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00584f
C7724 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C7725 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C7726 XThR.Tn[13] XA.XIR[14].XIC[6].icell.Ien 0.00338f
C7727 XA.XIR[10].XIC[10].icell.SM Vbias 0.00701f
C7728 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04031f
C7729 XA.XIR[6].XIC[0].icell.Ien VPWR 0.1903f
C7730 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PUM 0.00465f
C7731 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C7732 XThR.XTB5.A XThR.XTB7.B 0.30355f
C7733 XA.XIR[3].XIC[0].icell.SM Vbias 0.00675f
C7734 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.SM 0.0039f
C7735 a_n1319_6405# VPWR 0.00676f
C7736 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00584f
C7737 XThR.Tn[12] XA.XIR[13].XIC[14].icell.SM 0.00121f
C7738 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.25759f
C7739 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.15202f
C7740 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.SM 0.00168f
C7741 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02762f
C7742 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00214f
C7743 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00584f
C7744 XA.XIR[12].XIC[0].icell.Ien Vbias 0.20951f
C7745 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.03425f
C7746 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PUM 0.00465f
C7747 XA.XIR[7].XIC[14].icell.Ien Iout 0.06417f
C7748 a_6243_9615# XThC.Tn[6] 0.26142f
C7749 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.SM 0.00168f
C7750 XThR.Tn[0] XA.XIR[1].XIC[9].icell.Ien 0.00338f
C7751 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.SM 0.00168f
C7752 XA.XIR[11].XIC[4].icell.PDM VPWR 0.00799f
C7753 XThR.Tn[11] Vbias 3.74874f
C7754 XA.XIR[11].XIC[11].icell.Ien Iout 0.06417f
C7755 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.SM 0.00168f
C7756 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.SM 0.0039f
C7757 XA.XIR[4].XIC[0].icell.SM Iout 0.00388f
C7758 XThR.Tn[7] XA.XIR[8].XIC_15.icell.Ien 0.00117f
C7759 XA.XIR[10].XIC[8].icell.PDM VPWR 0.00799f
C7760 XA.XIR[7].XIC[9].icell.PDM Vbias 0.04261f
C7761 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00584f
C7762 XA.XIR[9].XIC[2].icell.PUM Vbias 0.0031f
C7763 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C7764 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00214f
C7765 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C7766 XA.XIR[13].XIC[1].icell.Ien Iout 0.06417f
C7767 XThR.Tn[5] XA.XIR[6].XIC[11].icell.Ien 0.00338f
C7768 XA.XIR[15].XIC[7].icell.PDM Vbias 0.04261f
C7769 XA.XIR[4].XIC[4].icell.PUM Vbias 0.0031f
C7770 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C7771 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00214f
C7772 XA.XIR[6].XIC[5].icell.Ien VPWR 0.1903f
C7773 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00584f
C7774 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.SM 0.00168f
C7775 XA.XIR[10].XIC[13].icell.PUM Vbias 0.0031f
C7776 XA.XIR[15].XIC[6].icell.SM VPWR 0.00158f
C7777 XA.XIR[5].XIC[8].icell.PUM VPWR 0.00937f
C7778 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02762f
C7779 XThR.XTB6.Y a_n997_2667# 0.00468f
C7780 XA.XIR[15].XIC[2].icell.SM Iout 0.00388f
C7781 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PUM 0.00465f
C7782 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02762f
C7783 a_8739_9569# Vbias 0.00278f
C7784 XA.XIR[9].XIC[5].icell.PDM Vbias 0.04261f
C7785 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00214f
C7786 XA.XIR[4].XIC[9].icell.SM VPWR 0.00158f
C7787 XThR.XTB7.B data[5] 0.00593f
C7788 XA.XIR[13].XIC[12].icell.SM Vbias 0.00701f
C7789 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02762f
C7790 XA.XIR[0].XIC[0].icell.SM VPWR 0.00158f
C7791 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.03425f
C7792 XThR.Tn[12] XA.XIR[13].XIC[11].icell.Ien 0.00338f
C7793 XThC.XTB5.A XThC.XTBN.A 0.06305f
C7794 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02762f
C7795 XA.XIR[2].XIC[0].icell.PDM VPWR 0.00799f
C7796 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.03425f
C7797 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.15202f
C7798 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.SM 0.0039f
C7799 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C7800 XA.XIR[4].XIC[5].icell.SM Iout 0.00388f
C7801 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C7802 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02762f
C7803 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00584f
C7804 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC[0].icell.Ien 0.00214f
C7805 XA.XIR[9].XIC[7].icell.PUM Vbias 0.0031f
C7806 XA.XIR[8].XIC[3].icell.SM VPWR 0.00158f
C7807 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Iout 0.00401f
C7808 XA.XIR[10].XIC[13].icell.PDM VPWR 0.00799f
C7809 XThC.XTB7.A XThC.Tn[2] 0.12602f
C7810 XThR.Tn[13] XA.XIR[14].XIC[0].icell.SM 0.00127f
C7811 XA.XIR[12].XIC[3].icell.PUM VPWR 0.00937f
C7812 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00584f
C7813 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C7814 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00584f
C7815 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.SM 0.00168f
C7816 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.SM 0.00168f
C7817 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C7818 XA.XIR[14].XIC[13].icell.Ien Iout 0.06417f
C7819 XA.XIR[11].XIC[4].icell.Ien VPWR 0.1903f
C7820 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.03425f
C7821 XA.XIR[9].XIC[12].icell.PDM Iout 0.00117f
C7822 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04037f
C7823 XA.XIR[3].XIC[8].icell.SM Vbias 0.00701f
C7824 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.SM 0.0039f
C7825 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.SM 0.0039f
C7826 XA.XIR[13].XIC[14].icell.PDM VPWR 0.00809f
C7827 XA.XIR[1].XIC[10].icell.PDM Vbias 0.04261f
C7828 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9] 0.00341f
C7829 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02762f
C7830 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00214f
C7831 XA.XIR[6].XIC[13].icell.Ien Vbias 0.21098f
C7832 XA.XIR[9].XIC[12].icell.SM VPWR 0.00158f
C7833 XA.XIR[10].XIC[14].icell.Ien Vbias 0.21098f
C7834 XA.XIR[10].XIC[6].icell.Ien VPWR 0.1903f
C7835 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11] 0.00341f
C7836 XThC.Tn[11] XThR.Tn[6] 0.28739f
C7837 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.15202f
C7838 XA.XIR[1].XIC[1].icell.Ien Iout 0.06417f
C7839 XA.XIR[9].XIC[8].icell.SM Iout 0.00388f
C7840 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00214f
C7841 XA.XIR[2].XIC[1].icell.SM Vbias 0.00701f
C7842 XA.XIR[10].XIC[2].icell.Ien Iout 0.06417f
C7843 XA.XIR[7].XIC[3].icell.PUM Vbias 0.0031f
C7844 XA.XIR[5].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7845 XA.XIR[4].XIC[10].icell.PDM Vbias 0.04261f
C7846 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00584f
C7847 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C7848 XThR.Tn[9] XA.XIR[10].XIC[2].icell.Ien 0.00338f
C7849 XA.XIR[0].XIC[5].icell.SM VPWR 0.00158f
C7850 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C7851 XThR.Tn[7] XA.XIR[8].XIC[0].icell.SM 0.00121f
C7852 XA.XIR[13].XIC_15.icell.PUM Vbias 0.0031f
C7853 XA.XIR[1].XIC[3].icell.SM Vbias 0.00704f
C7854 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00584f
C7855 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C7856 XA.XIR[0].XIC[1].icell.SM Iout 0.00367f
C7857 XA.XIR[3].XIC_15.icell.Ien VPWR 0.25566f
C7858 XA.XIR[14].XIC[7].icell.Ien Vbias 0.21098f
C7859 XThC.Tn[13] XThR.Tn[11] 0.2874f
C7860 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PUM 0.00465f
C7861 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C7862 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00584f
C7863 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12] 0.00341f
C7864 XA.XIR[13].XIC[9].icell.Ien Vbias 0.21098f
C7865 XA.XIR[3].XIC[11].icell.Ien Iout 0.06417f
C7866 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39036f
C7867 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8] 0.00341f
C7868 XA.XIR[2].XIC[8].icell.Ien VPWR 0.1903f
C7869 XA.XIR[8].XIC[11].icell.SM Vbias 0.00701f
C7870 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[8].icell.Ien 0.00214f
C7871 XThC.Tn[3] XThR.Tn[7] 0.28739f
C7872 XThC.Tn[11] Vbias 2.46509f
C7873 XA.XIR[7].XIC[8].icell.SM VPWR 0.00158f
C7874 XThC.XTB7.B XThC.Tn[1] 0.0014f
C7875 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C7876 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.3891f
C7877 XA.XIR[2].XIC[4].icell.Ien Iout 0.06417f
C7878 XA.XIR[14].XIC[14].icell.SM Iout 0.00388f
C7879 XA.XIR[7].XIC[4].icell.SM Iout 0.00388f
C7880 XA.XIR[1].XIC[10].icell.Ien VPWR 0.1903f
C7881 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.15202f
C7882 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04031f
C7883 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00214f
C7884 XA.XIR[1].XIC[6].icell.Ien Iout 0.06417f
C7885 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C7886 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PUM 0.00465f
C7887 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C7888 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02762f
C7889 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00214f
C7890 XThR.Tn[7] XA.XIR[8].XIC[5].icell.SM 0.00121f
C7891 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C7892 XThC.XTB3.Y a_5949_9615# 0.009f
C7893 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02809f
C7894 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.03425f
C7895 XThR.Tn[5] XA.XIR[6].XIC[1].icell.SM 0.00121f
C7896 XA.XIR[10].XIC[11].icell.PUM Vbias 0.0031f
C7897 XA.XIR[8].XIC[14].icell.Ien Iout 0.06417f
C7898 XThR.XTB5.A XThR.XTBN.Y 0.00282f
C7899 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.SM 0.0039f
C7900 XA.XIR[6].XIC_dummy_left.icell.SM VPWR 0.00269f
C7901 XThR.Tn[11] XA.XIR[12].XIC[3].icell.Ien 0.00338f
C7902 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PUM 0.00465f
C7903 XThR.Tn[8] XA.XIR[9].XIC[14].icell.Ien 0.00338f
C7904 XA.XIR[0].XIC[13].icell.SM Vbias 0.00716f
C7905 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.03425f
C7906 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C7907 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02762f
C7908 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C7909 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.15202f
C7910 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00214f
C7911 XThR.Tn[4] XA.XIR[4].XIC[10].icell.PDM 0.00341f
C7912 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04031f
C7913 XA.XIR[13].XIC[10].icell.SM Vbias 0.00701f
C7914 XThR.XTB7.B XThR.Tn[9] 0.0565f
C7915 XThR.Tn[10] XA.XIR[11].XIC[6].icell.SM 0.00121f
C7916 XA.XIR[10].XIC[0].icell.SM VPWR 0.00158f
C7917 XA.XIR[7].XIC[0].icell.PDM VPWR 0.00799f
C7918 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00584f
C7919 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.SM 0.0039f
C7920 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C7921 XThR.Tn[3] XA.XIR[3].XIC[11].icell.PDM 0.00341f
C7922 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C7923 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02762f
C7924 XA.XIR[6].XIC[7].icell.PDM VPWR 0.00799f
C7925 XThR.Tn[1] XA.XIR[2].XIC[7].icell.Ien 0.00338f
C7926 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.SM 0.00168f
C7927 XA.XIR[15].XIC[1].icell.PUM Vbias 0.0031f
C7928 XThC.Tn[2] XThR.Tn[3] 0.28739f
C7929 XA.XIR[5].XIC[1].icell.Ien Vbias 0.21098f
C7930 XA.XIR[0].XIC_dummy_right.icell.SM VPWR 0.00123f
C7931 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.15202f
C7932 XThC.XTBN.Y XThC.Tn[14] 0.50214f
C7933 XThR.Tn[14] Vbias 3.74893f
C7934 XA.XIR[5].XIC[14].icell.PDM VPWR 0.00809f
C7935 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.15202f
C7936 XA.XIR[14].XIC[4].icell.PDM VPWR 0.00799f
C7937 XThC.Tn[11] XThR.Tn[4] 0.28739f
C7938 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.03425f
C7939 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.03425f
C7940 XA.XIR[14].XIC[11].icell.Ien Iout 0.06417f
C7941 XA.XIR[11].XIC[0].icell.PDM Vbias 0.04207f
C7942 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.SM 0.0039f
C7943 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C7944 XA.XIR[5].XIC[2].icell.PDM Iout 0.00117f
C7945 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C7946 XA.XIR[13].XIC[8].icell.PDM VPWR 0.00799f
C7947 XA.XIR[10].XIC[4].icell.PDM Vbias 0.04261f
C7948 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C7949 Vbias data[0] 0.00282f
C7950 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PUM 0.00429f
C7951 XA.XIR[10].XIC[12].icell.Ien Vbias 0.21098f
C7952 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00584f
C7953 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.03023f
C7954 XThC.XTB7.Y a_10051_9569# 0.013f
C7955 XA.XIR[6].XIC[1].icell.Ien Iout 0.06417f
C7956 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.SM 0.00168f
C7957 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PUM 0.00465f
C7958 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.15202f
C7959 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.SM 0.00168f
C7960 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C7961 XThR.Tn[0] XA.XIR[1].XIC[14].icell.Ien 0.00338f
C7962 XThC.Tn[5] XThR.Tn[0] 0.28744f
C7963 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.15202f
C7964 XA.XIR[12].XIC[1].icell.PDM Iout 0.00117f
C7965 XThC.Tn[7] XThR.Tn[5] 0.28739f
C7966 XA.XIR[6].XIC[3].icell.SM Vbias 0.00701f
C7967 XA.XIR[9].XIC[4].icell.PUM VPWR 0.00937f
C7968 bias[1] Vbias 0.04991f
C7969 XA.XIR[13].XIC[13].icell.PUM Vbias 0.0031f
C7970 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PUM 0.00465f
C7971 XThR.Tn[2] Iout 1.16236f
C7972 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.SM 0.00168f
C7973 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.SM 0.00168f
C7974 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C7975 XThC.Tn[11] XThC.Tn[13] 0.00226f
C7976 XA.XIR[15].XIC[6].icell.PUM Vbias 0.0031f
C7977 XA.XIR[11].XIC[7].icell.PDM Iout 0.00117f
C7978 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.SM 0.0039f
C7979 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C7980 XA.XIR[5].XIC[6].icell.Ien Vbias 0.21098f
C7981 XA.XIR[11].XIC[12].icell.SM VPWR 0.00158f
C7982 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02762f
C7983 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.SM 0.0039f
C7984 XA.XIR[10].XIC[12].icell.PDM VPWR 0.00799f
C7985 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C7986 XA.XIR[4].XIC[9].icell.PUM Vbias 0.0031f
C7987 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00584f
C7988 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02762f
C7989 XA.XIR[3].XIC[5].icell.SM VPWR 0.00158f
C7990 XA.XIR[1].XIC[1].icell.PDM VPWR 0.00799f
C7991 data[7] VGND 0.49949f
C7992 data[6] VGND 0.47974f
C7993 data[4] VGND 0.59317f
C7994 data[5] VGND 1.17814f
C7995 Iout VGND 0.32054p
C7996 data[3] VGND 0.49912f
C7997 data[2] VGND 0.48064f
C7998 data[0] VGND 0.59421f
C7999 data[1] VGND 1.17844f
C8000 bias[2] VGND 0.77552f
C8001 bias[0] VGND 1.22004f
C8002 Vbias VGND 0.23111p
C8003 bias[1] VGND 0.62458f
C8004 VPWR VGND 0.34079p
C8005 a_n997_715# VGND 0.5638f
C8006 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.75246f
C8007 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C8008 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64516f
C8009 XA.XIR[15].XIC_15.icell.SM VGND 0.00474f
C8010 XA.XIR[15].XIC_dummy_right.icell.PUM VGND 0.00215f
C8011 XA.XIR[15].XIC_15.icell.Ien VGND 0.44292f
C8012 XA.XIR[15].XIC[14].icell.SM VGND 0.00502f
C8013 XA.XIR[15].XIC_15.icell.PUM VGND 0.00282f
C8014 XA.XIR[15].XIC[14].icell.Ien VGND 0.44322f
C8015 XA.XIR[15].XIC[13].icell.SM VGND 0.00502f
C8016 XA.XIR[15].XIC[14].icell.PUM VGND 0.00293f
C8017 XA.XIR[15].XIC[13].icell.Ien VGND 0.44322f
C8018 XA.XIR[15].XIC[12].icell.SM VGND 0.00502f
C8019 XA.XIR[15].XIC[13].icell.PUM VGND 0.00293f
C8020 XA.XIR[15].XIC[12].icell.Ien VGND 0.44322f
C8021 XA.XIR[15].XIC[11].icell.SM VGND 0.00502f
C8022 XA.XIR[15].XIC[12].icell.PUM VGND 0.00293f
C8023 XA.XIR[15].XIC[11].icell.Ien VGND 0.44322f
C8024 XA.XIR[15].XIC[10].icell.SM VGND 0.00502f
C8025 XA.XIR[15].XIC[11].icell.PUM VGND 0.00293f
C8026 XA.XIR[15].XIC[10].icell.Ien VGND 0.44322f
C8027 XA.XIR[15].XIC[9].icell.SM VGND 0.00502f
C8028 XA.XIR[15].XIC[10].icell.PUM VGND 0.00293f
C8029 XA.XIR[15].XIC[9].icell.Ien VGND 0.44322f
C8030 XA.XIR[15].XIC[8].icell.SM VGND 0.00502f
C8031 XA.XIR[15].XIC[9].icell.PUM VGND 0.00293f
C8032 XA.XIR[15].XIC[8].icell.Ien VGND 0.44322f
C8033 XA.XIR[15].XIC[7].icell.SM VGND 0.00502f
C8034 XA.XIR[15].XIC[8].icell.PUM VGND 0.00293f
C8035 XA.XIR[15].XIC[7].icell.Ien VGND 0.44322f
C8036 XA.XIR[15].XIC[6].icell.SM VGND 0.00502f
C8037 XA.XIR[15].XIC[7].icell.PUM VGND 0.00293f
C8038 XA.XIR[15].XIC[6].icell.Ien VGND 0.44322f
C8039 XA.XIR[15].XIC[5].icell.SM VGND 0.00502f
C8040 XA.XIR[15].XIC[6].icell.PUM VGND 0.00293f
C8041 XA.XIR[15].XIC[5].icell.Ien VGND 0.44322f
C8042 XA.XIR[15].XIC[4].icell.SM VGND 0.00502f
C8043 XA.XIR[15].XIC[5].icell.PUM VGND 0.00293f
C8044 XA.XIR[15].XIC[4].icell.Ien VGND 0.44322f
C8045 XA.XIR[15].XIC[3].icell.SM VGND 0.00502f
C8046 XA.XIR[15].XIC[4].icell.PUM VGND 0.00293f
C8047 XA.XIR[15].XIC[3].icell.Ien VGND 0.44322f
C8048 XA.XIR[15].XIC[2].icell.SM VGND 0.00502f
C8049 XA.XIR[15].XIC[3].icell.PUM VGND 0.00293f
C8050 XA.XIR[15].XIC[2].icell.Ien VGND 0.44322f
C8051 XA.XIR[15].XIC[1].icell.SM VGND 0.00502f
C8052 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70718f
C8053 XA.XIR[15].XIC[2].icell.PUM VGND 0.00293f
C8054 XA.XIR[15].XIC[1].icell.Ien VGND 0.44322f
C8055 XA.XIR[15].XIC[0].icell.SM VGND 0.00502f
C8056 XA.XIR[15].XIC[1].icell.PUM VGND 0.00293f
C8057 XA.XIR[15].XIC[0].icell.Ien VGND 0.44356f
C8058 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01044f
C8059 XA.XIR[15].XIC[0].icell.PUM VGND 0.00516f
C8060 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.61163f
C8061 XA.XIR[15].XIC_dummy_left.icell.PUM VGND 0.00215f
C8062 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23279f
C8063 XA.XIR[15].XIC_15.icell.PDM VGND 0.18779f
C8064 XA.XIR[15].XIC[14].icell.PDM VGND 0.18733f
C8065 XA.XIR[15].XIC[13].icell.PDM VGND 0.18733f
C8066 XA.XIR[15].XIC[12].icell.PDM VGND 0.18733f
C8067 XA.XIR[15].XIC[11].icell.PDM VGND 0.18733f
C8068 XA.XIR[15].XIC[10].icell.PDM VGND 0.18733f
C8069 XA.XIR[15].XIC[9].icell.PDM VGND 0.18733f
C8070 XA.XIR[15].XIC[8].icell.PDM VGND 0.18733f
C8071 XA.XIR[15].XIC[7].icell.PDM VGND 0.18733f
C8072 XA.XIR[15].XIC[6].icell.PDM VGND 0.18733f
C8073 XA.XIR[15].XIC[5].icell.PDM VGND 0.18733f
C8074 XA.XIR[15].XIC[4].icell.PDM VGND 0.18733f
C8075 XA.XIR[15].XIC[3].icell.PDM VGND 0.18733f
C8076 XA.XIR[15].XIC[2].icell.PDM VGND 0.18733f
C8077 XA.XIR[15].XIC[1].icell.PDM VGND 0.18733f
C8078 XA.XIR[15].XIC[0].icell.PDM VGND 0.18741f
C8079 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C8080 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85795f
C8081 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C8082 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60802f
C8083 XA.XIR[14].XIC_15.icell.SM VGND 0.00474f
C8084 XA.XIR[14].XIC_dummy_right.icell.PUM VGND 0.00215f
C8085 XA.XIR[14].XIC_15.icell.Ien VGND 0.37063f
C8086 XA.XIR[14].XIC[14].icell.SM VGND 0.00502f
C8087 XA.XIR[14].XIC_15.icell.PUM VGND 0.00282f
C8088 XA.XIR[14].XIC[14].icell.Ien VGND 0.37144f
C8089 XA.XIR[14].XIC[13].icell.SM VGND 0.00502f
C8090 XA.XIR[14].XIC[14].icell.PUM VGND 0.00293f
C8091 XA.XIR[14].XIC[13].icell.Ien VGND 0.37144f
C8092 XA.XIR[14].XIC[12].icell.SM VGND 0.00502f
C8093 XA.XIR[14].XIC[13].icell.PUM VGND 0.00293f
C8094 XA.XIR[14].XIC[12].icell.Ien VGND 0.37144f
C8095 XA.XIR[14].XIC[11].icell.SM VGND 0.00502f
C8096 XA.XIR[14].XIC[12].icell.PUM VGND 0.00293f
C8097 XA.XIR[14].XIC[11].icell.Ien VGND 0.37144f
C8098 XA.XIR[14].XIC[10].icell.SM VGND 0.00502f
C8099 XA.XIR[14].XIC[11].icell.PUM VGND 0.00293f
C8100 XA.XIR[14].XIC[10].icell.Ien VGND 0.37144f
C8101 XA.XIR[14].XIC[9].icell.SM VGND 0.00502f
C8102 XA.XIR[14].XIC[10].icell.PUM VGND 0.00293f
C8103 XA.XIR[14].XIC[9].icell.Ien VGND 0.37144f
C8104 XA.XIR[14].XIC[8].icell.SM VGND 0.00502f
C8105 XA.XIR[14].XIC[9].icell.PUM VGND 0.00293f
C8106 XA.XIR[14].XIC[8].icell.Ien VGND 0.37144f
C8107 XA.XIR[14].XIC[7].icell.SM VGND 0.00502f
C8108 XA.XIR[14].XIC[8].icell.PUM VGND 0.00293f
C8109 XA.XIR[14].XIC[7].icell.Ien VGND 0.37144f
C8110 XA.XIR[14].XIC[6].icell.SM VGND 0.00502f
C8111 XA.XIR[14].XIC[7].icell.PUM VGND 0.00293f
C8112 XA.XIR[14].XIC[6].icell.Ien VGND 0.37144f
C8113 XA.XIR[14].XIC[5].icell.SM VGND 0.00502f
C8114 XA.XIR[14].XIC[6].icell.PUM VGND 0.00293f
C8115 XA.XIR[14].XIC[5].icell.Ien VGND 0.37144f
C8116 XA.XIR[14].XIC[4].icell.SM VGND 0.00502f
C8117 XA.XIR[14].XIC[5].icell.PUM VGND 0.00293f
C8118 XA.XIR[14].XIC[4].icell.Ien VGND 0.37144f
C8119 XA.XIR[14].XIC[3].icell.SM VGND 0.00502f
C8120 XA.XIR[14].XIC[4].icell.PUM VGND 0.00293f
C8121 XA.XIR[14].XIC[3].icell.Ien VGND 0.37144f
C8122 XA.XIR[14].XIC[2].icell.SM VGND 0.00502f
C8123 XA.XIR[14].XIC[3].icell.PUM VGND 0.00293f
C8124 XA.XIR[14].XIC[2].icell.Ien VGND 0.37144f
C8125 XA.XIR[14].XIC[1].icell.SM VGND 0.00502f
C8126 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80696f
C8127 XThR.Tn[14] VGND 14.14128f
C8128 XA.XIR[14].XIC[2].icell.PUM VGND 0.00293f
C8129 XA.XIR[14].XIC[1].icell.Ien VGND 0.37144f
C8130 XA.XIR[14].XIC[0].icell.SM VGND 0.00502f
C8131 a_n997_1579# VGND 0.54776f
C8132 XA.XIR[14].XIC[1].icell.PUM VGND 0.00293f
C8133 XA.XIR[14].XIC[0].icell.Ien VGND 0.37178f
C8134 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01044f
C8135 XA.XIR[14].XIC[0].icell.PUM VGND 0.00516f
C8136 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57579f
C8137 XA.XIR[14].XIC_dummy_left.icell.PUM VGND 0.00215f
C8138 a_n997_1803# VGND 0.53619f
C8139 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C8140 XA.XIR[14].XIC_15.icell.PDM VGND 0.18855f
C8141 XA.XIR[14].XIC[14].icell.PDM VGND 0.18809f
C8142 XA.XIR[14].XIC[13].icell.PDM VGND 0.18809f
C8143 XA.XIR[14].XIC[12].icell.PDM VGND 0.18809f
C8144 XA.XIR[14].XIC[11].icell.PDM VGND 0.18809f
C8145 XA.XIR[14].XIC[10].icell.PDM VGND 0.18809f
C8146 XA.XIR[14].XIC[9].icell.PDM VGND 0.18809f
C8147 XA.XIR[14].XIC[8].icell.PDM VGND 0.18809f
C8148 XA.XIR[14].XIC[7].icell.PDM VGND 0.18809f
C8149 XA.XIR[14].XIC[6].icell.PDM VGND 0.18809f
C8150 XA.XIR[14].XIC[5].icell.PDM VGND 0.18809f
C8151 XA.XIR[14].XIC[4].icell.PDM VGND 0.18809f
C8152 XA.XIR[14].XIC[3].icell.PDM VGND 0.18809f
C8153 XA.XIR[14].XIC[2].icell.PDM VGND 0.18809f
C8154 XA.XIR[14].XIC[1].icell.PDM VGND 0.18809f
C8155 XA.XIR[14].XIC[0].icell.PDM VGND 0.18817f
C8156 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C8157 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85795f
C8158 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C8159 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60802f
C8160 XA.XIR[13].XIC_15.icell.SM VGND 0.00474f
C8161 XA.XIR[13].XIC_dummy_right.icell.PUM VGND 0.00215f
C8162 XA.XIR[13].XIC_15.icell.Ien VGND 0.37063f
C8163 XA.XIR[13].XIC[14].icell.SM VGND 0.00502f
C8164 XA.XIR[13].XIC_15.icell.PUM VGND 0.00282f
C8165 XA.XIR[13].XIC[14].icell.Ien VGND 0.37144f
C8166 XA.XIR[13].XIC[13].icell.SM VGND 0.00502f
C8167 XA.XIR[13].XIC[14].icell.PUM VGND 0.00293f
C8168 XA.XIR[13].XIC[13].icell.Ien VGND 0.37144f
C8169 XA.XIR[13].XIC[12].icell.SM VGND 0.00502f
C8170 XA.XIR[13].XIC[13].icell.PUM VGND 0.00293f
C8171 XA.XIR[13].XIC[12].icell.Ien VGND 0.37144f
C8172 XA.XIR[13].XIC[11].icell.SM VGND 0.00502f
C8173 XA.XIR[13].XIC[12].icell.PUM VGND 0.00293f
C8174 XA.XIR[13].XIC[11].icell.Ien VGND 0.37144f
C8175 XA.XIR[13].XIC[10].icell.SM VGND 0.00502f
C8176 XA.XIR[13].XIC[11].icell.PUM VGND 0.00293f
C8177 XA.XIR[13].XIC[10].icell.Ien VGND 0.37144f
C8178 XA.XIR[13].XIC[9].icell.SM VGND 0.00502f
C8179 XA.XIR[13].XIC[10].icell.PUM VGND 0.00293f
C8180 XA.XIR[13].XIC[9].icell.Ien VGND 0.37144f
C8181 XA.XIR[13].XIC[8].icell.SM VGND 0.00502f
C8182 XA.XIR[13].XIC[9].icell.PUM VGND 0.00293f
C8183 XA.XIR[13].XIC[8].icell.Ien VGND 0.37144f
C8184 XA.XIR[13].XIC[7].icell.SM VGND 0.00502f
C8185 XA.XIR[13].XIC[8].icell.PUM VGND 0.00293f
C8186 XA.XIR[13].XIC[7].icell.Ien VGND 0.37144f
C8187 XA.XIR[13].XIC[6].icell.SM VGND 0.00502f
C8188 XA.XIR[13].XIC[7].icell.PUM VGND 0.00293f
C8189 XA.XIR[13].XIC[6].icell.Ien VGND 0.37144f
C8190 XA.XIR[13].XIC[5].icell.SM VGND 0.00502f
C8191 XA.XIR[13].XIC[6].icell.PUM VGND 0.00293f
C8192 XA.XIR[13].XIC[5].icell.Ien VGND 0.37144f
C8193 XA.XIR[13].XIC[4].icell.SM VGND 0.00502f
C8194 XA.XIR[13].XIC[5].icell.PUM VGND 0.00293f
C8195 XA.XIR[13].XIC[4].icell.Ien VGND 0.37144f
C8196 XA.XIR[13].XIC[3].icell.SM VGND 0.00502f
C8197 XA.XIR[13].XIC[4].icell.PUM VGND 0.00293f
C8198 XA.XIR[13].XIC[3].icell.Ien VGND 0.37144f
C8199 XA.XIR[13].XIC[2].icell.SM VGND 0.00502f
C8200 XA.XIR[13].XIC[3].icell.PUM VGND 0.00293f
C8201 XA.XIR[13].XIC[2].icell.Ien VGND 0.37144f
C8202 XA.XIR[13].XIC[1].icell.SM VGND 0.00502f
C8203 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.807f
C8204 XThR.Tn[13] VGND 14.01892f
C8205 XA.XIR[13].XIC[2].icell.PUM VGND 0.00293f
C8206 XA.XIR[13].XIC[1].icell.Ien VGND 0.37144f
C8207 XA.XIR[13].XIC[0].icell.SM VGND 0.00502f
C8208 XA.XIR[13].XIC[1].icell.PUM VGND 0.00293f
C8209 XA.XIR[13].XIC[0].icell.Ien VGND 0.37178f
C8210 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01044f
C8211 XA.XIR[13].XIC[0].icell.PUM VGND 0.00516f
C8212 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57425f
C8213 XA.XIR[13].XIC_dummy_left.icell.PUM VGND 0.00215f
C8214 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C8215 XA.XIR[13].XIC_15.icell.PDM VGND 0.18855f
C8216 XA.XIR[13].XIC[14].icell.PDM VGND 0.18809f
C8217 XA.XIR[13].XIC[13].icell.PDM VGND 0.18809f
C8218 XA.XIR[13].XIC[12].icell.PDM VGND 0.18809f
C8219 XA.XIR[13].XIC[11].icell.PDM VGND 0.18809f
C8220 XA.XIR[13].XIC[10].icell.PDM VGND 0.18809f
C8221 XA.XIR[13].XIC[9].icell.PDM VGND 0.18809f
C8222 XA.XIR[13].XIC[8].icell.PDM VGND 0.18809f
C8223 XA.XIR[13].XIC[7].icell.PDM VGND 0.18809f
C8224 XA.XIR[13].XIC[6].icell.PDM VGND 0.18809f
C8225 XA.XIR[13].XIC[5].icell.PDM VGND 0.18809f
C8226 XA.XIR[13].XIC[4].icell.PDM VGND 0.18809f
C8227 XA.XIR[13].XIC[3].icell.PDM VGND 0.18809f
C8228 XA.XIR[13].XIC[2].icell.PDM VGND 0.18809f
C8229 XA.XIR[13].XIC[1].icell.PDM VGND 0.18809f
C8230 XA.XIR[13].XIC[0].icell.PDM VGND 0.18817f
C8231 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C8232 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85795f
C8233 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C8234 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60802f
C8235 XA.XIR[12].XIC_15.icell.SM VGND 0.00474f
C8236 XA.XIR[12].XIC_dummy_right.icell.PUM VGND 0.00215f
C8237 XA.XIR[12].XIC_15.icell.Ien VGND 0.37063f
C8238 XA.XIR[12].XIC[14].icell.SM VGND 0.00502f
C8239 XA.XIR[12].XIC_15.icell.PUM VGND 0.00282f
C8240 XA.XIR[12].XIC[14].icell.Ien VGND 0.37144f
C8241 XA.XIR[12].XIC[13].icell.SM VGND 0.00502f
C8242 XA.XIR[12].XIC[14].icell.PUM VGND 0.00293f
C8243 XA.XIR[12].XIC[13].icell.Ien VGND 0.37144f
C8244 XA.XIR[12].XIC[12].icell.SM VGND 0.00502f
C8245 XA.XIR[12].XIC[13].icell.PUM VGND 0.00293f
C8246 XA.XIR[12].XIC[12].icell.Ien VGND 0.37144f
C8247 XA.XIR[12].XIC[11].icell.SM VGND 0.00502f
C8248 XA.XIR[12].XIC[12].icell.PUM VGND 0.00293f
C8249 XA.XIR[12].XIC[11].icell.Ien VGND 0.37144f
C8250 XA.XIR[12].XIC[10].icell.SM VGND 0.00502f
C8251 XA.XIR[12].XIC[11].icell.PUM VGND 0.00293f
C8252 XA.XIR[12].XIC[10].icell.Ien VGND 0.37144f
C8253 XA.XIR[12].XIC[9].icell.SM VGND 0.00502f
C8254 XA.XIR[12].XIC[10].icell.PUM VGND 0.00293f
C8255 XA.XIR[12].XIC[9].icell.Ien VGND 0.37144f
C8256 XA.XIR[12].XIC[8].icell.SM VGND 0.00502f
C8257 XA.XIR[12].XIC[9].icell.PUM VGND 0.00293f
C8258 XA.XIR[12].XIC[8].icell.Ien VGND 0.37144f
C8259 XA.XIR[12].XIC[7].icell.SM VGND 0.00502f
C8260 XA.XIR[12].XIC[8].icell.PUM VGND 0.00293f
C8261 XA.XIR[12].XIC[7].icell.Ien VGND 0.37144f
C8262 XA.XIR[12].XIC[6].icell.SM VGND 0.00502f
C8263 XA.XIR[12].XIC[7].icell.PUM VGND 0.00293f
C8264 XA.XIR[12].XIC[6].icell.Ien VGND 0.37144f
C8265 XA.XIR[12].XIC[5].icell.SM VGND 0.00502f
C8266 XA.XIR[12].XIC[6].icell.PUM VGND 0.00293f
C8267 XA.XIR[12].XIC[5].icell.Ien VGND 0.37144f
C8268 XA.XIR[12].XIC[4].icell.SM VGND 0.00502f
C8269 XA.XIR[12].XIC[5].icell.PUM VGND 0.00293f
C8270 XA.XIR[12].XIC[4].icell.Ien VGND 0.37144f
C8271 XA.XIR[12].XIC[3].icell.SM VGND 0.00502f
C8272 XA.XIR[12].XIC[4].icell.PUM VGND 0.00293f
C8273 XA.XIR[12].XIC[3].icell.Ien VGND 0.37144f
C8274 XA.XIR[12].XIC[2].icell.SM VGND 0.00502f
C8275 XA.XIR[12].XIC[3].icell.PUM VGND 0.00293f
C8276 XA.XIR[12].XIC[2].icell.Ien VGND 0.37144f
C8277 XA.XIR[12].XIC[1].icell.SM VGND 0.00502f
C8278 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80565f
C8279 XThR.Tn[12] VGND 13.90987f
C8280 XA.XIR[12].XIC[2].icell.PUM VGND 0.00293f
C8281 XA.XIR[12].XIC[1].icell.Ien VGND 0.37144f
C8282 XA.XIR[12].XIC[0].icell.SM VGND 0.00502f
C8283 XA.XIR[12].XIC[1].icell.PUM VGND 0.00293f
C8284 XA.XIR[12].XIC[0].icell.Ien VGND 0.37178f
C8285 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01044f
C8286 XA.XIR[12].XIC[0].icell.PUM VGND 0.00516f
C8287 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.57283f
C8288 XA.XIR[12].XIC_dummy_left.icell.PUM VGND 0.00215f
C8289 a_n997_2667# VGND 0.5457f
C8290 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C8291 XA.XIR[12].XIC_15.icell.PDM VGND 0.18855f
C8292 XA.XIR[12].XIC[14].icell.PDM VGND 0.18809f
C8293 XA.XIR[12].XIC[13].icell.PDM VGND 0.18809f
C8294 XA.XIR[12].XIC[12].icell.PDM VGND 0.18809f
C8295 XA.XIR[12].XIC[11].icell.PDM VGND 0.18809f
C8296 XA.XIR[12].XIC[10].icell.PDM VGND 0.18809f
C8297 XA.XIR[12].XIC[9].icell.PDM VGND 0.18809f
C8298 XA.XIR[12].XIC[8].icell.PDM VGND 0.18809f
C8299 XA.XIR[12].XIC[7].icell.PDM VGND 0.18809f
C8300 XA.XIR[12].XIC[6].icell.PDM VGND 0.18809f
C8301 XA.XIR[12].XIC[5].icell.PDM VGND 0.18809f
C8302 XA.XIR[12].XIC[4].icell.PDM VGND 0.18809f
C8303 XA.XIR[12].XIC[3].icell.PDM VGND 0.18809f
C8304 XA.XIR[12].XIC[2].icell.PDM VGND 0.18809f
C8305 XA.XIR[12].XIC[1].icell.PDM VGND 0.18809f
C8306 XA.XIR[12].XIC[0].icell.PDM VGND 0.18817f
C8307 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C8308 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85795f
C8309 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C8310 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60802f
C8311 XA.XIR[11].XIC_15.icell.SM VGND 0.00474f
C8312 XA.XIR[11].XIC_dummy_right.icell.PUM VGND 0.00215f
C8313 XA.XIR[11].XIC_15.icell.Ien VGND 0.37063f
C8314 XA.XIR[11].XIC[14].icell.SM VGND 0.00502f
C8315 XA.XIR[11].XIC_15.icell.PUM VGND 0.00282f
C8316 XA.XIR[11].XIC[14].icell.Ien VGND 0.37144f
C8317 XA.XIR[11].XIC[13].icell.SM VGND 0.00502f
C8318 XA.XIR[11].XIC[14].icell.PUM VGND 0.00293f
C8319 XA.XIR[11].XIC[13].icell.Ien VGND 0.37144f
C8320 XA.XIR[11].XIC[12].icell.SM VGND 0.00502f
C8321 XA.XIR[11].XIC[13].icell.PUM VGND 0.00293f
C8322 XA.XIR[11].XIC[12].icell.Ien VGND 0.37144f
C8323 XA.XIR[11].XIC[11].icell.SM VGND 0.00502f
C8324 XA.XIR[11].XIC[12].icell.PUM VGND 0.00293f
C8325 XA.XIR[11].XIC[11].icell.Ien VGND 0.37144f
C8326 XA.XIR[11].XIC[10].icell.SM VGND 0.00502f
C8327 XA.XIR[11].XIC[11].icell.PUM VGND 0.00293f
C8328 XA.XIR[11].XIC[10].icell.Ien VGND 0.37144f
C8329 XA.XIR[11].XIC[9].icell.SM VGND 0.00502f
C8330 XA.XIR[11].XIC[10].icell.PUM VGND 0.00293f
C8331 XA.XIR[11].XIC[9].icell.Ien VGND 0.37144f
C8332 XA.XIR[11].XIC[8].icell.SM VGND 0.00502f
C8333 XA.XIR[11].XIC[9].icell.PUM VGND 0.00293f
C8334 XA.XIR[11].XIC[8].icell.Ien VGND 0.37144f
C8335 XA.XIR[11].XIC[7].icell.SM VGND 0.00502f
C8336 XA.XIR[11].XIC[8].icell.PUM VGND 0.00293f
C8337 XA.XIR[11].XIC[7].icell.Ien VGND 0.37144f
C8338 XA.XIR[11].XIC[6].icell.SM VGND 0.00502f
C8339 XA.XIR[11].XIC[7].icell.PUM VGND 0.00293f
C8340 XA.XIR[11].XIC[6].icell.Ien VGND 0.37144f
C8341 XA.XIR[11].XIC[5].icell.SM VGND 0.00502f
C8342 XA.XIR[11].XIC[6].icell.PUM VGND 0.00293f
C8343 XA.XIR[11].XIC[5].icell.Ien VGND 0.37144f
C8344 XA.XIR[11].XIC[4].icell.SM VGND 0.00502f
C8345 XA.XIR[11].XIC[5].icell.PUM VGND 0.00293f
C8346 XA.XIR[11].XIC[4].icell.Ien VGND 0.37144f
C8347 XA.XIR[11].XIC[3].icell.SM VGND 0.00502f
C8348 XA.XIR[11].XIC[4].icell.PUM VGND 0.00293f
C8349 XA.XIR[11].XIC[3].icell.Ien VGND 0.37144f
C8350 XA.XIR[11].XIC[2].icell.SM VGND 0.00502f
C8351 XA.XIR[11].XIC[3].icell.PUM VGND 0.00293f
C8352 XA.XIR[11].XIC[2].icell.Ien VGND 0.37144f
C8353 XA.XIR[11].XIC[1].icell.SM VGND 0.00502f
C8354 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.808f
C8355 XThR.Tn[11] VGND 13.97038f
C8356 XA.XIR[11].XIC[2].icell.PUM VGND 0.00293f
C8357 XA.XIR[11].XIC[1].icell.Ien VGND 0.37144f
C8358 XA.XIR[11].XIC[0].icell.SM VGND 0.00502f
C8359 a_n997_2891# VGND 0.54795f
C8360 a_n1331_2891# VGND 0.00194f
C8361 XA.XIR[11].XIC[1].icell.PUM VGND 0.00293f
C8362 XA.XIR[11].XIC[0].icell.Ien VGND 0.37178f
C8363 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01044f
C8364 XA.XIR[11].XIC[0].icell.PUM VGND 0.00516f
C8365 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57297f
C8366 XA.XIR[11].XIC_dummy_left.icell.PUM VGND 0.00215f
C8367 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C8368 XA.XIR[11].XIC_15.icell.PDM VGND 0.18855f
C8369 XA.XIR[11].XIC[14].icell.PDM VGND 0.18809f
C8370 XA.XIR[11].XIC[13].icell.PDM VGND 0.18809f
C8371 XA.XIR[11].XIC[12].icell.PDM VGND 0.18809f
C8372 XA.XIR[11].XIC[11].icell.PDM VGND 0.18809f
C8373 XA.XIR[11].XIC[10].icell.PDM VGND 0.18809f
C8374 XA.XIR[11].XIC[9].icell.PDM VGND 0.18809f
C8375 XA.XIR[11].XIC[8].icell.PDM VGND 0.18809f
C8376 XA.XIR[11].XIC[7].icell.PDM VGND 0.18809f
C8377 XA.XIR[11].XIC[6].icell.PDM VGND 0.18809f
C8378 XA.XIR[11].XIC[5].icell.PDM VGND 0.18809f
C8379 XA.XIR[11].XIC[4].icell.PDM VGND 0.18809f
C8380 XA.XIR[11].XIC[3].icell.PDM VGND 0.18809f
C8381 XA.XIR[11].XIC[2].icell.PDM VGND 0.18809f
C8382 XA.XIR[11].XIC[1].icell.PDM VGND 0.18809f
C8383 XA.XIR[11].XIC[0].icell.PDM VGND 0.18817f
C8384 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C8385 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85795f
C8386 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C8387 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60802f
C8388 XA.XIR[10].XIC_15.icell.SM VGND 0.00474f
C8389 XA.XIR[10].XIC_dummy_right.icell.PUM VGND 0.00215f
C8390 XA.XIR[10].XIC_15.icell.Ien VGND 0.37063f
C8391 XA.XIR[10].XIC[14].icell.SM VGND 0.00502f
C8392 XA.XIR[10].XIC_15.icell.PUM VGND 0.00282f
C8393 XA.XIR[10].XIC[14].icell.Ien VGND 0.37144f
C8394 XA.XIR[10].XIC[13].icell.SM VGND 0.00502f
C8395 XA.XIR[10].XIC[14].icell.PUM VGND 0.00293f
C8396 XA.XIR[10].XIC[13].icell.Ien VGND 0.37144f
C8397 XA.XIR[10].XIC[12].icell.SM VGND 0.00502f
C8398 XA.XIR[10].XIC[13].icell.PUM VGND 0.00293f
C8399 XA.XIR[10].XIC[12].icell.Ien VGND 0.37144f
C8400 XA.XIR[10].XIC[11].icell.SM VGND 0.00502f
C8401 XA.XIR[10].XIC[12].icell.PUM VGND 0.00293f
C8402 XA.XIR[10].XIC[11].icell.Ien VGND 0.37144f
C8403 XA.XIR[10].XIC[10].icell.SM VGND 0.00502f
C8404 XA.XIR[10].XIC[11].icell.PUM VGND 0.00293f
C8405 XA.XIR[10].XIC[10].icell.Ien VGND 0.37144f
C8406 XA.XIR[10].XIC[9].icell.SM VGND 0.00502f
C8407 XA.XIR[10].XIC[10].icell.PUM VGND 0.00293f
C8408 XA.XIR[10].XIC[9].icell.Ien VGND 0.37144f
C8409 XA.XIR[10].XIC[8].icell.SM VGND 0.00502f
C8410 XA.XIR[10].XIC[9].icell.PUM VGND 0.00293f
C8411 XA.XIR[10].XIC[8].icell.Ien VGND 0.37144f
C8412 XA.XIR[10].XIC[7].icell.SM VGND 0.00502f
C8413 XA.XIR[10].XIC[8].icell.PUM VGND 0.00293f
C8414 XA.XIR[10].XIC[7].icell.Ien VGND 0.37144f
C8415 XA.XIR[10].XIC[6].icell.SM VGND 0.00502f
C8416 XA.XIR[10].XIC[7].icell.PUM VGND 0.00293f
C8417 XA.XIR[10].XIC[6].icell.Ien VGND 0.37144f
C8418 XA.XIR[10].XIC[5].icell.SM VGND 0.00502f
C8419 XA.XIR[10].XIC[6].icell.PUM VGND 0.00293f
C8420 XA.XIR[10].XIC[5].icell.Ien VGND 0.37144f
C8421 XA.XIR[10].XIC[4].icell.SM VGND 0.00502f
C8422 XA.XIR[10].XIC[5].icell.PUM VGND 0.00293f
C8423 XA.XIR[10].XIC[4].icell.Ien VGND 0.37144f
C8424 XA.XIR[10].XIC[3].icell.SM VGND 0.00502f
C8425 XA.XIR[10].XIC[4].icell.PUM VGND 0.00293f
C8426 XA.XIR[10].XIC[3].icell.Ien VGND 0.37144f
C8427 XA.XIR[10].XIC[2].icell.SM VGND 0.00502f
C8428 XA.XIR[10].XIC[3].icell.PUM VGND 0.00293f
C8429 XA.XIR[10].XIC[2].icell.Ien VGND 0.37144f
C8430 XA.XIR[10].XIC[1].icell.SM VGND 0.00502f
C8431 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80684f
C8432 XThR.Tn[10] VGND 13.91105f
C8433 XA.XIR[10].XIC[2].icell.PUM VGND 0.00293f
C8434 XA.XIR[10].XIC[1].icell.Ien VGND 0.37144f
C8435 XA.XIR[10].XIC[0].icell.SM VGND 0.00502f
C8436 XA.XIR[10].XIC[1].icell.PUM VGND 0.00293f
C8437 XA.XIR[10].XIC[0].icell.Ien VGND 0.37178f
C8438 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01044f
C8439 XA.XIR[10].XIC[0].icell.PUM VGND 0.00516f
C8440 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57425f
C8441 XA.XIR[10].XIC_dummy_left.icell.PUM VGND 0.00215f
C8442 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C8443 XA.XIR[10].XIC_15.icell.PDM VGND 0.18855f
C8444 XA.XIR[10].XIC[14].icell.PDM VGND 0.18809f
C8445 XA.XIR[10].XIC[13].icell.PDM VGND 0.18809f
C8446 XA.XIR[10].XIC[12].icell.PDM VGND 0.18809f
C8447 XA.XIR[10].XIC[11].icell.PDM VGND 0.18809f
C8448 XA.XIR[10].XIC[10].icell.PDM VGND 0.18809f
C8449 XA.XIR[10].XIC[9].icell.PDM VGND 0.18809f
C8450 XA.XIR[10].XIC[8].icell.PDM VGND 0.18809f
C8451 XA.XIR[10].XIC[7].icell.PDM VGND 0.18809f
C8452 XA.XIR[10].XIC[6].icell.PDM VGND 0.18809f
C8453 XA.XIR[10].XIC[5].icell.PDM VGND 0.18809f
C8454 XA.XIR[10].XIC[4].icell.PDM VGND 0.18809f
C8455 XA.XIR[10].XIC[3].icell.PDM VGND 0.18809f
C8456 XA.XIR[10].XIC[2].icell.PDM VGND 0.18809f
C8457 XA.XIR[10].XIC[1].icell.PDM VGND 0.18809f
C8458 XA.XIR[10].XIC[0].icell.PDM VGND 0.18817f
C8459 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C8460 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85795f
C8461 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C8462 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60802f
C8463 XA.XIR[9].XIC_15.icell.SM VGND 0.00474f
C8464 XA.XIR[9].XIC_dummy_right.icell.PUM VGND 0.00215f
C8465 XA.XIR[9].XIC_15.icell.Ien VGND 0.37063f
C8466 XA.XIR[9].XIC[14].icell.SM VGND 0.00502f
C8467 XA.XIR[9].XIC_15.icell.PUM VGND 0.00282f
C8468 XA.XIR[9].XIC[14].icell.Ien VGND 0.37144f
C8469 XA.XIR[9].XIC[13].icell.SM VGND 0.00502f
C8470 XA.XIR[9].XIC[14].icell.PUM VGND 0.00293f
C8471 XA.XIR[9].XIC[13].icell.Ien VGND 0.37144f
C8472 XA.XIR[9].XIC[12].icell.SM VGND 0.00502f
C8473 XA.XIR[9].XIC[13].icell.PUM VGND 0.00293f
C8474 XA.XIR[9].XIC[12].icell.Ien VGND 0.37144f
C8475 XA.XIR[9].XIC[11].icell.SM VGND 0.00502f
C8476 XA.XIR[9].XIC[12].icell.PUM VGND 0.00293f
C8477 XA.XIR[9].XIC[11].icell.Ien VGND 0.37144f
C8478 XA.XIR[9].XIC[10].icell.SM VGND 0.00502f
C8479 XA.XIR[9].XIC[11].icell.PUM VGND 0.00293f
C8480 XA.XIR[9].XIC[10].icell.Ien VGND 0.37144f
C8481 XA.XIR[9].XIC[9].icell.SM VGND 0.00502f
C8482 XA.XIR[9].XIC[10].icell.PUM VGND 0.00293f
C8483 XA.XIR[9].XIC[9].icell.Ien VGND 0.37144f
C8484 XA.XIR[9].XIC[8].icell.SM VGND 0.00502f
C8485 XA.XIR[9].XIC[9].icell.PUM VGND 0.00293f
C8486 XA.XIR[9].XIC[8].icell.Ien VGND 0.37144f
C8487 XA.XIR[9].XIC[7].icell.SM VGND 0.00502f
C8488 XA.XIR[9].XIC[8].icell.PUM VGND 0.00293f
C8489 XA.XIR[9].XIC[7].icell.Ien VGND 0.37144f
C8490 XA.XIR[9].XIC[6].icell.SM VGND 0.00502f
C8491 XA.XIR[9].XIC[7].icell.PUM VGND 0.00293f
C8492 XA.XIR[9].XIC[6].icell.Ien VGND 0.37144f
C8493 XA.XIR[9].XIC[5].icell.SM VGND 0.00502f
C8494 XA.XIR[9].XIC[6].icell.PUM VGND 0.00293f
C8495 XA.XIR[9].XIC[5].icell.Ien VGND 0.37144f
C8496 XA.XIR[9].XIC[4].icell.SM VGND 0.00502f
C8497 XA.XIR[9].XIC[5].icell.PUM VGND 0.00293f
C8498 XA.XIR[9].XIC[4].icell.Ien VGND 0.37144f
C8499 XA.XIR[9].XIC[3].icell.SM VGND 0.00502f
C8500 XA.XIR[9].XIC[4].icell.PUM VGND 0.00293f
C8501 XA.XIR[9].XIC[3].icell.Ien VGND 0.37144f
C8502 XA.XIR[9].XIC[2].icell.SM VGND 0.00502f
C8503 XA.XIR[9].XIC[3].icell.PUM VGND 0.00293f
C8504 XA.XIR[9].XIC[2].icell.Ien VGND 0.37144f
C8505 XA.XIR[9].XIC[1].icell.SM VGND 0.00502f
C8506 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.8087f
C8507 XA.XIR[9].XIC[2].icell.PUM VGND 0.00293f
C8508 XA.XIR[9].XIC[1].icell.Ien VGND 0.37144f
C8509 XA.XIR[9].XIC[0].icell.SM VGND 0.00502f
C8510 XThR.Tn[9] VGND 13.95272f
C8511 a_n997_3755# VGND 0.54861f
C8512 XA.XIR[9].XIC[1].icell.PUM VGND 0.00293f
C8513 XA.XIR[9].XIC[0].icell.Ien VGND 0.37178f
C8514 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01044f
C8515 XA.XIR[9].XIC[0].icell.PUM VGND 0.00516f
C8516 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.57323f
C8517 a_n997_3979# VGND 0.54721f
C8518 XA.XIR[9].XIC_dummy_left.icell.PUM VGND 0.00215f
C8519 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C8520 XA.XIR[9].XIC_15.icell.PDM VGND 0.18855f
C8521 XA.XIR[9].XIC[14].icell.PDM VGND 0.18809f
C8522 XA.XIR[9].XIC[13].icell.PDM VGND 0.18809f
C8523 XA.XIR[9].XIC[12].icell.PDM VGND 0.18809f
C8524 XA.XIR[9].XIC[11].icell.PDM VGND 0.18809f
C8525 XA.XIR[9].XIC[10].icell.PDM VGND 0.18809f
C8526 XA.XIR[9].XIC[9].icell.PDM VGND 0.18809f
C8527 XA.XIR[9].XIC[8].icell.PDM VGND 0.18809f
C8528 XA.XIR[9].XIC[7].icell.PDM VGND 0.18809f
C8529 XA.XIR[9].XIC[6].icell.PDM VGND 0.18809f
C8530 XA.XIR[9].XIC[5].icell.PDM VGND 0.18809f
C8531 XA.XIR[9].XIC[4].icell.PDM VGND 0.18809f
C8532 XA.XIR[9].XIC[3].icell.PDM VGND 0.18809f
C8533 XA.XIR[9].XIC[2].icell.PDM VGND 0.18809f
C8534 XA.XIR[9].XIC[1].icell.PDM VGND 0.18809f
C8535 XA.XIR[9].XIC[0].icell.PDM VGND 0.18817f
C8536 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C8537 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85795f
C8538 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C8539 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60802f
C8540 XA.XIR[8].XIC_15.icell.SM VGND 0.00474f
C8541 XA.XIR[8].XIC_dummy_right.icell.PUM VGND 0.00215f
C8542 XA.XIR[8].XIC_15.icell.Ien VGND 0.37063f
C8543 XA.XIR[8].XIC[14].icell.SM VGND 0.00502f
C8544 XA.XIR[8].XIC_15.icell.PUM VGND 0.00282f
C8545 XA.XIR[8].XIC[14].icell.Ien VGND 0.37144f
C8546 XA.XIR[8].XIC[13].icell.SM VGND 0.00502f
C8547 XA.XIR[8].XIC[14].icell.PUM VGND 0.00293f
C8548 XA.XIR[8].XIC[13].icell.Ien VGND 0.37144f
C8549 XA.XIR[8].XIC[12].icell.SM VGND 0.00502f
C8550 XA.XIR[8].XIC[13].icell.PUM VGND 0.00293f
C8551 XA.XIR[8].XIC[12].icell.Ien VGND 0.37144f
C8552 XA.XIR[8].XIC[11].icell.SM VGND 0.00502f
C8553 XA.XIR[8].XIC[12].icell.PUM VGND 0.00293f
C8554 XA.XIR[8].XIC[11].icell.Ien VGND 0.37144f
C8555 XA.XIR[8].XIC[10].icell.SM VGND 0.00502f
C8556 XA.XIR[8].XIC[11].icell.PUM VGND 0.00293f
C8557 XA.XIR[8].XIC[10].icell.Ien VGND 0.37144f
C8558 XA.XIR[8].XIC[9].icell.SM VGND 0.00502f
C8559 XA.XIR[8].XIC[10].icell.PUM VGND 0.00293f
C8560 XA.XIR[8].XIC[9].icell.Ien VGND 0.37144f
C8561 XA.XIR[8].XIC[8].icell.SM VGND 0.00502f
C8562 XA.XIR[8].XIC[9].icell.PUM VGND 0.00293f
C8563 XA.XIR[8].XIC[8].icell.Ien VGND 0.37144f
C8564 XA.XIR[8].XIC[7].icell.SM VGND 0.00502f
C8565 XA.XIR[8].XIC[8].icell.PUM VGND 0.00293f
C8566 XA.XIR[8].XIC[7].icell.Ien VGND 0.37144f
C8567 XA.XIR[8].XIC[6].icell.SM VGND 0.00502f
C8568 XA.XIR[8].XIC[7].icell.PUM VGND 0.00293f
C8569 XA.XIR[8].XIC[6].icell.Ien VGND 0.37144f
C8570 XA.XIR[8].XIC[5].icell.SM VGND 0.00502f
C8571 XA.XIR[8].XIC[6].icell.PUM VGND 0.00293f
C8572 XA.XIR[8].XIC[5].icell.Ien VGND 0.37144f
C8573 XA.XIR[8].XIC[4].icell.SM VGND 0.00502f
C8574 XA.XIR[8].XIC[5].icell.PUM VGND 0.00293f
C8575 XA.XIR[8].XIC[4].icell.Ien VGND 0.37144f
C8576 XA.XIR[8].XIC[3].icell.SM VGND 0.00502f
C8577 XA.XIR[8].XIC[4].icell.PUM VGND 0.00293f
C8578 XA.XIR[8].XIC[3].icell.Ien VGND 0.37144f
C8579 XA.XIR[8].XIC[2].icell.SM VGND 0.00502f
C8580 XA.XIR[8].XIC[3].icell.PUM VGND 0.00293f
C8581 XA.XIR[8].XIC[2].icell.Ien VGND 0.37144f
C8582 XA.XIR[8].XIC[1].icell.SM VGND 0.00502f
C8583 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80602f
C8584 XA.XIR[8].XIC[2].icell.PUM VGND 0.00293f
C8585 XA.XIR[8].XIC[1].icell.Ien VGND 0.37144f
C8586 XA.XIR[8].XIC[0].icell.SM VGND 0.00502f
C8587 XThR.Tn[8] VGND 13.8971f
C8588 XA.XIR[8].XIC[1].icell.PUM VGND 0.00293f
C8589 XA.XIR[8].XIC[0].icell.Ien VGND 0.37178f
C8590 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01044f
C8591 XA.XIR[8].XIC[0].icell.PUM VGND 0.00516f
C8592 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57311f
C8593 XA.XIR[8].XIC_dummy_left.icell.PUM VGND 0.00215f
C8594 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C8595 XA.XIR[8].XIC_15.icell.PDM VGND 0.18855f
C8596 XA.XIR[8].XIC[14].icell.PDM VGND 0.18809f
C8597 XA.XIR[8].XIC[13].icell.PDM VGND 0.18809f
C8598 XA.XIR[8].XIC[12].icell.PDM VGND 0.18809f
C8599 XA.XIR[8].XIC[11].icell.PDM VGND 0.18809f
C8600 XA.XIR[8].XIC[10].icell.PDM VGND 0.18809f
C8601 XA.XIR[8].XIC[9].icell.PDM VGND 0.18809f
C8602 XA.XIR[8].XIC[8].icell.PDM VGND 0.18809f
C8603 XA.XIR[8].XIC[7].icell.PDM VGND 0.18809f
C8604 XA.XIR[8].XIC[6].icell.PDM VGND 0.18809f
C8605 XA.XIR[8].XIC[5].icell.PDM VGND 0.18809f
C8606 XA.XIR[8].XIC[4].icell.PDM VGND 0.18809f
C8607 XA.XIR[8].XIC[3].icell.PDM VGND 0.18809f
C8608 XA.XIR[8].XIC[2].icell.PDM VGND 0.18809f
C8609 XA.XIR[8].XIC[1].icell.PDM VGND 0.18809f
C8610 XA.XIR[8].XIC[0].icell.PDM VGND 0.18817f
C8611 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C8612 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85795f
C8613 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C8614 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60802f
C8615 XA.XIR[7].XIC_15.icell.SM VGND 0.00474f
C8616 XA.XIR[7].XIC_dummy_right.icell.PUM VGND 0.00215f
C8617 XA.XIR[7].XIC_15.icell.Ien VGND 0.37063f
C8618 XA.XIR[7].XIC[14].icell.SM VGND 0.00502f
C8619 XA.XIR[7].XIC_15.icell.PUM VGND 0.00282f
C8620 XA.XIR[7].XIC[14].icell.Ien VGND 0.37144f
C8621 XA.XIR[7].XIC[13].icell.SM VGND 0.00502f
C8622 XA.XIR[7].XIC[14].icell.PUM VGND 0.00293f
C8623 XA.XIR[7].XIC[13].icell.Ien VGND 0.37144f
C8624 XA.XIR[7].XIC[12].icell.SM VGND 0.00502f
C8625 XA.XIR[7].XIC[13].icell.PUM VGND 0.00293f
C8626 XA.XIR[7].XIC[12].icell.Ien VGND 0.37144f
C8627 XA.XIR[7].XIC[11].icell.SM VGND 0.00502f
C8628 XA.XIR[7].XIC[12].icell.PUM VGND 0.00293f
C8629 XA.XIR[7].XIC[11].icell.Ien VGND 0.37144f
C8630 XA.XIR[7].XIC[10].icell.SM VGND 0.00502f
C8631 XA.XIR[7].XIC[11].icell.PUM VGND 0.00293f
C8632 XA.XIR[7].XIC[10].icell.Ien VGND 0.37144f
C8633 XA.XIR[7].XIC[9].icell.SM VGND 0.00502f
C8634 XA.XIR[7].XIC[10].icell.PUM VGND 0.00293f
C8635 XA.XIR[7].XIC[9].icell.Ien VGND 0.37144f
C8636 XA.XIR[7].XIC[8].icell.SM VGND 0.00502f
C8637 XA.XIR[7].XIC[9].icell.PUM VGND 0.00293f
C8638 XA.XIR[7].XIC[8].icell.Ien VGND 0.37144f
C8639 XA.XIR[7].XIC[7].icell.SM VGND 0.00502f
C8640 XA.XIR[7].XIC[8].icell.PUM VGND 0.00293f
C8641 XA.XIR[7].XIC[7].icell.Ien VGND 0.37144f
C8642 XA.XIR[7].XIC[6].icell.SM VGND 0.00502f
C8643 XA.XIR[7].XIC[7].icell.PUM VGND 0.00293f
C8644 XA.XIR[7].XIC[6].icell.Ien VGND 0.37144f
C8645 XA.XIR[7].XIC[5].icell.SM VGND 0.00502f
C8646 XA.XIR[7].XIC[6].icell.PUM VGND 0.00293f
C8647 XA.XIR[7].XIC[5].icell.Ien VGND 0.37144f
C8648 XA.XIR[7].XIC[4].icell.SM VGND 0.00502f
C8649 XA.XIR[7].XIC[5].icell.PUM VGND 0.00293f
C8650 XA.XIR[7].XIC[4].icell.Ien VGND 0.37144f
C8651 XA.XIR[7].XIC[3].icell.SM VGND 0.00502f
C8652 XA.XIR[7].XIC[4].icell.PUM VGND 0.00293f
C8653 XA.XIR[7].XIC[3].icell.Ien VGND 0.37144f
C8654 XA.XIR[7].XIC[2].icell.SM VGND 0.00502f
C8655 XA.XIR[7].XIC[3].icell.PUM VGND 0.00293f
C8656 XA.XIR[7].XIC[2].icell.Ien VGND 0.37144f
C8657 XA.XIR[7].XIC[1].icell.SM VGND 0.00502f
C8658 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80634f
C8659 XA.XIR[7].XIC[2].icell.PUM VGND 0.00293f
C8660 XA.XIR[7].XIC[1].icell.Ien VGND 0.37144f
C8661 XA.XIR[7].XIC[0].icell.SM VGND 0.00502f
C8662 XA.XIR[7].XIC[1].icell.PUM VGND 0.00293f
C8663 XA.XIR[7].XIC[0].icell.Ien VGND 0.37178f
C8664 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01044f
C8665 XThR.Tn[7] VGND 14.38144f
C8666 XThR.XTBN.A VGND 1.22814f
C8667 XA.XIR[7].XIC[0].icell.PUM VGND 0.00516f
C8668 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57579f
C8669 XA.XIR[7].XIC_dummy_left.icell.PUM VGND 0.00222f
C8670 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C8671 XA.XIR[7].XIC_15.icell.PDM VGND 0.18855f
C8672 XA.XIR[7].XIC[14].icell.PDM VGND 0.18809f
C8673 XA.XIR[7].XIC[13].icell.PDM VGND 0.18809f
C8674 XA.XIR[7].XIC[12].icell.PDM VGND 0.18809f
C8675 XA.XIR[7].XIC[11].icell.PDM VGND 0.18809f
C8676 XA.XIR[7].XIC[10].icell.PDM VGND 0.18809f
C8677 XA.XIR[7].XIC[9].icell.PDM VGND 0.18809f
C8678 XA.XIR[7].XIC[8].icell.PDM VGND 0.18809f
C8679 XA.XIR[7].XIC[7].icell.PDM VGND 0.18809f
C8680 XA.XIR[7].XIC[6].icell.PDM VGND 0.18809f
C8681 XA.XIR[7].XIC[5].icell.PDM VGND 0.18809f
C8682 XA.XIR[7].XIC[4].icell.PDM VGND 0.18809f
C8683 XA.XIR[7].XIC[3].icell.PDM VGND 0.18809f
C8684 XA.XIR[7].XIC[2].icell.PDM VGND 0.18809f
C8685 XA.XIR[7].XIC[1].icell.PDM VGND 0.18809f
C8686 XA.XIR[7].XIC[0].icell.PDM VGND 0.18817f
C8687 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C8688 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85795f
C8689 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C8690 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60802f
C8691 XA.XIR[6].XIC_15.icell.SM VGND 0.00474f
C8692 XA.XIR[6].XIC_dummy_right.icell.PUM VGND 0.00215f
C8693 XA.XIR[6].XIC_15.icell.Ien VGND 0.37063f
C8694 XA.XIR[6].XIC[14].icell.SM VGND 0.00502f
C8695 XA.XIR[6].XIC_15.icell.PUM VGND 0.00282f
C8696 XA.XIR[6].XIC[14].icell.Ien VGND 0.37144f
C8697 XA.XIR[6].XIC[13].icell.SM VGND 0.00502f
C8698 XA.XIR[6].XIC[14].icell.PUM VGND 0.00293f
C8699 XA.XIR[6].XIC[13].icell.Ien VGND 0.37144f
C8700 XA.XIR[6].XIC[12].icell.SM VGND 0.00502f
C8701 XA.XIR[6].XIC[13].icell.PUM VGND 0.00293f
C8702 XA.XIR[6].XIC[12].icell.Ien VGND 0.37144f
C8703 XA.XIR[6].XIC[11].icell.SM VGND 0.00502f
C8704 XA.XIR[6].XIC[12].icell.PUM VGND 0.00293f
C8705 XA.XIR[6].XIC[11].icell.Ien VGND 0.37144f
C8706 XA.XIR[6].XIC[10].icell.SM VGND 0.00502f
C8707 XA.XIR[6].XIC[11].icell.PUM VGND 0.00293f
C8708 XA.XIR[6].XIC[10].icell.Ien VGND 0.37144f
C8709 XA.XIR[6].XIC[9].icell.SM VGND 0.00502f
C8710 XA.XIR[6].XIC[10].icell.PUM VGND 0.00293f
C8711 XA.XIR[6].XIC[9].icell.Ien VGND 0.37144f
C8712 XA.XIR[6].XIC[8].icell.SM VGND 0.00502f
C8713 XA.XIR[6].XIC[9].icell.PUM VGND 0.00293f
C8714 XA.XIR[6].XIC[8].icell.Ien VGND 0.37144f
C8715 XA.XIR[6].XIC[7].icell.SM VGND 0.00502f
C8716 XA.XIR[6].XIC[8].icell.PUM VGND 0.00293f
C8717 XA.XIR[6].XIC[7].icell.Ien VGND 0.37144f
C8718 XA.XIR[6].XIC[6].icell.SM VGND 0.00502f
C8719 XA.XIR[6].XIC[7].icell.PUM VGND 0.00293f
C8720 XA.XIR[6].XIC[6].icell.Ien VGND 0.37144f
C8721 XA.XIR[6].XIC[5].icell.SM VGND 0.00502f
C8722 XA.XIR[6].XIC[6].icell.PUM VGND 0.00293f
C8723 XA.XIR[6].XIC[5].icell.Ien VGND 0.37144f
C8724 XA.XIR[6].XIC[4].icell.SM VGND 0.00502f
C8725 XA.XIR[6].XIC[5].icell.PUM VGND 0.00293f
C8726 XA.XIR[6].XIC[4].icell.Ien VGND 0.37144f
C8727 XA.XIR[6].XIC[3].icell.SM VGND 0.00502f
C8728 XA.XIR[6].XIC[4].icell.PUM VGND 0.00293f
C8729 XA.XIR[6].XIC[3].icell.Ien VGND 0.37144f
C8730 XA.XIR[6].XIC[2].icell.SM VGND 0.00502f
C8731 XA.XIR[6].XIC[3].icell.PUM VGND 0.00293f
C8732 XA.XIR[6].XIC[2].icell.Ien VGND 0.37144f
C8733 XA.XIR[6].XIC[1].icell.SM VGND 0.00502f
C8734 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80729f
C8735 XA.XIR[6].XIC[2].icell.PUM VGND 0.00293f
C8736 XA.XIR[6].XIC[1].icell.Ien VGND 0.37144f
C8737 XA.XIR[6].XIC[0].icell.SM VGND 0.00502f
C8738 XA.XIR[6].XIC[1].icell.PUM VGND 0.00293f
C8739 XA.XIR[6].XIC[0].icell.Ien VGND 0.37178f
C8740 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01044f
C8741 XA.XIR[6].XIC[0].icell.PUM VGND 0.00516f
C8742 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57425f
C8743 XThR.Tn[6] VGND 13.98754f
C8744 a_n1049_5317# VGND 0.02283f
C8745 XA.XIR[6].XIC_dummy_left.icell.PUM VGND 0.00215f
C8746 XThR.XTB7.Y VGND 1.36132f
C8747 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C8748 XA.XIR[6].XIC_15.icell.PDM VGND 0.18855f
C8749 XA.XIR[6].XIC[14].icell.PDM VGND 0.18809f
C8750 XA.XIR[6].XIC[13].icell.PDM VGND 0.18809f
C8751 XA.XIR[6].XIC[12].icell.PDM VGND 0.18809f
C8752 XA.XIR[6].XIC[11].icell.PDM VGND 0.18809f
C8753 XA.XIR[6].XIC[10].icell.PDM VGND 0.18809f
C8754 XA.XIR[6].XIC[9].icell.PDM VGND 0.18809f
C8755 XA.XIR[6].XIC[8].icell.PDM VGND 0.18809f
C8756 XA.XIR[6].XIC[7].icell.PDM VGND 0.18809f
C8757 XA.XIR[6].XIC[6].icell.PDM VGND 0.18809f
C8758 XA.XIR[6].XIC[5].icell.PDM VGND 0.18809f
C8759 XA.XIR[6].XIC[4].icell.PDM VGND 0.18809f
C8760 XA.XIR[6].XIC[3].icell.PDM VGND 0.18809f
C8761 XA.XIR[6].XIC[2].icell.PDM VGND 0.18809f
C8762 XA.XIR[6].XIC[1].icell.PDM VGND 0.18809f
C8763 XA.XIR[6].XIC[0].icell.PDM VGND 0.18817f
C8764 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C8765 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85795f
C8766 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C8767 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60802f
C8768 XA.XIR[5].XIC_15.icell.SM VGND 0.00474f
C8769 XA.XIR[5].XIC_dummy_right.icell.PUM VGND 0.00215f
C8770 XA.XIR[5].XIC_15.icell.Ien VGND 0.37063f
C8771 XA.XIR[5].XIC[14].icell.SM VGND 0.00502f
C8772 XA.XIR[5].XIC_15.icell.PUM VGND 0.00282f
C8773 XA.XIR[5].XIC[14].icell.Ien VGND 0.37144f
C8774 XA.XIR[5].XIC[13].icell.SM VGND 0.00502f
C8775 XA.XIR[5].XIC[14].icell.PUM VGND 0.00293f
C8776 XA.XIR[5].XIC[13].icell.Ien VGND 0.37144f
C8777 XA.XIR[5].XIC[12].icell.SM VGND 0.00502f
C8778 XA.XIR[5].XIC[13].icell.PUM VGND 0.00293f
C8779 XA.XIR[5].XIC[12].icell.Ien VGND 0.37144f
C8780 XA.XIR[5].XIC[11].icell.SM VGND 0.00502f
C8781 XA.XIR[5].XIC[12].icell.PUM VGND 0.00293f
C8782 XA.XIR[5].XIC[11].icell.Ien VGND 0.37144f
C8783 XA.XIR[5].XIC[10].icell.SM VGND 0.00502f
C8784 XA.XIR[5].XIC[11].icell.PUM VGND 0.00293f
C8785 XA.XIR[5].XIC[10].icell.Ien VGND 0.37144f
C8786 XA.XIR[5].XIC[9].icell.SM VGND 0.00502f
C8787 XA.XIR[5].XIC[10].icell.PUM VGND 0.00293f
C8788 XA.XIR[5].XIC[9].icell.Ien VGND 0.37144f
C8789 XA.XIR[5].XIC[8].icell.SM VGND 0.00502f
C8790 XA.XIR[5].XIC[9].icell.PUM VGND 0.00293f
C8791 XA.XIR[5].XIC[8].icell.Ien VGND 0.37144f
C8792 XA.XIR[5].XIC[7].icell.SM VGND 0.00502f
C8793 XA.XIR[5].XIC[8].icell.PUM VGND 0.00293f
C8794 XA.XIR[5].XIC[7].icell.Ien VGND 0.37144f
C8795 XA.XIR[5].XIC[6].icell.SM VGND 0.00502f
C8796 XA.XIR[5].XIC[7].icell.PUM VGND 0.00293f
C8797 XA.XIR[5].XIC[6].icell.Ien VGND 0.37144f
C8798 XA.XIR[5].XIC[5].icell.SM VGND 0.00502f
C8799 XA.XIR[5].XIC[6].icell.PUM VGND 0.00293f
C8800 XA.XIR[5].XIC[5].icell.Ien VGND 0.37144f
C8801 XA.XIR[5].XIC[4].icell.SM VGND 0.00502f
C8802 XA.XIR[5].XIC[5].icell.PUM VGND 0.00293f
C8803 XA.XIR[5].XIC[4].icell.Ien VGND 0.37144f
C8804 XA.XIR[5].XIC[3].icell.SM VGND 0.00502f
C8805 XA.XIR[5].XIC[4].icell.PUM VGND 0.00293f
C8806 XA.XIR[5].XIC[3].icell.Ien VGND 0.37144f
C8807 XA.XIR[5].XIC[2].icell.SM VGND 0.00502f
C8808 XA.XIR[5].XIC[3].icell.PUM VGND 0.00293f
C8809 XA.XIR[5].XIC[2].icell.Ien VGND 0.37144f
C8810 XA.XIR[5].XIC[1].icell.SM VGND 0.00502f
C8811 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80598f
C8812 XA.XIR[5].XIC[2].icell.PUM VGND 0.00293f
C8813 XA.XIR[5].XIC[1].icell.Ien VGND 0.37144f
C8814 XA.XIR[5].XIC[0].icell.SM VGND 0.00502f
C8815 a_n1049_5611# VGND 0.02888f
C8816 XA.XIR[5].XIC[1].icell.PUM VGND 0.00293f
C8817 XA.XIR[5].XIC[0].icell.Ien VGND 0.37178f
C8818 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01044f
C8819 XA.XIR[5].XIC[0].icell.PUM VGND 0.00516f
C8820 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57291f
C8821 XA.XIR[5].XIC_dummy_left.icell.PUM VGND 0.00215f
C8822 XThR.Tn[5] VGND 13.96673f
C8823 XThR.XTB6.Y VGND 1.38212f
C8824 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C8825 XA.XIR[5].XIC_15.icell.PDM VGND 0.18855f
C8826 XA.XIR[5].XIC[14].icell.PDM VGND 0.18809f
C8827 XA.XIR[5].XIC[13].icell.PDM VGND 0.18809f
C8828 XA.XIR[5].XIC[12].icell.PDM VGND 0.18809f
C8829 XA.XIR[5].XIC[11].icell.PDM VGND 0.18809f
C8830 XA.XIR[5].XIC[10].icell.PDM VGND 0.18809f
C8831 XA.XIR[5].XIC[9].icell.PDM VGND 0.18809f
C8832 XA.XIR[5].XIC[8].icell.PDM VGND 0.18809f
C8833 XA.XIR[5].XIC[7].icell.PDM VGND 0.18809f
C8834 XA.XIR[5].XIC[6].icell.PDM VGND 0.18809f
C8835 XA.XIR[5].XIC[5].icell.PDM VGND 0.18809f
C8836 XA.XIR[5].XIC[4].icell.PDM VGND 0.18809f
C8837 XA.XIR[5].XIC[3].icell.PDM VGND 0.18809f
C8838 XA.XIR[5].XIC[2].icell.PDM VGND 0.18809f
C8839 XA.XIR[5].XIC[1].icell.PDM VGND 0.18809f
C8840 XA.XIR[5].XIC[0].icell.PDM VGND 0.18817f
C8841 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C8842 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85795f
C8843 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C8844 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60802f
C8845 XA.XIR[4].XIC_15.icell.SM VGND 0.00474f
C8846 XA.XIR[4].XIC_dummy_right.icell.PUM VGND 0.00215f
C8847 XA.XIR[4].XIC_15.icell.Ien VGND 0.37063f
C8848 XA.XIR[4].XIC[14].icell.SM VGND 0.00502f
C8849 XA.XIR[4].XIC_15.icell.PUM VGND 0.00282f
C8850 XA.XIR[4].XIC[14].icell.Ien VGND 0.37144f
C8851 XA.XIR[4].XIC[13].icell.SM VGND 0.00502f
C8852 XA.XIR[4].XIC[14].icell.PUM VGND 0.00293f
C8853 XA.XIR[4].XIC[13].icell.Ien VGND 0.37144f
C8854 XA.XIR[4].XIC[12].icell.SM VGND 0.00502f
C8855 XA.XIR[4].XIC[13].icell.PUM VGND 0.00293f
C8856 XA.XIR[4].XIC[12].icell.Ien VGND 0.37144f
C8857 XA.XIR[4].XIC[11].icell.SM VGND 0.00502f
C8858 XA.XIR[4].XIC[12].icell.PUM VGND 0.00293f
C8859 XA.XIR[4].XIC[11].icell.Ien VGND 0.37144f
C8860 XA.XIR[4].XIC[10].icell.SM VGND 0.00502f
C8861 XA.XIR[4].XIC[11].icell.PUM VGND 0.00293f
C8862 XA.XIR[4].XIC[10].icell.Ien VGND 0.37144f
C8863 XA.XIR[4].XIC[9].icell.SM VGND 0.00502f
C8864 XA.XIR[4].XIC[10].icell.PUM VGND 0.00293f
C8865 XA.XIR[4].XIC[9].icell.Ien VGND 0.37144f
C8866 XA.XIR[4].XIC[8].icell.SM VGND 0.00502f
C8867 XA.XIR[4].XIC[9].icell.PUM VGND 0.00293f
C8868 XA.XIR[4].XIC[8].icell.Ien VGND 0.37144f
C8869 XA.XIR[4].XIC[7].icell.SM VGND 0.00502f
C8870 XA.XIR[4].XIC[8].icell.PUM VGND 0.00293f
C8871 XA.XIR[4].XIC[7].icell.Ien VGND 0.37144f
C8872 XA.XIR[4].XIC[6].icell.SM VGND 0.00502f
C8873 XA.XIR[4].XIC[7].icell.PUM VGND 0.00293f
C8874 XA.XIR[4].XIC[6].icell.Ien VGND 0.37144f
C8875 XA.XIR[4].XIC[5].icell.SM VGND 0.00502f
C8876 XA.XIR[4].XIC[6].icell.PUM VGND 0.00293f
C8877 XA.XIR[4].XIC[5].icell.Ien VGND 0.37144f
C8878 XA.XIR[4].XIC[4].icell.SM VGND 0.00502f
C8879 XA.XIR[4].XIC[5].icell.PUM VGND 0.00293f
C8880 XA.XIR[4].XIC[4].icell.Ien VGND 0.37144f
C8881 XA.XIR[4].XIC[3].icell.SM VGND 0.00502f
C8882 XA.XIR[4].XIC[4].icell.PUM VGND 0.00293f
C8883 XA.XIR[4].XIC[3].icell.Ien VGND 0.37144f
C8884 XA.XIR[4].XIC[2].icell.SM VGND 0.00502f
C8885 XA.XIR[4].XIC[3].icell.PUM VGND 0.00293f
C8886 XA.XIR[4].XIC[2].icell.Ien VGND 0.37144f
C8887 XA.XIR[4].XIC[1].icell.SM VGND 0.00502f
C8888 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.8077f
C8889 XA.XIR[4].XIC[2].icell.PUM VGND 0.00293f
C8890 XA.XIR[4].XIC[1].icell.Ien VGND 0.37144f
C8891 XA.XIR[4].XIC[0].icell.SM VGND 0.00502f
C8892 XA.XIR[4].XIC[1].icell.PUM VGND 0.00293f
C8893 XA.XIR[4].XIC[0].icell.Ien VGND 0.37178f
C8894 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01044f
C8895 XA.XIR[4].XIC[0].icell.PUM VGND 0.00516f
C8896 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57336f
C8897 XA.XIR[4].XIC_dummy_left.icell.PUM VGND 0.00215f
C8898 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C8899 XA.XIR[4].XIC_15.icell.PDM VGND 0.18855f
C8900 XA.XIR[4].XIC[14].icell.PDM VGND 0.18809f
C8901 XA.XIR[4].XIC[13].icell.PDM VGND 0.18809f
C8902 XA.XIR[4].XIC[12].icell.PDM VGND 0.18809f
C8903 XA.XIR[4].XIC[11].icell.PDM VGND 0.18809f
C8904 XA.XIR[4].XIC[10].icell.PDM VGND 0.18809f
C8905 XA.XIR[4].XIC[9].icell.PDM VGND 0.18809f
C8906 XA.XIR[4].XIC[8].icell.PDM VGND 0.18809f
C8907 XA.XIR[4].XIC[7].icell.PDM VGND 0.18809f
C8908 XA.XIR[4].XIC[6].icell.PDM VGND 0.18809f
C8909 XA.XIR[4].XIC[5].icell.PDM VGND 0.18809f
C8910 XA.XIR[4].XIC[4].icell.PDM VGND 0.18809f
C8911 XA.XIR[4].XIC[3].icell.PDM VGND 0.18809f
C8912 XA.XIR[4].XIC[2].icell.PDM VGND 0.18809f
C8913 XA.XIR[4].XIC[1].icell.PDM VGND 0.18809f
C8914 XA.XIR[4].XIC[0].icell.PDM VGND 0.18817f
C8915 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C8916 XThR.Tn[4] VGND 14.03736f
C8917 a_n1049_6405# VGND 0.02935f
C8918 a_n1319_6405# VGND 0.00166f
C8919 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85795f
C8920 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C8921 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60802f
C8922 XA.XIR[3].XIC_15.icell.SM VGND 0.00474f
C8923 XA.XIR[3].XIC_dummy_right.icell.PUM VGND 0.00215f
C8924 XA.XIR[3].XIC_15.icell.Ien VGND 0.37063f
C8925 XA.XIR[3].XIC[14].icell.SM VGND 0.00502f
C8926 XA.XIR[3].XIC_15.icell.PUM VGND 0.00282f
C8927 XA.XIR[3].XIC[14].icell.Ien VGND 0.37144f
C8928 XA.XIR[3].XIC[13].icell.SM VGND 0.00502f
C8929 XA.XIR[3].XIC[14].icell.PUM VGND 0.00293f
C8930 XA.XIR[3].XIC[13].icell.Ien VGND 0.37144f
C8931 XA.XIR[3].XIC[12].icell.SM VGND 0.00502f
C8932 XA.XIR[3].XIC[13].icell.PUM VGND 0.00293f
C8933 XA.XIR[3].XIC[12].icell.Ien VGND 0.37144f
C8934 XA.XIR[3].XIC[11].icell.SM VGND 0.00502f
C8935 XA.XIR[3].XIC[12].icell.PUM VGND 0.00293f
C8936 XA.XIR[3].XIC[11].icell.Ien VGND 0.37144f
C8937 XA.XIR[3].XIC[10].icell.SM VGND 0.00502f
C8938 XA.XIR[3].XIC[11].icell.PUM VGND 0.00293f
C8939 XA.XIR[3].XIC[10].icell.Ien VGND 0.37144f
C8940 XA.XIR[3].XIC[9].icell.SM VGND 0.00502f
C8941 XA.XIR[3].XIC[10].icell.PUM VGND 0.00293f
C8942 XA.XIR[3].XIC[9].icell.Ien VGND 0.37144f
C8943 XA.XIR[3].XIC[8].icell.SM VGND 0.00502f
C8944 XA.XIR[3].XIC[9].icell.PUM VGND 0.00293f
C8945 XA.XIR[3].XIC[8].icell.Ien VGND 0.37144f
C8946 XA.XIR[3].XIC[7].icell.SM VGND 0.00502f
C8947 XA.XIR[3].XIC[8].icell.PUM VGND 0.00293f
C8948 XA.XIR[3].XIC[7].icell.Ien VGND 0.37144f
C8949 XA.XIR[3].XIC[6].icell.SM VGND 0.00502f
C8950 XA.XIR[3].XIC[7].icell.PUM VGND 0.00293f
C8951 XA.XIR[3].XIC[6].icell.Ien VGND 0.37144f
C8952 XA.XIR[3].XIC[5].icell.SM VGND 0.00502f
C8953 XA.XIR[3].XIC[6].icell.PUM VGND 0.00293f
C8954 XA.XIR[3].XIC[5].icell.Ien VGND 0.37144f
C8955 XA.XIR[3].XIC[4].icell.SM VGND 0.00502f
C8956 XA.XIR[3].XIC[5].icell.PUM VGND 0.00293f
C8957 XA.XIR[3].XIC[4].icell.Ien VGND 0.37144f
C8958 XA.XIR[3].XIC[3].icell.SM VGND 0.00502f
C8959 XA.XIR[3].XIC[4].icell.PUM VGND 0.00293f
C8960 XA.XIR[3].XIC[3].icell.Ien VGND 0.37144f
C8961 XA.XIR[3].XIC[2].icell.SM VGND 0.00502f
C8962 XA.XIR[3].XIC[3].icell.PUM VGND 0.00293f
C8963 XA.XIR[3].XIC[2].icell.Ien VGND 0.37144f
C8964 XA.XIR[3].XIC[1].icell.SM VGND 0.00502f
C8965 XThR.XTB5.Y VGND 1.32753f
C8966 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80611f
C8967 XA.XIR[3].XIC[2].icell.PUM VGND 0.00293f
C8968 XA.XIR[3].XIC[1].icell.Ien VGND 0.37144f
C8969 XA.XIR[3].XIC[0].icell.SM VGND 0.00502f
C8970 XA.XIR[3].XIC[1].icell.PUM VGND 0.00293f
C8971 XA.XIR[3].XIC[0].icell.Ien VGND 0.37178f
C8972 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01044f
C8973 XA.XIR[3].XIC[0].icell.PUM VGND 0.00516f
C8974 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57425f
C8975 a_n1049_6699# VGND 0.02979f
C8976 XA.XIR[3].XIC_dummy_left.icell.PUM VGND 0.00215f
C8977 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C8978 XA.XIR[3].XIC_15.icell.PDM VGND 0.18855f
C8979 XA.XIR[3].XIC[14].icell.PDM VGND 0.18809f
C8980 XA.XIR[3].XIC[13].icell.PDM VGND 0.18809f
C8981 XA.XIR[3].XIC[12].icell.PDM VGND 0.18809f
C8982 XA.XIR[3].XIC[11].icell.PDM VGND 0.18809f
C8983 XA.XIR[3].XIC[10].icell.PDM VGND 0.18809f
C8984 XA.XIR[3].XIC[9].icell.PDM VGND 0.18809f
C8985 XA.XIR[3].XIC[8].icell.PDM VGND 0.18809f
C8986 XA.XIR[3].XIC[7].icell.PDM VGND 0.18809f
C8987 XA.XIR[3].XIC[6].icell.PDM VGND 0.18809f
C8988 XA.XIR[3].XIC[5].icell.PDM VGND 0.18809f
C8989 XA.XIR[3].XIC[4].icell.PDM VGND 0.18809f
C8990 XA.XIR[3].XIC[3].icell.PDM VGND 0.18809f
C8991 XA.XIR[3].XIC[2].icell.PDM VGND 0.18809f
C8992 XA.XIR[3].XIC[1].icell.PDM VGND 0.18809f
C8993 XA.XIR[3].XIC[0].icell.PDM VGND 0.18817f
C8994 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C8995 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85795f
C8996 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C8997 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60802f
C8998 XA.XIR[2].XIC_15.icell.SM VGND 0.00474f
C8999 XA.XIR[2].XIC_dummy_right.icell.PUM VGND 0.00215f
C9000 XA.XIR[2].XIC_15.icell.Ien VGND 0.37063f
C9001 XA.XIR[2].XIC[14].icell.SM VGND 0.00502f
C9002 XA.XIR[2].XIC_15.icell.PUM VGND 0.00282f
C9003 XA.XIR[2].XIC[14].icell.Ien VGND 0.37144f
C9004 XA.XIR[2].XIC[13].icell.SM VGND 0.00502f
C9005 XA.XIR[2].XIC[14].icell.PUM VGND 0.00293f
C9006 XA.XIR[2].XIC[13].icell.Ien VGND 0.37144f
C9007 XA.XIR[2].XIC[12].icell.SM VGND 0.00502f
C9008 XA.XIR[2].XIC[13].icell.PUM VGND 0.00293f
C9009 XA.XIR[2].XIC[12].icell.Ien VGND 0.37144f
C9010 XA.XIR[2].XIC[11].icell.SM VGND 0.00502f
C9011 XA.XIR[2].XIC[12].icell.PUM VGND 0.00293f
C9012 XA.XIR[2].XIC[11].icell.Ien VGND 0.37144f
C9013 XA.XIR[2].XIC[10].icell.SM VGND 0.00502f
C9014 XA.XIR[2].XIC[11].icell.PUM VGND 0.00293f
C9015 XA.XIR[2].XIC[10].icell.Ien VGND 0.37144f
C9016 XA.XIR[2].XIC[9].icell.SM VGND 0.00502f
C9017 XA.XIR[2].XIC[10].icell.PUM VGND 0.00293f
C9018 XA.XIR[2].XIC[9].icell.Ien VGND 0.37144f
C9019 XA.XIR[2].XIC[8].icell.SM VGND 0.00502f
C9020 XA.XIR[2].XIC[9].icell.PUM VGND 0.00293f
C9021 XA.XIR[2].XIC[8].icell.Ien VGND 0.37144f
C9022 XA.XIR[2].XIC[7].icell.SM VGND 0.00502f
C9023 XA.XIR[2].XIC[8].icell.PUM VGND 0.00293f
C9024 XA.XIR[2].XIC[7].icell.Ien VGND 0.37144f
C9025 XA.XIR[2].XIC[6].icell.SM VGND 0.00502f
C9026 XA.XIR[2].XIC[7].icell.PUM VGND 0.00293f
C9027 XA.XIR[2].XIC[6].icell.Ien VGND 0.37144f
C9028 XA.XIR[2].XIC[5].icell.SM VGND 0.00502f
C9029 XA.XIR[2].XIC[6].icell.PUM VGND 0.00293f
C9030 XA.XIR[2].XIC[5].icell.Ien VGND 0.37144f
C9031 XA.XIR[2].XIC[4].icell.SM VGND 0.00502f
C9032 XA.XIR[2].XIC[5].icell.PUM VGND 0.00293f
C9033 XA.XIR[2].XIC[4].icell.Ien VGND 0.37144f
C9034 XA.XIR[2].XIC[3].icell.SM VGND 0.00502f
C9035 XA.XIR[2].XIC[4].icell.PUM VGND 0.00293f
C9036 XA.XIR[2].XIC[3].icell.Ien VGND 0.37144f
C9037 XA.XIR[2].XIC[2].icell.SM VGND 0.00502f
C9038 XA.XIR[2].XIC[3].icell.PUM VGND 0.00293f
C9039 XA.XIR[2].XIC[2].icell.Ien VGND 0.37144f
C9040 XA.XIR[2].XIC[1].icell.SM VGND 0.00502f
C9041 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80825f
C9042 XA.XIR[2].XIC[2].icell.PUM VGND 0.00293f
C9043 XA.XIR[2].XIC[1].icell.Ien VGND 0.37144f
C9044 XA.XIR[2].XIC[0].icell.SM VGND 0.00502f
C9045 XThR.Tn[3] VGND 13.98256f
C9046 XThR.XTB4.Y VGND 1.76953f
C9047 XA.XIR[2].XIC[1].icell.PUM VGND 0.00293f
C9048 XA.XIR[2].XIC[0].icell.Ien VGND 0.37178f
C9049 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01044f
C9050 XA.XIR[2].XIC[0].icell.PUM VGND 0.00516f
C9051 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57559f
C9052 a_n1335_7243# VGND 0.00179f
C9053 XA.XIR[2].XIC_dummy_left.icell.PUM VGND 0.00215f
C9054 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C9055 XA.XIR[2].XIC_15.icell.PDM VGND 0.18855f
C9056 XA.XIR[2].XIC[14].icell.PDM VGND 0.18809f
C9057 XA.XIR[2].XIC[13].icell.PDM VGND 0.18809f
C9058 XA.XIR[2].XIC[12].icell.PDM VGND 0.18809f
C9059 XA.XIR[2].XIC[11].icell.PDM VGND 0.18809f
C9060 XA.XIR[2].XIC[10].icell.PDM VGND 0.18809f
C9061 XA.XIR[2].XIC[9].icell.PDM VGND 0.18809f
C9062 XA.XIR[2].XIC[8].icell.PDM VGND 0.18809f
C9063 XA.XIR[2].XIC[7].icell.PDM VGND 0.18809f
C9064 XA.XIR[2].XIC[6].icell.PDM VGND 0.18809f
C9065 XA.XIR[2].XIC[5].icell.PDM VGND 0.18809f
C9066 XA.XIR[2].XIC[4].icell.PDM VGND 0.18809f
C9067 XA.XIR[2].XIC[3].icell.PDM VGND 0.18809f
C9068 XA.XIR[2].XIC[2].icell.PDM VGND 0.18809f
C9069 XA.XIR[2].XIC[1].icell.PDM VGND 0.18809f
C9070 XA.XIR[2].XIC[0].icell.PDM VGND 0.18817f
C9071 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C9072 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85795f
C9073 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C9074 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60802f
C9075 XA.XIR[1].XIC_15.icell.SM VGND 0.00474f
C9076 XA.XIR[1].XIC_dummy_right.icell.PUM VGND 0.00215f
C9077 XA.XIR[1].XIC_15.icell.Ien VGND 0.37063f
C9078 XA.XIR[1].XIC[14].icell.SM VGND 0.00502f
C9079 XA.XIR[1].XIC_15.icell.PUM VGND 0.00282f
C9080 XA.XIR[1].XIC[14].icell.Ien VGND 0.37144f
C9081 XA.XIR[1].XIC[13].icell.SM VGND 0.00502f
C9082 XA.XIR[1].XIC[14].icell.PUM VGND 0.00293f
C9083 XA.XIR[1].XIC[13].icell.Ien VGND 0.37144f
C9084 XA.XIR[1].XIC[12].icell.SM VGND 0.00502f
C9085 XA.XIR[1].XIC[13].icell.PUM VGND 0.00293f
C9086 XA.XIR[1].XIC[12].icell.Ien VGND 0.37144f
C9087 XA.XIR[1].XIC[11].icell.SM VGND 0.00502f
C9088 XA.XIR[1].XIC[12].icell.PUM VGND 0.00293f
C9089 XA.XIR[1].XIC[11].icell.Ien VGND 0.37144f
C9090 XA.XIR[1].XIC[10].icell.SM VGND 0.00502f
C9091 XA.XIR[1].XIC[11].icell.PUM VGND 0.00293f
C9092 XA.XIR[1].XIC[10].icell.Ien VGND 0.37144f
C9093 XA.XIR[1].XIC[9].icell.SM VGND 0.00502f
C9094 XA.XIR[1].XIC[10].icell.PUM VGND 0.00293f
C9095 XA.XIR[1].XIC[9].icell.Ien VGND 0.37144f
C9096 XA.XIR[1].XIC[8].icell.SM VGND 0.00502f
C9097 XA.XIR[1].XIC[9].icell.PUM VGND 0.00293f
C9098 XA.XIR[1].XIC[8].icell.Ien VGND 0.37144f
C9099 XA.XIR[1].XIC[7].icell.SM VGND 0.00502f
C9100 XA.XIR[1].XIC[8].icell.PUM VGND 0.00293f
C9101 XA.XIR[1].XIC[7].icell.Ien VGND 0.37144f
C9102 XA.XIR[1].XIC[6].icell.SM VGND 0.00502f
C9103 XA.XIR[1].XIC[7].icell.PUM VGND 0.00293f
C9104 XA.XIR[1].XIC[6].icell.Ien VGND 0.37144f
C9105 XA.XIR[1].XIC[5].icell.SM VGND 0.00502f
C9106 XA.XIR[1].XIC[6].icell.PUM VGND 0.00293f
C9107 XA.XIR[1].XIC[5].icell.Ien VGND 0.37144f
C9108 XA.XIR[1].XIC[4].icell.SM VGND 0.00502f
C9109 XA.XIR[1].XIC[5].icell.PUM VGND 0.00293f
C9110 XA.XIR[1].XIC[4].icell.Ien VGND 0.37144f
C9111 XA.XIR[1].XIC[3].icell.SM VGND 0.00502f
C9112 XA.XIR[1].XIC[4].icell.PUM VGND 0.00293f
C9113 XA.XIR[1].XIC[3].icell.Ien VGND 0.37144f
C9114 XA.XIR[1].XIC[2].icell.SM VGND 0.00502f
C9115 XA.XIR[1].XIC[3].icell.PUM VGND 0.00293f
C9116 XA.XIR[1].XIC[2].icell.Ien VGND 0.37144f
C9117 XA.XIR[1].XIC[1].icell.SM VGND 0.00502f
C9118 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80611f
C9119 XA.XIR[1].XIC[2].icell.PUM VGND 0.00293f
C9120 XA.XIR[1].XIC[1].icell.Ien VGND 0.37144f
C9121 XA.XIR[1].XIC[0].icell.SM VGND 0.00502f
C9122 XThR.Tn[2] VGND 14.03476f
C9123 a_n1049_7493# VGND 0.02484f
C9124 XThR.XTB3.Y VGND 2.09162f
C9125 XThR.XTB7.A VGND 1.95537f
C9126 XA.XIR[1].XIC[1].icell.PUM VGND 0.00293f
C9127 XA.XIR[1].XIC[0].icell.Ien VGND 0.37178f
C9128 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01044f
C9129 XA.XIR[1].XIC[0].icell.PUM VGND 0.00516f
C9130 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57378f
C9131 XA.XIR[1].XIC_dummy_left.icell.PUM VGND 0.00215f
C9132 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C9133 XA.XIR[1].XIC_15.icell.PDM VGND 0.18855f
C9134 XA.XIR[1].XIC[14].icell.PDM VGND 0.18809f
C9135 XA.XIR[1].XIC[13].icell.PDM VGND 0.18809f
C9136 XA.XIR[1].XIC[12].icell.PDM VGND 0.18809f
C9137 XA.XIR[1].XIC[11].icell.PDM VGND 0.18809f
C9138 XA.XIR[1].XIC[10].icell.PDM VGND 0.18809f
C9139 XA.XIR[1].XIC[9].icell.PDM VGND 0.18809f
C9140 XA.XIR[1].XIC[8].icell.PDM VGND 0.18809f
C9141 XA.XIR[1].XIC[7].icell.PDM VGND 0.18809f
C9142 XA.XIR[1].XIC[6].icell.PDM VGND 0.18809f
C9143 XA.XIR[1].XIC[5].icell.PDM VGND 0.18809f
C9144 XA.XIR[1].XIC[4].icell.PDM VGND 0.18809f
C9145 XA.XIR[1].XIC[3].icell.PDM VGND 0.18809f
C9146 XA.XIR[1].XIC[2].icell.PDM VGND 0.18809f
C9147 XA.XIR[1].XIC[1].icell.PDM VGND 0.18809f
C9148 XA.XIR[1].XIC[0].icell.PDM VGND 0.18817f
C9149 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C9150 a_n1049_7787# VGND 0.03396f
C9151 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87409f
C9152 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C9153 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61781f
C9154 XA.XIR[0].XIC_15.icell.SM VGND 0.00474f
C9155 XA.XIR[0].XIC_dummy_right.icell.PUM VGND 0.00207f
C9156 XA.XIR[0].XIC_15.icell.Ien VGND 0.37673f
C9157 XA.XIR[0].XIC[14].icell.SM VGND 0.00624f
C9158 XA.XIR[0].XIC_15.icell.PUM VGND 0.00468f
C9159 XA.XIR[0].XIC[14].icell.Ien VGND 0.38432f
C9160 XA.XIR[0].XIC[13].icell.SM VGND 0.00624f
C9161 XA.XIR[0].XIC[14].icell.PUM VGND 0.00392f
C9162 XA.XIR[0].XIC[13].icell.Ien VGND 0.38436f
C9163 XA.XIR[0].XIC[12].icell.SM VGND 0.00624f
C9164 XA.XIR[0].XIC[13].icell.PUM VGND 0.00397f
C9165 XA.XIR[0].XIC[12].icell.Ien VGND 0.381f
C9166 XA.XIR[0].XIC[11].icell.SM VGND 0.00624f
C9167 XA.XIR[0].XIC[12].icell.PUM VGND 0.00392f
C9168 XA.XIR[0].XIC[11].icell.Ien VGND 0.38167f
C9169 XA.XIR[0].XIC[10].icell.SM VGND 0.00624f
C9170 XA.XIR[0].XIC[11].icell.PUM VGND 0.00392f
C9171 XA.XIR[0].XIC[10].icell.Ien VGND 0.38301f
C9172 XA.XIR[0].XIC[9].icell.SM VGND 0.00624f
C9173 XA.XIR[0].XIC[10].icell.PUM VGND 0.00392f
C9174 XA.XIR[0].XIC[9].icell.Ien VGND 0.38128f
C9175 XA.XIR[0].XIC[8].icell.SM VGND 0.00624f
C9176 XA.XIR[0].XIC[9].icell.PUM VGND 0.00392f
C9177 XA.XIR[0].XIC[8].icell.Ien VGND 0.38176f
C9178 XA.XIR[0].XIC[7].icell.SM VGND 0.00624f
C9179 XA.XIR[0].XIC[8].icell.PUM VGND 0.00392f
C9180 XA.XIR[0].XIC[7].icell.Ien VGND 0.382f
C9181 XA.XIR[0].XIC[6].icell.SM VGND 0.00624f
C9182 XA.XIR[0].XIC[7].icell.PUM VGND 0.00392f
C9183 XA.XIR[0].XIC[6].icell.Ien VGND 0.38192f
C9184 XA.XIR[0].XIC[5].icell.SM VGND 0.00624f
C9185 XA.XIR[0].XIC[6].icell.PUM VGND 0.00403f
C9186 XA.XIR[0].XIC[5].icell.Ien VGND 0.38091f
C9187 XA.XIR[0].XIC[4].icell.SM VGND 0.00624f
C9188 XA.XIR[0].XIC[5].icell.PUM VGND 0.00392f
C9189 XA.XIR[0].XIC[4].icell.Ien VGND 0.38104f
C9190 XA.XIR[0].XIC[3].icell.SM VGND 0.00624f
C9191 XA.XIR[0].XIC[4].icell.PUM VGND 0.00392f
C9192 XA.XIR[0].XIC[3].icell.Ien VGND 0.38229f
C9193 XA.XIR[0].XIC[2].icell.SM VGND 0.00624f
C9194 XA.XIR[0].XIC[3].icell.PUM VGND 0.00392f
C9195 XA.XIR[0].XIC[2].icell.Ien VGND 0.38432f
C9196 XA.XIR[0].XIC[1].icell.SM VGND 0.00624f
C9197 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.841f
C9198 XA.XIR[0].XIC[2].icell.PUM VGND 0.00392f
C9199 XA.XIR[0].XIC[1].icell.Ien VGND 0.38432f
C9200 XA.XIR[0].XIC[0].icell.SM VGND 0.00624f
C9201 XA.XIR[0].XIC[1].icell.PUM VGND 0.00394f
C9202 XA.XIR[0].XIC[0].icell.Ien VGND 0.38446f
C9203 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01044f
C9204 XThR.Tn[1] VGND 14.06925f
C9205 a_n1335_8107# VGND 0.00163f
C9206 XThR.XTB2.Y VGND 1.47668f
C9207 XThR.XTB6.A VGND 0.95641f
C9208 XA.XIR[0].XIC[0].icell.PUM VGND 0.00623f
C9209 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58675f
C9210 XA.XIR[0].XIC_dummy_left.icell.PUM VGND 0.0035f
C9211 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.25101f
C9212 XA.XIR[0].XIC_15.icell.PDM VGND 0.20765f
C9213 XA.XIR[0].XIC[14].icell.PDM VGND 0.24599f
C9214 XA.XIR[0].XIC[13].icell.PDM VGND 0.24583f
C9215 XA.XIR[0].XIC[12].icell.PDM VGND 0.24144f
C9216 XA.XIR[0].XIC[11].icell.PDM VGND 0.24182f
C9217 XA.XIR[0].XIC[10].icell.PDM VGND 0.24172f
C9218 XA.XIR[0].XIC[9].icell.PDM VGND 0.24144f
C9219 XA.XIR[0].XIC[8].icell.PDM VGND 0.24144f
C9220 XA.XIR[0].XIC[7].icell.PDM VGND 0.24388f
C9221 XA.XIR[0].XIC[6].icell.PDM VGND 0.24108f
C9222 XA.XIR[0].XIC[5].icell.PDM VGND 0.24297f
C9223 XA.XIR[0].XIC[4].icell.PDM VGND 0.24156f
C9224 XA.XIR[0].XIC[3].icell.PDM VGND 0.24455f
C9225 XA.XIR[0].XIC[2].icell.PDM VGND 0.24578f
C9226 XA.XIR[0].XIC[1].icell.PDM VGND 0.24578f
C9227 XA.XIR[0].XIC[0].icell.PDM VGND 0.24491f
C9228 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24713f
C9229 a_n1335_8331# VGND 0.00203f
C9230 XThR.Tn[0] VGND 14.40644f
C9231 a_n1049_8581# VGND 0.04324f
C9232 XThR.XTBN.Y VGND 7.54172f
C9233 XThR.XTB1.Y VGND 1.81265f
C9234 XThR.XTB7.B VGND 2.61156f
C9235 XThR.XTB5.A VGND 1.76044f
C9236 XThC.Tn[14] VGND 9.98563f
C9237 XThC.Tn[13] VGND 9.79145f
C9238 XThC.Tn[12] VGND 9.63534f
C9239 XThC.Tn[11] VGND 9.46598f
C9240 XThC.Tn[10] VGND 9.29745f
C9241 XThC.Tn[9] VGND 9.27278f
C9242 XThC.Tn[8] VGND 9.24802f
C9243 a_10915_9569# VGND 0.55837f
C9244 a_10051_9569# VGND 0.55761f
C9245 a_9827_9569# VGND 0.54461f
C9246 a_8963_9569# VGND 0.55448f
C9247 a_8739_9569# VGND 0.55288f
C9248 a_7875_9569# VGND 0.55432f
C9249 a_7651_9569# VGND 0.55717f
C9250 XThC.Tn[7] VGND 10.56205f
C9251 XThC.Tn[6] VGND 10.35711f
C9252 XThC.Tn[5] VGND 10.62787f
C9253 XThC.Tn[4] VGND 10.6808f
C9254 XThC.Tn[3] VGND 9.9249f
C9255 XThC.Tn[2] VGND 10.4557f
C9256 XThC.Tn[1] VGND 10.33149f
C9257 XThC.Tn[0] VGND 10.74903f
C9258 a_6243_9615# VGND 0.0299f
C9259 a_5949_9615# VGND 0.03432f
C9260 a_5155_9615# VGND 0.03615f
C9261 a_4861_9615# VGND 0.03632f
C9262 a_4067_9615# VGND 0.03071f
C9263 a_3773_9615# VGND 0.03867f
C9264 a_2979_9615# VGND 0.04107f
C9265 a_8739_10571# VGND 0.00194f
C9266 XThC.XTBN.Y VGND 7.90394f
C9267 XThC.XTB7.Y VGND 1.36247f
C9268 XThC.XTB6.Y VGND 1.3829f
C9269 a_5155_10571# VGND 0.00165f
C9270 XThC.XTB7.B VGND 2.73083f
C9271 XThC.XTB5.Y VGND 1.32591f
C9272 XThC.XTBN.A VGND 1.23171f
C9273 a_4387_10575# VGND 0.00179f
C9274 a_3523_10575# VGND 0.00163f
C9275 a_3299_10575# VGND 0.00202f
C9276 XThC.XTB4.Y VGND 1.69875f
C9277 XThC.XTB3.Y VGND 1.96765f
C9278 XThC.XTB7.A VGND 1.96056f
C9279 XThC.XTB6.A VGND 0.95757f
C9280 XThC.XTB2.Y VGND 1.47589f
C9281 XThC.XTB1.Y VGND 1.77676f
C9282 XThC.XTB5.A VGND 1.75974f
C9283 XThR.XTB3.Y.t1 VGND 0.06176f
C9284 XThR.XTB3.Y.n0 VGND 0.01521f
C9285 XThR.XTB3.Y.t8 VGND 0.04903f
C9286 XThR.XTB3.Y.t15 VGND 0.02889f
C9287 XThR.XTB3.Y.t13 VGND 0.04903f
C9288 XThR.XTB3.Y.t6 VGND 0.02889f
C9289 XThR.XTB3.Y.t9 VGND 0.04903f
C9290 XThR.XTB3.Y.t17 VGND 0.02889f
C9291 XThR.XTB3.Y.n1 VGND 0.08226f
C9292 XThR.XTB3.Y.n2 VGND 0.08688f
C9293 XThR.XTB3.Y.n3 VGND 0.03573f
C9294 XThR.XTB3.Y.n4 VGND 0.0707f
C9295 XThR.XTB3.Y.t12 VGND 0.04903f
C9296 XThR.XTB3.Y.t4 VGND 0.02889f
C9297 XThR.XTB3.Y.n5 VGND 0.06608f
C9298 XThR.XTB3.Y.n6 VGND 0.03236f
C9299 XThR.XTB3.Y.n7 VGND 0.02685f
C9300 XThR.XTB3.Y.t18 VGND 0.04903f
C9301 XThR.XTB3.Y.t5 VGND 0.02889f
C9302 XThR.XTB3.Y.n8 VGND 0.03005f
C9303 XThR.XTB3.Y.t7 VGND 0.04903f
C9304 XThR.XTB3.Y.t10 VGND 0.02889f
C9305 XThR.XTB3.Y.n9 VGND 0.05992f
C9306 XThR.XTB3.Y.t11 VGND 0.04903f
C9307 XThR.XTB3.Y.t16 VGND 0.02889f
C9308 XThR.XTB3.Y.n10 VGND 0.06454f
C9309 XThR.XTB3.Y.n11 VGND 0.03645f
C9310 XThR.XTB3.Y.n12 VGND 0.06034f
C9311 XThR.XTB3.Y.n13 VGND 0.03128f
C9312 XThR.XTB3.Y.n14 VGND 0.02851f
C9313 XThR.XTB3.Y.n15 VGND 0.06454f
C9314 XThR.XTB3.Y.t14 VGND 0.04903f
C9315 XThR.XTB3.Y.t3 VGND 0.02889f
C9316 XThR.XTB3.Y.n16 VGND 0.05838f
C9317 XThR.XTB3.Y.n17 VGND 0.03236f
C9318 XThR.XTB3.Y.n18 VGND 0.04707f
C9319 XThR.XTB3.Y.n19 VGND 1.31347f
C9320 XThR.XTB3.Y.t2 VGND 0.03152f
C9321 XThR.XTB3.Y.t0 VGND 0.03152f
C9322 XThR.XTB3.Y.n20 VGND 0.06766f
C9323 XThR.XTB3.Y.n21 VGND 0.157f
C9324 XThR.XTB3.Y.n22 VGND 0.03296f
C9325 XThR.XTB1.Y.t1 VGND 0.03165f
C9326 XThR.XTB1.Y.n0 VGND 0.0078f
C9327 XThR.XTB1.Y.t8 VGND 0.02512f
C9328 XThR.XTB1.Y.t15 VGND 0.0148f
C9329 XThR.XTB1.Y.t14 VGND 0.02512f
C9330 XThR.XTB1.Y.t7 VGND 0.0148f
C9331 XThR.XTB1.Y.t10 VGND 0.02512f
C9332 XThR.XTB1.Y.t18 VGND 0.0148f
C9333 XThR.XTB1.Y.n1 VGND 0.04215f
C9334 XThR.XTB1.Y.n2 VGND 0.04452f
C9335 XThR.XTB1.Y.n3 VGND 0.01831f
C9336 XThR.XTB1.Y.n4 VGND 0.03623f
C9337 XThR.XTB1.Y.t13 VGND 0.02512f
C9338 XThR.XTB1.Y.t4 VGND 0.0148f
C9339 XThR.XTB1.Y.n5 VGND 0.03386f
C9340 XThR.XTB1.Y.n6 VGND 0.01658f
C9341 XThR.XTB1.Y.n7 VGND 0.01376f
C9342 XThR.XTB1.Y.t6 VGND 0.02512f
C9343 XThR.XTB1.Y.t11 VGND 0.0148f
C9344 XThR.XTB1.Y.n8 VGND 0.0154f
C9345 XThR.XTB1.Y.t12 VGND 0.02512f
C9346 XThR.XTB1.Y.t16 VGND 0.0148f
C9347 XThR.XTB1.Y.n9 VGND 0.0307f
C9348 XThR.XTB1.Y.t17 VGND 0.02512f
C9349 XThR.XTB1.Y.t5 VGND 0.0148f
C9350 XThR.XTB1.Y.n10 VGND 0.03307f
C9351 XThR.XTB1.Y.n11 VGND 0.01868f
C9352 XThR.XTB1.Y.n12 VGND 0.03092f
C9353 XThR.XTB1.Y.n13 VGND 0.01603f
C9354 XThR.XTB1.Y.n14 VGND 0.01461f
C9355 XThR.XTB1.Y.n15 VGND 0.03307f
C9356 XThR.XTB1.Y.t3 VGND 0.02512f
C9357 XThR.XTB1.Y.t9 VGND 0.0148f
C9358 XThR.XTB1.Y.n16 VGND 0.02991f
C9359 XThR.XTB1.Y.n17 VGND 0.01658f
C9360 XThR.XTB1.Y.n18 VGND 0.02412f
C9361 XThR.XTB1.Y.n19 VGND 0.75219f
C9362 XThR.XTB1.Y.t2 VGND 0.01615f
C9363 XThR.XTB1.Y.t0 VGND 0.01615f
C9364 XThR.XTB1.Y.n20 VGND 0.03467f
C9365 XThR.XTB1.Y.n21 VGND 0.08068f
C9366 XThR.XTB1.Y.n22 VGND 0.01689f
C9367 XThR.XTB4.Y.t8 VGND 0.02956f
C9368 XThR.XTB4.Y.t15 VGND 0.05016f
C9369 XThR.XTB4.Y.t16 VGND 0.02956f
C9370 XThR.XTB4.Y.t5 VGND 0.05016f
C9371 XThR.XTB4.Y.t10 VGND 0.02956f
C9372 XThR.XTB4.Y.t17 VGND 0.05016f
C9373 XThR.XTB4.Y.n0 VGND 0.08416f
C9374 XThR.XTB4.Y.n1 VGND 0.08889f
C9375 XThR.XTB4.Y.n2 VGND 0.03656f
C9376 XThR.XTB4.Y.n3 VGND 0.07234f
C9377 XThR.XTB4.Y.t13 VGND 0.02956f
C9378 XThR.XTB4.Y.t4 VGND 0.05016f
C9379 XThR.XTB4.Y.n4 VGND 0.06761f
C9380 XThR.XTB4.Y.n5 VGND 0.0331f
C9381 XThR.XTB4.Y.n6 VGND 0.01685f
C9382 XThR.XTB4.Y.n7 VGND 0.05355f
C9383 XThR.XTB4.Y.n8 VGND 0.64921f
C9384 XThR.XTB4.Y.t14 VGND 0.02956f
C9385 XThR.XTB4.Y.t7 VGND 0.05016f
C9386 XThR.XTB4.Y.n9 VGND 0.03074f
C9387 XThR.XTB4.Y.t3 VGND 0.02956f
C9388 XThR.XTB4.Y.t12 VGND 0.05016f
C9389 XThR.XTB4.Y.n10 VGND 0.0613f
C9390 XThR.XTB4.Y.t9 VGND 0.02956f
C9391 XThR.XTB4.Y.t2 VGND 0.05016f
C9392 XThR.XTB4.Y.n11 VGND 0.06603f
C9393 XThR.XTB4.Y.n12 VGND 0.03729f
C9394 XThR.XTB4.Y.n13 VGND 0.06174f
C9395 XThR.XTB4.Y.n14 VGND 0.03201f
C9396 XThR.XTB4.Y.n15 VGND 0.02916f
C9397 XThR.XTB4.Y.n16 VGND 0.06603f
C9398 XThR.XTB4.Y.t11 VGND 0.02956f
C9399 XThR.XTB4.Y.t6 VGND 0.05016f
C9400 XThR.XTB4.Y.n17 VGND 0.05972f
C9401 XThR.XTB4.Y.n18 VGND 0.0331f
C9402 XThR.XTB4.Y.n19 VGND 0.05647f
C9403 XThR.XTB4.Y.n20 VGND 1.3092f
C9404 XThR.XTB4.Y.t1 VGND 0.06491f
C9405 XThR.XTB4.Y.n21 VGND 0.12281f
C9406 XThR.XTB4.Y.n22 VGND 0.02892f
C9407 XThR.XTB4.Y.t0 VGND 0.11919f
C9408 XThR.Tn[13].t9 VGND 0.02397f
C9409 XThR.Tn[13].t11 VGND 0.02397f
C9410 XThR.Tn[13].n0 VGND 0.07277f
C9411 XThR.Tn[13].t10 VGND 0.02397f
C9412 XThR.Tn[13].t8 VGND 0.02397f
C9413 XThR.Tn[13].n1 VGND 0.05327f
C9414 XThR.Tn[13].n2 VGND 0.24224f
C9415 XThR.Tn[13].t7 VGND 0.01558f
C9416 XThR.Tn[13].t5 VGND 0.01558f
C9417 XThR.Tn[13].n3 VGND 0.03885f
C9418 XThR.Tn[13].t6 VGND 0.01558f
C9419 XThR.Tn[13].t4 VGND 0.01558f
C9420 XThR.Tn[13].n4 VGND 0.03116f
C9421 XThR.Tn[13].n5 VGND 0.07837f
C9422 XThR.Tn[13].t72 VGND 0.01873f
C9423 XThR.Tn[13].t64 VGND 0.02051f
C9424 XThR.Tn[13].n6 VGND 0.05008f
C9425 XThR.Tn[13].n7 VGND 0.09621f
C9426 XThR.Tn[13].t28 VGND 0.01873f
C9427 XThR.Tn[13].t21 VGND 0.02051f
C9428 XThR.Tn[13].n8 VGND 0.05008f
C9429 XThR.Tn[13].t44 VGND 0.01867f
C9430 XThR.Tn[13].t12 VGND 0.02044f
C9431 XThR.Tn[13].n9 VGND 0.05211f
C9432 XThR.Tn[13].n10 VGND 0.03661f
C9433 XThR.Tn[13].n11 VGND 0.00669f
C9434 XThR.Tn[13].n12 VGND 0.11748f
C9435 XThR.Tn[13].t65 VGND 0.01873f
C9436 XThR.Tn[13].t57 VGND 0.02051f
C9437 XThR.Tn[13].n13 VGND 0.05008f
C9438 XThR.Tn[13].t19 VGND 0.01867f
C9439 XThR.Tn[13].t52 VGND 0.02044f
C9440 XThR.Tn[13].n14 VGND 0.05211f
C9441 XThR.Tn[13].n15 VGND 0.03661f
C9442 XThR.Tn[13].n16 VGND 0.00669f
C9443 XThR.Tn[13].n17 VGND 0.11748f
C9444 XThR.Tn[13].t22 VGND 0.01873f
C9445 XThR.Tn[13].t14 VGND 0.02051f
C9446 XThR.Tn[13].n18 VGND 0.05008f
C9447 XThR.Tn[13].t34 VGND 0.01867f
C9448 XThR.Tn[13].t70 VGND 0.02044f
C9449 XThR.Tn[13].n19 VGND 0.05211f
C9450 XThR.Tn[13].n20 VGND 0.03661f
C9451 XThR.Tn[13].n21 VGND 0.00669f
C9452 XThR.Tn[13].n22 VGND 0.11748f
C9453 XThR.Tn[13].t49 VGND 0.01873f
C9454 XThR.Tn[13].t39 VGND 0.02051f
C9455 XThR.Tn[13].n23 VGND 0.05008f
C9456 XThR.Tn[13].t66 VGND 0.01867f
C9457 XThR.Tn[13].t35 VGND 0.02044f
C9458 XThR.Tn[13].n24 VGND 0.05211f
C9459 XThR.Tn[13].n25 VGND 0.03661f
C9460 XThR.Tn[13].n26 VGND 0.00669f
C9461 XThR.Tn[13].n27 VGND 0.11748f
C9462 XThR.Tn[13].t24 VGND 0.01873f
C9463 XThR.Tn[13].t16 VGND 0.02051f
C9464 XThR.Tn[13].n28 VGND 0.05008f
C9465 XThR.Tn[13].t37 VGND 0.01867f
C9466 XThR.Tn[13].t71 VGND 0.02044f
C9467 XThR.Tn[13].n29 VGND 0.05211f
C9468 XThR.Tn[13].n30 VGND 0.03661f
C9469 XThR.Tn[13].n31 VGND 0.00669f
C9470 XThR.Tn[13].n32 VGND 0.11748f
C9471 XThR.Tn[13].t60 VGND 0.01873f
C9472 XThR.Tn[13].t30 VGND 0.02051f
C9473 XThR.Tn[13].n33 VGND 0.05008f
C9474 XThR.Tn[13].t13 VGND 0.01867f
C9475 XThR.Tn[13].t26 VGND 0.02044f
C9476 XThR.Tn[13].n34 VGND 0.05211f
C9477 XThR.Tn[13].n35 VGND 0.03661f
C9478 XThR.Tn[13].n36 VGND 0.00669f
C9479 XThR.Tn[13].n37 VGND 0.11748f
C9480 XThR.Tn[13].t29 VGND 0.01873f
C9481 XThR.Tn[13].t25 VGND 0.02051f
C9482 XThR.Tn[13].n38 VGND 0.05008f
C9483 XThR.Tn[13].t43 VGND 0.01867f
C9484 XThR.Tn[13].t18 VGND 0.02044f
C9485 XThR.Tn[13].n39 VGND 0.05211f
C9486 XThR.Tn[13].n40 VGND 0.03661f
C9487 XThR.Tn[13].n41 VGND 0.00669f
C9488 XThR.Tn[13].n42 VGND 0.11748f
C9489 XThR.Tn[13].t32 VGND 0.01873f
C9490 XThR.Tn[13].t38 VGND 0.02051f
C9491 XThR.Tn[13].n43 VGND 0.05008f
C9492 XThR.Tn[13].t48 VGND 0.01867f
C9493 XThR.Tn[13].t33 VGND 0.02044f
C9494 XThR.Tn[13].n44 VGND 0.05211f
C9495 XThR.Tn[13].n45 VGND 0.03661f
C9496 XThR.Tn[13].n46 VGND 0.00669f
C9497 XThR.Tn[13].n47 VGND 0.11748f
C9498 XThR.Tn[13].t51 VGND 0.01873f
C9499 XThR.Tn[13].t59 VGND 0.02051f
C9500 XThR.Tn[13].n48 VGND 0.05008f
C9501 XThR.Tn[13].t68 VGND 0.01867f
C9502 XThR.Tn[13].t53 VGND 0.02044f
C9503 XThR.Tn[13].n49 VGND 0.05211f
C9504 XThR.Tn[13].n50 VGND 0.03661f
C9505 XThR.Tn[13].n51 VGND 0.00669f
C9506 XThR.Tn[13].n52 VGND 0.11748f
C9507 XThR.Tn[13].t41 VGND 0.01873f
C9508 XThR.Tn[13].t17 VGND 0.02051f
C9509 XThR.Tn[13].n53 VGND 0.05008f
C9510 XThR.Tn[13].t58 VGND 0.01867f
C9511 XThR.Tn[13].t73 VGND 0.02044f
C9512 XThR.Tn[13].n54 VGND 0.05211f
C9513 XThR.Tn[13].n55 VGND 0.03661f
C9514 XThR.Tn[13].n56 VGND 0.00669f
C9515 XThR.Tn[13].n57 VGND 0.11748f
C9516 XThR.Tn[13].t63 VGND 0.01873f
C9517 XThR.Tn[13].t55 VGND 0.02051f
C9518 XThR.Tn[13].n58 VGND 0.05008f
C9519 XThR.Tn[13].t15 VGND 0.01867f
C9520 XThR.Tn[13].t45 VGND 0.02044f
C9521 XThR.Tn[13].n59 VGND 0.05211f
C9522 XThR.Tn[13].n60 VGND 0.03661f
C9523 XThR.Tn[13].n61 VGND 0.00669f
C9524 XThR.Tn[13].n62 VGND 0.11748f
C9525 XThR.Tn[13].t31 VGND 0.01873f
C9526 XThR.Tn[13].t27 VGND 0.02051f
C9527 XThR.Tn[13].n63 VGND 0.05008f
C9528 XThR.Tn[13].t46 VGND 0.01867f
C9529 XThR.Tn[13].t20 VGND 0.02044f
C9530 XThR.Tn[13].n64 VGND 0.05211f
C9531 XThR.Tn[13].n65 VGND 0.03661f
C9532 XThR.Tn[13].n66 VGND 0.00669f
C9533 XThR.Tn[13].n67 VGND 0.11748f
C9534 XThR.Tn[13].t50 VGND 0.01873f
C9535 XThR.Tn[13].t40 VGND 0.02051f
C9536 XThR.Tn[13].n68 VGND 0.05008f
C9537 XThR.Tn[13].t67 VGND 0.01867f
C9538 XThR.Tn[13].t36 VGND 0.02044f
C9539 XThR.Tn[13].n69 VGND 0.05211f
C9540 XThR.Tn[13].n70 VGND 0.03661f
C9541 XThR.Tn[13].n71 VGND 0.00669f
C9542 XThR.Tn[13].n72 VGND 0.11748f
C9543 XThR.Tn[13].t69 VGND 0.01873f
C9544 XThR.Tn[13].t62 VGND 0.02051f
C9545 XThR.Tn[13].n73 VGND 0.05008f
C9546 XThR.Tn[13].t23 VGND 0.01867f
C9547 XThR.Tn[13].t54 VGND 0.02044f
C9548 XThR.Tn[13].n74 VGND 0.05211f
C9549 XThR.Tn[13].n75 VGND 0.03661f
C9550 XThR.Tn[13].n76 VGND 0.00669f
C9551 XThR.Tn[13].n77 VGND 0.11748f
C9552 XThR.Tn[13].t42 VGND 0.01873f
C9553 XThR.Tn[13].t56 VGND 0.02051f
C9554 XThR.Tn[13].n78 VGND 0.05008f
C9555 XThR.Tn[13].t61 VGND 0.01867f
C9556 XThR.Tn[13].t47 VGND 0.02044f
C9557 XThR.Tn[13].n79 VGND 0.05211f
C9558 XThR.Tn[13].n80 VGND 0.03661f
C9559 XThR.Tn[13].n81 VGND 0.00669f
C9560 XThR.Tn[13].n82 VGND 0.11748f
C9561 XThR.Tn[13].n83 VGND 0.10676f
C9562 XThR.Tn[13].n84 VGND 0.41858f
C9563 XThR.Tn[13].t2 VGND 0.02397f
C9564 XThR.Tn[13].t0 VGND 0.02397f
C9565 XThR.Tn[13].n85 VGND 0.05178f
C9566 XThR.Tn[13].t3 VGND 0.02397f
C9567 XThR.Tn[13].t1 VGND 0.02397f
C9568 XThR.Tn[13].n86 VGND 0.07881f
C9569 XThR.Tn[13].n87 VGND 0.21883f
C9570 XThR.Tn[13].n88 VGND 0.0293f
C9571 XThC.XTB3.Y.t2 VGND 0.06296f
C9572 XThC.XTB3.Y.n0 VGND 0.04069f
C9573 XThC.XTB3.Y.n1 VGND 0.05192f
C9574 XThC.XTB3.Y.t1 VGND 0.03159f
C9575 XThC.XTB3.Y.t0 VGND 0.03159f
C9576 XThC.XTB3.Y.n2 VGND 0.06782f
C9577 XThC.XTB3.Y.t10 VGND 0.04914f
C9578 XThC.XTB3.Y.t17 VGND 0.02896f
C9579 XThC.XTB3.Y.n3 VGND 0.05852f
C9580 XThC.XTB3.Y.t14 VGND 0.04914f
C9581 XThC.XTB3.Y.t5 VGND 0.02896f
C9582 XThC.XTB3.Y.n4 VGND 0.03012f
C9583 XThC.XTB3.Y.t15 VGND 0.04914f
C9584 XThC.XTB3.Y.t6 VGND 0.02896f
C9585 XThC.XTB3.Y.n5 VGND 0.06469f
C9586 XThC.XTB3.Y.t3 VGND 0.04914f
C9587 XThC.XTB3.Y.t9 VGND 0.02896f
C9588 XThC.XTB3.Y.n6 VGND 0.06006f
C9589 XThC.XTB3.Y.n7 VGND 0.03654f
C9590 XThC.XTB3.Y.n8 VGND 0.06049f
C9591 XThC.XTB3.Y.n9 VGND 0.0234f
C9592 XThC.XTB3.Y.n10 VGND 0.02857f
C9593 XThC.XTB3.Y.n11 VGND 0.06469f
C9594 XThC.XTB3.Y.n12 VGND 0.03243f
C9595 XThC.XTB3.Y.n13 VGND 0.05514f
C9596 XThC.XTB3.Y.t16 VGND 0.04914f
C9597 XThC.XTB3.Y.t7 VGND 0.02896f
C9598 XThC.XTB3.Y.n14 VGND 0.06624f
C9599 XThC.XTB3.Y.t4 VGND 0.04914f
C9600 XThC.XTB3.Y.t13 VGND 0.02896f
C9601 XThC.XTB3.Y.t12 VGND 0.04914f
C9602 XThC.XTB3.Y.t18 VGND 0.02896f
C9603 XThC.XTB3.Y.t11 VGND 0.04914f
C9604 XThC.XTB3.Y.t8 VGND 0.02896f
C9605 XThC.XTB3.Y.n15 VGND 0.08245f
C9606 XThC.XTB3.Y.n16 VGND 0.08709f
C9607 XThC.XTB3.Y.n17 VGND 0.03356f
C9608 XThC.XTB3.Y.n18 VGND 0.07087f
C9609 XThC.XTB3.Y.n19 VGND 0.03243f
C9610 XThC.XTB3.Y.n20 VGND 0.02691f
C9611 XThC.XTB3.Y.n21 VGND 1.39635f
C9612 XThC.XTB3.Y.n22 VGND 0.14933f
C9613 XThR.Tn[8].t6 VGND 0.02415f
C9614 XThR.Tn[8].t4 VGND 0.02415f
C9615 XThR.Tn[8].n0 VGND 0.07334f
C9616 XThR.Tn[8].t7 VGND 0.02415f
C9617 XThR.Tn[8].t5 VGND 0.02415f
C9618 XThR.Tn[8].n1 VGND 0.05369f
C9619 XThR.Tn[8].n2 VGND 0.24415f
C9620 XThR.Tn[8].t8 VGND 0.02415f
C9621 XThR.Tn[8].t10 VGND 0.02415f
C9622 XThR.Tn[8].n3 VGND 0.05219f
C9623 XThR.Tn[8].t1 VGND 0.02415f
C9624 XThR.Tn[8].t9 VGND 0.02415f
C9625 XThR.Tn[8].n4 VGND 0.07943f
C9626 XThR.Tn[8].n5 VGND 0.22055f
C9627 XThR.Tn[8].n6 VGND 0.01087f
C9628 XThR.Tn[8].t39 VGND 0.01888f
C9629 XThR.Tn[8].t33 VGND 0.02067f
C9630 XThR.Tn[8].n7 VGND 0.05048f
C9631 XThR.Tn[8].n8 VGND 0.09697f
C9632 XThR.Tn[8].t59 VGND 0.01888f
C9633 XThR.Tn[8].t49 VGND 0.02067f
C9634 XThR.Tn[8].n9 VGND 0.05048f
C9635 XThR.Tn[8].t13 VGND 0.01882f
C9636 XThR.Tn[8].t45 VGND 0.02061f
C9637 XThR.Tn[8].n10 VGND 0.05252f
C9638 XThR.Tn[8].n11 VGND 0.0369f
C9639 XThR.Tn[8].n12 VGND 0.00675f
C9640 XThR.Tn[8].n13 VGND 0.11841f
C9641 XThR.Tn[8].t34 VGND 0.01888f
C9642 XThR.Tn[8].t26 VGND 0.02067f
C9643 XThR.Tn[8].n14 VGND 0.05048f
C9644 XThR.Tn[8].t53 VGND 0.01882f
C9645 XThR.Tn[8].t22 VGND 0.02061f
C9646 XThR.Tn[8].n15 VGND 0.05252f
C9647 XThR.Tn[8].n16 VGND 0.0369f
C9648 XThR.Tn[8].n17 VGND 0.00675f
C9649 XThR.Tn[8].n18 VGND 0.11841f
C9650 XThR.Tn[8].t50 VGND 0.01888f
C9651 XThR.Tn[8].t43 VGND 0.02067f
C9652 XThR.Tn[8].n19 VGND 0.05048f
C9653 XThR.Tn[8].t65 VGND 0.01882f
C9654 XThR.Tn[8].t40 VGND 0.02061f
C9655 XThR.Tn[8].n20 VGND 0.05252f
C9656 XThR.Tn[8].n21 VGND 0.0369f
C9657 XThR.Tn[8].n22 VGND 0.00675f
C9658 XThR.Tn[8].n23 VGND 0.11841f
C9659 XThR.Tn[8].t12 VGND 0.01888f
C9660 XThR.Tn[8].t70 VGND 0.02067f
C9661 XThR.Tn[8].n24 VGND 0.05048f
C9662 XThR.Tn[8].t36 VGND 0.01882f
C9663 XThR.Tn[8].t66 VGND 0.02061f
C9664 XThR.Tn[8].n25 VGND 0.05252f
C9665 XThR.Tn[8].n26 VGND 0.0369f
C9666 XThR.Tn[8].n27 VGND 0.00675f
C9667 XThR.Tn[8].n28 VGND 0.11841f
C9668 XThR.Tn[8].t52 VGND 0.01888f
C9669 XThR.Tn[8].t44 VGND 0.02067f
C9670 XThR.Tn[8].n29 VGND 0.05048f
C9671 XThR.Tn[8].t68 VGND 0.01882f
C9672 XThR.Tn[8].t41 VGND 0.02061f
C9673 XThR.Tn[8].n30 VGND 0.05252f
C9674 XThR.Tn[8].n31 VGND 0.0369f
C9675 XThR.Tn[8].n32 VGND 0.00675f
C9676 XThR.Tn[8].n33 VGND 0.11841f
C9677 XThR.Tn[8].t28 VGND 0.01888f
C9678 XThR.Tn[8].t61 VGND 0.02067f
C9679 XThR.Tn[8].n34 VGND 0.05048f
C9680 XThR.Tn[8].t47 VGND 0.01882f
C9681 XThR.Tn[8].t58 VGND 0.02061f
C9682 XThR.Tn[8].n35 VGND 0.05252f
C9683 XThR.Tn[8].n36 VGND 0.0369f
C9684 XThR.Tn[8].n37 VGND 0.00675f
C9685 XThR.Tn[8].n38 VGND 0.11841f
C9686 XThR.Tn[8].t60 VGND 0.01888f
C9687 XThR.Tn[8].t56 VGND 0.02067f
C9688 XThR.Tn[8].n39 VGND 0.05048f
C9689 XThR.Tn[8].t14 VGND 0.01882f
C9690 XThR.Tn[8].t51 VGND 0.02061f
C9691 XThR.Tn[8].n40 VGND 0.05252f
C9692 XThR.Tn[8].n41 VGND 0.0369f
C9693 XThR.Tn[8].n42 VGND 0.00675f
C9694 XThR.Tn[8].n43 VGND 0.11841f
C9695 XThR.Tn[8].t63 VGND 0.01888f
C9696 XThR.Tn[8].t69 VGND 0.02067f
C9697 XThR.Tn[8].n44 VGND 0.05048f
C9698 XThR.Tn[8].t20 VGND 0.01882f
C9699 XThR.Tn[8].t64 VGND 0.02061f
C9700 XThR.Tn[8].n45 VGND 0.05252f
C9701 XThR.Tn[8].n46 VGND 0.0369f
C9702 XThR.Tn[8].n47 VGND 0.00675f
C9703 XThR.Tn[8].n48 VGND 0.11841f
C9704 XThR.Tn[8].t17 VGND 0.01888f
C9705 XThR.Tn[8].t27 VGND 0.02067f
C9706 XThR.Tn[8].n49 VGND 0.05048f
C9707 XThR.Tn[8].t38 VGND 0.01882f
C9708 XThR.Tn[8].t24 VGND 0.02061f
C9709 XThR.Tn[8].n50 VGND 0.05252f
C9710 XThR.Tn[8].n51 VGND 0.0369f
C9711 XThR.Tn[8].n52 VGND 0.00675f
C9712 XThR.Tn[8].n53 VGND 0.11841f
C9713 XThR.Tn[8].t72 VGND 0.01888f
C9714 XThR.Tn[8].t46 VGND 0.02067f
C9715 XThR.Tn[8].n54 VGND 0.05048f
C9716 XThR.Tn[8].t31 VGND 0.01882f
C9717 XThR.Tn[8].t42 VGND 0.02061f
C9718 XThR.Tn[8].n55 VGND 0.05252f
C9719 XThR.Tn[8].n56 VGND 0.0369f
C9720 XThR.Tn[8].n57 VGND 0.00675f
C9721 XThR.Tn[8].n58 VGND 0.11841f
C9722 XThR.Tn[8].t30 VGND 0.01888f
C9723 XThR.Tn[8].t21 VGND 0.02067f
C9724 XThR.Tn[8].n59 VGND 0.05048f
C9725 XThR.Tn[8].t48 VGND 0.01882f
C9726 XThR.Tn[8].t16 VGND 0.02061f
C9727 XThR.Tn[8].n60 VGND 0.05252f
C9728 XThR.Tn[8].n61 VGND 0.0369f
C9729 XThR.Tn[8].n62 VGND 0.00675f
C9730 XThR.Tn[8].n63 VGND 0.11841f
C9731 XThR.Tn[8].t62 VGND 0.01888f
C9732 XThR.Tn[8].t57 VGND 0.02067f
C9733 XThR.Tn[8].n64 VGND 0.05048f
C9734 XThR.Tn[8].t18 VGND 0.01882f
C9735 XThR.Tn[8].t54 VGND 0.02061f
C9736 XThR.Tn[8].n65 VGND 0.05252f
C9737 XThR.Tn[8].n66 VGND 0.0369f
C9738 XThR.Tn[8].n67 VGND 0.00675f
C9739 XThR.Tn[8].n68 VGND 0.11841f
C9740 XThR.Tn[8].t15 VGND 0.01888f
C9741 XThR.Tn[8].t71 VGND 0.02067f
C9742 XThR.Tn[8].n69 VGND 0.05048f
C9743 XThR.Tn[8].t37 VGND 0.01882f
C9744 XThR.Tn[8].t67 VGND 0.02061f
C9745 XThR.Tn[8].n70 VGND 0.05252f
C9746 XThR.Tn[8].n71 VGND 0.0369f
C9747 XThR.Tn[8].n72 VGND 0.00675f
C9748 XThR.Tn[8].n73 VGND 0.11841f
C9749 XThR.Tn[8].t35 VGND 0.01888f
C9750 XThR.Tn[8].t29 VGND 0.02067f
C9751 XThR.Tn[8].n74 VGND 0.05048f
C9752 XThR.Tn[8].t55 VGND 0.01882f
C9753 XThR.Tn[8].t25 VGND 0.02061f
C9754 XThR.Tn[8].n75 VGND 0.05252f
C9755 XThR.Tn[8].n76 VGND 0.0369f
C9756 XThR.Tn[8].n77 VGND 0.00675f
C9757 XThR.Tn[8].n78 VGND 0.11841f
C9758 XThR.Tn[8].t73 VGND 0.01888f
C9759 XThR.Tn[8].t23 VGND 0.02067f
C9760 XThR.Tn[8].n79 VGND 0.05048f
C9761 XThR.Tn[8].t32 VGND 0.01882f
C9762 XThR.Tn[8].t19 VGND 0.02061f
C9763 XThR.Tn[8].n80 VGND 0.05252f
C9764 XThR.Tn[8].n81 VGND 0.0369f
C9765 XThR.Tn[8].n82 VGND 0.00675f
C9766 XThR.Tn[8].n83 VGND 0.11841f
C9767 XThR.Tn[8].n84 VGND 0.10761f
C9768 XThR.Tn[8].n85 VGND 0.32972f
C9769 XThR.Tn[8].t11 VGND 0.0157f
C9770 XThR.Tn[8].t3 VGND 0.0157f
C9771 XThR.Tn[8].n86 VGND 0.03916f
C9772 XThR.Tn[8].t2 VGND 0.0157f
C9773 XThR.Tn[8].t0 VGND 0.0157f
C9774 XThR.Tn[8].n87 VGND 0.0314f
C9775 XThR.Tn[8].n88 VGND 0.07241f
C9776 XThR.Tn[0].t5 VGND 0.02293f
C9777 XThR.Tn[0].t6 VGND 0.02293f
C9778 XThR.Tn[0].n0 VGND 0.04628f
C9779 XThR.Tn[0].t4 VGND 0.02293f
C9780 XThR.Tn[0].t3 VGND 0.02293f
C9781 XThR.Tn[0].n1 VGND 0.05416f
C9782 XThR.Tn[0].n2 VGND 0.16245f
C9783 XThR.Tn[0].t8 VGND 0.0149f
C9784 XThR.Tn[0].t9 VGND 0.0149f
C9785 XThR.Tn[0].n3 VGND 0.03394f
C9786 XThR.Tn[0].t7 VGND 0.0149f
C9787 XThR.Tn[0].t10 VGND 0.0149f
C9788 XThR.Tn[0].n4 VGND 0.03394f
C9789 XThR.Tn[0].t11 VGND 0.0149f
C9790 XThR.Tn[0].t1 VGND 0.0149f
C9791 XThR.Tn[0].n5 VGND 0.05655f
C9792 XThR.Tn[0].t2 VGND 0.0149f
C9793 XThR.Tn[0].t0 VGND 0.0149f
C9794 XThR.Tn[0].n6 VGND 0.03394f
C9795 XThR.Tn[0].n7 VGND 0.16164f
C9796 XThR.Tn[0].n8 VGND 0.09992f
C9797 XThR.Tn[0].n9 VGND 0.11277f
C9798 XThR.Tn[0].t48 VGND 0.01792f
C9799 XThR.Tn[0].t40 VGND 0.01962f
C9800 XThR.Tn[0].n10 VGND 0.04792f
C9801 XThR.Tn[0].n11 VGND 0.09205f
C9802 XThR.Tn[0].t67 VGND 0.01792f
C9803 XThR.Tn[0].t58 VGND 0.01962f
C9804 XThR.Tn[0].n12 VGND 0.04792f
C9805 XThR.Tn[0].t24 VGND 0.01786f
C9806 XThR.Tn[0].t50 VGND 0.01956f
C9807 XThR.Tn[0].n13 VGND 0.04986f
C9808 XThR.Tn[0].n14 VGND 0.03503f
C9809 XThR.Tn[0].n15 VGND 0.0064f
C9810 XThR.Tn[0].n16 VGND 0.11241f
C9811 XThR.Tn[0].t41 VGND 0.01792f
C9812 XThR.Tn[0].t33 VGND 0.01962f
C9813 XThR.Tn[0].n17 VGND 0.04792f
C9814 XThR.Tn[0].t61 VGND 0.01786f
C9815 XThR.Tn[0].t26 VGND 0.01956f
C9816 XThR.Tn[0].n18 VGND 0.04986f
C9817 XThR.Tn[0].n19 VGND 0.03503f
C9818 XThR.Tn[0].n20 VGND 0.0064f
C9819 XThR.Tn[0].n21 VGND 0.11241f
C9820 XThR.Tn[0].t59 VGND 0.01792f
C9821 XThR.Tn[0].t51 VGND 0.01962f
C9822 XThR.Tn[0].n22 VGND 0.04792f
C9823 XThR.Tn[0].t12 VGND 0.01786f
C9824 XThR.Tn[0].t44 VGND 0.01956f
C9825 XThR.Tn[0].n23 VGND 0.04986f
C9826 XThR.Tn[0].n24 VGND 0.03503f
C9827 XThR.Tn[0].n25 VGND 0.0064f
C9828 XThR.Tn[0].n26 VGND 0.11241f
C9829 XThR.Tn[0].t21 VGND 0.01792f
C9830 XThR.Tn[0].t15 VGND 0.01962f
C9831 XThR.Tn[0].n27 VGND 0.04792f
C9832 XThR.Tn[0].t43 VGND 0.01786f
C9833 XThR.Tn[0].t72 VGND 0.01956f
C9834 XThR.Tn[0].n28 VGND 0.04986f
C9835 XThR.Tn[0].n29 VGND 0.03503f
C9836 XThR.Tn[0].n30 VGND 0.0064f
C9837 XThR.Tn[0].n31 VGND 0.11241f
C9838 XThR.Tn[0].t60 VGND 0.01792f
C9839 XThR.Tn[0].t52 VGND 0.01962f
C9840 XThR.Tn[0].n32 VGND 0.04792f
C9841 XThR.Tn[0].t13 VGND 0.01786f
C9842 XThR.Tn[0].t46 VGND 0.01956f
C9843 XThR.Tn[0].n33 VGND 0.04986f
C9844 XThR.Tn[0].n34 VGND 0.03503f
C9845 XThR.Tn[0].n35 VGND 0.0064f
C9846 XThR.Tn[0].n36 VGND 0.11241f
C9847 XThR.Tn[0].t35 VGND 0.01792f
C9848 XThR.Tn[0].t68 VGND 0.01962f
C9849 XThR.Tn[0].n37 VGND 0.04792f
C9850 XThR.Tn[0].t54 VGND 0.01786f
C9851 XThR.Tn[0].t64 VGND 0.01956f
C9852 XThR.Tn[0].n38 VGND 0.04986f
C9853 XThR.Tn[0].n39 VGND 0.03503f
C9854 XThR.Tn[0].n40 VGND 0.0064f
C9855 XThR.Tn[0].n41 VGND 0.11241f
C9856 XThR.Tn[0].t66 VGND 0.01792f
C9857 XThR.Tn[0].t63 VGND 0.01962f
C9858 XThR.Tn[0].n42 VGND 0.04792f
C9859 XThR.Tn[0].t23 VGND 0.01786f
C9860 XThR.Tn[0].t55 VGND 0.01956f
C9861 XThR.Tn[0].n43 VGND 0.04986f
C9862 XThR.Tn[0].n44 VGND 0.03503f
C9863 XThR.Tn[0].n45 VGND 0.0064f
C9864 XThR.Tn[0].n46 VGND 0.11241f
C9865 XThR.Tn[0].t70 VGND 0.01792f
C9866 XThR.Tn[0].t14 VGND 0.01962f
C9867 XThR.Tn[0].n47 VGND 0.04792f
C9868 XThR.Tn[0].t28 VGND 0.01786f
C9869 XThR.Tn[0].t71 VGND 0.01956f
C9870 XThR.Tn[0].n48 VGND 0.04986f
C9871 XThR.Tn[0].n49 VGND 0.03503f
C9872 XThR.Tn[0].n50 VGND 0.0064f
C9873 XThR.Tn[0].n51 VGND 0.11241f
C9874 XThR.Tn[0].t25 VGND 0.01792f
C9875 XThR.Tn[0].t34 VGND 0.01962f
C9876 XThR.Tn[0].n52 VGND 0.04792f
C9877 XThR.Tn[0].t47 VGND 0.01786f
C9878 XThR.Tn[0].t29 VGND 0.01956f
C9879 XThR.Tn[0].n53 VGND 0.04986f
C9880 XThR.Tn[0].n54 VGND 0.03503f
C9881 XThR.Tn[0].n55 VGND 0.0064f
C9882 XThR.Tn[0].n56 VGND 0.11241f
C9883 XThR.Tn[0].t17 VGND 0.01792f
C9884 XThR.Tn[0].t53 VGND 0.01962f
C9885 XThR.Tn[0].n57 VGND 0.04792f
C9886 XThR.Tn[0].t38 VGND 0.01786f
C9887 XThR.Tn[0].t49 VGND 0.01956f
C9888 XThR.Tn[0].n58 VGND 0.04986f
C9889 XThR.Tn[0].n59 VGND 0.03503f
C9890 XThR.Tn[0].n60 VGND 0.0064f
C9891 XThR.Tn[0].n61 VGND 0.11241f
C9892 XThR.Tn[0].t37 VGND 0.01792f
C9893 XThR.Tn[0].t31 VGND 0.01962f
C9894 XThR.Tn[0].n62 VGND 0.04792f
C9895 XThR.Tn[0].t56 VGND 0.01786f
C9896 XThR.Tn[0].t19 VGND 0.01956f
C9897 XThR.Tn[0].n63 VGND 0.04986f
C9898 XThR.Tn[0].n64 VGND 0.03503f
C9899 XThR.Tn[0].n65 VGND 0.0064f
C9900 XThR.Tn[0].n66 VGND 0.11241f
C9901 XThR.Tn[0].t69 VGND 0.01792f
C9902 XThR.Tn[0].t65 VGND 0.01962f
C9903 XThR.Tn[0].n67 VGND 0.04792f
C9904 XThR.Tn[0].t27 VGND 0.01786f
C9905 XThR.Tn[0].t57 VGND 0.01956f
C9906 XThR.Tn[0].n68 VGND 0.04986f
C9907 XThR.Tn[0].n69 VGND 0.03503f
C9908 XThR.Tn[0].n70 VGND 0.0064f
C9909 XThR.Tn[0].n71 VGND 0.11241f
C9910 XThR.Tn[0].t22 VGND 0.01792f
C9911 XThR.Tn[0].t16 VGND 0.01962f
C9912 XThR.Tn[0].n72 VGND 0.04792f
C9913 XThR.Tn[0].t45 VGND 0.01786f
C9914 XThR.Tn[0].t73 VGND 0.01956f
C9915 XThR.Tn[0].n73 VGND 0.04986f
C9916 XThR.Tn[0].n74 VGND 0.03503f
C9917 XThR.Tn[0].n75 VGND 0.0064f
C9918 XThR.Tn[0].n76 VGND 0.11241f
C9919 XThR.Tn[0].t42 VGND 0.01792f
C9920 XThR.Tn[0].t36 VGND 0.01962f
C9921 XThR.Tn[0].n77 VGND 0.04792f
C9922 XThR.Tn[0].t62 VGND 0.01786f
C9923 XThR.Tn[0].t30 VGND 0.01956f
C9924 XThR.Tn[0].n78 VGND 0.04986f
C9925 XThR.Tn[0].n79 VGND 0.03503f
C9926 XThR.Tn[0].n80 VGND 0.0064f
C9927 XThR.Tn[0].n81 VGND 0.11241f
C9928 XThR.Tn[0].t18 VGND 0.01792f
C9929 XThR.Tn[0].t32 VGND 0.01962f
C9930 XThR.Tn[0].n82 VGND 0.04792f
C9931 XThR.Tn[0].t39 VGND 0.01786f
C9932 XThR.Tn[0].t20 VGND 0.01956f
C9933 XThR.Tn[0].n83 VGND 0.04986f
C9934 XThR.Tn[0].n84 VGND 0.03503f
C9935 XThR.Tn[0].n85 VGND 0.0064f
C9936 XThR.Tn[0].n86 VGND 0.11241f
C9937 XThR.Tn[0].n87 VGND 0.10215f
C9938 XThR.Tn[0].n88 VGND 0.29249f
C9939 XThR.Tn[7].t7 VGND 0.01503f
C9940 XThR.Tn[7].t4 VGND 0.01503f
C9941 XThR.Tn[7].n0 VGND 0.04638f
C9942 XThR.Tn[7].t6 VGND 0.01503f
C9943 XThR.Tn[7].t5 VGND 0.01503f
C9944 XThR.Tn[7].n1 VGND 0.03319f
C9945 XThR.Tn[7].n2 VGND 0.17022f
C9946 XThR.Tn[7].t2 VGND 0.02312f
C9947 XThR.Tn[7].t3 VGND 0.02312f
C9948 XThR.Tn[7].n3 VGND 0.0704f
C9949 XThR.Tn[7].t1 VGND 0.02312f
C9950 XThR.Tn[7].t0 VGND 0.02312f
C9951 XThR.Tn[7].n4 VGND 0.05122f
C9952 XThR.Tn[7].n5 VGND 0.22538f
C9953 XThR.Tn[7].n6 VGND 0.02809f
C9954 XThR.Tn[7].t53 VGND 0.01807f
C9955 XThR.Tn[7].t45 VGND 0.01979f
C9956 XThR.Tn[7].n7 VGND 0.04832f
C9957 XThR.Tn[7].n8 VGND 0.09282f
C9958 XThR.Tn[7].t8 VGND 0.01807f
C9959 XThR.Tn[7].t60 VGND 0.01979f
C9960 XThR.Tn[7].n9 VGND 0.04832f
C9961 XThR.Tn[7].t26 VGND 0.01801f
C9962 XThR.Tn[7].t38 VGND 0.01972f
C9963 XThR.Tn[7].n10 VGND 0.05027f
C9964 XThR.Tn[7].n11 VGND 0.03532f
C9965 XThR.Tn[7].n12 VGND 0.00646f
C9966 XThR.Tn[7].n13 VGND 0.11334f
C9967 XThR.Tn[7].t47 VGND 0.01807f
C9968 XThR.Tn[7].t37 VGND 0.01979f
C9969 XThR.Tn[7].n14 VGND 0.04832f
C9970 XThR.Tn[7].t66 VGND 0.01801f
C9971 XThR.Tn[7].t15 VGND 0.01972f
C9972 XThR.Tn[7].n15 VGND 0.05027f
C9973 XThR.Tn[7].n16 VGND 0.03532f
C9974 XThR.Tn[7].n17 VGND 0.00646f
C9975 XThR.Tn[7].n18 VGND 0.11334f
C9976 XThR.Tn[7].t62 VGND 0.01807f
C9977 XThR.Tn[7].t55 VGND 0.01979f
C9978 XThR.Tn[7].n19 VGND 0.04832f
C9979 XThR.Tn[7].t18 VGND 0.01801f
C9980 XThR.Tn[7].t32 VGND 0.01972f
C9981 XThR.Tn[7].n20 VGND 0.05027f
C9982 XThR.Tn[7].n21 VGND 0.03532f
C9983 XThR.Tn[7].n22 VGND 0.00646f
C9984 XThR.Tn[7].n23 VGND 0.11334f
C9985 XThR.Tn[7].t25 VGND 0.01807f
C9986 XThR.Tn[7].t21 VGND 0.01979f
C9987 XThR.Tn[7].n24 VGND 0.04832f
C9988 XThR.Tn[7].t50 VGND 0.01801f
C9989 XThR.Tn[7].t63 VGND 0.01972f
C9990 XThR.Tn[7].n25 VGND 0.05027f
C9991 XThR.Tn[7].n26 VGND 0.03532f
C9992 XThR.Tn[7].n27 VGND 0.00646f
C9993 XThR.Tn[7].n28 VGND 0.11334f
C9994 XThR.Tn[7].t65 VGND 0.01807f
C9995 XThR.Tn[7].t56 VGND 0.01979f
C9996 XThR.Tn[7].n29 VGND 0.04832f
C9997 XThR.Tn[7].t19 VGND 0.01801f
C9998 XThR.Tn[7].t34 VGND 0.01972f
C9999 XThR.Tn[7].n30 VGND 0.05027f
C10000 XThR.Tn[7].n31 VGND 0.03532f
C10001 XThR.Tn[7].n32 VGND 0.00646f
C10002 XThR.Tn[7].n33 VGND 0.11334f
C10003 XThR.Tn[7].t40 VGND 0.01807f
C10004 XThR.Tn[7].t11 VGND 0.01979f
C10005 XThR.Tn[7].n34 VGND 0.04832f
C10006 XThR.Tn[7].t58 VGND 0.01801f
C10007 XThR.Tn[7].t54 VGND 0.01972f
C10008 XThR.Tn[7].n35 VGND 0.05027f
C10009 XThR.Tn[7].n36 VGND 0.03532f
C10010 XThR.Tn[7].n37 VGND 0.00646f
C10011 XThR.Tn[7].n38 VGND 0.11334f
C10012 XThR.Tn[7].t9 VGND 0.01807f
C10013 XThR.Tn[7].t68 VGND 0.01979f
C10014 XThR.Tn[7].n39 VGND 0.04832f
C10015 XThR.Tn[7].t27 VGND 0.01801f
C10016 XThR.Tn[7].t46 VGND 0.01972f
C10017 XThR.Tn[7].n40 VGND 0.05027f
C10018 XThR.Tn[7].n41 VGND 0.03532f
C10019 XThR.Tn[7].n42 VGND 0.00646f
C10020 XThR.Tn[7].n43 VGND 0.11334f
C10021 XThR.Tn[7].t14 VGND 0.01807f
C10022 XThR.Tn[7].t20 VGND 0.01979f
C10023 XThR.Tn[7].n44 VGND 0.04832f
C10024 XThR.Tn[7].t31 VGND 0.01801f
C10025 XThR.Tn[7].t61 VGND 0.01972f
C10026 XThR.Tn[7].n45 VGND 0.05027f
C10027 XThR.Tn[7].n46 VGND 0.03532f
C10028 XThR.Tn[7].n47 VGND 0.00646f
C10029 XThR.Tn[7].n48 VGND 0.11334f
C10030 XThR.Tn[7].t29 VGND 0.01807f
C10031 XThR.Tn[7].t39 VGND 0.01979f
C10032 XThR.Tn[7].n49 VGND 0.04832f
C10033 XThR.Tn[7].t52 VGND 0.01801f
C10034 XThR.Tn[7].t16 VGND 0.01972f
C10035 XThR.Tn[7].n50 VGND 0.05027f
C10036 XThR.Tn[7].n51 VGND 0.03532f
C10037 XThR.Tn[7].n52 VGND 0.00646f
C10038 XThR.Tn[7].n53 VGND 0.11334f
C10039 XThR.Tn[7].t23 VGND 0.01807f
C10040 XThR.Tn[7].t57 VGND 0.01979f
C10041 XThR.Tn[7].n54 VGND 0.04832f
C10042 XThR.Tn[7].t43 VGND 0.01801f
C10043 XThR.Tn[7].t36 VGND 0.01972f
C10044 XThR.Tn[7].n55 VGND 0.05027f
C10045 XThR.Tn[7].n56 VGND 0.03532f
C10046 XThR.Tn[7].n57 VGND 0.00646f
C10047 XThR.Tn[7].n58 VGND 0.11334f
C10048 XThR.Tn[7].t42 VGND 0.01807f
C10049 XThR.Tn[7].t33 VGND 0.01979f
C10050 XThR.Tn[7].n59 VGND 0.04832f
C10051 XThR.Tn[7].t59 VGND 0.01801f
C10052 XThR.Tn[7].t10 VGND 0.01972f
C10053 XThR.Tn[7].n60 VGND 0.05027f
C10054 XThR.Tn[7].n61 VGND 0.03532f
C10055 XThR.Tn[7].n62 VGND 0.00646f
C10056 XThR.Tn[7].n63 VGND 0.11334f
C10057 XThR.Tn[7].t12 VGND 0.01807f
C10058 XThR.Tn[7].t69 VGND 0.01979f
C10059 XThR.Tn[7].n64 VGND 0.04832f
C10060 XThR.Tn[7].t30 VGND 0.01801f
C10061 XThR.Tn[7].t48 VGND 0.01972f
C10062 XThR.Tn[7].n65 VGND 0.05027f
C10063 XThR.Tn[7].n66 VGND 0.03532f
C10064 XThR.Tn[7].n67 VGND 0.00646f
C10065 XThR.Tn[7].n68 VGND 0.11334f
C10066 XThR.Tn[7].t28 VGND 0.01807f
C10067 XThR.Tn[7].t22 VGND 0.01979f
C10068 XThR.Tn[7].n69 VGND 0.04832f
C10069 XThR.Tn[7].t51 VGND 0.01801f
C10070 XThR.Tn[7].t64 VGND 0.01972f
C10071 XThR.Tn[7].n70 VGND 0.05027f
C10072 XThR.Tn[7].n71 VGND 0.03532f
C10073 XThR.Tn[7].n72 VGND 0.00646f
C10074 XThR.Tn[7].n73 VGND 0.11334f
C10075 XThR.Tn[7].t49 VGND 0.01807f
C10076 XThR.Tn[7].t41 VGND 0.01979f
C10077 XThR.Tn[7].n74 VGND 0.04832f
C10078 XThR.Tn[7].t67 VGND 0.01801f
C10079 XThR.Tn[7].t17 VGND 0.01972f
C10080 XThR.Tn[7].n75 VGND 0.05027f
C10081 XThR.Tn[7].n76 VGND 0.03532f
C10082 XThR.Tn[7].n77 VGND 0.00646f
C10083 XThR.Tn[7].n78 VGND 0.11334f
C10084 XThR.Tn[7].t24 VGND 0.01807f
C10085 XThR.Tn[7].t35 VGND 0.01979f
C10086 XThR.Tn[7].n79 VGND 0.04832f
C10087 XThR.Tn[7].t44 VGND 0.01801f
C10088 XThR.Tn[7].t13 VGND 0.01972f
C10089 XThR.Tn[7].n80 VGND 0.05027f
C10090 XThR.Tn[7].n81 VGND 0.03532f
C10091 XThR.Tn[7].n82 VGND 0.00646f
C10092 XThR.Tn[7].n83 VGND 0.11334f
C10093 XThR.Tn[7].n84 VGND 0.103f
C10094 XThR.Tn[7].n85 VGND 0.41812f
C10095 XThR.Tn[11].t5 VGND 0.01567f
C10096 XThR.Tn[11].t2 VGND 0.01567f
C10097 XThR.Tn[11].n0 VGND 0.03134f
C10098 XThR.Tn[11].t4 VGND 0.01567f
C10099 XThR.Tn[11].t0 VGND 0.01567f
C10100 XThR.Tn[11].n1 VGND 0.03908f
C10101 XThR.Tn[11].n2 VGND 0.07883f
C10102 XThR.Tn[11].t6 VGND 0.0241f
C10103 XThR.Tn[11].t8 VGND 0.0241f
C10104 XThR.Tn[11].n3 VGND 0.07319f
C10105 XThR.Tn[11].t7 VGND 0.0241f
C10106 XThR.Tn[11].t9 VGND 0.0241f
C10107 XThR.Tn[11].n4 VGND 0.05358f
C10108 XThR.Tn[11].n5 VGND 0.24365f
C10109 XThR.Tn[11].t3 VGND 0.0241f
C10110 XThR.Tn[11].t11 VGND 0.0241f
C10111 XThR.Tn[11].n6 VGND 0.05208f
C10112 XThR.Tn[11].t1 VGND 0.0241f
C10113 XThR.Tn[11].t10 VGND 0.0241f
C10114 XThR.Tn[11].n7 VGND 0.07927f
C10115 XThR.Tn[11].n8 VGND 0.2201f
C10116 XThR.Tn[11].n9 VGND 0.02947f
C10117 XThR.Tn[11].t56 VGND 0.01884f
C10118 XThR.Tn[11].t48 VGND 0.02063f
C10119 XThR.Tn[11].n10 VGND 0.05037f
C10120 XThR.Tn[11].n11 VGND 0.09677f
C10121 XThR.Tn[11].t12 VGND 0.01884f
C10122 XThR.Tn[11].t67 VGND 0.02063f
C10123 XThR.Tn[11].n12 VGND 0.05037f
C10124 XThR.Tn[11].t27 VGND 0.01878f
C10125 XThR.Tn[11].t58 VGND 0.02056f
C10126 XThR.Tn[11].n13 VGND 0.05241f
C10127 XThR.Tn[11].n14 VGND 0.03682f
C10128 XThR.Tn[11].n15 VGND 0.00673f
C10129 XThR.Tn[11].n16 VGND 0.11816f
C10130 XThR.Tn[11].t49 VGND 0.01884f
C10131 XThR.Tn[11].t41 VGND 0.02063f
C10132 XThR.Tn[11].n17 VGND 0.05037f
C10133 XThR.Tn[11].t65 VGND 0.01878f
C10134 XThR.Tn[11].t36 VGND 0.02056f
C10135 XThR.Tn[11].n18 VGND 0.05241f
C10136 XThR.Tn[11].n19 VGND 0.03682f
C10137 XThR.Tn[11].n20 VGND 0.00673f
C10138 XThR.Tn[11].n21 VGND 0.11816f
C10139 XThR.Tn[11].t68 VGND 0.01884f
C10140 XThR.Tn[11].t60 VGND 0.02063f
C10141 XThR.Tn[11].n22 VGND 0.05037f
C10142 XThR.Tn[11].t18 VGND 0.01878f
C10143 XThR.Tn[11].t54 VGND 0.02056f
C10144 XThR.Tn[11].n23 VGND 0.05241f
C10145 XThR.Tn[11].n24 VGND 0.03682f
C10146 XThR.Tn[11].n25 VGND 0.00673f
C10147 XThR.Tn[11].n26 VGND 0.11816f
C10148 XThR.Tn[11].t33 VGND 0.01884f
C10149 XThR.Tn[11].t23 VGND 0.02063f
C10150 XThR.Tn[11].n27 VGND 0.05037f
C10151 XThR.Tn[11].t50 VGND 0.01878f
C10152 XThR.Tn[11].t19 VGND 0.02056f
C10153 XThR.Tn[11].n28 VGND 0.05241f
C10154 XThR.Tn[11].n29 VGND 0.03682f
C10155 XThR.Tn[11].n30 VGND 0.00673f
C10156 XThR.Tn[11].n31 VGND 0.11816f
C10157 XThR.Tn[11].t70 VGND 0.01884f
C10158 XThR.Tn[11].t62 VGND 0.02063f
C10159 XThR.Tn[11].n32 VGND 0.05037f
C10160 XThR.Tn[11].t21 VGND 0.01878f
C10161 XThR.Tn[11].t55 VGND 0.02056f
C10162 XThR.Tn[11].n33 VGND 0.05241f
C10163 XThR.Tn[11].n34 VGND 0.03682f
C10164 XThR.Tn[11].n35 VGND 0.00673f
C10165 XThR.Tn[11].n36 VGND 0.11816f
C10166 XThR.Tn[11].t44 VGND 0.01884f
C10167 XThR.Tn[11].t14 VGND 0.02063f
C10168 XThR.Tn[11].n37 VGND 0.05037f
C10169 XThR.Tn[11].t59 VGND 0.01878f
C10170 XThR.Tn[11].t72 VGND 0.02056f
C10171 XThR.Tn[11].n38 VGND 0.05241f
C10172 XThR.Tn[11].n39 VGND 0.03682f
C10173 XThR.Tn[11].n40 VGND 0.00673f
C10174 XThR.Tn[11].n41 VGND 0.11816f
C10175 XThR.Tn[11].t13 VGND 0.01884f
C10176 XThR.Tn[11].t71 VGND 0.02063f
C10177 XThR.Tn[11].n42 VGND 0.05037f
C10178 XThR.Tn[11].t28 VGND 0.01878f
C10179 XThR.Tn[11].t64 VGND 0.02056f
C10180 XThR.Tn[11].n43 VGND 0.05241f
C10181 XThR.Tn[11].n44 VGND 0.03682f
C10182 XThR.Tn[11].n45 VGND 0.00673f
C10183 XThR.Tn[11].n46 VGND 0.11816f
C10184 XThR.Tn[11].t16 VGND 0.01884f
C10185 XThR.Tn[11].t22 VGND 0.02063f
C10186 XThR.Tn[11].n47 VGND 0.05037f
C10187 XThR.Tn[11].t32 VGND 0.01878f
C10188 XThR.Tn[11].t17 VGND 0.02056f
C10189 XThR.Tn[11].n48 VGND 0.05241f
C10190 XThR.Tn[11].n49 VGND 0.03682f
C10191 XThR.Tn[11].n50 VGND 0.00673f
C10192 XThR.Tn[11].n51 VGND 0.11816f
C10193 XThR.Tn[11].t35 VGND 0.01884f
C10194 XThR.Tn[11].t43 VGND 0.02063f
C10195 XThR.Tn[11].n52 VGND 0.05037f
C10196 XThR.Tn[11].t52 VGND 0.01878f
C10197 XThR.Tn[11].t37 VGND 0.02056f
C10198 XThR.Tn[11].n53 VGND 0.05241f
C10199 XThR.Tn[11].n54 VGND 0.03682f
C10200 XThR.Tn[11].n55 VGND 0.00673f
C10201 XThR.Tn[11].n56 VGND 0.11816f
C10202 XThR.Tn[11].t25 VGND 0.01884f
C10203 XThR.Tn[11].t63 VGND 0.02063f
C10204 XThR.Tn[11].n57 VGND 0.05037f
C10205 XThR.Tn[11].t42 VGND 0.01878f
C10206 XThR.Tn[11].t57 VGND 0.02056f
C10207 XThR.Tn[11].n58 VGND 0.05241f
C10208 XThR.Tn[11].n59 VGND 0.03682f
C10209 XThR.Tn[11].n60 VGND 0.00673f
C10210 XThR.Tn[11].n61 VGND 0.11816f
C10211 XThR.Tn[11].t47 VGND 0.01884f
C10212 XThR.Tn[11].t39 VGND 0.02063f
C10213 XThR.Tn[11].n62 VGND 0.05037f
C10214 XThR.Tn[11].t61 VGND 0.01878f
C10215 XThR.Tn[11].t29 VGND 0.02056f
C10216 XThR.Tn[11].n63 VGND 0.05241f
C10217 XThR.Tn[11].n64 VGND 0.03682f
C10218 XThR.Tn[11].n65 VGND 0.00673f
C10219 XThR.Tn[11].n66 VGND 0.11816f
C10220 XThR.Tn[11].t15 VGND 0.01884f
C10221 XThR.Tn[11].t73 VGND 0.02063f
C10222 XThR.Tn[11].n67 VGND 0.05037f
C10223 XThR.Tn[11].t30 VGND 0.01878f
C10224 XThR.Tn[11].t66 VGND 0.02056f
C10225 XThR.Tn[11].n68 VGND 0.05241f
C10226 XThR.Tn[11].n69 VGND 0.03682f
C10227 XThR.Tn[11].n70 VGND 0.00673f
C10228 XThR.Tn[11].n71 VGND 0.11816f
C10229 XThR.Tn[11].t34 VGND 0.01884f
C10230 XThR.Tn[11].t24 VGND 0.02063f
C10231 XThR.Tn[11].n72 VGND 0.05037f
C10232 XThR.Tn[11].t51 VGND 0.01878f
C10233 XThR.Tn[11].t20 VGND 0.02056f
C10234 XThR.Tn[11].n73 VGND 0.05241f
C10235 XThR.Tn[11].n74 VGND 0.03682f
C10236 XThR.Tn[11].n75 VGND 0.00673f
C10237 XThR.Tn[11].n76 VGND 0.11816f
C10238 XThR.Tn[11].t53 VGND 0.01884f
C10239 XThR.Tn[11].t46 VGND 0.02063f
C10240 XThR.Tn[11].n77 VGND 0.05037f
C10241 XThR.Tn[11].t69 VGND 0.01878f
C10242 XThR.Tn[11].t38 VGND 0.02056f
C10243 XThR.Tn[11].n78 VGND 0.05241f
C10244 XThR.Tn[11].n79 VGND 0.03682f
C10245 XThR.Tn[11].n80 VGND 0.00673f
C10246 XThR.Tn[11].n81 VGND 0.11816f
C10247 XThR.Tn[11].t26 VGND 0.01884f
C10248 XThR.Tn[11].t40 VGND 0.02063f
C10249 XThR.Tn[11].n82 VGND 0.05037f
C10250 XThR.Tn[11].t45 VGND 0.01878f
C10251 XThR.Tn[11].t31 VGND 0.02056f
C10252 XThR.Tn[11].n83 VGND 0.05241f
C10253 XThR.Tn[11].n84 VGND 0.03682f
C10254 XThR.Tn[11].n85 VGND 0.00673f
C10255 XThR.Tn[11].n86 VGND 0.11816f
C10256 XThR.Tn[11].n87 VGND 0.10738f
C10257 XThR.Tn[11].n88 VGND 0.38486f
C10258 XThR.Tn[4].t9 VGND 0.02325f
C10259 XThR.Tn[4].t10 VGND 0.02325f
C10260 XThR.Tn[4].n0 VGND 0.04693f
C10261 XThR.Tn[4].t8 VGND 0.02325f
C10262 XThR.Tn[4].t11 VGND 0.02325f
C10263 XThR.Tn[4].n1 VGND 0.05491f
C10264 XThR.Tn[4].n2 VGND 0.16472f
C10265 XThR.Tn[4].t7 VGND 0.01511f
C10266 XThR.Tn[4].t4 VGND 0.01511f
C10267 XThR.Tn[4].n3 VGND 0.03442f
C10268 XThR.Tn[4].t6 VGND 0.01511f
C10269 XThR.Tn[4].t5 VGND 0.01511f
C10270 XThR.Tn[4].n4 VGND 0.03442f
C10271 XThR.Tn[4].t0 VGND 0.01511f
C10272 XThR.Tn[4].t1 VGND 0.01511f
C10273 XThR.Tn[4].n5 VGND 0.05735f
C10274 XThR.Tn[4].t3 VGND 0.01511f
C10275 XThR.Tn[4].t2 VGND 0.01511f
C10276 XThR.Tn[4].n6 VGND 0.03442f
C10277 XThR.Tn[4].n7 VGND 0.1639f
C10278 XThR.Tn[4].n8 VGND 0.10132f
C10279 XThR.Tn[4].n9 VGND 0.11435f
C10280 XThR.Tn[4].t44 VGND 0.01817f
C10281 XThR.Tn[4].t38 VGND 0.0199f
C10282 XThR.Tn[4].n10 VGND 0.04859f
C10283 XThR.Tn[4].n11 VGND 0.09334f
C10284 XThR.Tn[4].t65 VGND 0.01817f
C10285 XThR.Tn[4].t54 VGND 0.0199f
C10286 XThR.Tn[4].n12 VGND 0.04859f
C10287 XThR.Tn[4].t19 VGND 0.01811f
C10288 XThR.Tn[4].t50 VGND 0.01983f
C10289 XThR.Tn[4].n13 VGND 0.05056f
C10290 XThR.Tn[4].n14 VGND 0.03552f
C10291 XThR.Tn[4].n15 VGND 0.00649f
C10292 XThR.Tn[4].n16 VGND 0.11398f
C10293 XThR.Tn[4].t39 VGND 0.01817f
C10294 XThR.Tn[4].t31 VGND 0.0199f
C10295 XThR.Tn[4].n17 VGND 0.04859f
C10296 XThR.Tn[4].t58 VGND 0.01811f
C10297 XThR.Tn[4].t27 VGND 0.01983f
C10298 XThR.Tn[4].n18 VGND 0.05056f
C10299 XThR.Tn[4].n19 VGND 0.03552f
C10300 XThR.Tn[4].n20 VGND 0.00649f
C10301 XThR.Tn[4].n21 VGND 0.11398f
C10302 XThR.Tn[4].t55 VGND 0.01817f
C10303 XThR.Tn[4].t48 VGND 0.0199f
C10304 XThR.Tn[4].n22 VGND 0.04859f
C10305 XThR.Tn[4].t70 VGND 0.01811f
C10306 XThR.Tn[4].t45 VGND 0.01983f
C10307 XThR.Tn[4].n23 VGND 0.05056f
C10308 XThR.Tn[4].n24 VGND 0.03552f
C10309 XThR.Tn[4].n25 VGND 0.00649f
C10310 XThR.Tn[4].n26 VGND 0.11398f
C10311 XThR.Tn[4].t17 VGND 0.01817f
C10312 XThR.Tn[4].t13 VGND 0.0199f
C10313 XThR.Tn[4].n27 VGND 0.04859f
C10314 XThR.Tn[4].t41 VGND 0.01811f
C10315 XThR.Tn[4].t71 VGND 0.01983f
C10316 XThR.Tn[4].n28 VGND 0.05056f
C10317 XThR.Tn[4].n29 VGND 0.03552f
C10318 XThR.Tn[4].n30 VGND 0.00649f
C10319 XThR.Tn[4].n31 VGND 0.11398f
C10320 XThR.Tn[4].t57 VGND 0.01817f
C10321 XThR.Tn[4].t49 VGND 0.0199f
C10322 XThR.Tn[4].n32 VGND 0.04859f
C10323 XThR.Tn[4].t73 VGND 0.01811f
C10324 XThR.Tn[4].t46 VGND 0.01983f
C10325 XThR.Tn[4].n33 VGND 0.05056f
C10326 XThR.Tn[4].n34 VGND 0.03552f
C10327 XThR.Tn[4].n35 VGND 0.00649f
C10328 XThR.Tn[4].n36 VGND 0.11398f
C10329 XThR.Tn[4].t33 VGND 0.01817f
C10330 XThR.Tn[4].t66 VGND 0.0199f
C10331 XThR.Tn[4].n37 VGND 0.04859f
C10332 XThR.Tn[4].t52 VGND 0.01811f
C10333 XThR.Tn[4].t63 VGND 0.01983f
C10334 XThR.Tn[4].n38 VGND 0.05056f
C10335 XThR.Tn[4].n39 VGND 0.03552f
C10336 XThR.Tn[4].n40 VGND 0.00649f
C10337 XThR.Tn[4].n41 VGND 0.11398f
C10338 XThR.Tn[4].t64 VGND 0.01817f
C10339 XThR.Tn[4].t61 VGND 0.0199f
C10340 XThR.Tn[4].n42 VGND 0.04859f
C10341 XThR.Tn[4].t18 VGND 0.01811f
C10342 XThR.Tn[4].t56 VGND 0.01983f
C10343 XThR.Tn[4].n43 VGND 0.05056f
C10344 XThR.Tn[4].n44 VGND 0.03552f
C10345 XThR.Tn[4].n45 VGND 0.00649f
C10346 XThR.Tn[4].n46 VGND 0.11398f
C10347 XThR.Tn[4].t68 VGND 0.01817f
C10348 XThR.Tn[4].t12 VGND 0.0199f
C10349 XThR.Tn[4].n47 VGND 0.04859f
C10350 XThR.Tn[4].t25 VGND 0.01811f
C10351 XThR.Tn[4].t69 VGND 0.01983f
C10352 XThR.Tn[4].n48 VGND 0.05056f
C10353 XThR.Tn[4].n49 VGND 0.03552f
C10354 XThR.Tn[4].n50 VGND 0.00649f
C10355 XThR.Tn[4].n51 VGND 0.11398f
C10356 XThR.Tn[4].t22 VGND 0.01817f
C10357 XThR.Tn[4].t32 VGND 0.0199f
C10358 XThR.Tn[4].n52 VGND 0.04859f
C10359 XThR.Tn[4].t43 VGND 0.01811f
C10360 XThR.Tn[4].t29 VGND 0.01983f
C10361 XThR.Tn[4].n53 VGND 0.05056f
C10362 XThR.Tn[4].n54 VGND 0.03552f
C10363 XThR.Tn[4].n55 VGND 0.00649f
C10364 XThR.Tn[4].n56 VGND 0.11398f
C10365 XThR.Tn[4].t15 VGND 0.01817f
C10366 XThR.Tn[4].t51 VGND 0.0199f
C10367 XThR.Tn[4].n57 VGND 0.04859f
C10368 XThR.Tn[4].t36 VGND 0.01811f
C10369 XThR.Tn[4].t47 VGND 0.01983f
C10370 XThR.Tn[4].n58 VGND 0.05056f
C10371 XThR.Tn[4].n59 VGND 0.03552f
C10372 XThR.Tn[4].n60 VGND 0.00649f
C10373 XThR.Tn[4].n61 VGND 0.11398f
C10374 XThR.Tn[4].t35 VGND 0.01817f
C10375 XThR.Tn[4].t26 VGND 0.0199f
C10376 XThR.Tn[4].n62 VGND 0.04859f
C10377 XThR.Tn[4].t53 VGND 0.01811f
C10378 XThR.Tn[4].t21 VGND 0.01983f
C10379 XThR.Tn[4].n63 VGND 0.05056f
C10380 XThR.Tn[4].n64 VGND 0.03552f
C10381 XThR.Tn[4].n65 VGND 0.00649f
C10382 XThR.Tn[4].n66 VGND 0.11398f
C10383 XThR.Tn[4].t67 VGND 0.01817f
C10384 XThR.Tn[4].t62 VGND 0.0199f
C10385 XThR.Tn[4].n67 VGND 0.04859f
C10386 XThR.Tn[4].t23 VGND 0.01811f
C10387 XThR.Tn[4].t59 VGND 0.01983f
C10388 XThR.Tn[4].n68 VGND 0.05056f
C10389 XThR.Tn[4].n69 VGND 0.03552f
C10390 XThR.Tn[4].n70 VGND 0.00649f
C10391 XThR.Tn[4].n71 VGND 0.11398f
C10392 XThR.Tn[4].t20 VGND 0.01817f
C10393 XThR.Tn[4].t14 VGND 0.0199f
C10394 XThR.Tn[4].n72 VGND 0.04859f
C10395 XThR.Tn[4].t42 VGND 0.01811f
C10396 XThR.Tn[4].t72 VGND 0.01983f
C10397 XThR.Tn[4].n73 VGND 0.05056f
C10398 XThR.Tn[4].n74 VGND 0.03552f
C10399 XThR.Tn[4].n75 VGND 0.00649f
C10400 XThR.Tn[4].n76 VGND 0.11398f
C10401 XThR.Tn[4].t40 VGND 0.01817f
C10402 XThR.Tn[4].t34 VGND 0.0199f
C10403 XThR.Tn[4].n77 VGND 0.04859f
C10404 XThR.Tn[4].t60 VGND 0.01811f
C10405 XThR.Tn[4].t30 VGND 0.01983f
C10406 XThR.Tn[4].n78 VGND 0.05056f
C10407 XThR.Tn[4].n79 VGND 0.03552f
C10408 XThR.Tn[4].n80 VGND 0.00649f
C10409 XThR.Tn[4].n81 VGND 0.11398f
C10410 XThR.Tn[4].t16 VGND 0.01817f
C10411 XThR.Tn[4].t28 VGND 0.0199f
C10412 XThR.Tn[4].n82 VGND 0.04859f
C10413 XThR.Tn[4].t37 VGND 0.01811f
C10414 XThR.Tn[4].t24 VGND 0.01983f
C10415 XThR.Tn[4].n83 VGND 0.05056f
C10416 XThR.Tn[4].n84 VGND 0.03552f
C10417 XThR.Tn[4].n85 VGND 0.00649f
C10418 XThR.Tn[4].n86 VGND 0.11398f
C10419 XThR.Tn[4].n87 VGND 0.10358f
C10420 XThR.Tn[4].n88 VGND 0.19569f
C10421 XThC.Tn[7].t6 VGND 0.01228f
C10422 XThC.Tn[7].t5 VGND 0.01228f
C10423 XThC.Tn[7].n0 VGND 0.03791f
C10424 XThC.Tn[7].t4 VGND 0.01228f
C10425 XThC.Tn[7].t7 VGND 0.01228f
C10426 XThC.Tn[7].n1 VGND 0.02713f
C10427 XThC.Tn[7].n2 VGND 0.13418f
C10428 XThC.Tn[7].t0 VGND 0.0189f
C10429 XThC.Tn[7].t3 VGND 0.0189f
C10430 XThC.Tn[7].n3 VGND 0.0407f
C10431 XThC.Tn[7].t2 VGND 0.0189f
C10432 XThC.Tn[7].t1 VGND 0.0189f
C10433 XThC.Tn[7].n4 VGND 0.06179f
C10434 XThC.Tn[7].n5 VGND 0.18167f
C10435 XThC.Tn[7].t8 VGND 0.01498f
C10436 XThC.Tn[7].t11 VGND 0.01636f
C10437 XThC.Tn[7].n6 VGND 0.03652f
C10438 XThC.Tn[7].n7 VGND 0.02502f
C10439 XThC.Tn[7].n8 VGND 0.08213f
C10440 XThC.Tn[7].t25 VGND 0.01498f
C10441 XThC.Tn[7].t30 VGND 0.01636f
C10442 XThC.Tn[7].n9 VGND 0.03652f
C10443 XThC.Tn[7].n10 VGND 0.02502f
C10444 XThC.Tn[7].n11 VGND 0.08235f
C10445 XThC.Tn[7].n12 VGND 0.13573f
C10446 XThC.Tn[7].t27 VGND 0.01498f
C10447 XThC.Tn[7].t34 VGND 0.01636f
C10448 XThC.Tn[7].n13 VGND 0.03652f
C10449 XThC.Tn[7].n14 VGND 0.02502f
C10450 XThC.Tn[7].n15 VGND 0.08235f
C10451 XThC.Tn[7].n16 VGND 0.13573f
C10452 XThC.Tn[7].t29 VGND 0.01498f
C10453 XThC.Tn[7].t35 VGND 0.01636f
C10454 XThC.Tn[7].n17 VGND 0.03652f
C10455 XThC.Tn[7].n18 VGND 0.02502f
C10456 XThC.Tn[7].n19 VGND 0.08235f
C10457 XThC.Tn[7].n20 VGND 0.13573f
C10458 XThC.Tn[7].t18 VGND 0.01498f
C10459 XThC.Tn[7].t22 VGND 0.01636f
C10460 XThC.Tn[7].n21 VGND 0.03652f
C10461 XThC.Tn[7].n22 VGND 0.02502f
C10462 XThC.Tn[7].n23 VGND 0.08235f
C10463 XThC.Tn[7].n24 VGND 0.13573f
C10464 XThC.Tn[7].t20 VGND 0.01498f
C10465 XThC.Tn[7].t23 VGND 0.01636f
C10466 XThC.Tn[7].n25 VGND 0.03652f
C10467 XThC.Tn[7].n26 VGND 0.02502f
C10468 XThC.Tn[7].n27 VGND 0.08235f
C10469 XThC.Tn[7].n28 VGND 0.13573f
C10470 XThC.Tn[7].t33 VGND 0.01498f
C10471 XThC.Tn[7].t39 VGND 0.01636f
C10472 XThC.Tn[7].n29 VGND 0.03652f
C10473 XThC.Tn[7].n30 VGND 0.02502f
C10474 XThC.Tn[7].n31 VGND 0.08235f
C10475 XThC.Tn[7].n32 VGND 0.13573f
C10476 XThC.Tn[7].t10 VGND 0.01498f
C10477 XThC.Tn[7].t14 VGND 0.01636f
C10478 XThC.Tn[7].n33 VGND 0.03652f
C10479 XThC.Tn[7].n34 VGND 0.02502f
C10480 XThC.Tn[7].n35 VGND 0.08235f
C10481 XThC.Tn[7].n36 VGND 0.13573f
C10482 XThC.Tn[7].t12 VGND 0.01498f
C10483 XThC.Tn[7].t16 VGND 0.01636f
C10484 XThC.Tn[7].n37 VGND 0.03652f
C10485 XThC.Tn[7].n38 VGND 0.02502f
C10486 XThC.Tn[7].n39 VGND 0.08235f
C10487 XThC.Tn[7].n40 VGND 0.13573f
C10488 XThC.Tn[7].t31 VGND 0.01498f
C10489 XThC.Tn[7].t36 VGND 0.01636f
C10490 XThC.Tn[7].n41 VGND 0.03652f
C10491 XThC.Tn[7].n42 VGND 0.02502f
C10492 XThC.Tn[7].n43 VGND 0.08235f
C10493 XThC.Tn[7].n44 VGND 0.13573f
C10494 XThC.Tn[7].t32 VGND 0.01498f
C10495 XThC.Tn[7].t38 VGND 0.01636f
C10496 XThC.Tn[7].n45 VGND 0.03652f
C10497 XThC.Tn[7].n46 VGND 0.02502f
C10498 XThC.Tn[7].n47 VGND 0.08235f
C10499 XThC.Tn[7].n48 VGND 0.13573f
C10500 XThC.Tn[7].t13 VGND 0.01498f
C10501 XThC.Tn[7].t17 VGND 0.01636f
C10502 XThC.Tn[7].n49 VGND 0.03652f
C10503 XThC.Tn[7].n50 VGND 0.02502f
C10504 XThC.Tn[7].n51 VGND 0.08235f
C10505 XThC.Tn[7].n52 VGND 0.13573f
C10506 XThC.Tn[7].t21 VGND 0.01498f
C10507 XThC.Tn[7].t26 VGND 0.01636f
C10508 XThC.Tn[7].n53 VGND 0.03652f
C10509 XThC.Tn[7].n54 VGND 0.02502f
C10510 XThC.Tn[7].n55 VGND 0.08235f
C10511 XThC.Tn[7].n56 VGND 0.13573f
C10512 XThC.Tn[7].t24 VGND 0.01498f
C10513 XThC.Tn[7].t28 VGND 0.01636f
C10514 XThC.Tn[7].n57 VGND 0.03652f
C10515 XThC.Tn[7].n58 VGND 0.02502f
C10516 XThC.Tn[7].n59 VGND 0.08235f
C10517 XThC.Tn[7].n60 VGND 0.13573f
C10518 XThC.Tn[7].t37 VGND 0.01498f
C10519 XThC.Tn[7].t9 VGND 0.01636f
C10520 XThC.Tn[7].n61 VGND 0.03652f
C10521 XThC.Tn[7].n62 VGND 0.02502f
C10522 XThC.Tn[7].n63 VGND 0.08235f
C10523 XThC.Tn[7].n64 VGND 0.13573f
C10524 XThC.Tn[7].t15 VGND 0.01498f
C10525 XThC.Tn[7].t19 VGND 0.01636f
C10526 XThC.Tn[7].n65 VGND 0.03652f
C10527 XThC.Tn[7].n66 VGND 0.02502f
C10528 XThC.Tn[7].n67 VGND 0.08235f
C10529 XThC.Tn[7].n68 VGND 0.13573f
C10530 XThC.Tn[7].n69 VGND 0.34086f
C10531 XThC.Tn[7].n70 VGND 0.02261f
C10532 XThR.Tn[1].t4 VGND 0.02304f
C10533 XThR.Tn[1].t5 VGND 0.02304f
C10534 XThR.Tn[1].n0 VGND 0.0465f
C10535 XThR.Tn[1].t7 VGND 0.02304f
C10536 XThR.Tn[1].t6 VGND 0.02304f
C10537 XThR.Tn[1].n1 VGND 0.05441f
C10538 XThR.Tn[1].n2 VGND 0.15232f
C10539 XThR.Tn[1].t11 VGND 0.01497f
C10540 XThR.Tn[1].t8 VGND 0.01497f
C10541 XThR.Tn[1].n3 VGND 0.0341f
C10542 XThR.Tn[1].t10 VGND 0.01497f
C10543 XThR.Tn[1].t9 VGND 0.01497f
C10544 XThR.Tn[1].n4 VGND 0.0341f
C10545 XThR.Tn[1].t2 VGND 0.01497f
C10546 XThR.Tn[1].t1 VGND 0.01497f
C10547 XThR.Tn[1].n5 VGND 0.0341f
C10548 XThR.Tn[1].t3 VGND 0.01497f
C10549 XThR.Tn[1].t0 VGND 0.01497f
C10550 XThR.Tn[1].n6 VGND 0.05682f
C10551 XThR.Tn[1].n7 VGND 0.16239f
C10552 XThR.Tn[1].n8 VGND 0.10039f
C10553 XThR.Tn[1].n9 VGND 0.11329f
C10554 XThR.Tn[1].t24 VGND 0.01801f
C10555 XThR.Tn[1].t18 VGND 0.01972f
C10556 XThR.Tn[1].n10 VGND 0.04814f
C10557 XThR.Tn[1].n11 VGND 0.09248f
C10558 XThR.Tn[1].t44 VGND 0.01801f
C10559 XThR.Tn[1].t34 VGND 0.01972f
C10560 XThR.Tn[1].n12 VGND 0.04814f
C10561 XThR.Tn[1].t61 VGND 0.01795f
C10562 XThR.Tn[1].t30 VGND 0.01965f
C10563 XThR.Tn[1].n13 VGND 0.05009f
C10564 XThR.Tn[1].n14 VGND 0.03519f
C10565 XThR.Tn[1].n15 VGND 0.00643f
C10566 XThR.Tn[1].n16 VGND 0.11293f
C10567 XThR.Tn[1].t19 VGND 0.01801f
C10568 XThR.Tn[1].t73 VGND 0.01972f
C10569 XThR.Tn[1].n17 VGND 0.04814f
C10570 XThR.Tn[1].t38 VGND 0.01795f
C10571 XThR.Tn[1].t69 VGND 0.01965f
C10572 XThR.Tn[1].n18 VGND 0.05009f
C10573 XThR.Tn[1].n19 VGND 0.03519f
C10574 XThR.Tn[1].n20 VGND 0.00643f
C10575 XThR.Tn[1].n21 VGND 0.11293f
C10576 XThR.Tn[1].t35 VGND 0.01801f
C10577 XThR.Tn[1].t28 VGND 0.01972f
C10578 XThR.Tn[1].n22 VGND 0.04814f
C10579 XThR.Tn[1].t50 VGND 0.01795f
C10580 XThR.Tn[1].t25 VGND 0.01965f
C10581 XThR.Tn[1].n23 VGND 0.05009f
C10582 XThR.Tn[1].n24 VGND 0.03519f
C10583 XThR.Tn[1].n25 VGND 0.00643f
C10584 XThR.Tn[1].n26 VGND 0.11293f
C10585 XThR.Tn[1].t59 VGND 0.01801f
C10586 XThR.Tn[1].t55 VGND 0.01972f
C10587 XThR.Tn[1].n27 VGND 0.04814f
C10588 XThR.Tn[1].t21 VGND 0.01795f
C10589 XThR.Tn[1].t51 VGND 0.01965f
C10590 XThR.Tn[1].n28 VGND 0.05009f
C10591 XThR.Tn[1].n29 VGND 0.03519f
C10592 XThR.Tn[1].n30 VGND 0.00643f
C10593 XThR.Tn[1].n31 VGND 0.11293f
C10594 XThR.Tn[1].t37 VGND 0.01801f
C10595 XThR.Tn[1].t29 VGND 0.01972f
C10596 XThR.Tn[1].n32 VGND 0.04814f
C10597 XThR.Tn[1].t53 VGND 0.01795f
C10598 XThR.Tn[1].t26 VGND 0.01965f
C10599 XThR.Tn[1].n33 VGND 0.05009f
C10600 XThR.Tn[1].n34 VGND 0.03519f
C10601 XThR.Tn[1].n35 VGND 0.00643f
C10602 XThR.Tn[1].n36 VGND 0.11293f
C10603 XThR.Tn[1].t13 VGND 0.01801f
C10604 XThR.Tn[1].t46 VGND 0.01972f
C10605 XThR.Tn[1].n37 VGND 0.04814f
C10606 XThR.Tn[1].t32 VGND 0.01795f
C10607 XThR.Tn[1].t43 VGND 0.01965f
C10608 XThR.Tn[1].n38 VGND 0.05009f
C10609 XThR.Tn[1].n39 VGND 0.03519f
C10610 XThR.Tn[1].n40 VGND 0.00643f
C10611 XThR.Tn[1].n41 VGND 0.11293f
C10612 XThR.Tn[1].t45 VGND 0.01801f
C10613 XThR.Tn[1].t41 VGND 0.01972f
C10614 XThR.Tn[1].n42 VGND 0.04814f
C10615 XThR.Tn[1].t60 VGND 0.01795f
C10616 XThR.Tn[1].t36 VGND 0.01965f
C10617 XThR.Tn[1].n43 VGND 0.05009f
C10618 XThR.Tn[1].n44 VGND 0.03519f
C10619 XThR.Tn[1].n45 VGND 0.00643f
C10620 XThR.Tn[1].n46 VGND 0.11293f
C10621 XThR.Tn[1].t48 VGND 0.01801f
C10622 XThR.Tn[1].t54 VGND 0.01972f
C10623 XThR.Tn[1].n47 VGND 0.04814f
C10624 XThR.Tn[1].t67 VGND 0.01795f
C10625 XThR.Tn[1].t49 VGND 0.01965f
C10626 XThR.Tn[1].n48 VGND 0.05009f
C10627 XThR.Tn[1].n49 VGND 0.03519f
C10628 XThR.Tn[1].n50 VGND 0.00643f
C10629 XThR.Tn[1].n51 VGND 0.11293f
C10630 XThR.Tn[1].t64 VGND 0.01801f
C10631 XThR.Tn[1].t12 VGND 0.01972f
C10632 XThR.Tn[1].n52 VGND 0.04814f
C10633 XThR.Tn[1].t23 VGND 0.01795f
C10634 XThR.Tn[1].t71 VGND 0.01965f
C10635 XThR.Tn[1].n53 VGND 0.05009f
C10636 XThR.Tn[1].n54 VGND 0.03519f
C10637 XThR.Tn[1].n55 VGND 0.00643f
C10638 XThR.Tn[1].n56 VGND 0.11293f
C10639 XThR.Tn[1].t57 VGND 0.01801f
C10640 XThR.Tn[1].t31 VGND 0.01972f
C10641 XThR.Tn[1].n57 VGND 0.04814f
C10642 XThR.Tn[1].t16 VGND 0.01795f
C10643 XThR.Tn[1].t27 VGND 0.01965f
C10644 XThR.Tn[1].n58 VGND 0.05009f
C10645 XThR.Tn[1].n59 VGND 0.03519f
C10646 XThR.Tn[1].n60 VGND 0.00643f
C10647 XThR.Tn[1].n61 VGND 0.11293f
C10648 XThR.Tn[1].t15 VGND 0.01801f
C10649 XThR.Tn[1].t68 VGND 0.01972f
C10650 XThR.Tn[1].n62 VGND 0.04814f
C10651 XThR.Tn[1].t33 VGND 0.01795f
C10652 XThR.Tn[1].t63 VGND 0.01965f
C10653 XThR.Tn[1].n63 VGND 0.05009f
C10654 XThR.Tn[1].n64 VGND 0.03519f
C10655 XThR.Tn[1].n65 VGND 0.00643f
C10656 XThR.Tn[1].n66 VGND 0.11293f
C10657 XThR.Tn[1].t47 VGND 0.01801f
C10658 XThR.Tn[1].t42 VGND 0.01972f
C10659 XThR.Tn[1].n67 VGND 0.04814f
C10660 XThR.Tn[1].t65 VGND 0.01795f
C10661 XThR.Tn[1].t39 VGND 0.01965f
C10662 XThR.Tn[1].n68 VGND 0.05009f
C10663 XThR.Tn[1].n69 VGND 0.03519f
C10664 XThR.Tn[1].n70 VGND 0.00643f
C10665 XThR.Tn[1].n71 VGND 0.11293f
C10666 XThR.Tn[1].t62 VGND 0.01801f
C10667 XThR.Tn[1].t56 VGND 0.01972f
C10668 XThR.Tn[1].n72 VGND 0.04814f
C10669 XThR.Tn[1].t22 VGND 0.01795f
C10670 XThR.Tn[1].t52 VGND 0.01965f
C10671 XThR.Tn[1].n73 VGND 0.05009f
C10672 XThR.Tn[1].n74 VGND 0.03519f
C10673 XThR.Tn[1].n75 VGND 0.00643f
C10674 XThR.Tn[1].n76 VGND 0.11293f
C10675 XThR.Tn[1].t20 VGND 0.01801f
C10676 XThR.Tn[1].t14 VGND 0.01972f
C10677 XThR.Tn[1].n77 VGND 0.04814f
C10678 XThR.Tn[1].t40 VGND 0.01795f
C10679 XThR.Tn[1].t72 VGND 0.01965f
C10680 XThR.Tn[1].n78 VGND 0.05009f
C10681 XThR.Tn[1].n79 VGND 0.03519f
C10682 XThR.Tn[1].n80 VGND 0.00643f
C10683 XThR.Tn[1].n81 VGND 0.11293f
C10684 XThR.Tn[1].t58 VGND 0.01801f
C10685 XThR.Tn[1].t70 VGND 0.01972f
C10686 XThR.Tn[1].n82 VGND 0.04814f
C10687 XThR.Tn[1].t17 VGND 0.01795f
C10688 XThR.Tn[1].t66 VGND 0.01965f
C10689 XThR.Tn[1].n83 VGND 0.05009f
C10690 XThR.Tn[1].n84 VGND 0.03519f
C10691 XThR.Tn[1].n85 VGND 0.00643f
C10692 XThR.Tn[1].n86 VGND 0.11293f
C10693 XThR.Tn[1].n87 VGND 0.10263f
C10694 XThR.Tn[1].n88 VGND 0.29541f
C10695 XThR.Tn[1].n89 VGND 0.04821f
C10696 XThC.Tn[8].t9 VGND 0.01304f
C10697 XThC.Tn[8].t8 VGND 0.01304f
C10698 XThC.Tn[8].n0 VGND 0.03253f
C10699 XThC.Tn[8].t11 VGND 0.01304f
C10700 XThC.Tn[8].t10 VGND 0.01304f
C10701 XThC.Tn[8].n1 VGND 0.02608f
C10702 XThC.Tn[8].n2 VGND 0.06561f
C10703 XThC.Tn[8].n3 VGND 0.02453f
C10704 XThC.Tn[8].t43 VGND 0.0159f
C10705 XThC.Tn[8].t41 VGND 0.01737f
C10706 XThC.Tn[8].n4 VGND 0.03878f
C10707 XThC.Tn[8].n5 VGND 0.02657f
C10708 XThC.Tn[8].n6 VGND 0.0872f
C10709 XThC.Tn[8].t29 VGND 0.0159f
C10710 XThC.Tn[8].t26 VGND 0.01737f
C10711 XThC.Tn[8].n7 VGND 0.03878f
C10712 XThC.Tn[8].n8 VGND 0.02657f
C10713 XThC.Tn[8].n9 VGND 0.08744f
C10714 XThC.Tn[8].n10 VGND 0.1441f
C10715 XThC.Tn[8].t34 VGND 0.0159f
C10716 XThC.Tn[8].t28 VGND 0.01737f
C10717 XThC.Tn[8].n11 VGND 0.03878f
C10718 XThC.Tn[8].n12 VGND 0.02657f
C10719 XThC.Tn[8].n13 VGND 0.08744f
C10720 XThC.Tn[8].n14 VGND 0.1441f
C10721 XThC.Tn[8].t35 VGND 0.0159f
C10722 XThC.Tn[8].t30 VGND 0.01737f
C10723 XThC.Tn[8].n15 VGND 0.03878f
C10724 XThC.Tn[8].n16 VGND 0.02657f
C10725 XThC.Tn[8].n17 VGND 0.08744f
C10726 XThC.Tn[8].n18 VGND 0.1441f
C10727 XThC.Tn[8].t22 VGND 0.0159f
C10728 XThC.Tn[8].t19 VGND 0.01737f
C10729 XThC.Tn[8].n19 VGND 0.03878f
C10730 XThC.Tn[8].n20 VGND 0.02657f
C10731 XThC.Tn[8].n21 VGND 0.08744f
C10732 XThC.Tn[8].n22 VGND 0.1441f
C10733 XThC.Tn[8].t23 VGND 0.0159f
C10734 XThC.Tn[8].t20 VGND 0.01737f
C10735 XThC.Tn[8].n23 VGND 0.03878f
C10736 XThC.Tn[8].n24 VGND 0.02657f
C10737 XThC.Tn[8].n25 VGND 0.08744f
C10738 XThC.Tn[8].n26 VGND 0.1441f
C10739 XThC.Tn[8].t39 VGND 0.0159f
C10740 XThC.Tn[8].t33 VGND 0.01737f
C10741 XThC.Tn[8].n27 VGND 0.03878f
C10742 XThC.Tn[8].n28 VGND 0.02657f
C10743 XThC.Tn[8].n29 VGND 0.08744f
C10744 XThC.Tn[8].n30 VGND 0.1441f
C10745 XThC.Tn[8].t14 VGND 0.0159f
C10746 XThC.Tn[8].t42 VGND 0.01737f
C10747 XThC.Tn[8].n31 VGND 0.03878f
C10748 XThC.Tn[8].n32 VGND 0.02657f
C10749 XThC.Tn[8].n33 VGND 0.08744f
C10750 XThC.Tn[8].n34 VGND 0.1441f
C10751 XThC.Tn[8].t16 VGND 0.0159f
C10752 XThC.Tn[8].t12 VGND 0.01737f
C10753 XThC.Tn[8].n35 VGND 0.03878f
C10754 XThC.Tn[8].n36 VGND 0.02657f
C10755 XThC.Tn[8].n37 VGND 0.08744f
C10756 XThC.Tn[8].n38 VGND 0.1441f
C10757 XThC.Tn[8].t36 VGND 0.0159f
C10758 XThC.Tn[8].t31 VGND 0.01737f
C10759 XThC.Tn[8].n39 VGND 0.03878f
C10760 XThC.Tn[8].n40 VGND 0.02657f
C10761 XThC.Tn[8].n41 VGND 0.08744f
C10762 XThC.Tn[8].n42 VGND 0.1441f
C10763 XThC.Tn[8].t38 VGND 0.0159f
C10764 XThC.Tn[8].t32 VGND 0.01737f
C10765 XThC.Tn[8].n43 VGND 0.03878f
C10766 XThC.Tn[8].n44 VGND 0.02657f
C10767 XThC.Tn[8].n45 VGND 0.08744f
C10768 XThC.Tn[8].n46 VGND 0.1441f
C10769 XThC.Tn[8].t17 VGND 0.0159f
C10770 XThC.Tn[8].t13 VGND 0.01737f
C10771 XThC.Tn[8].n47 VGND 0.03878f
C10772 XThC.Tn[8].n48 VGND 0.02657f
C10773 XThC.Tn[8].n49 VGND 0.08744f
C10774 XThC.Tn[8].n50 VGND 0.1441f
C10775 XThC.Tn[8].t25 VGND 0.0159f
C10776 XThC.Tn[8].t21 VGND 0.01737f
C10777 XThC.Tn[8].n51 VGND 0.03878f
C10778 XThC.Tn[8].n52 VGND 0.02657f
C10779 XThC.Tn[8].n53 VGND 0.08744f
C10780 XThC.Tn[8].n54 VGND 0.1441f
C10781 XThC.Tn[8].t27 VGND 0.0159f
C10782 XThC.Tn[8].t24 VGND 0.01737f
C10783 XThC.Tn[8].n55 VGND 0.03878f
C10784 XThC.Tn[8].n56 VGND 0.02657f
C10785 XThC.Tn[8].n57 VGND 0.08744f
C10786 XThC.Tn[8].n58 VGND 0.1441f
C10787 XThC.Tn[8].t40 VGND 0.0159f
C10788 XThC.Tn[8].t37 VGND 0.01737f
C10789 XThC.Tn[8].n59 VGND 0.03878f
C10790 XThC.Tn[8].n60 VGND 0.02657f
C10791 XThC.Tn[8].n61 VGND 0.08744f
C10792 XThC.Tn[8].n62 VGND 0.1441f
C10793 XThC.Tn[8].t18 VGND 0.0159f
C10794 XThC.Tn[8].t15 VGND 0.01737f
C10795 XThC.Tn[8].n63 VGND 0.03878f
C10796 XThC.Tn[8].n64 VGND 0.02657f
C10797 XThC.Tn[8].n65 VGND 0.08744f
C10798 XThC.Tn[8].n66 VGND 0.1441f
C10799 XThC.Tn[8].n67 VGND 0.60346f
C10800 XThC.Tn[8].n68 VGND 0.23618f
C10801 XThC.Tn[8].t5 VGND 0.02006f
C10802 XThC.Tn[8].t6 VGND 0.02006f
C10803 XThC.Tn[8].n69 VGND 0.04335f
C10804 XThC.Tn[8].t4 VGND 0.02006f
C10805 XThC.Tn[8].t7 VGND 0.02006f
C10806 XThC.Tn[8].n70 VGND 0.06598f
C10807 XThC.Tn[8].n71 VGND 0.18333f
C10808 XThC.Tn[8].n72 VGND 0.02883f
C10809 XThC.Tn[8].t2 VGND 0.02006f
C10810 XThC.Tn[8].t1 VGND 0.02006f
C10811 XThC.Tn[8].n73 VGND 0.0446f
C10812 XThC.Tn[8].t0 VGND 0.02006f
C10813 XThC.Tn[8].t3 VGND 0.02006f
C10814 XThC.Tn[8].n74 VGND 0.06092f
C10815 XThC.Tn[8].n75 VGND 0.1985f
C10816 XThC.XTB1.Y.t2 VGND 0.03224f
C10817 XThC.XTB1.Y.n0 VGND 0.02084f
C10818 XThC.XTB1.Y.n1 VGND 0.02659f
C10819 XThC.XTB1.Y.t1 VGND 0.01618f
C10820 XThC.XTB1.Y.t0 VGND 0.01618f
C10821 XThC.XTB1.Y.n2 VGND 0.03473f
C10822 XThC.XTB1.Y.t17 VGND 0.02517f
C10823 XThC.XTB1.Y.t5 VGND 0.01483f
C10824 XThC.XTB1.Y.n3 VGND 0.02997f
C10825 XThC.XTB1.Y.t6 VGND 0.02517f
C10826 XThC.XTB1.Y.t12 VGND 0.01483f
C10827 XThC.XTB1.Y.n4 VGND 0.01542f
C10828 XThC.XTB1.Y.t8 VGND 0.02517f
C10829 XThC.XTB1.Y.t13 VGND 0.01483f
C10830 XThC.XTB1.Y.n5 VGND 0.03313f
C10831 XThC.XTB1.Y.t11 VGND 0.02517f
C10832 XThC.XTB1.Y.t16 VGND 0.01483f
C10833 XThC.XTB1.Y.n6 VGND 0.03076f
C10834 XThC.XTB1.Y.n7 VGND 0.01871f
C10835 XThC.XTB1.Y.n8 VGND 0.03098f
C10836 XThC.XTB1.Y.n9 VGND 0.01198f
C10837 XThC.XTB1.Y.n10 VGND 0.01463f
C10838 XThC.XTB1.Y.n11 VGND 0.03313f
C10839 XThC.XTB1.Y.n12 VGND 0.01661f
C10840 XThC.XTB1.Y.n13 VGND 0.02824f
C10841 XThC.XTB1.Y.t18 VGND 0.02517f
C10842 XThC.XTB1.Y.t9 VGND 0.01483f
C10843 XThC.XTB1.Y.n14 VGND 0.03392f
C10844 XThC.XTB1.Y.t7 VGND 0.02517f
C10845 XThC.XTB1.Y.t15 VGND 0.01483f
C10846 XThC.XTB1.Y.t14 VGND 0.02517f
C10847 XThC.XTB1.Y.t3 VGND 0.01483f
C10848 XThC.XTB1.Y.t10 VGND 0.02517f
C10849 XThC.XTB1.Y.t4 VGND 0.01483f
C10850 XThC.XTB1.Y.n15 VGND 0.04223f
C10851 XThC.XTB1.Y.n16 VGND 0.0446f
C10852 XThC.XTB1.Y.n17 VGND 0.01719f
C10853 XThC.XTB1.Y.n18 VGND 0.0363f
C10854 XThC.XTB1.Y.n19 VGND 0.01661f
C10855 XThC.XTB1.Y.n20 VGND 0.01378f
C10856 XThC.XTB1.Y.n21 VGND 0.77148f
C10857 XThC.XTB1.Y.n22 VGND 0.07634f
C10858 XThC.Tn[14].t4 VGND 0.01262f
C10859 XThC.Tn[14].t6 VGND 0.01262f
C10860 XThC.Tn[14].n0 VGND 0.03148f
C10861 XThC.Tn[14].t5 VGND 0.01262f
C10862 XThC.Tn[14].t7 VGND 0.01262f
C10863 XThC.Tn[14].n1 VGND 0.02524f
C10864 XThC.Tn[14].n2 VGND 0.06349f
C10865 XThC.Tn[14].t43 VGND 0.01539f
C10866 XThC.Tn[14].t38 VGND 0.01681f
C10867 XThC.Tn[14].n3 VGND 0.03752f
C10868 XThC.Tn[14].n4 VGND 0.02571f
C10869 XThC.Tn[14].n5 VGND 0.08438f
C10870 XThC.Tn[14].t29 VGND 0.01539f
C10871 XThC.Tn[14].t22 VGND 0.01681f
C10872 XThC.Tn[14].n6 VGND 0.03752f
C10873 XThC.Tn[14].n7 VGND 0.02571f
C10874 XThC.Tn[14].n8 VGND 0.08461f
C10875 XThC.Tn[14].n9 VGND 0.13945f
C10876 XThC.Tn[14].t32 VGND 0.01539f
C10877 XThC.Tn[14].t25 VGND 0.01681f
C10878 XThC.Tn[14].n10 VGND 0.03752f
C10879 XThC.Tn[14].n11 VGND 0.02571f
C10880 XThC.Tn[14].n12 VGND 0.08461f
C10881 XThC.Tn[14].n13 VGND 0.13945f
C10882 XThC.Tn[14].t34 VGND 0.01539f
C10883 XThC.Tn[14].t26 VGND 0.01681f
C10884 XThC.Tn[14].n14 VGND 0.03752f
C10885 XThC.Tn[14].n15 VGND 0.02571f
C10886 XThC.Tn[14].n16 VGND 0.08461f
C10887 XThC.Tn[14].n17 VGND 0.13945f
C10888 XThC.Tn[14].t20 VGND 0.01539f
C10889 XThC.Tn[14].t14 VGND 0.01681f
C10890 XThC.Tn[14].n18 VGND 0.03752f
C10891 XThC.Tn[14].n19 VGND 0.02571f
C10892 XThC.Tn[14].n20 VGND 0.08461f
C10893 XThC.Tn[14].n21 VGND 0.13945f
C10894 XThC.Tn[14].t23 VGND 0.01539f
C10895 XThC.Tn[14].t17 VGND 0.01681f
C10896 XThC.Tn[14].n22 VGND 0.03752f
C10897 XThC.Tn[14].n23 VGND 0.02571f
C10898 XThC.Tn[14].n24 VGND 0.08461f
C10899 XThC.Tn[14].n25 VGND 0.13945f
C10900 XThC.Tn[14].t37 VGND 0.01539f
C10901 XThC.Tn[14].t31 VGND 0.01681f
C10902 XThC.Tn[14].n26 VGND 0.03752f
C10903 XThC.Tn[14].n27 VGND 0.02571f
C10904 XThC.Tn[14].n28 VGND 0.08461f
C10905 XThC.Tn[14].n29 VGND 0.13945f
C10906 XThC.Tn[14].t13 VGND 0.01539f
C10907 XThC.Tn[14].t39 VGND 0.01681f
C10908 XThC.Tn[14].n30 VGND 0.03752f
C10909 XThC.Tn[14].n31 VGND 0.02571f
C10910 XThC.Tn[14].n32 VGND 0.08461f
C10911 XThC.Tn[14].n33 VGND 0.13945f
C10912 XThC.Tn[14].t15 VGND 0.01539f
C10913 XThC.Tn[14].t41 VGND 0.01681f
C10914 XThC.Tn[14].n34 VGND 0.03752f
C10915 XThC.Tn[14].n35 VGND 0.02571f
C10916 XThC.Tn[14].n36 VGND 0.08461f
C10917 XThC.Tn[14].n37 VGND 0.13945f
C10918 XThC.Tn[14].t35 VGND 0.01539f
C10919 XThC.Tn[14].t27 VGND 0.01681f
C10920 XThC.Tn[14].n38 VGND 0.03752f
C10921 XThC.Tn[14].n39 VGND 0.02571f
C10922 XThC.Tn[14].n40 VGND 0.08461f
C10923 XThC.Tn[14].n41 VGND 0.13945f
C10924 XThC.Tn[14].t36 VGND 0.01539f
C10925 XThC.Tn[14].t30 VGND 0.01681f
C10926 XThC.Tn[14].n42 VGND 0.03752f
C10927 XThC.Tn[14].n43 VGND 0.02571f
C10928 XThC.Tn[14].n44 VGND 0.08461f
C10929 XThC.Tn[14].n45 VGND 0.13945f
C10930 XThC.Tn[14].t16 VGND 0.01539f
C10931 XThC.Tn[14].t42 VGND 0.01681f
C10932 XThC.Tn[14].n46 VGND 0.03752f
C10933 XThC.Tn[14].n47 VGND 0.02571f
C10934 XThC.Tn[14].n48 VGND 0.08461f
C10935 XThC.Tn[14].n49 VGND 0.13945f
C10936 XThC.Tn[14].t24 VGND 0.01539f
C10937 XThC.Tn[14].t19 VGND 0.01681f
C10938 XThC.Tn[14].n50 VGND 0.03752f
C10939 XThC.Tn[14].n51 VGND 0.02571f
C10940 XThC.Tn[14].n52 VGND 0.08461f
C10941 XThC.Tn[14].n53 VGND 0.13945f
C10942 XThC.Tn[14].t28 VGND 0.01539f
C10943 XThC.Tn[14].t21 VGND 0.01681f
C10944 XThC.Tn[14].n54 VGND 0.03752f
C10945 XThC.Tn[14].n55 VGND 0.02571f
C10946 XThC.Tn[14].n56 VGND 0.08461f
C10947 XThC.Tn[14].n57 VGND 0.13945f
C10948 XThC.Tn[14].t40 VGND 0.01539f
C10949 XThC.Tn[14].t33 VGND 0.01681f
C10950 XThC.Tn[14].n58 VGND 0.03752f
C10951 XThC.Tn[14].n59 VGND 0.02571f
C10952 XThC.Tn[14].n60 VGND 0.08461f
C10953 XThC.Tn[14].n61 VGND 0.13945f
C10954 XThC.Tn[14].t18 VGND 0.01539f
C10955 XThC.Tn[14].t12 VGND 0.01681f
C10956 XThC.Tn[14].n62 VGND 0.03752f
C10957 XThC.Tn[14].n63 VGND 0.02571f
C10958 XThC.Tn[14].n64 VGND 0.08461f
C10959 XThC.Tn[14].n65 VGND 0.13945f
C10960 XThC.Tn[14].n66 VGND 0.91462f
C10961 XThC.Tn[14].n67 VGND 0.26906f
C10962 XThC.Tn[14].t0 VGND 0.01942f
C10963 XThC.Tn[14].t1 VGND 0.01942f
C10964 XThC.Tn[14].n68 VGND 0.04195f
C10965 XThC.Tn[14].t3 VGND 0.01942f
C10966 XThC.Tn[14].t2 VGND 0.01942f
C10967 XThC.Tn[14].n69 VGND 0.06385f
C10968 XThC.Tn[14].n70 VGND 0.1774f
C10969 XThC.Tn[14].n71 VGND 0.02789f
C10970 XThC.Tn[14].t11 VGND 0.01942f
C10971 XThC.Tn[14].t10 VGND 0.01942f
C10972 XThC.Tn[14].n72 VGND 0.05895f
C10973 XThC.Tn[14].t9 VGND 0.01942f
C10974 XThC.Tn[14].t8 VGND 0.01942f
C10975 XThC.Tn[14].n73 VGND 0.04316f
C10976 XThC.Tn[14].n74 VGND 0.19209f
C10977 XThR.Tn[10].t9 VGND 0.02415f
C10978 XThR.Tn[10].t7 VGND 0.02415f
C10979 XThR.Tn[10].n0 VGND 0.07333f
C10980 XThR.Tn[10].t10 VGND 0.02415f
C10981 XThR.Tn[10].t8 VGND 0.02415f
C10982 XThR.Tn[10].n1 VGND 0.05368f
C10983 XThR.Tn[10].n2 VGND 0.2441f
C10984 XThR.Tn[10].t2 VGND 0.0157f
C10985 XThR.Tn[10].t6 VGND 0.0157f
C10986 XThR.Tn[10].n3 VGND 0.03915f
C10987 XThR.Tn[10].t4 VGND 0.0157f
C10988 XThR.Tn[10].t11 VGND 0.0157f
C10989 XThR.Tn[10].n4 VGND 0.0314f
C10990 XThR.Tn[10].n5 VGND 0.07239f
C10991 XThR.Tn[10].t54 VGND 0.01887f
C10992 XThR.Tn[10].t47 VGND 0.02067f
C10993 XThR.Tn[10].n6 VGND 0.05047f
C10994 XThR.Tn[10].n7 VGND 0.09695f
C10995 XThR.Tn[10].t13 VGND 0.01887f
C10996 XThR.Tn[10].t63 VGND 0.02067f
C10997 XThR.Tn[10].n8 VGND 0.05047f
C10998 XThR.Tn[10].t50 VGND 0.01881f
C10999 XThR.Tn[10].t60 VGND 0.0206f
C11000 XThR.Tn[10].n9 VGND 0.05251f
C11001 XThR.Tn[10].n10 VGND 0.03689f
C11002 XThR.Tn[10].n11 VGND 0.00674f
C11003 XThR.Tn[10].n12 VGND 0.11838f
C11004 XThR.Tn[10].t48 VGND 0.01887f
C11005 XThR.Tn[10].t41 VGND 0.02067f
C11006 XThR.Tn[10].n13 VGND 0.05047f
C11007 XThR.Tn[10].t23 VGND 0.01881f
C11008 XThR.Tn[10].t36 VGND 0.0206f
C11009 XThR.Tn[10].n14 VGND 0.05251f
C11010 XThR.Tn[10].n15 VGND 0.03689f
C11011 XThR.Tn[10].n16 VGND 0.00674f
C11012 XThR.Tn[10].n17 VGND 0.11838f
C11013 XThR.Tn[10].t65 VGND 0.01887f
C11014 XThR.Tn[10].t58 VGND 0.02067f
C11015 XThR.Tn[10].n18 VGND 0.05047f
C11016 XThR.Tn[10].t40 VGND 0.01881f
C11017 XThR.Tn[10].t55 VGND 0.0206f
C11018 XThR.Tn[10].n19 VGND 0.05251f
C11019 XThR.Tn[10].n20 VGND 0.03689f
C11020 XThR.Tn[10].n21 VGND 0.00674f
C11021 XThR.Tn[10].n22 VGND 0.11838f
C11022 XThR.Tn[10].t30 VGND 0.01887f
C11023 XThR.Tn[10].t26 VGND 0.02067f
C11024 XThR.Tn[10].n23 VGND 0.05047f
C11025 XThR.Tn[10].t70 VGND 0.01881f
C11026 XThR.Tn[10].t21 VGND 0.0206f
C11027 XThR.Tn[10].n24 VGND 0.05251f
C11028 XThR.Tn[10].n25 VGND 0.03689f
C11029 XThR.Tn[10].n26 VGND 0.00674f
C11030 XThR.Tn[10].n27 VGND 0.11838f
C11031 XThR.Tn[10].t67 VGND 0.01887f
C11032 XThR.Tn[10].t59 VGND 0.02067f
C11033 XThR.Tn[10].n28 VGND 0.05047f
C11034 XThR.Tn[10].t42 VGND 0.01881f
C11035 XThR.Tn[10].t56 VGND 0.0206f
C11036 XThR.Tn[10].n29 VGND 0.05251f
C11037 XThR.Tn[10].n30 VGND 0.03689f
C11038 XThR.Tn[10].n31 VGND 0.00674f
C11039 XThR.Tn[10].n32 VGND 0.11838f
C11040 XThR.Tn[10].t44 VGND 0.01887f
C11041 XThR.Tn[10].t15 VGND 0.02067f
C11042 XThR.Tn[10].n33 VGND 0.05047f
C11043 XThR.Tn[10].t18 VGND 0.01881f
C11044 XThR.Tn[10].t12 VGND 0.0206f
C11045 XThR.Tn[10].n34 VGND 0.05251f
C11046 XThR.Tn[10].n35 VGND 0.03689f
C11047 XThR.Tn[10].n36 VGND 0.00674f
C11048 XThR.Tn[10].n37 VGND 0.11838f
C11049 XThR.Tn[10].t14 VGND 0.01887f
C11050 XThR.Tn[10].t69 VGND 0.02067f
C11051 XThR.Tn[10].n38 VGND 0.05047f
C11052 XThR.Tn[10].t51 VGND 0.01881f
C11053 XThR.Tn[10].t66 VGND 0.0206f
C11054 XThR.Tn[10].n39 VGND 0.05251f
C11055 XThR.Tn[10].n40 VGND 0.03689f
C11056 XThR.Tn[10].n41 VGND 0.00674f
C11057 XThR.Tn[10].n42 VGND 0.11838f
C11058 XThR.Tn[10].t17 VGND 0.01887f
C11059 XThR.Tn[10].t24 VGND 0.02067f
C11060 XThR.Tn[10].n43 VGND 0.05047f
C11061 XThR.Tn[10].t53 VGND 0.01881f
C11062 XThR.Tn[10].t20 VGND 0.0206f
C11063 XThR.Tn[10].n44 VGND 0.05251f
C11064 XThR.Tn[10].n45 VGND 0.03689f
C11065 XThR.Tn[10].n46 VGND 0.00674f
C11066 XThR.Tn[10].n47 VGND 0.11838f
C11067 XThR.Tn[10].t33 VGND 0.01887f
C11068 XThR.Tn[10].t43 VGND 0.02067f
C11069 XThR.Tn[10].n48 VGND 0.05047f
C11070 XThR.Tn[10].t73 VGND 0.01881f
C11071 XThR.Tn[10].t38 VGND 0.0206f
C11072 XThR.Tn[10].n49 VGND 0.05251f
C11073 XThR.Tn[10].n50 VGND 0.03689f
C11074 XThR.Tn[10].n51 VGND 0.00674f
C11075 XThR.Tn[10].n52 VGND 0.11838f
C11076 XThR.Tn[10].t28 VGND 0.01887f
C11077 XThR.Tn[10].t61 VGND 0.02067f
C11078 XThR.Tn[10].n53 VGND 0.05047f
C11079 XThR.Tn[10].t62 VGND 0.01881f
C11080 XThR.Tn[10].t57 VGND 0.0206f
C11081 XThR.Tn[10].n54 VGND 0.05251f
C11082 XThR.Tn[10].n55 VGND 0.03689f
C11083 XThR.Tn[10].n56 VGND 0.00674f
C11084 XThR.Tn[10].n57 VGND 0.11838f
C11085 XThR.Tn[10].t46 VGND 0.01887f
C11086 XThR.Tn[10].t35 VGND 0.02067f
C11087 XThR.Tn[10].n58 VGND 0.05047f
C11088 XThR.Tn[10].t19 VGND 0.01881f
C11089 XThR.Tn[10].t32 VGND 0.0206f
C11090 XThR.Tn[10].n59 VGND 0.05251f
C11091 XThR.Tn[10].n60 VGND 0.03689f
C11092 XThR.Tn[10].n61 VGND 0.00674f
C11093 XThR.Tn[10].n62 VGND 0.11838f
C11094 XThR.Tn[10].t16 VGND 0.01887f
C11095 XThR.Tn[10].t72 VGND 0.02067f
C11096 XThR.Tn[10].n63 VGND 0.05047f
C11097 XThR.Tn[10].t52 VGND 0.01881f
C11098 XThR.Tn[10].t68 VGND 0.0206f
C11099 XThR.Tn[10].n64 VGND 0.05251f
C11100 XThR.Tn[10].n65 VGND 0.03689f
C11101 XThR.Tn[10].n66 VGND 0.00674f
C11102 XThR.Tn[10].n67 VGND 0.11838f
C11103 XThR.Tn[10].t31 VGND 0.01887f
C11104 XThR.Tn[10].t27 VGND 0.02067f
C11105 XThR.Tn[10].n68 VGND 0.05047f
C11106 XThR.Tn[10].t71 VGND 0.01881f
C11107 XThR.Tn[10].t22 VGND 0.0206f
C11108 XThR.Tn[10].n69 VGND 0.05251f
C11109 XThR.Tn[10].n70 VGND 0.03689f
C11110 XThR.Tn[10].n71 VGND 0.00674f
C11111 XThR.Tn[10].n72 VGND 0.11838f
C11112 XThR.Tn[10].t49 VGND 0.01887f
C11113 XThR.Tn[10].t45 VGND 0.02067f
C11114 XThR.Tn[10].n73 VGND 0.05047f
C11115 XThR.Tn[10].t25 VGND 0.01881f
C11116 XThR.Tn[10].t39 VGND 0.0206f
C11117 XThR.Tn[10].n74 VGND 0.05251f
C11118 XThR.Tn[10].n75 VGND 0.03689f
C11119 XThR.Tn[10].n76 VGND 0.00674f
C11120 XThR.Tn[10].n77 VGND 0.11838f
C11121 XThR.Tn[10].t29 VGND 0.01887f
C11122 XThR.Tn[10].t37 VGND 0.02067f
C11123 XThR.Tn[10].n78 VGND 0.05047f
C11124 XThR.Tn[10].t64 VGND 0.01881f
C11125 XThR.Tn[10].t34 VGND 0.0206f
C11126 XThR.Tn[10].n79 VGND 0.05251f
C11127 XThR.Tn[10].n80 VGND 0.03689f
C11128 XThR.Tn[10].n81 VGND 0.00674f
C11129 XThR.Tn[10].n82 VGND 0.11838f
C11130 XThR.Tn[10].n83 VGND 0.10758f
C11131 XThR.Tn[10].n84 VGND 0.3312f
C11132 XThR.Tn[10].t3 VGND 0.02415f
C11133 XThR.Tn[10].t0 VGND 0.02415f
C11134 XThR.Tn[10].n85 VGND 0.05218f
C11135 XThR.Tn[10].t1 VGND 0.02415f
C11136 XThR.Tn[10].t5 VGND 0.02415f
C11137 XThR.Tn[10].n86 VGND 0.07942f
C11138 XThR.Tn[10].n87 VGND 0.22051f
C11139 XThR.Tn[10].n88 VGND 0.01087f
C11140 XThC.Tn[3].t1 VGND 0.01826f
C11141 XThC.Tn[3].t0 VGND 0.01826f
C11142 XThC.Tn[3].n0 VGND 0.03685f
C11143 XThC.Tn[3].t3 VGND 0.01826f
C11144 XThC.Tn[3].t2 VGND 0.01826f
C11145 XThC.Tn[3].n1 VGND 0.04312f
C11146 XThC.Tn[3].n2 VGND 0.12934f
C11147 XThC.Tn[3].t11 VGND 0.01187f
C11148 XThC.Tn[3].t10 VGND 0.01187f
C11149 XThC.Tn[3].n3 VGND 0.04503f
C11150 XThC.Tn[3].t9 VGND 0.01187f
C11151 XThC.Tn[3].t8 VGND 0.01187f
C11152 XThC.Tn[3].n4 VGND 0.02703f
C11153 XThC.Tn[3].n5 VGND 0.1287f
C11154 XThC.Tn[3].t7 VGND 0.01187f
C11155 XThC.Tn[3].t6 VGND 0.01187f
C11156 XThC.Tn[3].n6 VGND 0.02703f
C11157 XThC.Tn[3].n7 VGND 0.07956f
C11158 XThC.Tn[3].t5 VGND 0.01187f
C11159 XThC.Tn[3].t4 VGND 0.01187f
C11160 XThC.Tn[3].n8 VGND 0.02703f
C11161 XThC.Tn[3].n9 VGND 0.08979f
C11162 XThC.Tn[3].t12 VGND 0.01447f
C11163 XThC.Tn[3].t42 VGND 0.01581f
C11164 XThC.Tn[3].n10 VGND 0.03529f
C11165 XThC.Tn[3].n11 VGND 0.02417f
C11166 XThC.Tn[3].n12 VGND 0.07935f
C11167 XThC.Tn[3].t30 VGND 0.01447f
C11168 XThC.Tn[3].t27 VGND 0.01581f
C11169 XThC.Tn[3].n13 VGND 0.03529f
C11170 XThC.Tn[3].n14 VGND 0.02417f
C11171 XThC.Tn[3].n15 VGND 0.07957f
C11172 XThC.Tn[3].n16 VGND 0.13113f
C11173 XThC.Tn[3].t35 VGND 0.01447f
C11174 XThC.Tn[3].t29 VGND 0.01581f
C11175 XThC.Tn[3].n17 VGND 0.03529f
C11176 XThC.Tn[3].n18 VGND 0.02417f
C11177 XThC.Tn[3].n19 VGND 0.07957f
C11178 XThC.Tn[3].n20 VGND 0.13113f
C11179 XThC.Tn[3].t36 VGND 0.01447f
C11180 XThC.Tn[3].t31 VGND 0.01581f
C11181 XThC.Tn[3].n21 VGND 0.03529f
C11182 XThC.Tn[3].n22 VGND 0.02417f
C11183 XThC.Tn[3].n23 VGND 0.07957f
C11184 XThC.Tn[3].n24 VGND 0.13113f
C11185 XThC.Tn[3].t23 VGND 0.01447f
C11186 XThC.Tn[3].t20 VGND 0.01581f
C11187 XThC.Tn[3].n25 VGND 0.03529f
C11188 XThC.Tn[3].n26 VGND 0.02417f
C11189 XThC.Tn[3].n27 VGND 0.07957f
C11190 XThC.Tn[3].n28 VGND 0.13113f
C11191 XThC.Tn[3].t24 VGND 0.01447f
C11192 XThC.Tn[3].t21 VGND 0.01581f
C11193 XThC.Tn[3].n29 VGND 0.03529f
C11194 XThC.Tn[3].n30 VGND 0.02417f
C11195 XThC.Tn[3].n31 VGND 0.07957f
C11196 XThC.Tn[3].n32 VGND 0.13113f
C11197 XThC.Tn[3].t40 VGND 0.01447f
C11198 XThC.Tn[3].t34 VGND 0.01581f
C11199 XThC.Tn[3].n33 VGND 0.03529f
C11200 XThC.Tn[3].n34 VGND 0.02417f
C11201 XThC.Tn[3].n35 VGND 0.07957f
C11202 XThC.Tn[3].n36 VGND 0.13113f
C11203 XThC.Tn[3].t15 VGND 0.01447f
C11204 XThC.Tn[3].t43 VGND 0.01581f
C11205 XThC.Tn[3].n37 VGND 0.03529f
C11206 XThC.Tn[3].n38 VGND 0.02417f
C11207 XThC.Tn[3].n39 VGND 0.07957f
C11208 XThC.Tn[3].n40 VGND 0.13113f
C11209 XThC.Tn[3].t17 VGND 0.01447f
C11210 XThC.Tn[3].t13 VGND 0.01581f
C11211 XThC.Tn[3].n41 VGND 0.03529f
C11212 XThC.Tn[3].n42 VGND 0.02417f
C11213 XThC.Tn[3].n43 VGND 0.07957f
C11214 XThC.Tn[3].n44 VGND 0.13113f
C11215 XThC.Tn[3].t37 VGND 0.01447f
C11216 XThC.Tn[3].t32 VGND 0.01581f
C11217 XThC.Tn[3].n45 VGND 0.03529f
C11218 XThC.Tn[3].n46 VGND 0.02417f
C11219 XThC.Tn[3].n47 VGND 0.07957f
C11220 XThC.Tn[3].n48 VGND 0.13113f
C11221 XThC.Tn[3].t39 VGND 0.01447f
C11222 XThC.Tn[3].t33 VGND 0.01581f
C11223 XThC.Tn[3].n49 VGND 0.03529f
C11224 XThC.Tn[3].n50 VGND 0.02417f
C11225 XThC.Tn[3].n51 VGND 0.07957f
C11226 XThC.Tn[3].n52 VGND 0.13113f
C11227 XThC.Tn[3].t18 VGND 0.01447f
C11228 XThC.Tn[3].t14 VGND 0.01581f
C11229 XThC.Tn[3].n53 VGND 0.03529f
C11230 XThC.Tn[3].n54 VGND 0.02417f
C11231 XThC.Tn[3].n55 VGND 0.07957f
C11232 XThC.Tn[3].n56 VGND 0.13113f
C11233 XThC.Tn[3].t26 VGND 0.01447f
C11234 XThC.Tn[3].t22 VGND 0.01581f
C11235 XThC.Tn[3].n57 VGND 0.03529f
C11236 XThC.Tn[3].n58 VGND 0.02417f
C11237 XThC.Tn[3].n59 VGND 0.07957f
C11238 XThC.Tn[3].n60 VGND 0.13113f
C11239 XThC.Tn[3].t28 VGND 0.01447f
C11240 XThC.Tn[3].t25 VGND 0.01581f
C11241 XThC.Tn[3].n61 VGND 0.03529f
C11242 XThC.Tn[3].n62 VGND 0.02417f
C11243 XThC.Tn[3].n63 VGND 0.07957f
C11244 XThC.Tn[3].n64 VGND 0.13113f
C11245 XThC.Tn[3].t41 VGND 0.01447f
C11246 XThC.Tn[3].t38 VGND 0.01581f
C11247 XThC.Tn[3].n65 VGND 0.03529f
C11248 XThC.Tn[3].n66 VGND 0.02417f
C11249 XThC.Tn[3].n67 VGND 0.07957f
C11250 XThC.Tn[3].n68 VGND 0.13113f
C11251 XThC.Tn[3].t19 VGND 0.01447f
C11252 XThC.Tn[3].t16 VGND 0.01581f
C11253 XThC.Tn[3].n69 VGND 0.03529f
C11254 XThC.Tn[3].n70 VGND 0.02417f
C11255 XThC.Tn[3].n71 VGND 0.07957f
C11256 XThC.Tn[3].n72 VGND 0.13113f
C11257 XThC.Tn[3].n73 VGND 0.77119f
C11258 XThC.Tn[3].n74 VGND 0.1112f
C11259 XThC.Tn[1].t3 VGND 0.01715f
C11260 XThC.Tn[1].t2 VGND 0.01715f
C11261 XThC.Tn[1].n0 VGND 0.03462f
C11262 XThC.Tn[1].t1 VGND 0.01715f
C11263 XThC.Tn[1].t0 VGND 0.01715f
C11264 XThC.Tn[1].n1 VGND 0.04051f
C11265 XThC.Tn[1].n2 VGND 0.12152f
C11266 XThC.Tn[1].t11 VGND 0.01115f
C11267 XThC.Tn[1].t10 VGND 0.01115f
C11268 XThC.Tn[1].n3 VGND 0.04231f
C11269 XThC.Tn[1].t9 VGND 0.01115f
C11270 XThC.Tn[1].t8 VGND 0.01115f
C11271 XThC.Tn[1].n4 VGND 0.02539f
C11272 XThC.Tn[1].n5 VGND 0.12091f
C11273 XThC.Tn[1].t7 VGND 0.01115f
C11274 XThC.Tn[1].t6 VGND 0.01115f
C11275 XThC.Tn[1].n6 VGND 0.02539f
C11276 XThC.Tn[1].n7 VGND 0.07475f
C11277 XThC.Tn[1].t5 VGND 0.01115f
C11278 XThC.Tn[1].t4 VGND 0.01115f
C11279 XThC.Tn[1].n8 VGND 0.02539f
C11280 XThC.Tn[1].n9 VGND 0.08436f
C11281 XThC.Tn[1].t31 VGND 0.0136f
C11282 XThC.Tn[1].t29 VGND 0.01485f
C11283 XThC.Tn[1].n10 VGND 0.03315f
C11284 XThC.Tn[1].n11 VGND 0.02271f
C11285 XThC.Tn[1].n12 VGND 0.07455f
C11286 XThC.Tn[1].t17 VGND 0.0136f
C11287 XThC.Tn[1].t14 VGND 0.01485f
C11288 XThC.Tn[1].n13 VGND 0.03315f
C11289 XThC.Tn[1].n14 VGND 0.02271f
C11290 XThC.Tn[1].n15 VGND 0.07475f
C11291 XThC.Tn[1].n16 VGND 0.1232f
C11292 XThC.Tn[1].t22 VGND 0.0136f
C11293 XThC.Tn[1].t16 VGND 0.01485f
C11294 XThC.Tn[1].n17 VGND 0.03315f
C11295 XThC.Tn[1].n18 VGND 0.02271f
C11296 XThC.Tn[1].n19 VGND 0.07475f
C11297 XThC.Tn[1].n20 VGND 0.1232f
C11298 XThC.Tn[1].t23 VGND 0.0136f
C11299 XThC.Tn[1].t18 VGND 0.01485f
C11300 XThC.Tn[1].n21 VGND 0.03315f
C11301 XThC.Tn[1].n22 VGND 0.02271f
C11302 XThC.Tn[1].n23 VGND 0.07475f
C11303 XThC.Tn[1].n24 VGND 0.1232f
C11304 XThC.Tn[1].t42 VGND 0.0136f
C11305 XThC.Tn[1].t39 VGND 0.01485f
C11306 XThC.Tn[1].n25 VGND 0.03315f
C11307 XThC.Tn[1].n26 VGND 0.02271f
C11308 XThC.Tn[1].n27 VGND 0.07475f
C11309 XThC.Tn[1].n28 VGND 0.1232f
C11310 XThC.Tn[1].t43 VGND 0.0136f
C11311 XThC.Tn[1].t40 VGND 0.01485f
C11312 XThC.Tn[1].n29 VGND 0.03315f
C11313 XThC.Tn[1].n30 VGND 0.02271f
C11314 XThC.Tn[1].n31 VGND 0.07475f
C11315 XThC.Tn[1].n32 VGND 0.1232f
C11316 XThC.Tn[1].t27 VGND 0.0136f
C11317 XThC.Tn[1].t21 VGND 0.01485f
C11318 XThC.Tn[1].n33 VGND 0.03315f
C11319 XThC.Tn[1].n34 VGND 0.02271f
C11320 XThC.Tn[1].n35 VGND 0.07475f
C11321 XThC.Tn[1].n36 VGND 0.1232f
C11322 XThC.Tn[1].t34 VGND 0.0136f
C11323 XThC.Tn[1].t30 VGND 0.01485f
C11324 XThC.Tn[1].n37 VGND 0.03315f
C11325 XThC.Tn[1].n38 VGND 0.02271f
C11326 XThC.Tn[1].n39 VGND 0.07475f
C11327 XThC.Tn[1].n40 VGND 0.1232f
C11328 XThC.Tn[1].t36 VGND 0.0136f
C11329 XThC.Tn[1].t32 VGND 0.01485f
C11330 XThC.Tn[1].n41 VGND 0.03315f
C11331 XThC.Tn[1].n42 VGND 0.02271f
C11332 XThC.Tn[1].n43 VGND 0.07475f
C11333 XThC.Tn[1].n44 VGND 0.1232f
C11334 XThC.Tn[1].t24 VGND 0.0136f
C11335 XThC.Tn[1].t19 VGND 0.01485f
C11336 XThC.Tn[1].n45 VGND 0.03315f
C11337 XThC.Tn[1].n46 VGND 0.02271f
C11338 XThC.Tn[1].n47 VGND 0.07475f
C11339 XThC.Tn[1].n48 VGND 0.1232f
C11340 XThC.Tn[1].t26 VGND 0.0136f
C11341 XThC.Tn[1].t20 VGND 0.01485f
C11342 XThC.Tn[1].n49 VGND 0.03315f
C11343 XThC.Tn[1].n50 VGND 0.02271f
C11344 XThC.Tn[1].n51 VGND 0.07475f
C11345 XThC.Tn[1].n52 VGND 0.1232f
C11346 XThC.Tn[1].t37 VGND 0.0136f
C11347 XThC.Tn[1].t33 VGND 0.01485f
C11348 XThC.Tn[1].n53 VGND 0.03315f
C11349 XThC.Tn[1].n54 VGND 0.02271f
C11350 XThC.Tn[1].n55 VGND 0.07475f
C11351 XThC.Tn[1].n56 VGND 0.1232f
C11352 XThC.Tn[1].t13 VGND 0.0136f
C11353 XThC.Tn[1].t41 VGND 0.01485f
C11354 XThC.Tn[1].n57 VGND 0.03315f
C11355 XThC.Tn[1].n58 VGND 0.02271f
C11356 XThC.Tn[1].n59 VGND 0.07475f
C11357 XThC.Tn[1].n60 VGND 0.1232f
C11358 XThC.Tn[1].t15 VGND 0.0136f
C11359 XThC.Tn[1].t12 VGND 0.01485f
C11360 XThC.Tn[1].n61 VGND 0.03315f
C11361 XThC.Tn[1].n62 VGND 0.02271f
C11362 XThC.Tn[1].n63 VGND 0.07475f
C11363 XThC.Tn[1].n64 VGND 0.1232f
C11364 XThC.Tn[1].t28 VGND 0.0136f
C11365 XThC.Tn[1].t25 VGND 0.01485f
C11366 XThC.Tn[1].n65 VGND 0.03315f
C11367 XThC.Tn[1].n66 VGND 0.02271f
C11368 XThC.Tn[1].n67 VGND 0.07475f
C11369 XThC.Tn[1].n68 VGND 0.1232f
C11370 XThC.Tn[1].t38 VGND 0.0136f
C11371 XThC.Tn[1].t35 VGND 0.01485f
C11372 XThC.Tn[1].n69 VGND 0.03315f
C11373 XThC.Tn[1].n70 VGND 0.02271f
C11374 XThC.Tn[1].n71 VGND 0.07475f
C11375 XThC.Tn[1].n72 VGND 0.1232f
C11376 XThC.Tn[1].n73 VGND 0.62603f
C11377 XThC.Tn[1].n74 VGND 0.11896f
C11378 Vbias.t2 VGND 0.30464f
C11379 Vbias.t1 VGND 1.19882f
C11380 Vbias.n0 VGND 2.23968f
C11381 Vbias.t4 VGND 0.06536f
C11382 Vbias.t3 VGND 0.06536f
C11383 Vbias.n1 VGND 0.44035f
C11384 Vbias.t5 VGND 0.06536f
C11385 Vbias.t0 VGND 0.06536f
C11386 Vbias.n2 VGND 0.44035f
C11387 Vbias.n3 VGND 1.32031f
C11388 Vbias.n4 VGND 0.92467f
C11389 Vbias.n5 VGND 0.99869f
C11390 Vbias.t181 VGND 0.31986f
C11391 Vbias.n6 VGND 0.3159f
C11392 Vbias.t110 VGND 0.31986f
C11393 Vbias.n7 VGND 0.3159f
C11394 Vbias.n8 VGND 0.08895f
C11395 Vbias.n9 VGND 0.33621f
C11396 Vbias.t146 VGND 0.31986f
C11397 Vbias.n10 VGND 0.3159f
C11398 Vbias.t238 VGND 0.31986f
C11399 Vbias.n11 VGND 0.3159f
C11400 Vbias.n12 VGND 0.33621f
C11401 Vbias.t210 VGND 0.31986f
C11402 Vbias.n13 VGND 0.3159f
C11403 Vbias.n14 VGND 0.08895f
C11404 Vbias.t24 VGND 0.31986f
C11405 Vbias.n15 VGND 0.3159f
C11406 Vbias.t12 VGND 0.31986f
C11407 Vbias.n16 VGND 0.3159f
C11408 Vbias.n17 VGND 0.33621f
C11409 Vbias.t193 VGND 0.31986f
C11410 Vbias.n18 VGND 0.3159f
C11411 Vbias.n19 VGND 0.18787f
C11412 Vbias.n20 VGND 0.18787f
C11413 Vbias.t173 VGND 0.31986f
C11414 Vbias.n21 VGND 0.3159f
C11415 Vbias.n22 VGND 0.33621f
C11416 Vbias.t248 VGND 0.31986f
C11417 Vbias.n23 VGND 0.3159f
C11418 Vbias.t95 VGND 0.31986f
C11419 Vbias.n24 VGND 0.3159f
C11420 Vbias.n25 VGND 0.33621f
C11421 Vbias.t25 VGND 0.31986f
C11422 Vbias.n26 VGND 0.3159f
C11423 Vbias.t258 VGND 0.31986f
C11424 Vbias.n27 VGND 0.3159f
C11425 Vbias.n28 VGND 0.33621f
C11426 Vbias.t75 VGND 0.31986f
C11427 Vbias.n29 VGND 0.3159f
C11428 Vbias.t246 VGND 0.31986f
C11429 Vbias.n30 VGND 0.3159f
C11430 Vbias.n31 VGND 0.33621f
C11431 Vbias.t171 VGND 0.31986f
C11432 Vbias.n32 VGND 0.3159f
C11433 Vbias.t96 VGND 0.31986f
C11434 Vbias.n33 VGND 0.3159f
C11435 Vbias.n34 VGND 0.33621f
C11436 Vbias.t169 VGND 0.31986f
C11437 Vbias.n35 VGND 0.3159f
C11438 Vbias.t147 VGND 0.31986f
C11439 Vbias.n36 VGND 0.3159f
C11440 Vbias.n37 VGND 0.33621f
C11441 Vbias.t76 VGND 0.31986f
C11442 Vbias.n38 VGND 0.3159f
C11443 Vbias.t247 VGND 0.31986f
C11444 Vbias.n39 VGND 0.3159f
C11445 Vbias.n40 VGND 0.33621f
C11446 Vbias.t60 VGND 0.31986f
C11447 Vbias.n41 VGND 0.3159f
C11448 Vbias.t227 VGND 0.31986f
C11449 Vbias.n42 VGND 0.3159f
C11450 Vbias.n43 VGND 0.33621f
C11451 Vbias.t156 VGND 0.31986f
C11452 Vbias.n44 VGND 0.3159f
C11453 Vbias.t69 VGND 0.31986f
C11454 Vbias.n45 VGND 0.3159f
C11455 Vbias.n46 VGND 0.33621f
C11456 Vbias.t141 VGND 0.31986f
C11457 Vbias.n47 VGND 0.3159f
C11458 Vbias.t56 VGND 0.31986f
C11459 Vbias.n48 VGND 0.3159f
C11460 Vbias.n49 VGND 0.33621f
C11461 Vbias.t242 VGND 0.31986f
C11462 Vbias.n50 VGND 0.3159f
C11463 Vbias.t229 VGND 0.31986f
C11464 Vbias.n51 VGND 0.3159f
C11465 Vbias.n52 VGND 0.33621f
C11466 Vbias.t41 VGND 0.31986f
C11467 Vbias.n53 VGND 0.3159f
C11468 Vbias.t201 VGND 0.31986f
C11469 Vbias.n54 VGND 0.3159f
C11470 Vbias.n55 VGND 0.33621f
C11471 Vbias.t130 VGND 0.31986f
C11472 Vbias.n56 VGND 0.3159f
C11473 Vbias.t57 VGND 0.31986f
C11474 Vbias.n57 VGND 0.3159f
C11475 Vbias.t129 VGND 0.31986f
C11476 Vbias.n58 VGND 0.3159f
C11477 Vbias.n59 VGND 0.04244f
C11478 Vbias.t87 VGND 0.31986f
C11479 Vbias.n60 VGND 0.3159f
C11480 Vbias.t225 VGND 0.31986f
C11481 Vbias.n61 VGND 0.3159f
C11482 Vbias.n62 VGND 0.08895f
C11483 Vbias.n63 VGND 0.18787f
C11484 Vbias.t205 VGND 0.31986f
C11485 Vbias.n64 VGND 0.3159f
C11486 Vbias.n65 VGND 0.08895f
C11487 Vbias.n66 VGND 0.18787f
C11488 Vbias.t52 VGND 0.31986f
C11489 Vbias.n67 VGND 0.3159f
C11490 Vbias.n68 VGND 0.08895f
C11491 Vbias.n69 VGND 0.18787f
C11492 Vbias.t32 VGND 0.31986f
C11493 Vbias.n70 VGND 0.3159f
C11494 Vbias.n71 VGND 0.08895f
C11495 Vbias.n72 VGND 0.18787f
C11496 Vbias.t199 VGND 0.31986f
C11497 Vbias.n73 VGND 0.3159f
C11498 Vbias.n74 VGND 0.08895f
C11499 Vbias.n75 VGND 0.18787f
C11500 Vbias.t125 VGND 0.31986f
C11501 Vbias.n76 VGND 0.3159f
C11502 Vbias.n77 VGND 0.08895f
C11503 Vbias.n78 VGND 0.18787f
C11504 Vbias.t102 VGND 0.31986f
C11505 Vbias.n79 VGND 0.3159f
C11506 Vbias.n80 VGND 0.08895f
C11507 Vbias.n81 VGND 0.18787f
C11508 Vbias.t18 VGND 0.31986f
C11509 Vbias.n82 VGND 0.3159f
C11510 Vbias.n83 VGND 0.08895f
C11511 Vbias.n84 VGND 0.18787f
C11512 Vbias.t183 VGND 0.31986f
C11513 Vbias.n85 VGND 0.3159f
C11514 Vbias.n86 VGND 0.08895f
C11515 Vbias.n87 VGND 0.18787f
C11516 Vbias.t99 VGND 0.31986f
C11517 Vbias.n88 VGND 0.3159f
C11518 Vbias.n89 VGND 0.08895f
C11519 Vbias.n90 VGND 0.18787f
C11520 Vbias.t14 VGND 0.31986f
C11521 Vbias.n91 VGND 0.3159f
C11522 Vbias.n92 VGND 0.08895f
C11523 Vbias.n93 VGND 0.18787f
C11524 Vbias.t261 VGND 0.31986f
C11525 Vbias.n94 VGND 0.3159f
C11526 Vbias.n95 VGND 0.08895f
C11527 Vbias.n96 VGND 0.18787f
C11528 Vbias.t160 VGND 0.31986f
C11529 Vbias.n97 VGND 0.3159f
C11530 Vbias.n98 VGND 0.08895f
C11531 Vbias.n99 VGND 0.18787f
C11532 Vbias.n100 VGND 0.08634f
C11533 Vbias.n101 VGND 0.33621f
C11534 Vbias.t16 VGND 0.31986f
C11535 Vbias.n102 VGND 0.3159f
C11536 Vbias.t88 VGND 0.31986f
C11537 Vbias.n103 VGND 0.3159f
C11538 Vbias.n104 VGND 0.33621f
C11539 Vbias.t17 VGND 0.31986f
C11540 Vbias.n105 VGND 0.3159f
C11541 Vbias.t113 VGND 0.31986f
C11542 Vbias.n106 VGND 0.3159f
C11543 Vbias.n107 VGND 0.33621f
C11544 Vbias.t185 VGND 0.31986f
C11545 Vbias.n108 VGND 0.3159f
C11546 Vbias.t196 VGND 0.31986f
C11547 Vbias.n109 VGND 0.3159f
C11548 Vbias.n110 VGND 0.33621f
C11549 Vbias.t124 VGND 0.31986f
C11550 Vbias.n111 VGND 0.3159f
C11551 Vbias.t213 VGND 0.31986f
C11552 Vbias.n112 VGND 0.3159f
C11553 Vbias.n113 VGND 0.33621f
C11554 Vbias.t29 VGND 0.31986f
C11555 Vbias.n114 VGND 0.3159f
C11556 Vbias.t112 VGND 0.31986f
C11557 Vbias.n115 VGND 0.3159f
C11558 Vbias.n116 VGND 0.33621f
C11559 Vbias.t40 VGND 0.31986f
C11560 Vbias.n117 VGND 0.3159f
C11561 Vbias.t127 VGND 0.31986f
C11562 Vbias.n118 VGND 0.3159f
C11563 Vbias.n119 VGND 0.33621f
C11564 Vbias.t200 VGND 0.31986f
C11565 Vbias.n120 VGND 0.3159f
C11566 Vbias.t33 VGND 0.31986f
C11567 Vbias.n121 VGND 0.3159f
C11568 Vbias.n122 VGND 0.33621f
C11569 Vbias.t219 VGND 0.31986f
C11570 Vbias.n123 VGND 0.3159f
C11571 Vbias.t240 VGND 0.31986f
C11572 Vbias.n124 VGND 0.3159f
C11573 Vbias.n125 VGND 0.33621f
C11574 Vbias.t53 VGND 0.31986f
C11575 Vbias.n126 VGND 0.3159f
C11576 Vbias.t126 VGND 0.31986f
C11577 Vbias.n127 VGND 0.3159f
C11578 Vbias.n128 VGND 0.33621f
C11579 Vbias.t54 VGND 0.31986f
C11580 Vbias.n129 VGND 0.3159f
C11581 Vbias.t144 VGND 0.31986f
C11582 Vbias.n130 VGND 0.3159f
C11583 Vbias.n131 VGND 0.33621f
C11584 Vbias.t217 VGND 0.31986f
C11585 Vbias.n132 VGND 0.3159f
C11586 Vbias.t239 VGND 0.31986f
C11587 Vbias.n133 VGND 0.3159f
C11588 Vbias.n134 VGND 0.33621f
C11589 Vbias.t166 VGND 0.31986f
C11590 Vbias.n135 VGND 0.3159f
C11591 Vbias.t62 VGND 0.31986f
C11592 Vbias.n136 VGND 0.3159f
C11593 Vbias.n137 VGND 0.33621f
C11594 Vbias.t133 VGND 0.31986f
C11595 Vbias.n138 VGND 0.3159f
C11596 Vbias.t153 VGND 0.31986f
C11597 Vbias.n139 VGND 0.3159f
C11598 Vbias.n140 VGND 0.33621f
C11599 Vbias.t81 VGND 0.31986f
C11600 Vbias.n141 VGND 0.3159f
C11601 Vbias.t92 VGND 0.31986f
C11602 Vbias.n142 VGND 0.3159f
C11603 Vbias.n143 VGND 0.33621f
C11604 Vbias.t20 VGND 0.31986f
C11605 Vbias.n144 VGND 0.3159f
C11606 Vbias.t121 VGND 0.31986f
C11607 Vbias.n145 VGND 0.3159f
C11608 Vbias.t49 VGND 0.31986f
C11609 Vbias.n146 VGND 0.3159f
C11610 Vbias.n147 VGND 0.08634f
C11611 Vbias.n148 VGND 0.33621f
C11612 Vbias.t82 VGND 0.31986f
C11613 Vbias.n149 VGND 0.3159f
C11614 Vbias.t154 VGND 0.31986f
C11615 Vbias.n150 VGND 0.3159f
C11616 Vbias.n151 VGND 0.33621f
C11617 Vbias.t122 VGND 0.31986f
C11618 Vbias.n152 VGND 0.3159f
C11619 Vbias.t222 VGND 0.31986f
C11620 Vbias.n153 VGND 0.3159f
C11621 Vbias.n154 VGND 0.33621f
C11622 Vbias.t257 VGND 0.31986f
C11623 Vbias.n155 VGND 0.3159f
C11624 Vbias.t8 VGND 0.31986f
C11625 Vbias.n156 VGND 0.3159f
C11626 Vbias.n157 VGND 0.33621f
C11627 Vbias.t235 VGND 0.31986f
C11628 Vbias.n158 VGND 0.3159f
C11629 Vbias.t63 VGND 0.31986f
C11630 Vbias.n159 VGND 0.3159f
C11631 Vbias.n160 VGND 0.33621f
C11632 Vbias.t93 VGND 0.31986f
C11633 Vbias.n161 VGND 0.3159f
C11634 Vbias.t179 VGND 0.31986f
C11635 Vbias.n162 VGND 0.3159f
C11636 Vbias.n163 VGND 0.33621f
C11637 Vbias.t150 VGND 0.31986f
C11638 Vbias.n164 VGND 0.3159f
C11639 Vbias.t237 VGND 0.31986f
C11640 Vbias.n165 VGND 0.3159f
C11641 Vbias.n166 VGND 0.33621f
C11642 Vbias.t11 VGND 0.31986f
C11643 Vbias.n167 VGND 0.3159f
C11644 Vbias.t98 VGND 0.31986f
C11645 Vbias.n168 VGND 0.3159f
C11646 Vbias.n169 VGND 0.33621f
C11647 Vbias.t68 VGND 0.31986f
C11648 Vbias.n170 VGND 0.3159f
C11649 Vbias.t91 VGND 0.31986f
C11650 Vbias.n171 VGND 0.3159f
C11651 Vbias.n172 VGND 0.33621f
C11652 Vbias.t118 VGND 0.31986f
C11653 Vbias.n173 VGND 0.3159f
C11654 Vbias.t190 VGND 0.31986f
C11655 Vbias.n174 VGND 0.3159f
C11656 Vbias.n175 VGND 0.33621f
C11657 Vbias.t164 VGND 0.31986f
C11658 Vbias.n176 VGND 0.3159f
C11659 Vbias.t251 VGND 0.31986f
C11660 Vbias.n177 VGND 0.3159f
C11661 Vbias.n178 VGND 0.33621f
C11662 Vbias.t27 VGND 0.31986f
C11663 Vbias.n179 VGND 0.3159f
C11664 Vbias.t44 VGND 0.31986f
C11665 Vbias.n180 VGND 0.3159f
C11666 Vbias.n181 VGND 0.33621f
C11667 Vbias.t21 VGND 0.31986f
C11668 Vbias.n182 VGND 0.3159f
C11669 Vbias.t168 VGND 0.31986f
C11670 Vbias.n183 VGND 0.3159f
C11671 Vbias.n184 VGND 0.33621f
C11672 Vbias.t197 VGND 0.31986f
C11673 Vbias.n185 VGND 0.3159f
C11674 Vbias.t220 VGND 0.31986f
C11675 Vbias.n186 VGND 0.3159f
C11676 Vbias.n187 VGND 0.33621f
C11677 Vbias.t187 VGND 0.31986f
C11678 Vbias.n188 VGND 0.3159f
C11679 Vbias.t105 VGND 0.31986f
C11680 Vbias.n189 VGND 0.3159f
C11681 Vbias.n190 VGND 0.33621f
C11682 Vbias.t137 VGND 0.31986f
C11683 Vbias.n191 VGND 0.3159f
C11684 Vbias.n192 VGND 0.08895f
C11685 Vbias.n193 VGND 0.33621f
C11686 Vbias.t64 VGND 0.31986f
C11687 Vbias.n194 VGND 0.3159f
C11688 Vbias.t9 VGND 0.31986f
C11689 Vbias.n195 VGND 0.3159f
C11690 Vbias.n196 VGND 0.08634f
C11691 Vbias.t83 VGND 0.31986f
C11692 Vbias.n197 VGND 0.3159f
C11693 Vbias.n198 VGND 0.08895f
C11694 Vbias.n199 VGND 0.18787f
C11695 Vbias.t180 VGND 0.31986f
C11696 Vbias.n200 VGND 0.3159f
C11697 Vbias.n201 VGND 0.08895f
C11698 Vbias.n202 VGND 0.18787f
C11699 Vbias.t188 VGND 0.31986f
C11700 Vbias.n203 VGND 0.3159f
C11701 Vbias.n204 VGND 0.08895f
C11702 Vbias.n205 VGND 0.18787f
C11703 Vbias.t23 VGND 0.31986f
C11704 Vbias.n206 VGND 0.3159f
C11705 Vbias.n207 VGND 0.08895f
C11706 Vbias.n208 VGND 0.18787f
C11707 Vbias.t107 VGND 0.31986f
C11708 Vbias.n209 VGND 0.3159f
C11709 Vbias.n210 VGND 0.08895f
C11710 Vbias.n211 VGND 0.18787f
C11711 Vbias.t192 VGND 0.31986f
C11712 Vbias.n212 VGND 0.3159f
C11713 Vbias.n213 VGND 0.08895f
C11714 Vbias.n214 VGND 0.18787f
C11715 Vbias.t28 VGND 0.31986f
C11716 Vbias.n215 VGND 0.3159f
C11717 Vbias.n216 VGND 0.08895f
C11718 Vbias.n217 VGND 0.18787f
C11719 Vbias.t45 VGND 0.31986f
C11720 Vbias.n218 VGND 0.3159f
C11721 Vbias.n219 VGND 0.08895f
C11722 Vbias.n220 VGND 0.18787f
C11723 Vbias.t119 VGND 0.31986f
C11724 Vbias.n221 VGND 0.3159f
C11725 Vbias.n222 VGND 0.08895f
C11726 Vbias.n223 VGND 0.18787f
C11727 Vbias.t211 VGND 0.31986f
C11728 Vbias.n224 VGND 0.3159f
C11729 Vbias.n225 VGND 0.08895f
C11730 Vbias.n226 VGND 0.18787f
C11731 Vbias.t233 VGND 0.31986f
C11732 Vbias.n227 VGND 0.3159f
C11733 Vbias.n228 VGND 0.08895f
C11734 Vbias.n229 VGND 0.18787f
C11735 Vbias.t123 VGND 0.31986f
C11736 Vbias.n230 VGND 0.3159f
C11737 Vbias.n231 VGND 0.08895f
C11738 Vbias.n232 VGND 0.18787f
C11739 Vbias.t149 VGND 0.31986f
C11740 Vbias.n233 VGND 0.3159f
C11741 Vbias.n234 VGND 0.08895f
C11742 Vbias.n235 VGND 0.18787f
C11743 Vbias.t161 VGND 0.31986f
C11744 Vbias.n236 VGND 0.3159f
C11745 Vbias.n237 VGND 0.33621f
C11746 Vbias.t232 VGND 0.31986f
C11747 Vbias.n238 VGND 0.3159f
C11748 Vbias.n239 VGND 0.99869f
C11749 Vbias.t80 VGND 0.31986f
C11750 Vbias.n240 VGND 0.3159f
C11751 Vbias.n241 VGND 0.33621f
C11752 Vbias.t191 VGND 0.31986f
C11753 Vbias.n242 VGND 0.3159f
C11754 Vbias.t172 VGND 0.31986f
C11755 Vbias.n243 VGND 0.3159f
C11756 Vbias.n244 VGND 0.33621f
C11757 Vbias.t51 VGND 0.31986f
C11758 Vbias.n245 VGND 0.3159f
C11759 Vbias.t162 VGND 0.31986f
C11760 Vbias.n246 VGND 0.3159f
C11761 Vbias.n247 VGND 0.33621f
C11762 Vbias.t22 VGND 0.31986f
C11763 Vbias.n248 VGND 0.3159f
C11764 Vbias.t256 VGND 0.31986f
C11765 Vbias.n249 VGND 0.3159f
C11766 Vbias.n250 VGND 0.33621f
C11767 Vbias.t136 VGND 0.31986f
C11768 Vbias.n251 VGND 0.3159f
C11769 Vbias.t46 VGND 0.31986f
C11770 Vbias.n252 VGND 0.3159f
C11771 Vbias.n253 VGND 0.33621f
C11772 Vbias.t167 VGND 0.31986f
C11773 Vbias.n254 VGND 0.3159f
C11774 Vbias.t94 VGND 0.31986f
C11775 Vbias.n255 VGND 0.3159f
C11776 Vbias.n256 VGND 0.33621f
C11777 Vbias.t234 VGND 0.31986f
C11778 Vbias.n257 VGND 0.3159f
C11779 Vbias.t212 VGND 0.31986f
C11780 Vbias.n258 VGND 0.3159f
C11781 Vbias.n259 VGND 0.33621f
C11782 Vbias.t74 VGND 0.31986f
C11783 Vbias.n260 VGND 0.3159f
C11784 Vbias.t244 VGND 0.31986f
C11785 Vbias.n261 VGND 0.3159f
C11786 Vbias.n262 VGND 0.33621f
C11787 Vbias.t120 VGND 0.31986f
C11788 Vbias.n263 VGND 0.3159f
C11789 Vbias.t36 VGND 0.31986f
C11790 Vbias.n264 VGND 0.3159f
C11791 Vbias.n265 VGND 0.33621f
C11792 Vbias.t155 VGND 0.31986f
C11793 Vbias.n266 VGND 0.3159f
C11794 Vbias.t66 VGND 0.31986f
C11795 Vbias.n267 VGND 0.3159f
C11796 Vbias.n268 VGND 0.33621f
C11797 Vbias.t208 VGND 0.31986f
C11798 Vbias.n269 VGND 0.3159f
C11799 Vbias.t117 VGND 0.31986f
C11800 Vbias.n270 VGND 0.3159f
C11801 Vbias.n271 VGND 0.33621f
C11802 Vbias.t241 VGND 0.31986f
C11803 Vbias.n272 VGND 0.3159f
C11804 Vbias.t226 VGND 0.31986f
C11805 Vbias.n273 VGND 0.3159f
C11806 Vbias.n274 VGND 0.33621f
C11807 Vbias.t108 VGND 0.31986f
C11808 Vbias.n275 VGND 0.3159f
C11809 Vbias.t10 VGND 0.31986f
C11810 Vbias.n276 VGND 0.3159f
C11811 Vbias.n277 VGND 0.33621f
C11812 Vbias.t128 VGND 0.31986f
C11813 Vbias.n278 VGND 0.3159f
C11814 Vbias.t55 VGND 0.31986f
C11815 Vbias.n279 VGND 0.3159f
C11816 Vbias.t189 VGND 0.31986f
C11817 Vbias.n280 VGND 0.3159f
C11818 Vbias.n281 VGND 0.08634f
C11819 Vbias.n282 VGND 0.33621f
C11820 Vbias.n283 VGND 0.33621f
C11821 Vbias.t186 VGND 0.31986f
C11822 Vbias.n284 VGND 0.3159f
C11823 Vbias.t85 VGND 0.31986f
C11824 Vbias.n285 VGND 0.3159f
C11825 Vbias.n286 VGND 0.33621f
C11826 Vbias.t207 VGND 0.31986f
C11827 Vbias.n287 VGND 0.3159f
C11828 Vbias.t109 VGND 0.31986f
C11829 Vbias.n288 VGND 0.3159f
C11830 Vbias.t249 VGND 0.31986f
C11831 Vbias.n289 VGND 0.3159f
C11832 Vbias.n290 VGND 0.08895f
C11833 Vbias.n291 VGND 0.33621f
C11834 Vbias.t86 VGND 0.31986f
C11835 Vbias.n292 VGND 0.3159f
C11836 Vbias.t170 VGND 0.31986f
C11837 Vbias.n293 VGND 0.3159f
C11838 Vbias.n294 VGND 0.34679f
C11839 Vbias.t97 VGND 0.31986f
C11840 Vbias.n295 VGND 0.3159f
C11841 Vbias.t77 VGND 0.31986f
C11842 Vbias.n296 VGND 0.3159f
C11843 Vbias.n297 VGND 0.34679f
C11844 Vbias.t148 VGND 0.31986f
C11845 Vbias.n298 VGND 0.3159f
C11846 Vbias.t252 VGND 0.31986f
C11847 Vbias.n299 VGND 0.3159f
C11848 Vbias.n300 VGND 0.34679f
C11849 Vbias.t177 VGND 0.31986f
C11850 Vbias.n301 VGND 0.3159f
C11851 Vbias.t157 VGND 0.31986f
C11852 Vbias.n302 VGND 0.3159f
C11853 Vbias.n303 VGND 0.34679f
C11854 Vbias.t228 VGND 0.31986f
C11855 Vbias.n304 VGND 0.3159f
C11856 Vbias.t143 VGND 0.31986f
C11857 Vbias.n305 VGND 0.3159f
C11858 Vbias.n306 VGND 0.34679f
C11859 Vbias.t71 VGND 0.31986f
C11860 Vbias.n307 VGND 0.3159f
C11861 Vbias.t253 VGND 0.31986f
C11862 Vbias.n308 VGND 0.3159f
C11863 Vbias.n309 VGND 0.34679f
C11864 Vbias.t70 VGND 0.31986f
C11865 Vbias.n310 VGND 0.3159f
C11866 Vbias.t42 VGND 0.31986f
C11867 Vbias.n311 VGND 0.3159f
C11868 Vbias.n312 VGND 0.34679f
C11869 Vbias.t230 VGND 0.31986f
C11870 Vbias.n313 VGND 0.3159f
C11871 Vbias.t145 VGND 0.31986f
C11872 Vbias.n314 VGND 0.3159f
C11873 Vbias.n315 VGND 0.34679f
C11874 Vbias.t218 VGND 0.31986f
C11875 Vbias.n316 VGND 0.3159f
C11876 Vbias.t131 VGND 0.31986f
C11877 Vbias.n317 VGND 0.3159f
C11878 Vbias.n318 VGND 0.34679f
C11879 Vbias.t58 VGND 0.31986f
C11880 Vbias.n319 VGND 0.3159f
C11881 Vbias.t224 VGND 0.31986f
C11882 Vbias.n320 VGND 0.3159f
C11883 Vbias.n321 VGND 0.34679f
C11884 Vbias.t38 VGND 0.31986f
C11885 Vbias.n322 VGND 0.3159f
C11886 Vbias.t214 VGND 0.31986f
C11887 Vbias.n323 VGND 0.3159f
C11888 Vbias.n324 VGND 0.34679f
C11889 Vbias.t139 VGND 0.31986f
C11890 Vbias.n325 VGND 0.3159f
C11891 Vbias.t132 VGND 0.31986f
C11892 Vbias.n326 VGND 0.3159f
C11893 Vbias.n327 VGND 0.34679f
C11894 Vbias.t203 VGND 0.31986f
C11895 Vbias.n328 VGND 0.3159f
C11896 Vbias.t30 VGND 0.31986f
C11897 Vbias.n329 VGND 0.3159f
C11898 Vbias.n330 VGND 0.08634f
C11899 Vbias.t100 VGND 0.31986f
C11900 Vbias.n331 VGND 0.3159f
C11901 Vbias.n332 VGND 0.34679f
C11902 Vbias.t31 VGND 0.31986f
C11903 Vbias.n333 VGND 0.3159f
C11904 Vbias.t215 VGND 0.31986f
C11905 Vbias.n334 VGND 0.3159f
C11906 Vbias.t140 VGND 0.31986f
C11907 Vbias.n335 VGND 0.3159f
C11908 Vbias.n336 VGND 0.08634f
C11909 Vbias.t260 VGND 0.31986f
C11910 Vbias.n337 VGND 0.3159f
C11911 Vbias.t151 VGND 0.31986f
C11912 Vbias.n338 VGND 0.3159f
C11913 Vbias.t35 VGND 0.31986f
C11914 Vbias.n339 VGND 0.3159f
C11915 Vbias.n340 VGND 0.08895f
C11916 Vbias.t104 VGND 0.31986f
C11917 Vbias.n341 VGND 0.3159f
C11918 Vbias.n342 VGND 0.97075f
C11919 Vbias.t216 VGND 0.31986f
C11920 Vbias.n343 VGND 0.3159f
C11921 Vbias.n344 VGND 0.08895f
C11922 Vbias.n345 VGND 0.18787f
C11923 Vbias.t59 VGND 0.31986f
C11924 Vbias.n346 VGND 0.3159f
C11925 Vbias.n347 VGND 0.08895f
C11926 Vbias.n348 VGND 0.18787f
C11927 Vbias.t67 VGND 0.31986f
C11928 Vbias.n349 VGND 0.3159f
C11929 Vbias.n350 VGND 0.08895f
C11930 Vbias.n351 VGND 0.18787f
C11931 Vbias.t152 VGND 0.31986f
C11932 Vbias.n352 VGND 0.3159f
C11933 Vbias.n353 VGND 0.08895f
C11934 Vbias.n354 VGND 0.18787f
C11935 Vbias.t245 VGND 0.31986f
C11936 Vbias.n355 VGND 0.3159f
C11937 Vbias.n356 VGND 0.08895f
C11938 Vbias.n357 VGND 0.18787f
C11939 Vbias.t72 VGND 0.31986f
C11940 Vbias.n358 VGND 0.3159f
C11941 Vbias.n359 VGND 0.08895f
C11942 Vbias.n360 VGND 0.18787f
C11943 Vbias.t158 VGND 0.31986f
C11944 Vbias.n361 VGND 0.3159f
C11945 Vbias.n362 VGND 0.08895f
C11946 Vbias.n363 VGND 0.18787f
C11947 Vbias.t178 VGND 0.31986f
C11948 Vbias.n364 VGND 0.3159f
C11949 Vbias.n365 VGND 0.08895f
C11950 Vbias.n366 VGND 0.18787f
C11951 Vbias.t254 VGND 0.31986f
C11952 Vbias.n367 VGND 0.3159f
C11953 Vbias.n368 VGND 0.08895f
C11954 Vbias.n369 VGND 0.18787f
C11955 Vbias.t84 VGND 0.31986f
C11956 Vbias.n370 VGND 0.3159f
C11957 Vbias.n371 VGND 0.08895f
C11958 Vbias.n372 VGND 0.18787f
C11959 Vbias.t106 VGND 0.31986f
C11960 Vbias.n373 VGND 0.3159f
C11961 Vbias.n374 VGND 0.08895f
C11962 Vbias.n375 VGND 0.18787f
C11963 Vbias.t259 VGND 0.31986f
C11964 Vbias.n376 VGND 0.3159f
C11965 Vbias.n377 VGND 0.08895f
C11966 Vbias.n378 VGND 0.18787f
C11967 Vbias.t26 VGND 0.31986f
C11968 Vbias.n379 VGND 0.3159f
C11969 Vbias.n380 VGND 0.08895f
C11970 Vbias.n381 VGND 0.18787f
C11971 Vbias.n382 VGND 0.18787f
C11972 Vbias.t194 VGND 0.31986f
C11973 Vbias.n383 VGND 0.3159f
C11974 Vbias.t61 VGND 0.31986f
C11975 Vbias.n384 VGND 0.3159f
C11976 Vbias.n385 VGND 0.18787f
C11977 Vbias.n386 VGND 0.25639f
C11978 Vbias.n387 VGND 0.34679f
C11979 Vbias.n388 VGND 0.08895f
C11980 Vbias.n389 VGND 0.18787f
C11981 Vbias.n390 VGND 0.99869f
C11982 Vbias.n391 VGND 0.18787f
C11983 Vbias.n392 VGND 0.99869f
C11984 Vbias.n393 VGND 0.99869f
C11985 Vbias.n394 VGND 0.99869f
C11986 Vbias.t13 VGND 0.31986f
C11987 Vbias.n395 VGND 0.3159f
C11988 Vbias.n396 VGND 0.08895f
C11989 Vbias.n397 VGND 0.18787f
C11990 Vbias.n398 VGND 0.18787f
C11991 Vbias.n399 VGND 0.08895f
C11992 Vbias.n400 VGND 0.33621f
C11993 Vbias.n401 VGND 0.34679f
C11994 Vbias.n402 VGND 0.25639f
C11995 Vbias.n403 VGND 0.18787f
C11996 Vbias.t142 VGND 0.31986f
C11997 Vbias.n404 VGND 0.3159f
C11998 Vbias.n405 VGND 0.25639f
C11999 Vbias.n406 VGND 0.18787f
C12000 Vbias.t114 VGND 0.31986f
C12001 Vbias.n407 VGND 0.3159f
C12002 Vbias.n408 VGND 0.25639f
C12003 Vbias.n409 VGND 0.18787f
C12004 Vbias.t223 VGND 0.31986f
C12005 Vbias.n410 VGND 0.3159f
C12006 Vbias.n411 VGND 0.25639f
C12007 Vbias.n412 VGND 0.18787f
C12008 Vbias.t202 VGND 0.31986f
C12009 Vbias.n413 VGND 0.3159f
C12010 Vbias.n414 VGND 0.25639f
C12011 Vbias.n415 VGND 0.18787f
C12012 Vbias.t111 VGND 0.31986f
C12013 Vbias.n416 VGND 0.3159f
C12014 Vbias.n417 VGND 0.25639f
C12015 Vbias.n418 VGND 0.18787f
C12016 Vbias.t39 VGND 0.31986f
C12017 Vbias.n419 VGND 0.3159f
C12018 Vbias.n420 VGND 0.25639f
C12019 Vbias.n421 VGND 0.18787f
C12020 Vbias.t19 VGND 0.31986f
C12021 Vbias.n422 VGND 0.3159f
C12022 Vbias.n423 VGND 0.25639f
C12023 Vbias.n424 VGND 0.18787f
C12024 Vbias.t184 VGND 0.31986f
C12025 Vbias.n425 VGND 0.3159f
C12026 Vbias.n426 VGND 0.25639f
C12027 Vbias.n427 VGND 0.18787f
C12028 Vbias.t101 VGND 0.31986f
C12029 Vbias.n428 VGND 0.3159f
C12030 Vbias.n429 VGND 0.25639f
C12031 Vbias.n430 VGND 0.18787f
C12032 Vbias.t15 VGND 0.31986f
C12033 Vbias.n431 VGND 0.3159f
C12034 Vbias.n432 VGND 0.25639f
C12035 Vbias.n433 VGND 0.18787f
C12036 Vbias.t182 VGND 0.31986f
C12037 Vbias.n434 VGND 0.3159f
C12038 Vbias.n435 VGND 0.25639f
C12039 Vbias.n436 VGND 0.18787f
C12040 Vbias.t174 VGND 0.31986f
C12041 Vbias.n437 VGND 0.3159f
C12042 Vbias.n438 VGND 0.25639f
C12043 Vbias.n439 VGND 0.18787f
C12044 Vbias.t79 VGND 0.31986f
C12045 Vbias.n440 VGND 0.3159f
C12046 Vbias.n441 VGND 0.25639f
C12047 Vbias.n442 VGND 0.18787f
C12048 Vbias.n443 VGND 0.25378f
C12049 Vbias.n444 VGND 0.34679f
C12050 Vbias.n445 VGND 0.33621f
C12051 Vbias.n446 VGND 0.08634f
C12052 Vbias.n447 VGND 0.18787f
C12053 Vbias.n448 VGND 0.08895f
C12054 Vbias.n449 VGND 0.33621f
C12055 Vbias.n450 VGND 0.33621f
C12056 Vbias.n451 VGND 0.08895f
C12057 Vbias.n452 VGND 0.18787f
C12058 Vbias.n453 VGND 0.18787f
C12059 Vbias.n454 VGND 0.08895f
C12060 Vbias.n455 VGND 0.33621f
C12061 Vbias.n456 VGND 0.33621f
C12062 Vbias.n457 VGND 0.08895f
C12063 Vbias.n458 VGND 0.18787f
C12064 Vbias.n459 VGND 0.18787f
C12065 Vbias.n460 VGND 0.08895f
C12066 Vbias.n461 VGND 0.33621f
C12067 Vbias.n462 VGND 0.33621f
C12068 Vbias.n463 VGND 0.08895f
C12069 Vbias.n464 VGND 0.18787f
C12070 Vbias.n465 VGND 0.18787f
C12071 Vbias.n466 VGND 0.08895f
C12072 Vbias.n467 VGND 0.33621f
C12073 Vbias.n468 VGND 0.33621f
C12074 Vbias.n469 VGND 0.08895f
C12075 Vbias.n470 VGND 0.18787f
C12076 Vbias.n471 VGND 0.18787f
C12077 Vbias.n472 VGND 0.08895f
C12078 Vbias.n473 VGND 0.33621f
C12079 Vbias.n474 VGND 0.33621f
C12080 Vbias.n475 VGND 0.08895f
C12081 Vbias.n476 VGND 0.18787f
C12082 Vbias.n477 VGND 0.18787f
C12083 Vbias.n478 VGND 0.08895f
C12084 Vbias.n479 VGND 0.33621f
C12085 Vbias.n480 VGND 0.33621f
C12086 Vbias.n481 VGND 0.08895f
C12087 Vbias.n482 VGND 0.18787f
C12088 Vbias.n483 VGND 0.18787f
C12089 Vbias.n484 VGND 0.08895f
C12090 Vbias.n485 VGND 0.33621f
C12091 Vbias.n486 VGND 0.33621f
C12092 Vbias.n487 VGND 0.08895f
C12093 Vbias.n488 VGND 0.18787f
C12094 Vbias.n489 VGND 0.18787f
C12095 Vbias.n490 VGND 0.08895f
C12096 Vbias.n491 VGND 0.33621f
C12097 Vbias.n492 VGND 0.33621f
C12098 Vbias.n493 VGND 0.08895f
C12099 Vbias.n494 VGND 0.18787f
C12100 Vbias.n495 VGND 0.18787f
C12101 Vbias.n496 VGND 0.08895f
C12102 Vbias.n497 VGND 0.33621f
C12103 Vbias.n498 VGND 0.33621f
C12104 Vbias.n499 VGND 0.08895f
C12105 Vbias.n500 VGND 0.18787f
C12106 Vbias.n501 VGND 0.18787f
C12107 Vbias.n502 VGND 0.08895f
C12108 Vbias.n503 VGND 0.33621f
C12109 Vbias.n504 VGND 0.33621f
C12110 Vbias.n505 VGND 0.08895f
C12111 Vbias.n506 VGND 0.18787f
C12112 Vbias.n507 VGND 0.18787f
C12113 Vbias.n508 VGND 0.08895f
C12114 Vbias.n509 VGND 0.33621f
C12115 Vbias.n510 VGND 0.33621f
C12116 Vbias.n511 VGND 0.08895f
C12117 Vbias.n512 VGND 0.18787f
C12118 Vbias.n513 VGND 0.18787f
C12119 Vbias.n514 VGND 0.08895f
C12120 Vbias.n515 VGND 0.33621f
C12121 Vbias.n516 VGND 0.33621f
C12122 Vbias.n517 VGND 0.08895f
C12123 Vbias.n518 VGND 0.18787f
C12124 Vbias.n519 VGND 0.18787f
C12125 Vbias.n520 VGND 0.08895f
C12126 Vbias.n521 VGND 0.33621f
C12127 Vbias.n522 VGND 0.33621f
C12128 Vbias.n523 VGND 0.08895f
C12129 Vbias.n524 VGND 0.18787f
C12130 Vbias.t175 VGND 0.31986f
C12131 Vbias.n525 VGND 0.3159f
C12132 Vbias.n526 VGND 0.08895f
C12133 Vbias.n527 VGND 0.18787f
C12134 Vbias.n528 VGND 0.18787f
C12135 Vbias.n529 VGND 0.08895f
C12136 Vbias.n530 VGND 0.33621f
C12137 Vbias.n531 VGND 0.33621f
C12138 Vbias.n532 VGND 0.33621f
C12139 Vbias.n533 VGND 0.08895f
C12140 Vbias.n534 VGND 0.18787f
C12141 Vbias.n535 VGND 0.18787f
C12142 Vbias.n536 VGND 0.08895f
C12143 Vbias.n537 VGND 0.33621f
C12144 Vbias.n538 VGND 0.33621f
C12145 Vbias.n539 VGND 0.08895f
C12146 Vbias.n540 VGND 0.18787f
C12147 Vbias.t78 VGND 0.31986f
C12148 Vbias.n541 VGND 0.3159f
C12149 Vbias.n542 VGND 0.08895f
C12150 Vbias.n543 VGND 0.18787f
C12151 Vbias.t47 VGND 0.31986f
C12152 Vbias.n544 VGND 0.3159f
C12153 Vbias.n545 VGND 0.08895f
C12154 Vbias.n546 VGND 0.18787f
C12155 Vbias.t159 VGND 0.31986f
C12156 Vbias.n547 VGND 0.3159f
C12157 Vbias.n548 VGND 0.08895f
C12158 Vbias.n549 VGND 0.18787f
C12159 Vbias.t134 VGND 0.31986f
C12160 Vbias.n550 VGND 0.3159f
C12161 Vbias.n551 VGND 0.08895f
C12162 Vbias.n552 VGND 0.18787f
C12163 Vbias.t43 VGND 0.31986f
C12164 Vbias.n553 VGND 0.3159f
C12165 Vbias.n554 VGND 0.08895f
C12166 Vbias.n555 VGND 0.18787f
C12167 Vbias.t231 VGND 0.31986f
C12168 Vbias.n556 VGND 0.3159f
C12169 Vbias.n557 VGND 0.08895f
C12170 Vbias.n558 VGND 0.18787f
C12171 Vbias.t209 VGND 0.31986f
C12172 Vbias.n559 VGND 0.3159f
C12173 Vbias.n560 VGND 0.08895f
C12174 Vbias.n561 VGND 0.18787f
C12175 Vbias.t116 VGND 0.31986f
C12176 Vbias.n562 VGND 0.3159f
C12177 Vbias.n563 VGND 0.08895f
C12178 Vbias.n564 VGND 0.18787f
C12179 Vbias.t34 VGND 0.31986f
C12180 Vbias.n565 VGND 0.3159f
C12181 Vbias.n566 VGND 0.08895f
C12182 Vbias.n567 VGND 0.18787f
C12183 Vbias.t206 VGND 0.31986f
C12184 Vbias.n568 VGND 0.3159f
C12185 Vbias.n569 VGND 0.08895f
C12186 Vbias.n570 VGND 0.18787f
C12187 Vbias.t115 VGND 0.31986f
C12188 Vbias.n571 VGND 0.3159f
C12189 Vbias.n572 VGND 0.08895f
C12190 Vbias.n573 VGND 0.18787f
C12191 Vbias.t103 VGND 0.31986f
C12192 Vbias.n574 VGND 0.3159f
C12193 Vbias.n575 VGND 0.08895f
C12194 Vbias.n576 VGND 0.18787f
C12195 Vbias.t6 VGND 0.31986f
C12196 Vbias.n577 VGND 0.3159f
C12197 Vbias.n578 VGND 0.08895f
C12198 Vbias.n579 VGND 0.18787f
C12199 Vbias.n580 VGND 0.08634f
C12200 Vbias.n581 VGND 0.33621f
C12201 Vbias.n582 VGND 0.33621f
C12202 Vbias.n583 VGND 0.08634f
C12203 Vbias.n584 VGND 0.18787f
C12204 Vbias.n585 VGND 0.08895f
C12205 Vbias.n586 VGND 0.33621f
C12206 Vbias.n587 VGND 0.33621f
C12207 Vbias.n588 VGND 0.08895f
C12208 Vbias.n589 VGND 0.18787f
C12209 Vbias.n590 VGND 0.18787f
C12210 Vbias.n591 VGND 0.08895f
C12211 Vbias.n592 VGND 0.33621f
C12212 Vbias.n593 VGND 0.33621f
C12213 Vbias.n594 VGND 0.08895f
C12214 Vbias.n595 VGND 0.18787f
C12215 Vbias.n596 VGND 0.18787f
C12216 Vbias.n597 VGND 0.08895f
C12217 Vbias.n598 VGND 0.33621f
C12218 Vbias.n599 VGND 0.33621f
C12219 Vbias.n600 VGND 0.08895f
C12220 Vbias.n601 VGND 0.18787f
C12221 Vbias.n602 VGND 0.18787f
C12222 Vbias.n603 VGND 0.08895f
C12223 Vbias.n604 VGND 0.33621f
C12224 Vbias.n605 VGND 0.33621f
C12225 Vbias.n606 VGND 0.08895f
C12226 Vbias.n607 VGND 0.18787f
C12227 Vbias.n608 VGND 0.18787f
C12228 Vbias.n609 VGND 0.08895f
C12229 Vbias.n610 VGND 0.33621f
C12230 Vbias.n611 VGND 0.33621f
C12231 Vbias.n612 VGND 0.08895f
C12232 Vbias.n613 VGND 0.18787f
C12233 Vbias.n614 VGND 0.18787f
C12234 Vbias.n615 VGND 0.08895f
C12235 Vbias.n616 VGND 0.33621f
C12236 Vbias.n617 VGND 0.33621f
C12237 Vbias.n618 VGND 0.08895f
C12238 Vbias.n619 VGND 0.18787f
C12239 Vbias.n620 VGND 0.18787f
C12240 Vbias.n621 VGND 0.08895f
C12241 Vbias.n622 VGND 0.33621f
C12242 Vbias.n623 VGND 0.33621f
C12243 Vbias.n624 VGND 0.08895f
C12244 Vbias.n625 VGND 0.18787f
C12245 Vbias.n626 VGND 0.18787f
C12246 Vbias.n627 VGND 0.08895f
C12247 Vbias.n628 VGND 0.33621f
C12248 Vbias.n629 VGND 0.33621f
C12249 Vbias.n630 VGND 0.08895f
C12250 Vbias.n631 VGND 0.18787f
C12251 Vbias.n632 VGND 0.18787f
C12252 Vbias.n633 VGND 0.08895f
C12253 Vbias.n634 VGND 0.33621f
C12254 Vbias.n635 VGND 0.33621f
C12255 Vbias.n636 VGND 0.08895f
C12256 Vbias.n637 VGND 0.18787f
C12257 Vbias.n638 VGND 0.18787f
C12258 Vbias.n639 VGND 0.08895f
C12259 Vbias.n640 VGND 0.33621f
C12260 Vbias.n641 VGND 0.33621f
C12261 Vbias.n642 VGND 0.08895f
C12262 Vbias.n643 VGND 0.18787f
C12263 Vbias.n644 VGND 0.18787f
C12264 Vbias.n645 VGND 0.08895f
C12265 Vbias.n646 VGND 0.33621f
C12266 Vbias.n647 VGND 0.33621f
C12267 Vbias.n648 VGND 0.08895f
C12268 Vbias.n649 VGND 0.18787f
C12269 Vbias.n650 VGND 0.18787f
C12270 Vbias.n651 VGND 0.08895f
C12271 Vbias.n652 VGND 0.33621f
C12272 Vbias.n653 VGND 0.33621f
C12273 Vbias.n654 VGND 0.08895f
C12274 Vbias.n655 VGND 0.18787f
C12275 Vbias.n656 VGND 0.18787f
C12276 Vbias.n657 VGND 0.08895f
C12277 Vbias.n658 VGND 0.33621f
C12278 Vbias.n659 VGND 0.33621f
C12279 Vbias.n660 VGND 0.08895f
C12280 Vbias.n661 VGND 0.18787f
C12281 Vbias.t89 VGND 0.31986f
C12282 Vbias.n662 VGND 0.3159f
C12283 Vbias.n663 VGND 0.08895f
C12284 Vbias.n664 VGND 0.18787f
C12285 Vbias.t250 VGND 0.31986f
C12286 Vbias.n665 VGND 0.3159f
C12287 Vbias.n666 VGND 0.08895f
C12288 Vbias.n667 VGND 0.18787f
C12289 Vbias.n668 VGND 0.99869f
C12290 Vbias.n669 VGND 0.99869f
C12291 Vbias.n670 VGND 0.99869f
C12292 Vbias.t165 VGND 0.31986f
C12293 Vbias.n671 VGND 0.3159f
C12294 Vbias.n672 VGND 0.08895f
C12295 Vbias.n673 VGND 0.18787f
C12296 Vbias.t73 VGND 0.31986f
C12297 Vbias.n674 VGND 0.3159f
C12298 Vbias.n675 VGND 0.08895f
C12299 Vbias.n676 VGND 0.18787f
C12300 Vbias.n677 VGND 0.99869f
C12301 Vbias.t255 VGND 0.31986f
C12302 Vbias.n678 VGND 0.3159f
C12303 Vbias.n679 VGND 0.33621f
C12304 Vbias.n680 VGND 0.08895f
C12305 Vbias.n681 VGND 0.18787f
C12306 Vbias.n682 VGND 0.99869f
C12307 Vbias.t176 VGND 0.31986f
C12308 Vbias.n683 VGND 0.3159f
C12309 Vbias.n684 VGND 0.08895f
C12310 Vbias.n685 VGND 0.18787f
C12311 Vbias.n686 VGND 0.99869f
C12312 Vbias.n687 VGND 0.99869f
C12313 Vbias.n688 VGND 0.99869f
C12314 Vbias.n689 VGND 0.18787f
C12315 Vbias.n690 VGND 0.18787f
C12316 Vbias.n691 VGND 0.08895f
C12317 Vbias.n692 VGND 0.33621f
C12318 Vbias.n693 VGND 0.33621f
C12319 Vbias.n694 VGND 0.08895f
C12320 Vbias.n695 VGND 0.18787f
C12321 Vbias.n696 VGND 0.18787f
C12322 Vbias.n697 VGND 0.08895f
C12323 Vbias.n698 VGND 0.33621f
C12324 Vbias.n699 VGND 0.33621f
C12325 Vbias.n700 VGND 0.33621f
C12326 Vbias.n701 VGND 0.08895f
C12327 Vbias.n702 VGND 0.18787f
C12328 Vbias.t204 VGND 0.31986f
C12329 Vbias.n703 VGND 0.3159f
C12330 Vbias.n704 VGND 0.08895f
C12331 Vbias.n705 VGND 0.18787f
C12332 Vbias.n706 VGND 0.18787f
C12333 Vbias.n707 VGND 0.08895f
C12334 Vbias.n708 VGND 0.33621f
C12335 Vbias.n709 VGND 0.33621f
C12336 Vbias.n710 VGND 0.08895f
C12337 Vbias.n711 VGND 0.18787f
C12338 Vbias.n712 VGND 0.18787f
C12339 Vbias.n713 VGND 0.08895f
C12340 Vbias.n714 VGND 0.33621f
C12341 Vbias.n715 VGND 0.33621f
C12342 Vbias.n716 VGND 0.08895f
C12343 Vbias.n717 VGND 0.18787f
C12344 Vbias.n718 VGND 0.18787f
C12345 Vbias.n719 VGND 0.08895f
C12346 Vbias.n720 VGND 0.33621f
C12347 Vbias.n721 VGND 0.33621f
C12348 Vbias.n722 VGND 0.08895f
C12349 Vbias.n723 VGND 0.18787f
C12350 Vbias.n724 VGND 0.18787f
C12351 Vbias.n725 VGND 0.08895f
C12352 Vbias.n726 VGND 0.33621f
C12353 Vbias.n727 VGND 0.33621f
C12354 Vbias.n728 VGND 0.08895f
C12355 Vbias.n729 VGND 0.18787f
C12356 Vbias.n730 VGND 0.18787f
C12357 Vbias.n731 VGND 0.08895f
C12358 Vbias.n732 VGND 0.33621f
C12359 Vbias.n733 VGND 0.33621f
C12360 Vbias.n734 VGND 0.08895f
C12361 Vbias.n735 VGND 0.18787f
C12362 Vbias.n736 VGND 0.18787f
C12363 Vbias.n737 VGND 0.08895f
C12364 Vbias.n738 VGND 0.33621f
C12365 Vbias.n739 VGND 0.33621f
C12366 Vbias.n740 VGND 0.08895f
C12367 Vbias.n741 VGND 0.18787f
C12368 Vbias.n742 VGND 0.18787f
C12369 Vbias.n743 VGND 0.08895f
C12370 Vbias.n744 VGND 0.33621f
C12371 Vbias.n745 VGND 0.33621f
C12372 Vbias.n746 VGND 0.08895f
C12373 Vbias.n747 VGND 0.18787f
C12374 Vbias.n748 VGND 0.18787f
C12375 Vbias.n749 VGND 0.08895f
C12376 Vbias.n750 VGND 0.33621f
C12377 Vbias.n751 VGND 0.33621f
C12378 Vbias.n752 VGND 0.08895f
C12379 Vbias.n753 VGND 0.18787f
C12380 Vbias.n754 VGND 0.18787f
C12381 Vbias.n755 VGND 0.08895f
C12382 Vbias.n756 VGND 0.33621f
C12383 Vbias.n757 VGND 0.33621f
C12384 Vbias.n758 VGND 0.08895f
C12385 Vbias.n759 VGND 0.18787f
C12386 Vbias.n760 VGND 0.18787f
C12387 Vbias.n761 VGND 0.08895f
C12388 Vbias.n762 VGND 0.33621f
C12389 Vbias.n763 VGND 0.33621f
C12390 Vbias.n764 VGND 0.08895f
C12391 Vbias.n765 VGND 0.18787f
C12392 Vbias.n766 VGND 0.18787f
C12393 Vbias.n767 VGND 0.08895f
C12394 Vbias.n768 VGND 0.33621f
C12395 Vbias.n769 VGND 0.33621f
C12396 Vbias.n770 VGND 0.08895f
C12397 Vbias.n771 VGND 0.18787f
C12398 Vbias.n772 VGND 0.18787f
C12399 Vbias.n773 VGND 0.08895f
C12400 Vbias.n774 VGND 0.33621f
C12401 Vbias.n775 VGND 0.33621f
C12402 Vbias.n776 VGND 0.08895f
C12403 Vbias.n777 VGND 0.18787f
C12404 Vbias.n778 VGND 0.18787f
C12405 Vbias.n779 VGND 0.08895f
C12406 Vbias.n780 VGND 0.33621f
C12407 Vbias.n781 VGND 0.33621f
C12408 Vbias.n782 VGND 0.08895f
C12409 Vbias.n783 VGND 0.18787f
C12410 Vbias.n784 VGND 0.08634f
C12411 Vbias.n785 VGND 0.33621f
C12412 Vbias.n786 VGND 0.33621f
C12413 Vbias.n787 VGND 0.33621f
C12414 Vbias.n788 VGND 0.08634f
C12415 Vbias.t195 VGND 0.31986f
C12416 Vbias.n789 VGND 0.3159f
C12417 Vbias.n790 VGND 0.08895f
C12418 Vbias.n791 VGND 0.18787f
C12419 Vbias.t37 VGND 0.31986f
C12420 Vbias.n792 VGND 0.3159f
C12421 Vbias.n793 VGND 0.08895f
C12422 Vbias.n794 VGND 0.18787f
C12423 Vbias.t48 VGND 0.31986f
C12424 Vbias.n795 VGND 0.3159f
C12425 Vbias.n796 VGND 0.08895f
C12426 Vbias.n797 VGND 0.18787f
C12427 Vbias.t135 VGND 0.31986f
C12428 Vbias.n798 VGND 0.3159f
C12429 Vbias.n799 VGND 0.08895f
C12430 Vbias.n800 VGND 0.18787f
C12431 Vbias.t221 VGND 0.31986f
C12432 Vbias.n801 VGND 0.3159f
C12433 Vbias.n802 VGND 0.08895f
C12434 Vbias.n803 VGND 0.18787f
C12435 Vbias.t50 VGND 0.31986f
C12436 Vbias.n804 VGND 0.3159f
C12437 Vbias.n805 VGND 0.08895f
C12438 Vbias.n806 VGND 0.18787f
C12439 Vbias.t138 VGND 0.31986f
C12440 Vbias.n807 VGND 0.3159f
C12441 Vbias.n808 VGND 0.08895f
C12442 Vbias.n809 VGND 0.18787f
C12443 Vbias.t163 VGND 0.31986f
C12444 Vbias.n810 VGND 0.3159f
C12445 Vbias.n811 VGND 0.08895f
C12446 Vbias.n812 VGND 0.18787f
C12447 Vbias.t236 VGND 0.31986f
C12448 Vbias.n813 VGND 0.3159f
C12449 Vbias.n814 VGND 0.08895f
C12450 Vbias.n815 VGND 0.18787f
C12451 Vbias.t65 VGND 0.31986f
C12452 Vbias.n816 VGND 0.3159f
C12453 Vbias.n817 VGND 0.08895f
C12454 Vbias.n818 VGND 0.18787f
C12455 Vbias.t90 VGND 0.31986f
C12456 Vbias.n819 VGND 0.3159f
C12457 Vbias.n820 VGND 0.08895f
C12458 Vbias.n821 VGND 0.18787f
C12459 Vbias.t243 VGND 0.31986f
C12460 Vbias.n822 VGND 0.3159f
C12461 Vbias.n823 VGND 0.08895f
C12462 Vbias.n824 VGND 0.18787f
C12463 Vbias.t7 VGND 0.31986f
C12464 Vbias.n825 VGND 0.3159f
C12465 Vbias.n826 VGND 0.08895f
C12466 Vbias.n827 VGND 0.18787f
C12467 Vbias.n828 VGND 0.18787f
C12468 Vbias.n829 VGND 0.08895f
C12469 Vbias.n830 VGND 0.33621f
C12470 Vbias.n831 VGND 0.33621f
C12471 Vbias.n832 VGND 0.08895f
C12472 Vbias.n833 VGND 0.18787f
C12473 Vbias.n834 VGND 0.18787f
C12474 Vbias.n835 VGND 0.08895f
C12475 Vbias.n836 VGND 0.33621f
C12476 Vbias.n837 VGND 0.33621f
C12477 Vbias.n838 VGND 0.08895f
C12478 Vbias.n839 VGND 0.18787f
C12479 Vbias.n840 VGND 0.18787f
C12480 Vbias.n841 VGND 0.08895f
C12481 Vbias.n842 VGND 0.33621f
C12482 Vbias.n843 VGND 0.33621f
C12483 Vbias.n844 VGND 0.08895f
C12484 Vbias.n845 VGND 0.18787f
C12485 Vbias.n846 VGND 0.18787f
C12486 Vbias.n847 VGND 0.08895f
C12487 Vbias.n848 VGND 0.33621f
C12488 Vbias.n849 VGND 0.33621f
C12489 Vbias.n850 VGND 0.08895f
C12490 Vbias.n851 VGND 0.18787f
C12491 Vbias.n852 VGND 0.18787f
C12492 Vbias.n853 VGND 0.08895f
C12493 Vbias.n854 VGND 0.33621f
C12494 Vbias.n855 VGND 0.33621f
C12495 Vbias.n856 VGND 0.08895f
C12496 Vbias.n857 VGND 0.18787f
C12497 Vbias.n858 VGND 0.18787f
C12498 Vbias.n859 VGND 0.08895f
C12499 Vbias.n860 VGND 0.33621f
C12500 Vbias.n861 VGND 0.33621f
C12501 Vbias.n862 VGND 0.08895f
C12502 Vbias.n863 VGND 0.18787f
C12503 Vbias.n864 VGND 0.18787f
C12504 Vbias.n865 VGND 0.08895f
C12505 Vbias.n866 VGND 0.33621f
C12506 Vbias.n867 VGND 0.33621f
C12507 Vbias.n868 VGND 0.08895f
C12508 Vbias.n869 VGND 0.18787f
C12509 Vbias.n870 VGND 0.18787f
C12510 Vbias.n871 VGND 0.08895f
C12511 Vbias.n872 VGND 0.33621f
C12512 Vbias.n873 VGND 0.33621f
C12513 Vbias.n874 VGND 0.08895f
C12514 Vbias.n875 VGND 0.18787f
C12515 Vbias.n876 VGND 0.18787f
C12516 Vbias.n877 VGND 0.08895f
C12517 Vbias.n878 VGND 0.33621f
C12518 Vbias.n879 VGND 0.33621f
C12519 Vbias.n880 VGND 0.08895f
C12520 Vbias.n881 VGND 0.18787f
C12521 Vbias.n882 VGND 0.18787f
C12522 Vbias.n883 VGND 0.08895f
C12523 Vbias.n884 VGND 0.33621f
C12524 Vbias.n885 VGND 0.33621f
C12525 Vbias.n886 VGND 0.08895f
C12526 Vbias.n887 VGND 0.18787f
C12527 Vbias.n888 VGND 0.18787f
C12528 Vbias.n889 VGND 0.08895f
C12529 Vbias.n890 VGND 0.33621f
C12530 Vbias.n891 VGND 0.33621f
C12531 Vbias.n892 VGND 0.08895f
C12532 Vbias.n893 VGND 0.18787f
C12533 Vbias.n894 VGND 0.18787f
C12534 Vbias.n895 VGND 0.08895f
C12535 Vbias.n896 VGND 0.33621f
C12536 Vbias.n897 VGND 0.33621f
C12537 Vbias.n898 VGND 0.08895f
C12538 Vbias.n899 VGND 0.18787f
C12539 Vbias.n900 VGND 0.18787f
C12540 Vbias.n901 VGND 0.08895f
C12541 Vbias.n902 VGND 0.33621f
C12542 Vbias.n903 VGND 0.33621f
C12543 Vbias.n904 VGND 0.08895f
C12544 Vbias.n905 VGND 0.18787f
C12545 Vbias.t198 VGND 0.31986f
C12546 Vbias.n906 VGND 0.3159f
C12547 Vbias.n907 VGND 0.08634f
C12548 Vbias.n908 VGND 0.18787f
C12549 Vbias.n909 VGND 0.08895f
C12550 Vbias.n910 VGND 0.33621f
C12551 Vbias.n911 VGND 0.33621f
C12552 Vbias.n912 VGND 0.08895f
C12553 Vbias.n913 VGND 0.18787f
C12554 Vbias.n914 VGND 0.08634f
C12555 Vbias.n915 VGND 0.33621f
C12556 Vbias.n916 VGND 0.33621f
C12557 Vbias.n917 VGND 0.33344f
C12558 Vbias.n918 VGND 0.08634f
C12559 Vbias.n919 VGND 0.18787f
C12560 Vbias.n920 VGND 0.08895f
C12561 Vbias.n921 VGND 0.33344f
C12562 Vbias.n922 VGND 0.04505f
C12563 Vbias.n923 VGND 0.18787f
C12564 Vbias.n924 VGND 0.18787f
C12565 Vbias.n925 VGND 0.04505f
C12566 Vbias.n926 VGND 0.33344f
C12567 Vbias.n927 VGND 0.08895f
C12568 Vbias.n928 VGND 0.18787f
C12569 Vbias.n929 VGND 0.18787f
C12570 Vbias.n930 VGND 0.08895f
C12571 Vbias.n931 VGND 0.33344f
C12572 Vbias.n932 VGND 0.04505f
C12573 Vbias.n933 VGND 0.18787f
C12574 Vbias.n934 VGND 0.18787f
C12575 Vbias.n935 VGND 0.04505f
C12576 Vbias.n936 VGND 0.33344f
C12577 Vbias.n937 VGND 0.08895f
C12578 Vbias.n938 VGND 0.18787f
C12579 Vbias.n939 VGND 0.18787f
C12580 Vbias.n940 VGND 0.08895f
C12581 Vbias.n941 VGND 0.33344f
C12582 Vbias.n942 VGND 0.04505f
C12583 Vbias.n943 VGND 0.18787f
C12584 Vbias.n944 VGND 0.18787f
C12585 Vbias.n945 VGND 0.04505f
C12586 Vbias.n946 VGND 0.33344f
C12587 Vbias.n947 VGND 0.08895f
C12588 Vbias.n948 VGND 0.18787f
C12589 Vbias.n949 VGND 0.18787f
C12590 Vbias.n950 VGND 0.08895f
C12591 Vbias.n951 VGND 0.33344f
C12592 Vbias.n952 VGND 0.04505f
C12593 Vbias.n953 VGND 0.18787f
C12594 Vbias.n954 VGND 0.18787f
C12595 Vbias.n955 VGND 0.04505f
C12596 Vbias.n956 VGND 0.33344f
C12597 Vbias.n957 VGND 0.08895f
C12598 Vbias.n958 VGND 0.18787f
C12599 Vbias.n959 VGND 0.18787f
C12600 Vbias.n960 VGND 0.08895f
C12601 Vbias.n961 VGND 0.33344f
C12602 Vbias.n962 VGND 0.04505f
C12603 Vbias.n963 VGND 0.18787f
C12604 Vbias.n964 VGND 0.18787f
C12605 Vbias.n965 VGND 0.04505f
C12606 Vbias.n966 VGND 0.33344f
C12607 Vbias.n967 VGND 0.08895f
C12608 Vbias.n968 VGND 0.18787f
C12609 Vbias.n969 VGND 0.18787f
C12610 Vbias.n970 VGND 0.08895f
C12611 Vbias.n971 VGND 0.33344f
C12612 Vbias.n972 VGND 0.04505f
C12613 Vbias.n973 VGND 0.18787f
C12614 Vbias.n974 VGND 0.18787f
C12615 Vbias.n975 VGND 0.04505f
C12616 Vbias.n976 VGND 0.33344f
C12617 Vbias.n977 VGND 0.08895f
C12618 Vbias.n978 VGND 0.18787f
C12619 Vbias.n979 VGND 0.18787f
C12620 Vbias.n980 VGND 0.08895f
C12621 Vbias.n981 VGND 0.33344f
C12622 Vbias.n982 VGND 0.04505f
C12623 Vbias.n983 VGND 0.18787f
C12624 Vbias.n984 VGND 0.18787f
C12625 Vbias.n985 VGND 0.04505f
C12626 Vbias.n986 VGND 0.33344f
C12627 Vbias.n987 VGND 0.33621f
C12628 Vbias.n988 VGND 0.08895f
C12629 Vbias.n989 VGND 0.18787f
C12630 Vbias.n990 VGND 0.18787f
C12631 Vbias.n991 VGND 0.08895f
C12632 Vbias.n992 VGND 0.33621f
C12633 Vbias.n993 VGND 0.33344f
C12634 Vbias.n994 VGND 0.04505f
C12635 Vbias.n995 VGND 0.18787f
C12636 Vbias.n996 VGND 0.91809f
C12637 Vbias.n997 VGND 2.07913f
C12638 XThC.Tn[2].t8 VGND 0.0117f
C12639 XThC.Tn[2].t10 VGND 0.0117f
C12640 XThC.Tn[2].n0 VGND 0.04439f
C12641 XThC.Tn[2].t11 VGND 0.0117f
C12642 XThC.Tn[2].t9 VGND 0.0117f
C12643 XThC.Tn[2].n1 VGND 0.02664f
C12644 XThC.Tn[2].n2 VGND 0.12687f
C12645 XThC.Tn[2].t5 VGND 0.0117f
C12646 XThC.Tn[2].t4 VGND 0.0117f
C12647 XThC.Tn[2].n3 VGND 0.02664f
C12648 XThC.Tn[2].n4 VGND 0.07843f
C12649 XThC.Tn[2].t7 VGND 0.0117f
C12650 XThC.Tn[2].t6 VGND 0.0117f
C12651 XThC.Tn[2].n5 VGND 0.02664f
C12652 XThC.Tn[2].n6 VGND 0.08852f
C12653 XThC.Tn[2].t20 VGND 0.01427f
C12654 XThC.Tn[2].t18 VGND 0.01558f
C12655 XThC.Tn[2].n7 VGND 0.03478f
C12656 XThC.Tn[2].n8 VGND 0.02383f
C12657 XThC.Tn[2].n9 VGND 0.07822f
C12658 XThC.Tn[2].t38 VGND 0.01427f
C12659 XThC.Tn[2].t35 VGND 0.01558f
C12660 XThC.Tn[2].n10 VGND 0.03478f
C12661 XThC.Tn[2].n11 VGND 0.02383f
C12662 XThC.Tn[2].n12 VGND 0.07844f
C12663 XThC.Tn[2].n13 VGND 0.12927f
C12664 XThC.Tn[2].t43 VGND 0.01427f
C12665 XThC.Tn[2].t37 VGND 0.01558f
C12666 XThC.Tn[2].n14 VGND 0.03478f
C12667 XThC.Tn[2].n15 VGND 0.02383f
C12668 XThC.Tn[2].n16 VGND 0.07844f
C12669 XThC.Tn[2].n17 VGND 0.12927f
C12670 XThC.Tn[2].t12 VGND 0.01427f
C12671 XThC.Tn[2].t39 VGND 0.01558f
C12672 XThC.Tn[2].n18 VGND 0.03478f
C12673 XThC.Tn[2].n19 VGND 0.02383f
C12674 XThC.Tn[2].n20 VGND 0.07844f
C12675 XThC.Tn[2].n21 VGND 0.12927f
C12676 XThC.Tn[2].t31 VGND 0.01427f
C12677 XThC.Tn[2].t28 VGND 0.01558f
C12678 XThC.Tn[2].n22 VGND 0.03478f
C12679 XThC.Tn[2].n23 VGND 0.02383f
C12680 XThC.Tn[2].n24 VGND 0.07844f
C12681 XThC.Tn[2].n25 VGND 0.12927f
C12682 XThC.Tn[2].t32 VGND 0.01427f
C12683 XThC.Tn[2].t29 VGND 0.01558f
C12684 XThC.Tn[2].n26 VGND 0.03478f
C12685 XThC.Tn[2].n27 VGND 0.02383f
C12686 XThC.Tn[2].n28 VGND 0.07844f
C12687 XThC.Tn[2].n29 VGND 0.12927f
C12688 XThC.Tn[2].t16 VGND 0.01427f
C12689 XThC.Tn[2].t42 VGND 0.01558f
C12690 XThC.Tn[2].n30 VGND 0.03478f
C12691 XThC.Tn[2].n31 VGND 0.02383f
C12692 XThC.Tn[2].n32 VGND 0.07844f
C12693 XThC.Tn[2].n33 VGND 0.12927f
C12694 XThC.Tn[2].t23 VGND 0.01427f
C12695 XThC.Tn[2].t19 VGND 0.01558f
C12696 XThC.Tn[2].n34 VGND 0.03478f
C12697 XThC.Tn[2].n35 VGND 0.02383f
C12698 XThC.Tn[2].n36 VGND 0.07844f
C12699 XThC.Tn[2].n37 VGND 0.12927f
C12700 XThC.Tn[2].t25 VGND 0.01427f
C12701 XThC.Tn[2].t21 VGND 0.01558f
C12702 XThC.Tn[2].n38 VGND 0.03478f
C12703 XThC.Tn[2].n39 VGND 0.02383f
C12704 XThC.Tn[2].n40 VGND 0.07844f
C12705 XThC.Tn[2].n41 VGND 0.12927f
C12706 XThC.Tn[2].t13 VGND 0.01427f
C12707 XThC.Tn[2].t40 VGND 0.01558f
C12708 XThC.Tn[2].n42 VGND 0.03478f
C12709 XThC.Tn[2].n43 VGND 0.02383f
C12710 XThC.Tn[2].n44 VGND 0.07844f
C12711 XThC.Tn[2].n45 VGND 0.12927f
C12712 XThC.Tn[2].t15 VGND 0.01427f
C12713 XThC.Tn[2].t41 VGND 0.01558f
C12714 XThC.Tn[2].n46 VGND 0.03478f
C12715 XThC.Tn[2].n47 VGND 0.02383f
C12716 XThC.Tn[2].n48 VGND 0.07844f
C12717 XThC.Tn[2].n49 VGND 0.12927f
C12718 XThC.Tn[2].t26 VGND 0.01427f
C12719 XThC.Tn[2].t22 VGND 0.01558f
C12720 XThC.Tn[2].n50 VGND 0.03478f
C12721 XThC.Tn[2].n51 VGND 0.02383f
C12722 XThC.Tn[2].n52 VGND 0.07844f
C12723 XThC.Tn[2].n53 VGND 0.12927f
C12724 XThC.Tn[2].t34 VGND 0.01427f
C12725 XThC.Tn[2].t30 VGND 0.01558f
C12726 XThC.Tn[2].n54 VGND 0.03478f
C12727 XThC.Tn[2].n55 VGND 0.02383f
C12728 XThC.Tn[2].n56 VGND 0.07844f
C12729 XThC.Tn[2].n57 VGND 0.12927f
C12730 XThC.Tn[2].t36 VGND 0.01427f
C12731 XThC.Tn[2].t33 VGND 0.01558f
C12732 XThC.Tn[2].n58 VGND 0.03478f
C12733 XThC.Tn[2].n59 VGND 0.02383f
C12734 XThC.Tn[2].n60 VGND 0.07844f
C12735 XThC.Tn[2].n61 VGND 0.12927f
C12736 XThC.Tn[2].t17 VGND 0.01427f
C12737 XThC.Tn[2].t14 VGND 0.01558f
C12738 XThC.Tn[2].n62 VGND 0.03478f
C12739 XThC.Tn[2].n63 VGND 0.02383f
C12740 XThC.Tn[2].n64 VGND 0.07844f
C12741 XThC.Tn[2].n65 VGND 0.12927f
C12742 XThC.Tn[2].t27 VGND 0.01427f
C12743 XThC.Tn[2].t24 VGND 0.01558f
C12744 XThC.Tn[2].n66 VGND 0.03478f
C12745 XThC.Tn[2].n67 VGND 0.02383f
C12746 XThC.Tn[2].n68 VGND 0.07844f
C12747 XThC.Tn[2].n69 VGND 0.12927f
C12748 XThC.Tn[2].n70 VGND 0.50031f
C12749 XThC.Tn[2].n71 VGND 0.1061f
C12750 XThC.Tn[2].t1 VGND 0.018f
C12751 XThC.Tn[2].t0 VGND 0.018f
C12752 XThC.Tn[2].n72 VGND 0.04251f
C12753 XThC.Tn[2].t3 VGND 0.018f
C12754 XThC.Tn[2].t2 VGND 0.018f
C12755 XThC.Tn[2].n73 VGND 0.03633f
C12756 XThC.Tn[2].n74 VGND 0.119f
C12757 XThC.Tn[2].n75 VGND 0.03766f
C12758 XThC.Tn[4].t5 VGND 0.01821f
C12759 XThC.Tn[4].t4 VGND 0.01821f
C12760 XThC.Tn[4].n0 VGND 0.03675f
C12761 XThC.Tn[4].t7 VGND 0.01821f
C12762 XThC.Tn[4].t6 VGND 0.01821f
C12763 XThC.Tn[4].n1 VGND 0.043f
C12764 XThC.Tn[4].n2 VGND 0.12038f
C12765 XThC.Tn[4].t9 VGND 0.01183f
C12766 XThC.Tn[4].t8 VGND 0.01183f
C12767 XThC.Tn[4].n3 VGND 0.02695f
C12768 XThC.Tn[4].t11 VGND 0.01183f
C12769 XThC.Tn[4].t10 VGND 0.01183f
C12770 XThC.Tn[4].n4 VGND 0.02695f
C12771 XThC.Tn[4].t2 VGND 0.01183f
C12772 XThC.Tn[4].t1 VGND 0.01183f
C12773 XThC.Tn[4].n5 VGND 0.02695f
C12774 XThC.Tn[4].t0 VGND 0.01183f
C12775 XThC.Tn[4].t3 VGND 0.01183f
C12776 XThC.Tn[4].n6 VGND 0.0449f
C12777 XThC.Tn[4].n7 VGND 0.12834f
C12778 XThC.Tn[4].n8 VGND 0.07934f
C12779 XThC.Tn[4].n9 VGND 0.08954f
C12780 XThC.Tn[4].t28 VGND 0.01443f
C12781 XThC.Tn[4].t26 VGND 0.01576f
C12782 XThC.Tn[4].n10 VGND 0.03519f
C12783 XThC.Tn[4].n11 VGND 0.02411f
C12784 XThC.Tn[4].n12 VGND 0.07913f
C12785 XThC.Tn[4].t14 VGND 0.01443f
C12786 XThC.Tn[4].t43 VGND 0.01576f
C12787 XThC.Tn[4].n13 VGND 0.03519f
C12788 XThC.Tn[4].n14 VGND 0.02411f
C12789 XThC.Tn[4].n15 VGND 0.07935f
C12790 XThC.Tn[4].n16 VGND 0.13077f
C12791 XThC.Tn[4].t19 VGND 0.01443f
C12792 XThC.Tn[4].t13 VGND 0.01576f
C12793 XThC.Tn[4].n17 VGND 0.03519f
C12794 XThC.Tn[4].n18 VGND 0.02411f
C12795 XThC.Tn[4].n19 VGND 0.07935f
C12796 XThC.Tn[4].n20 VGND 0.13077f
C12797 XThC.Tn[4].t20 VGND 0.01443f
C12798 XThC.Tn[4].t15 VGND 0.01576f
C12799 XThC.Tn[4].n21 VGND 0.03519f
C12800 XThC.Tn[4].n22 VGND 0.02411f
C12801 XThC.Tn[4].n23 VGND 0.07935f
C12802 XThC.Tn[4].n24 VGND 0.13077f
C12803 XThC.Tn[4].t39 VGND 0.01443f
C12804 XThC.Tn[4].t36 VGND 0.01576f
C12805 XThC.Tn[4].n25 VGND 0.03519f
C12806 XThC.Tn[4].n26 VGND 0.02411f
C12807 XThC.Tn[4].n27 VGND 0.07935f
C12808 XThC.Tn[4].n28 VGND 0.13077f
C12809 XThC.Tn[4].t40 VGND 0.01443f
C12810 XThC.Tn[4].t37 VGND 0.01576f
C12811 XThC.Tn[4].n29 VGND 0.03519f
C12812 XThC.Tn[4].n30 VGND 0.02411f
C12813 XThC.Tn[4].n31 VGND 0.07935f
C12814 XThC.Tn[4].n32 VGND 0.13077f
C12815 XThC.Tn[4].t24 VGND 0.01443f
C12816 XThC.Tn[4].t18 VGND 0.01576f
C12817 XThC.Tn[4].n33 VGND 0.03519f
C12818 XThC.Tn[4].n34 VGND 0.02411f
C12819 XThC.Tn[4].n35 VGND 0.07935f
C12820 XThC.Tn[4].n36 VGND 0.13077f
C12821 XThC.Tn[4].t31 VGND 0.01443f
C12822 XThC.Tn[4].t27 VGND 0.01576f
C12823 XThC.Tn[4].n37 VGND 0.03519f
C12824 XThC.Tn[4].n38 VGND 0.02411f
C12825 XThC.Tn[4].n39 VGND 0.07935f
C12826 XThC.Tn[4].n40 VGND 0.13077f
C12827 XThC.Tn[4].t33 VGND 0.01443f
C12828 XThC.Tn[4].t29 VGND 0.01576f
C12829 XThC.Tn[4].n41 VGND 0.03519f
C12830 XThC.Tn[4].n42 VGND 0.02411f
C12831 XThC.Tn[4].n43 VGND 0.07935f
C12832 XThC.Tn[4].n44 VGND 0.13077f
C12833 XThC.Tn[4].t21 VGND 0.01443f
C12834 XThC.Tn[4].t16 VGND 0.01576f
C12835 XThC.Tn[4].n45 VGND 0.03519f
C12836 XThC.Tn[4].n46 VGND 0.02411f
C12837 XThC.Tn[4].n47 VGND 0.07935f
C12838 XThC.Tn[4].n48 VGND 0.13077f
C12839 XThC.Tn[4].t23 VGND 0.01443f
C12840 XThC.Tn[4].t17 VGND 0.01576f
C12841 XThC.Tn[4].n49 VGND 0.03519f
C12842 XThC.Tn[4].n50 VGND 0.02411f
C12843 XThC.Tn[4].n51 VGND 0.07935f
C12844 XThC.Tn[4].n52 VGND 0.13077f
C12845 XThC.Tn[4].t34 VGND 0.01443f
C12846 XThC.Tn[4].t30 VGND 0.01576f
C12847 XThC.Tn[4].n53 VGND 0.03519f
C12848 XThC.Tn[4].n54 VGND 0.02411f
C12849 XThC.Tn[4].n55 VGND 0.07935f
C12850 XThC.Tn[4].n56 VGND 0.13077f
C12851 XThC.Tn[4].t42 VGND 0.01443f
C12852 XThC.Tn[4].t38 VGND 0.01576f
C12853 XThC.Tn[4].n57 VGND 0.03519f
C12854 XThC.Tn[4].n58 VGND 0.02411f
C12855 XThC.Tn[4].n59 VGND 0.07935f
C12856 XThC.Tn[4].n60 VGND 0.13077f
C12857 XThC.Tn[4].t12 VGND 0.01443f
C12858 XThC.Tn[4].t41 VGND 0.01576f
C12859 XThC.Tn[4].n61 VGND 0.03519f
C12860 XThC.Tn[4].n62 VGND 0.02411f
C12861 XThC.Tn[4].n63 VGND 0.07935f
C12862 XThC.Tn[4].n64 VGND 0.13077f
C12863 XThC.Tn[4].t25 VGND 0.01443f
C12864 XThC.Tn[4].t22 VGND 0.01576f
C12865 XThC.Tn[4].n65 VGND 0.03519f
C12866 XThC.Tn[4].n66 VGND 0.02411f
C12867 XThC.Tn[4].n67 VGND 0.07935f
C12868 XThC.Tn[4].n68 VGND 0.13077f
C12869 XThC.Tn[4].t35 VGND 0.01443f
C12870 XThC.Tn[4].t32 VGND 0.01576f
C12871 XThC.Tn[4].n69 VGND 0.03519f
C12872 XThC.Tn[4].n70 VGND 0.02411f
C12873 XThC.Tn[4].n71 VGND 0.07935f
C12874 XThC.Tn[4].n72 VGND 0.13077f
C12875 XThC.Tn[4].n73 VGND 0.16028f
C12876 XThC.Tn[4].n74 VGND 0.0381f
C12877 XThR.Tn[5].t6 VGND 0.02327f
C12878 XThR.Tn[5].t7 VGND 0.02327f
C12879 XThR.Tn[5].n0 VGND 0.04698f
C12880 XThR.Tn[5].t5 VGND 0.02327f
C12881 XThR.Tn[5].t4 VGND 0.02327f
C12882 XThR.Tn[5].n1 VGND 0.05497f
C12883 XThR.Tn[5].n2 VGND 0.15388f
C12884 XThR.Tn[5].t11 VGND 0.01513f
C12885 XThR.Tn[5].t8 VGND 0.01513f
C12886 XThR.Tn[5].n3 VGND 0.03445f
C12887 XThR.Tn[5].t10 VGND 0.01513f
C12888 XThR.Tn[5].t9 VGND 0.01513f
C12889 XThR.Tn[5].n4 VGND 0.03445f
C12890 XThR.Tn[5].t0 VGND 0.01513f
C12891 XThR.Tn[5].t1 VGND 0.01513f
C12892 XThR.Tn[5].n5 VGND 0.0574f
C12893 XThR.Tn[5].t3 VGND 0.01513f
C12894 XThR.Tn[5].t2 VGND 0.01513f
C12895 XThR.Tn[5].n6 VGND 0.03445f
C12896 XThR.Tn[5].n7 VGND 0.16407f
C12897 XThR.Tn[5].n8 VGND 0.10142f
C12898 XThR.Tn[5].n9 VGND 0.11446f
C12899 XThR.Tn[5].t17 VGND 0.01819f
C12900 XThR.Tn[5].t72 VGND 0.01992f
C12901 XThR.Tn[5].n10 VGND 0.04864f
C12902 XThR.Tn[5].n11 VGND 0.09344f
C12903 XThR.Tn[5].t39 VGND 0.01819f
C12904 XThR.Tn[5].t26 VGND 0.01992f
C12905 XThR.Tn[5].n12 VGND 0.04864f
C12906 XThR.Tn[5].t13 VGND 0.01813f
C12907 XThR.Tn[5].t23 VGND 0.01985f
C12908 XThR.Tn[5].n13 VGND 0.05061f
C12909 XThR.Tn[5].n14 VGND 0.03555f
C12910 XThR.Tn[5].n15 VGND 0.0065f
C12911 XThR.Tn[5].n16 VGND 0.11409f
C12912 XThR.Tn[5].t73 VGND 0.01819f
C12913 XThR.Tn[5].t66 VGND 0.01992f
C12914 XThR.Tn[5].n17 VGND 0.04864f
C12915 XThR.Tn[5].t48 VGND 0.01813f
C12916 XThR.Tn[5].t61 VGND 0.01985f
C12917 XThR.Tn[5].n18 VGND 0.05061f
C12918 XThR.Tn[5].n19 VGND 0.03555f
C12919 XThR.Tn[5].n20 VGND 0.0065f
C12920 XThR.Tn[5].n21 VGND 0.11409f
C12921 XThR.Tn[5].t28 VGND 0.01819f
C12922 XThR.Tn[5].t21 VGND 0.01992f
C12923 XThR.Tn[5].n22 VGND 0.04864f
C12924 XThR.Tn[5].t65 VGND 0.01813f
C12925 XThR.Tn[5].t18 VGND 0.01985f
C12926 XThR.Tn[5].n23 VGND 0.05061f
C12927 XThR.Tn[5].n24 VGND 0.03555f
C12928 XThR.Tn[5].n25 VGND 0.0065f
C12929 XThR.Tn[5].n26 VGND 0.11409f
C12930 XThR.Tn[5].t55 VGND 0.01819f
C12931 XThR.Tn[5].t51 VGND 0.01992f
C12932 XThR.Tn[5].n27 VGND 0.04864f
C12933 XThR.Tn[5].t33 VGND 0.01813f
C12934 XThR.Tn[5].t46 VGND 0.01985f
C12935 XThR.Tn[5].n28 VGND 0.05061f
C12936 XThR.Tn[5].n29 VGND 0.03555f
C12937 XThR.Tn[5].n30 VGND 0.0065f
C12938 XThR.Tn[5].n31 VGND 0.11409f
C12939 XThR.Tn[5].t30 VGND 0.01819f
C12940 XThR.Tn[5].t22 VGND 0.01992f
C12941 XThR.Tn[5].n32 VGND 0.04864f
C12942 XThR.Tn[5].t67 VGND 0.01813f
C12943 XThR.Tn[5].t19 VGND 0.01985f
C12944 XThR.Tn[5].n33 VGND 0.05061f
C12945 XThR.Tn[5].n34 VGND 0.03555f
C12946 XThR.Tn[5].n35 VGND 0.0065f
C12947 XThR.Tn[5].n36 VGND 0.11409f
C12948 XThR.Tn[5].t69 VGND 0.01819f
C12949 XThR.Tn[5].t40 VGND 0.01992f
C12950 XThR.Tn[5].n37 VGND 0.04864f
C12951 XThR.Tn[5].t43 VGND 0.01813f
C12952 XThR.Tn[5].t37 VGND 0.01985f
C12953 XThR.Tn[5].n38 VGND 0.05061f
C12954 XThR.Tn[5].n39 VGND 0.03555f
C12955 XThR.Tn[5].n40 VGND 0.0065f
C12956 XThR.Tn[5].n41 VGND 0.11409f
C12957 XThR.Tn[5].t38 VGND 0.01819f
C12958 XThR.Tn[5].t32 VGND 0.01992f
C12959 XThR.Tn[5].n42 VGND 0.04864f
C12960 XThR.Tn[5].t14 VGND 0.01813f
C12961 XThR.Tn[5].t29 VGND 0.01985f
C12962 XThR.Tn[5].n43 VGND 0.05061f
C12963 XThR.Tn[5].n44 VGND 0.03555f
C12964 XThR.Tn[5].n45 VGND 0.0065f
C12965 XThR.Tn[5].n46 VGND 0.11409f
C12966 XThR.Tn[5].t42 VGND 0.01819f
C12967 XThR.Tn[5].t49 VGND 0.01992f
C12968 XThR.Tn[5].n47 VGND 0.04864f
C12969 XThR.Tn[5].t16 VGND 0.01813f
C12970 XThR.Tn[5].t45 VGND 0.01985f
C12971 XThR.Tn[5].n48 VGND 0.05061f
C12972 XThR.Tn[5].n49 VGND 0.03555f
C12973 XThR.Tn[5].n50 VGND 0.0065f
C12974 XThR.Tn[5].n51 VGND 0.11409f
C12975 XThR.Tn[5].t58 VGND 0.01819f
C12976 XThR.Tn[5].t68 VGND 0.01992f
C12977 XThR.Tn[5].n52 VGND 0.04864f
C12978 XThR.Tn[5].t36 VGND 0.01813f
C12979 XThR.Tn[5].t63 VGND 0.01985f
C12980 XThR.Tn[5].n53 VGND 0.05061f
C12981 XThR.Tn[5].n54 VGND 0.03555f
C12982 XThR.Tn[5].n55 VGND 0.0065f
C12983 XThR.Tn[5].n56 VGND 0.11409f
C12984 XThR.Tn[5].t53 VGND 0.01819f
C12985 XThR.Tn[5].t24 VGND 0.01992f
C12986 XThR.Tn[5].n57 VGND 0.04864f
C12987 XThR.Tn[5].t25 VGND 0.01813f
C12988 XThR.Tn[5].t20 VGND 0.01985f
C12989 XThR.Tn[5].n58 VGND 0.05061f
C12990 XThR.Tn[5].n59 VGND 0.03555f
C12991 XThR.Tn[5].n60 VGND 0.0065f
C12992 XThR.Tn[5].n61 VGND 0.11409f
C12993 XThR.Tn[5].t71 VGND 0.01819f
C12994 XThR.Tn[5].t60 VGND 0.01992f
C12995 XThR.Tn[5].n62 VGND 0.04864f
C12996 XThR.Tn[5].t44 VGND 0.01813f
C12997 XThR.Tn[5].t57 VGND 0.01985f
C12998 XThR.Tn[5].n63 VGND 0.05061f
C12999 XThR.Tn[5].n64 VGND 0.03555f
C13000 XThR.Tn[5].n65 VGND 0.0065f
C13001 XThR.Tn[5].n66 VGND 0.11409f
C13002 XThR.Tn[5].t41 VGND 0.01819f
C13003 XThR.Tn[5].t35 VGND 0.01992f
C13004 XThR.Tn[5].n67 VGND 0.04864f
C13005 XThR.Tn[5].t15 VGND 0.01813f
C13006 XThR.Tn[5].t31 VGND 0.01985f
C13007 XThR.Tn[5].n68 VGND 0.05061f
C13008 XThR.Tn[5].n69 VGND 0.03555f
C13009 XThR.Tn[5].n70 VGND 0.0065f
C13010 XThR.Tn[5].n71 VGND 0.11409f
C13011 XThR.Tn[5].t56 VGND 0.01819f
C13012 XThR.Tn[5].t52 VGND 0.01992f
C13013 XThR.Tn[5].n72 VGND 0.04864f
C13014 XThR.Tn[5].t34 VGND 0.01813f
C13015 XThR.Tn[5].t47 VGND 0.01985f
C13016 XThR.Tn[5].n73 VGND 0.05061f
C13017 XThR.Tn[5].n74 VGND 0.03555f
C13018 XThR.Tn[5].n75 VGND 0.0065f
C13019 XThR.Tn[5].n76 VGND 0.11409f
C13020 XThR.Tn[5].t12 VGND 0.01819f
C13021 XThR.Tn[5].t70 VGND 0.01992f
C13022 XThR.Tn[5].n77 VGND 0.04864f
C13023 XThR.Tn[5].t50 VGND 0.01813f
C13024 XThR.Tn[5].t64 VGND 0.01985f
C13025 XThR.Tn[5].n78 VGND 0.05061f
C13026 XThR.Tn[5].n79 VGND 0.03555f
C13027 XThR.Tn[5].n80 VGND 0.0065f
C13028 XThR.Tn[5].n81 VGND 0.11409f
C13029 XThR.Tn[5].t54 VGND 0.01819f
C13030 XThR.Tn[5].t62 VGND 0.01992f
C13031 XThR.Tn[5].n82 VGND 0.04864f
C13032 XThR.Tn[5].t27 VGND 0.01813f
C13033 XThR.Tn[5].t59 VGND 0.01985f
C13034 XThR.Tn[5].n83 VGND 0.05061f
C13035 XThR.Tn[5].n84 VGND 0.03555f
C13036 XThR.Tn[5].n85 VGND 0.0065f
C13037 XThR.Tn[5].n86 VGND 0.11409f
C13038 XThR.Tn[5].n87 VGND 0.10368f
C13039 XThR.Tn[5].n88 VGND 0.20081f
C13040 XThR.Tn[5].n89 VGND 0.0487f
C13041 XThR.Tn[3].t8 VGND 0.02315f
C13042 XThR.Tn[3].t9 VGND 0.02315f
C13043 XThR.Tn[3].n0 VGND 0.04673f
C13044 XThR.Tn[3].t7 VGND 0.02315f
C13045 XThR.Tn[3].t10 VGND 0.02315f
C13046 XThR.Tn[3].n1 VGND 0.05468f
C13047 XThR.Tn[3].n2 VGND 0.15307f
C13048 XThR.Tn[3].t6 VGND 0.01505f
C13049 XThR.Tn[3].t3 VGND 0.01505f
C13050 XThR.Tn[3].n3 VGND 0.03427f
C13051 XThR.Tn[3].t5 VGND 0.01505f
C13052 XThR.Tn[3].t4 VGND 0.01505f
C13053 XThR.Tn[3].n4 VGND 0.03427f
C13054 XThR.Tn[3].t11 VGND 0.01505f
C13055 XThR.Tn[3].t1 VGND 0.01505f
C13056 XThR.Tn[3].n5 VGND 0.03427f
C13057 XThR.Tn[3].t0 VGND 0.01505f
C13058 XThR.Tn[3].t2 VGND 0.01505f
C13059 XThR.Tn[3].n6 VGND 0.0571f
C13060 XThR.Tn[3].n7 VGND 0.16319f
C13061 XThR.Tn[3].n8 VGND 0.10088f
C13062 XThR.Tn[3].n9 VGND 0.11385f
C13063 XThR.Tn[3].t64 VGND 0.01809f
C13064 XThR.Tn[3].t57 VGND 0.01981f
C13065 XThR.Tn[3].n10 VGND 0.04838f
C13066 XThR.Tn[3].n11 VGND 0.09294f
C13067 XThR.Tn[3].t18 VGND 0.01809f
C13068 XThR.Tn[3].t70 VGND 0.01981f
C13069 XThR.Tn[3].n12 VGND 0.04838f
C13070 XThR.Tn[3].t24 VGND 0.01803f
C13071 XThR.Tn[3].t55 VGND 0.01975f
C13072 XThR.Tn[3].n13 VGND 0.05034f
C13073 XThR.Tn[3].n14 VGND 0.03536f
C13074 XThR.Tn[3].n15 VGND 0.00647f
C13075 XThR.Tn[3].n16 VGND 0.11349f
C13076 XThR.Tn[3].t59 VGND 0.01809f
C13077 XThR.Tn[3].t49 VGND 0.01981f
C13078 XThR.Tn[3].n17 VGND 0.04838f
C13079 XThR.Tn[3].t62 VGND 0.01803f
C13080 XThR.Tn[3].t29 VGND 0.01975f
C13081 XThR.Tn[3].n18 VGND 0.05034f
C13082 XThR.Tn[3].n19 VGND 0.03536f
C13083 XThR.Tn[3].n20 VGND 0.00647f
C13084 XThR.Tn[3].n21 VGND 0.11349f
C13085 XThR.Tn[3].t71 VGND 0.01809f
C13086 XThR.Tn[3].t67 VGND 0.01981f
C13087 XThR.Tn[3].n22 VGND 0.04838f
C13088 XThR.Tn[3].t12 VGND 0.01803f
C13089 XThR.Tn[3].t47 VGND 0.01975f
C13090 XThR.Tn[3].n23 VGND 0.05034f
C13091 XThR.Tn[3].n24 VGND 0.03536f
C13092 XThR.Tn[3].n25 VGND 0.00647f
C13093 XThR.Tn[3].n26 VGND 0.11349f
C13094 XThR.Tn[3].t39 VGND 0.01809f
C13095 XThR.Tn[3].t33 VGND 0.01981f
C13096 XThR.Tn[3].n27 VGND 0.04838f
C13097 XThR.Tn[3].t42 VGND 0.01803f
C13098 XThR.Tn[3].t13 VGND 0.01975f
C13099 XThR.Tn[3].n28 VGND 0.05034f
C13100 XThR.Tn[3].n29 VGND 0.03536f
C13101 XThR.Tn[3].n30 VGND 0.00647f
C13102 XThR.Tn[3].n31 VGND 0.11349f
C13103 XThR.Tn[3].t72 VGND 0.01809f
C13104 XThR.Tn[3].t68 VGND 0.01981f
C13105 XThR.Tn[3].n32 VGND 0.04838f
C13106 XThR.Tn[3].t16 VGND 0.01803f
C13107 XThR.Tn[3].t48 VGND 0.01975f
C13108 XThR.Tn[3].n33 VGND 0.05034f
C13109 XThR.Tn[3].n34 VGND 0.03536f
C13110 XThR.Tn[3].n35 VGND 0.00647f
C13111 XThR.Tn[3].n36 VGND 0.11349f
C13112 XThR.Tn[3].t52 VGND 0.01809f
C13113 XThR.Tn[3].t20 VGND 0.01981f
C13114 XThR.Tn[3].n37 VGND 0.04838f
C13115 XThR.Tn[3].t56 VGND 0.01803f
C13116 XThR.Tn[3].t66 VGND 0.01975f
C13117 XThR.Tn[3].n38 VGND 0.05034f
C13118 XThR.Tn[3].n39 VGND 0.03536f
C13119 XThR.Tn[3].n40 VGND 0.00647f
C13120 XThR.Tn[3].n41 VGND 0.11349f
C13121 XThR.Tn[3].t19 VGND 0.01809f
C13122 XThR.Tn[3].t14 VGND 0.01981f
C13123 XThR.Tn[3].n42 VGND 0.04838f
C13124 XThR.Tn[3].t23 VGND 0.01803f
C13125 XThR.Tn[3].t61 VGND 0.01975f
C13126 XThR.Tn[3].n43 VGND 0.05034f
C13127 XThR.Tn[3].n44 VGND 0.03536f
C13128 XThR.Tn[3].n45 VGND 0.00647f
C13129 XThR.Tn[3].n46 VGND 0.11349f
C13130 XThR.Tn[3].t22 VGND 0.01809f
C13131 XThR.Tn[3].t31 VGND 0.01981f
C13132 XThR.Tn[3].n47 VGND 0.04838f
C13133 XThR.Tn[3].t28 VGND 0.01803f
C13134 XThR.Tn[3].t73 VGND 0.01975f
C13135 XThR.Tn[3].n48 VGND 0.05034f
C13136 XThR.Tn[3].n49 VGND 0.03536f
C13137 XThR.Tn[3].n50 VGND 0.00647f
C13138 XThR.Tn[3].n51 VGND 0.11349f
C13139 XThR.Tn[3].t41 VGND 0.01809f
C13140 XThR.Tn[3].t51 VGND 0.01981f
C13141 XThR.Tn[3].n52 VGND 0.04838f
C13142 XThR.Tn[3].t45 VGND 0.01803f
C13143 XThR.Tn[3].t30 VGND 0.01975f
C13144 XThR.Tn[3].n53 VGND 0.05034f
C13145 XThR.Tn[3].n54 VGND 0.03536f
C13146 XThR.Tn[3].n55 VGND 0.00647f
C13147 XThR.Tn[3].n56 VGND 0.11349f
C13148 XThR.Tn[3].t35 VGND 0.01809f
C13149 XThR.Tn[3].t69 VGND 0.01981f
C13150 XThR.Tn[3].n57 VGND 0.04838f
C13151 XThR.Tn[3].t37 VGND 0.01803f
C13152 XThR.Tn[3].t50 VGND 0.01975f
C13153 XThR.Tn[3].n58 VGND 0.05034f
C13154 XThR.Tn[3].n59 VGND 0.03536f
C13155 XThR.Tn[3].n60 VGND 0.00647f
C13156 XThR.Tn[3].n61 VGND 0.11349f
C13157 XThR.Tn[3].t54 VGND 0.01809f
C13158 XThR.Tn[3].t44 VGND 0.01981f
C13159 XThR.Tn[3].n62 VGND 0.04838f
C13160 XThR.Tn[3].t58 VGND 0.01803f
C13161 XThR.Tn[3].t25 VGND 0.01975f
C13162 XThR.Tn[3].n63 VGND 0.05034f
C13163 XThR.Tn[3].n64 VGND 0.03536f
C13164 XThR.Tn[3].n65 VGND 0.00647f
C13165 XThR.Tn[3].n66 VGND 0.11349f
C13166 XThR.Tn[3].t21 VGND 0.01809f
C13167 XThR.Tn[3].t17 VGND 0.01981f
C13168 XThR.Tn[3].n67 VGND 0.04838f
C13169 XThR.Tn[3].t26 VGND 0.01803f
C13170 XThR.Tn[3].t63 VGND 0.01975f
C13171 XThR.Tn[3].n68 VGND 0.05034f
C13172 XThR.Tn[3].n69 VGND 0.03536f
C13173 XThR.Tn[3].n70 VGND 0.00647f
C13174 XThR.Tn[3].n71 VGND 0.11349f
C13175 XThR.Tn[3].t40 VGND 0.01809f
C13176 XThR.Tn[3].t34 VGND 0.01981f
C13177 XThR.Tn[3].n72 VGND 0.04838f
C13178 XThR.Tn[3].t43 VGND 0.01803f
C13179 XThR.Tn[3].t15 VGND 0.01975f
C13180 XThR.Tn[3].n73 VGND 0.05034f
C13181 XThR.Tn[3].n74 VGND 0.03536f
C13182 XThR.Tn[3].n75 VGND 0.00647f
C13183 XThR.Tn[3].n76 VGND 0.11349f
C13184 XThR.Tn[3].t60 VGND 0.01809f
C13185 XThR.Tn[3].t53 VGND 0.01981f
C13186 XThR.Tn[3].n77 VGND 0.04838f
C13187 XThR.Tn[3].t65 VGND 0.01803f
C13188 XThR.Tn[3].t32 VGND 0.01975f
C13189 XThR.Tn[3].n78 VGND 0.05034f
C13190 XThR.Tn[3].n79 VGND 0.03536f
C13191 XThR.Tn[3].n80 VGND 0.00647f
C13192 XThR.Tn[3].n81 VGND 0.11349f
C13193 XThR.Tn[3].t36 VGND 0.01809f
C13194 XThR.Tn[3].t46 VGND 0.01981f
C13195 XThR.Tn[3].n82 VGND 0.04838f
C13196 XThR.Tn[3].t38 VGND 0.01803f
C13197 XThR.Tn[3].t27 VGND 0.01975f
C13198 XThR.Tn[3].n83 VGND 0.05034f
C13199 XThR.Tn[3].n84 VGND 0.03536f
C13200 XThR.Tn[3].n85 VGND 0.00647f
C13201 XThR.Tn[3].n86 VGND 0.11349f
C13202 XThR.Tn[3].n87 VGND 0.10313f
C13203 XThR.Tn[3].n88 VGND 0.22842f
C13204 XThR.Tn[3].n89 VGND 0.04845f
C13205 XThC.XTB4.Y.t4 VGND 0.02956f
C13206 XThC.XTB4.Y.t13 VGND 0.05016f
C13207 XThC.XTB4.Y.n0 VGND 0.05972f
C13208 XThC.XTB4.Y.t7 VGND 0.02956f
C13209 XThC.XTB4.Y.t17 VGND 0.05016f
C13210 XThC.XTB4.Y.n1 VGND 0.03074f
C13211 XThC.XTB4.Y.t10 VGND 0.02956f
C13212 XThC.XTB4.Y.t2 VGND 0.05016f
C13213 XThC.XTB4.Y.n2 VGND 0.06603f
C13214 XThC.XTB4.Y.t14 VGND 0.02956f
C13215 XThC.XTB4.Y.t3 VGND 0.05016f
C13216 XThC.XTB4.Y.n3 VGND 0.0613f
C13217 XThC.XTB4.Y.n4 VGND 0.03729f
C13218 XThC.XTB4.Y.n5 VGND 0.06174f
C13219 XThC.XTB4.Y.n6 VGND 0.02389f
C13220 XThC.XTB4.Y.n7 VGND 0.02916f
C13221 XThC.XTB4.Y.n8 VGND 0.06603f
C13222 XThC.XTB4.Y.n9 VGND 0.0331f
C13223 XThC.XTB4.Y.n10 VGND 0.06459f
C13224 XThC.XTB4.Y.t5 VGND 0.02956f
C13225 XThC.XTB4.Y.t16 VGND 0.05016f
C13226 XThC.XTB4.Y.n11 VGND 0.06761f
C13227 XThC.XTB4.Y.t9 VGND 0.02956f
C13228 XThC.XTB4.Y.t6 VGND 0.05016f
C13229 XThC.XTB4.Y.t15 VGND 0.02956f
C13230 XThC.XTB4.Y.t12 VGND 0.05016f
C13231 XThC.XTB4.Y.t11 VGND 0.02956f
C13232 XThC.XTB4.Y.t8 VGND 0.05016f
C13233 XThC.XTB4.Y.n12 VGND 0.08416f
C13234 XThC.XTB4.Y.n13 VGND 0.08889f
C13235 XThC.XTB4.Y.n14 VGND 0.03426f
C13236 XThC.XTB4.Y.n15 VGND 0.07234f
C13237 XThC.XTB4.Y.n16 VGND 0.0331f
C13238 XThC.XTB4.Y.n17 VGND 0.02701f
C13239 XThC.XTB4.Y.n18 VGND 0.63971f
C13240 XThC.XTB4.Y.n19 VGND 1.30917f
C13241 XThC.XTB4.Y.t1 VGND 0.06491f
C13242 XThC.XTB4.Y.n20 VGND 0.11223f
C13243 XThC.XTB4.Y.t0 VGND 0.12238f
C13244 XThC.XTB4.Y.n21 VGND 0.16166f
C13245 XThC.Tn[0].t11 VGND 0.00786f
C13246 XThC.Tn[0].t8 VGND 0.00786f
C13247 XThC.Tn[0].n0 VGND 0.02982f
C13248 XThC.Tn[0].t9 VGND 0.00786f
C13249 XThC.Tn[0].t10 VGND 0.00786f
C13250 XThC.Tn[0].n1 VGND 0.01789f
C13251 XThC.Tn[0].n2 VGND 0.08522f
C13252 XThC.Tn[0].t7 VGND 0.00786f
C13253 XThC.Tn[0].t6 VGND 0.00786f
C13254 XThC.Tn[0].n3 VGND 0.01789f
C13255 XThC.Tn[0].n4 VGND 0.05268f
C13256 XThC.Tn[0].t5 VGND 0.00786f
C13257 XThC.Tn[0].t4 VGND 0.00786f
C13258 XThC.Tn[0].n5 VGND 0.01789f
C13259 XThC.Tn[0].n6 VGND 0.05945f
C13260 XThC.Tn[0].t18 VGND 0.00958f
C13261 XThC.Tn[0].t22 VGND 0.01047f
C13262 XThC.Tn[0].n7 VGND 0.02336f
C13263 XThC.Tn[0].n8 VGND 0.01601f
C13264 XThC.Tn[0].n9 VGND 0.05254f
C13265 XThC.Tn[0].t35 VGND 0.00958f
C13266 XThC.Tn[0].t41 VGND 0.01047f
C13267 XThC.Tn[0].n10 VGND 0.02336f
C13268 XThC.Tn[0].n11 VGND 0.01601f
C13269 XThC.Tn[0].n12 VGND 0.05268f
C13270 XThC.Tn[0].n13 VGND 0.08683f
C13271 XThC.Tn[0].t37 VGND 0.00958f
C13272 XThC.Tn[0].t12 VGND 0.01047f
C13273 XThC.Tn[0].n14 VGND 0.02336f
C13274 XThC.Tn[0].n15 VGND 0.01601f
C13275 XThC.Tn[0].n16 VGND 0.05268f
C13276 XThC.Tn[0].n17 VGND 0.08683f
C13277 XThC.Tn[0].t39 VGND 0.00958f
C13278 XThC.Tn[0].t13 VGND 0.01047f
C13279 XThC.Tn[0].n18 VGND 0.02336f
C13280 XThC.Tn[0].n19 VGND 0.01601f
C13281 XThC.Tn[0].n20 VGND 0.05268f
C13282 XThC.Tn[0].n21 VGND 0.08683f
C13283 XThC.Tn[0].t28 VGND 0.00958f
C13284 XThC.Tn[0].t32 VGND 0.01047f
C13285 XThC.Tn[0].n22 VGND 0.02336f
C13286 XThC.Tn[0].n23 VGND 0.01601f
C13287 XThC.Tn[0].n24 VGND 0.05268f
C13288 XThC.Tn[0].n25 VGND 0.08683f
C13289 XThC.Tn[0].t30 VGND 0.00958f
C13290 XThC.Tn[0].t34 VGND 0.01047f
C13291 XThC.Tn[0].n26 VGND 0.02336f
C13292 XThC.Tn[0].n27 VGND 0.01601f
C13293 XThC.Tn[0].n28 VGND 0.05268f
C13294 XThC.Tn[0].n29 VGND 0.08683f
C13295 XThC.Tn[0].t43 VGND 0.00958f
C13296 XThC.Tn[0].t17 VGND 0.01047f
C13297 XThC.Tn[0].n30 VGND 0.02336f
C13298 XThC.Tn[0].n31 VGND 0.01601f
C13299 XThC.Tn[0].n32 VGND 0.05268f
C13300 XThC.Tn[0].n33 VGND 0.08683f
C13301 XThC.Tn[0].t20 VGND 0.00958f
C13302 XThC.Tn[0].t25 VGND 0.01047f
C13303 XThC.Tn[0].n34 VGND 0.02336f
C13304 XThC.Tn[0].n35 VGND 0.01601f
C13305 XThC.Tn[0].n36 VGND 0.05268f
C13306 XThC.Tn[0].n37 VGND 0.08683f
C13307 XThC.Tn[0].t21 VGND 0.00958f
C13308 XThC.Tn[0].t26 VGND 0.01047f
C13309 XThC.Tn[0].n38 VGND 0.02336f
C13310 XThC.Tn[0].n39 VGND 0.01601f
C13311 XThC.Tn[0].n40 VGND 0.05268f
C13312 XThC.Tn[0].n41 VGND 0.08683f
C13313 XThC.Tn[0].t40 VGND 0.00958f
C13314 XThC.Tn[0].t15 VGND 0.01047f
C13315 XThC.Tn[0].n42 VGND 0.02336f
C13316 XThC.Tn[0].n43 VGND 0.01601f
C13317 XThC.Tn[0].n44 VGND 0.05268f
C13318 XThC.Tn[0].n45 VGND 0.08683f
C13319 XThC.Tn[0].t42 VGND 0.00958f
C13320 XThC.Tn[0].t16 VGND 0.01047f
C13321 XThC.Tn[0].n46 VGND 0.02336f
C13322 XThC.Tn[0].n47 VGND 0.01601f
C13323 XThC.Tn[0].n48 VGND 0.05268f
C13324 XThC.Tn[0].n49 VGND 0.08683f
C13325 XThC.Tn[0].t23 VGND 0.00958f
C13326 XThC.Tn[0].t27 VGND 0.01047f
C13327 XThC.Tn[0].n50 VGND 0.02336f
C13328 XThC.Tn[0].n51 VGND 0.01601f
C13329 XThC.Tn[0].n52 VGND 0.05268f
C13330 XThC.Tn[0].n53 VGND 0.08683f
C13331 XThC.Tn[0].t31 VGND 0.00958f
C13332 XThC.Tn[0].t36 VGND 0.01047f
C13333 XThC.Tn[0].n54 VGND 0.02336f
C13334 XThC.Tn[0].n55 VGND 0.01601f
C13335 XThC.Tn[0].n56 VGND 0.05268f
C13336 XThC.Tn[0].n57 VGND 0.08683f
C13337 XThC.Tn[0].t33 VGND 0.00958f
C13338 XThC.Tn[0].t38 VGND 0.01047f
C13339 XThC.Tn[0].n58 VGND 0.02336f
C13340 XThC.Tn[0].n59 VGND 0.01601f
C13341 XThC.Tn[0].n60 VGND 0.05268f
C13342 XThC.Tn[0].n61 VGND 0.08683f
C13343 XThC.Tn[0].t14 VGND 0.00958f
C13344 XThC.Tn[0].t19 VGND 0.01047f
C13345 XThC.Tn[0].n62 VGND 0.02336f
C13346 XThC.Tn[0].n63 VGND 0.01601f
C13347 XThC.Tn[0].n64 VGND 0.05268f
C13348 XThC.Tn[0].n65 VGND 0.08683f
C13349 XThC.Tn[0].t24 VGND 0.00958f
C13350 XThC.Tn[0].t29 VGND 0.01047f
C13351 XThC.Tn[0].n66 VGND 0.02336f
C13352 XThC.Tn[0].n67 VGND 0.01601f
C13353 XThC.Tn[0].n68 VGND 0.05268f
C13354 XThC.Tn[0].n69 VGND 0.08683f
C13355 XThC.Tn[0].n70 VGND 0.53669f
C13356 XThC.Tn[0].n71 VGND 0.06506f
C13357 XThC.Tn[0].t1 VGND 0.01209f
C13358 XThC.Tn[0].t0 VGND 0.01209f
C13359 XThC.Tn[0].n72 VGND 0.0244f
C13360 XThC.Tn[0].t3 VGND 0.01209f
C13361 XThC.Tn[0].t2 VGND 0.01209f
C13362 XThC.Tn[0].n73 VGND 0.02855f
C13363 XThC.Tn[0].n74 VGND 0.07993f
C13364 XThC.Tn[0].n75 VGND 0.0253f
C13365 XThC.Tn[13].t7 VGND 0.01267f
C13366 XThC.Tn[13].t5 VGND 0.01267f
C13367 XThC.Tn[13].n0 VGND 0.03161f
C13368 XThC.Tn[13].t4 VGND 0.01267f
C13369 XThC.Tn[13].t6 VGND 0.01267f
C13370 XThC.Tn[13].n1 VGND 0.02535f
C13371 XThC.Tn[13].n2 VGND 0.05845f
C13372 XThC.Tn[13].t29 VGND 0.01546f
C13373 XThC.Tn[13].t27 VGND 0.01688f
C13374 XThC.Tn[13].n3 VGND 0.03768f
C13375 XThC.Tn[13].n4 VGND 0.02582f
C13376 XThC.Tn[13].n5 VGND 0.08475f
C13377 XThC.Tn[13].t15 VGND 0.01546f
C13378 XThC.Tn[13].t12 VGND 0.01688f
C13379 XThC.Tn[13].n6 VGND 0.03768f
C13380 XThC.Tn[13].n7 VGND 0.02582f
C13381 XThC.Tn[13].n8 VGND 0.08498f
C13382 XThC.Tn[13].n9 VGND 0.14005f
C13383 XThC.Tn[13].t20 VGND 0.01546f
C13384 XThC.Tn[13].t14 VGND 0.01688f
C13385 XThC.Tn[13].n10 VGND 0.03768f
C13386 XThC.Tn[13].n11 VGND 0.02582f
C13387 XThC.Tn[13].n12 VGND 0.08498f
C13388 XThC.Tn[13].n13 VGND 0.14005f
C13389 XThC.Tn[13].t21 VGND 0.01546f
C13390 XThC.Tn[13].t16 VGND 0.01688f
C13391 XThC.Tn[13].n14 VGND 0.03768f
C13392 XThC.Tn[13].n15 VGND 0.02582f
C13393 XThC.Tn[13].n16 VGND 0.08498f
C13394 XThC.Tn[13].n17 VGND 0.14005f
C13395 XThC.Tn[13].t40 VGND 0.01546f
C13396 XThC.Tn[13].t37 VGND 0.01688f
C13397 XThC.Tn[13].n18 VGND 0.03768f
C13398 XThC.Tn[13].n19 VGND 0.02582f
C13399 XThC.Tn[13].n20 VGND 0.08498f
C13400 XThC.Tn[13].n21 VGND 0.14005f
C13401 XThC.Tn[13].t41 VGND 0.01546f
C13402 XThC.Tn[13].t38 VGND 0.01688f
C13403 XThC.Tn[13].n22 VGND 0.03768f
C13404 XThC.Tn[13].n23 VGND 0.02582f
C13405 XThC.Tn[13].n24 VGND 0.08498f
C13406 XThC.Tn[13].n25 VGND 0.14005f
C13407 XThC.Tn[13].t25 VGND 0.01546f
C13408 XThC.Tn[13].t19 VGND 0.01688f
C13409 XThC.Tn[13].n26 VGND 0.03768f
C13410 XThC.Tn[13].n27 VGND 0.02582f
C13411 XThC.Tn[13].n28 VGND 0.08498f
C13412 XThC.Tn[13].n29 VGND 0.14005f
C13413 XThC.Tn[13].t32 VGND 0.01546f
C13414 XThC.Tn[13].t28 VGND 0.01688f
C13415 XThC.Tn[13].n30 VGND 0.03768f
C13416 XThC.Tn[13].n31 VGND 0.02582f
C13417 XThC.Tn[13].n32 VGND 0.08498f
C13418 XThC.Tn[13].n33 VGND 0.14005f
C13419 XThC.Tn[13].t34 VGND 0.01546f
C13420 XThC.Tn[13].t30 VGND 0.01688f
C13421 XThC.Tn[13].n34 VGND 0.03768f
C13422 XThC.Tn[13].n35 VGND 0.02582f
C13423 XThC.Tn[13].n36 VGND 0.08498f
C13424 XThC.Tn[13].n37 VGND 0.14005f
C13425 XThC.Tn[13].t22 VGND 0.01546f
C13426 XThC.Tn[13].t17 VGND 0.01688f
C13427 XThC.Tn[13].n38 VGND 0.03768f
C13428 XThC.Tn[13].n39 VGND 0.02582f
C13429 XThC.Tn[13].n40 VGND 0.08498f
C13430 XThC.Tn[13].n41 VGND 0.14005f
C13431 XThC.Tn[13].t24 VGND 0.01546f
C13432 XThC.Tn[13].t18 VGND 0.01688f
C13433 XThC.Tn[13].n42 VGND 0.03768f
C13434 XThC.Tn[13].n43 VGND 0.02582f
C13435 XThC.Tn[13].n44 VGND 0.08498f
C13436 XThC.Tn[13].n45 VGND 0.14005f
C13437 XThC.Tn[13].t35 VGND 0.01546f
C13438 XThC.Tn[13].t31 VGND 0.01688f
C13439 XThC.Tn[13].n46 VGND 0.03768f
C13440 XThC.Tn[13].n47 VGND 0.02582f
C13441 XThC.Tn[13].n48 VGND 0.08498f
C13442 XThC.Tn[13].n49 VGND 0.14005f
C13443 XThC.Tn[13].t43 VGND 0.01546f
C13444 XThC.Tn[13].t39 VGND 0.01688f
C13445 XThC.Tn[13].n50 VGND 0.03768f
C13446 XThC.Tn[13].n51 VGND 0.02582f
C13447 XThC.Tn[13].n52 VGND 0.08498f
C13448 XThC.Tn[13].n53 VGND 0.14005f
C13449 XThC.Tn[13].t13 VGND 0.01546f
C13450 XThC.Tn[13].t42 VGND 0.01688f
C13451 XThC.Tn[13].n54 VGND 0.03768f
C13452 XThC.Tn[13].n55 VGND 0.02582f
C13453 XThC.Tn[13].n56 VGND 0.08498f
C13454 XThC.Tn[13].n57 VGND 0.14005f
C13455 XThC.Tn[13].t26 VGND 0.01546f
C13456 XThC.Tn[13].t23 VGND 0.01688f
C13457 XThC.Tn[13].n58 VGND 0.03768f
C13458 XThC.Tn[13].n59 VGND 0.02582f
C13459 XThC.Tn[13].n60 VGND 0.08498f
C13460 XThC.Tn[13].n61 VGND 0.14005f
C13461 XThC.Tn[13].t36 VGND 0.01546f
C13462 XThC.Tn[13].t33 VGND 0.01688f
C13463 XThC.Tn[13].n62 VGND 0.03768f
C13464 XThC.Tn[13].n63 VGND 0.02582f
C13465 XThC.Tn[13].n64 VGND 0.08498f
C13466 XThC.Tn[13].n65 VGND 0.14005f
C13467 XThC.Tn[13].n66 VGND 0.72631f
C13468 XThC.Tn[13].n67 VGND 0.25541f
C13469 XThC.Tn[13].t2 VGND 0.0195f
C13470 XThC.Tn[13].t1 VGND 0.0195f
C13471 XThC.Tn[13].n68 VGND 0.04213f
C13472 XThC.Tn[13].t0 VGND 0.0195f
C13473 XThC.Tn[13].t3 VGND 0.0195f
C13474 XThC.Tn[13].n69 VGND 0.06641f
C13475 XThC.Tn[13].n70 VGND 0.17588f
C13476 XThC.Tn[13].n71 VGND 0.01295f
C13477 XThC.Tn[13].t9 VGND 0.0195f
C13478 XThC.Tn[13].t8 VGND 0.0195f
C13479 XThC.Tn[13].n72 VGND 0.05921f
C13480 XThC.Tn[13].t11 VGND 0.0195f
C13481 XThC.Tn[13].t10 VGND 0.0195f
C13482 XThC.Tn[13].n73 VGND 0.04335f
C13483 XThC.Tn[13].n74 VGND 0.19292f
C13484 XThC.Tn[12].t7 VGND 0.01298f
C13485 XThC.Tn[12].t6 VGND 0.01298f
C13486 XThC.Tn[12].n0 VGND 0.03236f
C13487 XThC.Tn[12].t5 VGND 0.01298f
C13488 XThC.Tn[12].t4 VGND 0.01298f
C13489 XThC.Tn[12].n1 VGND 0.02595f
C13490 XThC.Tn[12].n2 VGND 0.06529f
C13491 XThC.Tn[12].t37 VGND 0.01582f
C13492 XThC.Tn[12].t35 VGND 0.01728f
C13493 XThC.Tn[12].n3 VGND 0.03858f
C13494 XThC.Tn[12].n4 VGND 0.02643f
C13495 XThC.Tn[12].n5 VGND 0.08676f
C13496 XThC.Tn[12].t23 VGND 0.01582f
C13497 XThC.Tn[12].t20 VGND 0.01728f
C13498 XThC.Tn[12].n6 VGND 0.03858f
C13499 XThC.Tn[12].n7 VGND 0.02643f
C13500 XThC.Tn[12].n8 VGND 0.087f
C13501 XThC.Tn[12].n9 VGND 0.14339f
C13502 XThC.Tn[12].t28 VGND 0.01582f
C13503 XThC.Tn[12].t22 VGND 0.01728f
C13504 XThC.Tn[12].n10 VGND 0.03858f
C13505 XThC.Tn[12].n11 VGND 0.02643f
C13506 XThC.Tn[12].n12 VGND 0.087f
C13507 XThC.Tn[12].n13 VGND 0.14339f
C13508 XThC.Tn[12].t29 VGND 0.01582f
C13509 XThC.Tn[12].t24 VGND 0.01728f
C13510 XThC.Tn[12].n14 VGND 0.03858f
C13511 XThC.Tn[12].n15 VGND 0.02643f
C13512 XThC.Tn[12].n16 VGND 0.087f
C13513 XThC.Tn[12].n17 VGND 0.14339f
C13514 XThC.Tn[12].t16 VGND 0.01582f
C13515 XThC.Tn[12].t13 VGND 0.01728f
C13516 XThC.Tn[12].n18 VGND 0.03858f
C13517 XThC.Tn[12].n19 VGND 0.02643f
C13518 XThC.Tn[12].n20 VGND 0.087f
C13519 XThC.Tn[12].n21 VGND 0.14339f
C13520 XThC.Tn[12].t17 VGND 0.01582f
C13521 XThC.Tn[12].t14 VGND 0.01728f
C13522 XThC.Tn[12].n22 VGND 0.03858f
C13523 XThC.Tn[12].n23 VGND 0.02643f
C13524 XThC.Tn[12].n24 VGND 0.087f
C13525 XThC.Tn[12].n25 VGND 0.14339f
C13526 XThC.Tn[12].t33 VGND 0.01582f
C13527 XThC.Tn[12].t27 VGND 0.01728f
C13528 XThC.Tn[12].n26 VGND 0.03858f
C13529 XThC.Tn[12].n27 VGND 0.02643f
C13530 XThC.Tn[12].n28 VGND 0.087f
C13531 XThC.Tn[12].n29 VGND 0.14339f
C13532 XThC.Tn[12].t40 VGND 0.01582f
C13533 XThC.Tn[12].t36 VGND 0.01728f
C13534 XThC.Tn[12].n30 VGND 0.03858f
C13535 XThC.Tn[12].n31 VGND 0.02643f
C13536 XThC.Tn[12].n32 VGND 0.087f
C13537 XThC.Tn[12].n33 VGND 0.14339f
C13538 XThC.Tn[12].t42 VGND 0.01582f
C13539 XThC.Tn[12].t38 VGND 0.01728f
C13540 XThC.Tn[12].n34 VGND 0.03858f
C13541 XThC.Tn[12].n35 VGND 0.02643f
C13542 XThC.Tn[12].n36 VGND 0.087f
C13543 XThC.Tn[12].n37 VGND 0.14339f
C13544 XThC.Tn[12].t30 VGND 0.01582f
C13545 XThC.Tn[12].t25 VGND 0.01728f
C13546 XThC.Tn[12].n38 VGND 0.03858f
C13547 XThC.Tn[12].n39 VGND 0.02643f
C13548 XThC.Tn[12].n40 VGND 0.087f
C13549 XThC.Tn[12].n41 VGND 0.14339f
C13550 XThC.Tn[12].t32 VGND 0.01582f
C13551 XThC.Tn[12].t26 VGND 0.01728f
C13552 XThC.Tn[12].n42 VGND 0.03858f
C13553 XThC.Tn[12].n43 VGND 0.02643f
C13554 XThC.Tn[12].n44 VGND 0.087f
C13555 XThC.Tn[12].n45 VGND 0.14339f
C13556 XThC.Tn[12].t43 VGND 0.01582f
C13557 XThC.Tn[12].t39 VGND 0.01728f
C13558 XThC.Tn[12].n46 VGND 0.03858f
C13559 XThC.Tn[12].n47 VGND 0.02643f
C13560 XThC.Tn[12].n48 VGND 0.087f
C13561 XThC.Tn[12].n49 VGND 0.14339f
C13562 XThC.Tn[12].t19 VGND 0.01582f
C13563 XThC.Tn[12].t15 VGND 0.01728f
C13564 XThC.Tn[12].n50 VGND 0.03858f
C13565 XThC.Tn[12].n51 VGND 0.02643f
C13566 XThC.Tn[12].n52 VGND 0.087f
C13567 XThC.Tn[12].n53 VGND 0.14339f
C13568 XThC.Tn[12].t21 VGND 0.01582f
C13569 XThC.Tn[12].t18 VGND 0.01728f
C13570 XThC.Tn[12].n54 VGND 0.03858f
C13571 XThC.Tn[12].n55 VGND 0.02643f
C13572 XThC.Tn[12].n56 VGND 0.087f
C13573 XThC.Tn[12].n57 VGND 0.14339f
C13574 XThC.Tn[12].t34 VGND 0.01582f
C13575 XThC.Tn[12].t31 VGND 0.01728f
C13576 XThC.Tn[12].n58 VGND 0.03858f
C13577 XThC.Tn[12].n59 VGND 0.02643f
C13578 XThC.Tn[12].n60 VGND 0.087f
C13579 XThC.Tn[12].n61 VGND 0.14339f
C13580 XThC.Tn[12].t12 VGND 0.01582f
C13581 XThC.Tn[12].t41 VGND 0.01728f
C13582 XThC.Tn[12].n62 VGND 0.03858f
C13583 XThC.Tn[12].n63 VGND 0.02643f
C13584 XThC.Tn[12].n64 VGND 0.087f
C13585 XThC.Tn[12].n65 VGND 0.14339f
C13586 XThC.Tn[12].n66 VGND 0.68185f
C13587 XThC.Tn[12].n67 VGND 0.24221f
C13588 XThC.Tn[12].t1 VGND 0.01996f
C13589 XThC.Tn[12].t2 VGND 0.01996f
C13590 XThC.Tn[12].n68 VGND 0.04313f
C13591 XThC.Tn[12].t0 VGND 0.01996f
C13592 XThC.Tn[12].t3 VGND 0.01996f
C13593 XThC.Tn[12].n69 VGND 0.06565f
C13594 XThC.Tn[12].n70 VGND 0.18241f
C13595 XThC.Tn[12].n71 VGND 0.02868f
C13596 XThC.Tn[12].t9 VGND 0.01996f
C13597 XThC.Tn[12].t8 VGND 0.01996f
C13598 XThC.Tn[12].n72 VGND 0.06062f
C13599 XThC.Tn[12].t11 VGND 0.01996f
C13600 XThC.Tn[12].t10 VGND 0.01996f
C13601 XThC.Tn[12].n73 VGND 0.04438f
C13602 XThC.Tn[12].n74 VGND 0.19752f
C13603 XThC.Tn[11].t7 VGND 0.01319f
C13604 XThC.Tn[11].t10 VGND 0.01319f
C13605 XThC.Tn[11].n0 VGND 0.0329f
C13606 XThC.Tn[11].t5 VGND 0.01319f
C13607 XThC.Tn[11].t11 VGND 0.01319f
C13608 XThC.Tn[11].n1 VGND 0.02638f
C13609 XThC.Tn[11].n2 VGND 0.06083f
C13610 XThC.Tn[11].t20 VGND 0.01608f
C13611 XThC.Tn[11].t18 VGND 0.01757f
C13612 XThC.Tn[11].n3 VGND 0.03922f
C13613 XThC.Tn[11].n4 VGND 0.02687f
C13614 XThC.Tn[11].n5 VGND 0.08819f
C13615 XThC.Tn[11].t38 VGND 0.01608f
C13616 XThC.Tn[11].t35 VGND 0.01757f
C13617 XThC.Tn[11].n6 VGND 0.03922f
C13618 XThC.Tn[11].n7 VGND 0.02687f
C13619 XThC.Tn[11].n8 VGND 0.08843f
C13620 XThC.Tn[11].n9 VGND 0.14574f
C13621 XThC.Tn[11].t43 VGND 0.01608f
C13622 XThC.Tn[11].t37 VGND 0.01757f
C13623 XThC.Tn[11].n10 VGND 0.03922f
C13624 XThC.Tn[11].n11 VGND 0.02687f
C13625 XThC.Tn[11].n12 VGND 0.08843f
C13626 XThC.Tn[11].n13 VGND 0.14574f
C13627 XThC.Tn[11].t12 VGND 0.01608f
C13628 XThC.Tn[11].t39 VGND 0.01757f
C13629 XThC.Tn[11].n14 VGND 0.03922f
C13630 XThC.Tn[11].n15 VGND 0.02687f
C13631 XThC.Tn[11].n16 VGND 0.08843f
C13632 XThC.Tn[11].n17 VGND 0.14574f
C13633 XThC.Tn[11].t31 VGND 0.01608f
C13634 XThC.Tn[11].t28 VGND 0.01757f
C13635 XThC.Tn[11].n18 VGND 0.03922f
C13636 XThC.Tn[11].n19 VGND 0.02687f
C13637 XThC.Tn[11].n20 VGND 0.08843f
C13638 XThC.Tn[11].n21 VGND 0.14574f
C13639 XThC.Tn[11].t32 VGND 0.01608f
C13640 XThC.Tn[11].t29 VGND 0.01757f
C13641 XThC.Tn[11].n22 VGND 0.03922f
C13642 XThC.Tn[11].n23 VGND 0.02687f
C13643 XThC.Tn[11].n24 VGND 0.08843f
C13644 XThC.Tn[11].n25 VGND 0.14574f
C13645 XThC.Tn[11].t16 VGND 0.01608f
C13646 XThC.Tn[11].t42 VGND 0.01757f
C13647 XThC.Tn[11].n26 VGND 0.03922f
C13648 XThC.Tn[11].n27 VGND 0.02687f
C13649 XThC.Tn[11].n28 VGND 0.08843f
C13650 XThC.Tn[11].n29 VGND 0.14574f
C13651 XThC.Tn[11].t23 VGND 0.01608f
C13652 XThC.Tn[11].t19 VGND 0.01757f
C13653 XThC.Tn[11].n30 VGND 0.03922f
C13654 XThC.Tn[11].n31 VGND 0.02687f
C13655 XThC.Tn[11].n32 VGND 0.08843f
C13656 XThC.Tn[11].n33 VGND 0.14574f
C13657 XThC.Tn[11].t25 VGND 0.01608f
C13658 XThC.Tn[11].t21 VGND 0.01757f
C13659 XThC.Tn[11].n34 VGND 0.03922f
C13660 XThC.Tn[11].n35 VGND 0.02687f
C13661 XThC.Tn[11].n36 VGND 0.08843f
C13662 XThC.Tn[11].n37 VGND 0.14574f
C13663 XThC.Tn[11].t13 VGND 0.01608f
C13664 XThC.Tn[11].t40 VGND 0.01757f
C13665 XThC.Tn[11].n38 VGND 0.03922f
C13666 XThC.Tn[11].n39 VGND 0.02687f
C13667 XThC.Tn[11].n40 VGND 0.08843f
C13668 XThC.Tn[11].n41 VGND 0.14574f
C13669 XThC.Tn[11].t15 VGND 0.01608f
C13670 XThC.Tn[11].t41 VGND 0.01757f
C13671 XThC.Tn[11].n42 VGND 0.03922f
C13672 XThC.Tn[11].n43 VGND 0.02687f
C13673 XThC.Tn[11].n44 VGND 0.08843f
C13674 XThC.Tn[11].n45 VGND 0.14574f
C13675 XThC.Tn[11].t26 VGND 0.01608f
C13676 XThC.Tn[11].t22 VGND 0.01757f
C13677 XThC.Tn[11].n46 VGND 0.03922f
C13678 XThC.Tn[11].n47 VGND 0.02687f
C13679 XThC.Tn[11].n48 VGND 0.08843f
C13680 XThC.Tn[11].n49 VGND 0.14574f
C13681 XThC.Tn[11].t34 VGND 0.01608f
C13682 XThC.Tn[11].t30 VGND 0.01757f
C13683 XThC.Tn[11].n50 VGND 0.03922f
C13684 XThC.Tn[11].n51 VGND 0.02687f
C13685 XThC.Tn[11].n52 VGND 0.08843f
C13686 XThC.Tn[11].n53 VGND 0.14574f
C13687 XThC.Tn[11].t36 VGND 0.01608f
C13688 XThC.Tn[11].t33 VGND 0.01757f
C13689 XThC.Tn[11].n54 VGND 0.03922f
C13690 XThC.Tn[11].n55 VGND 0.02687f
C13691 XThC.Tn[11].n56 VGND 0.08843f
C13692 XThC.Tn[11].n57 VGND 0.14574f
C13693 XThC.Tn[11].t17 VGND 0.01608f
C13694 XThC.Tn[11].t14 VGND 0.01757f
C13695 XThC.Tn[11].n58 VGND 0.03922f
C13696 XThC.Tn[11].n59 VGND 0.02687f
C13697 XThC.Tn[11].n60 VGND 0.08843f
C13698 XThC.Tn[11].n61 VGND 0.14574f
C13699 XThC.Tn[11].t27 VGND 0.01608f
C13700 XThC.Tn[11].t24 VGND 0.01757f
C13701 XThC.Tn[11].n62 VGND 0.03922f
C13702 XThC.Tn[11].n63 VGND 0.02687f
C13703 XThC.Tn[11].n64 VGND 0.08843f
C13704 XThC.Tn[11].n65 VGND 0.14574f
C13705 XThC.Tn[11].n66 VGND 0.6764f
C13706 XThC.Tn[11].n67 VGND 0.26496f
C13707 XThC.Tn[11].t4 VGND 0.02029f
C13708 XThC.Tn[11].t9 VGND 0.02029f
C13709 XThC.Tn[11].n68 VGND 0.04384f
C13710 XThC.Tn[11].t6 VGND 0.02029f
C13711 XThC.Tn[11].t8 VGND 0.02029f
C13712 XThC.Tn[11].n69 VGND 0.06911f
C13713 XThC.Tn[11].n70 VGND 0.18303f
C13714 XThC.Tn[11].n71 VGND 0.01348f
C13715 XThC.Tn[11].t2 VGND 0.02029f
C13716 XThC.Tn[11].t1 VGND 0.02029f
C13717 XThC.Tn[11].n72 VGND 0.04511f
C13718 XThC.Tn[11].t0 VGND 0.02029f
C13719 XThC.Tn[11].t3 VGND 0.02029f
C13720 XThC.Tn[11].n73 VGND 0.06161f
C13721 XThC.Tn[11].n74 VGND 0.20076f
C13722 XThC.Tn[9].t9 VGND 0.013f
C13723 XThC.Tn[9].t8 VGND 0.013f
C13724 XThC.Tn[9].n0 VGND 0.03242f
C13725 XThC.Tn[9].t10 VGND 0.013f
C13726 XThC.Tn[9].t11 VGND 0.013f
C13727 XThC.Tn[9].n1 VGND 0.026f
C13728 XThC.Tn[9].n2 VGND 0.05995f
C13729 XThC.Tn[9].t26 VGND 0.01585f
C13730 XThC.Tn[9].t12 VGND 0.01732f
C13731 XThC.Tn[9].n3 VGND 0.03865f
C13732 XThC.Tn[9].n4 VGND 0.02648f
C13733 XThC.Tn[9].n5 VGND 0.08692f
C13734 XThC.Tn[9].t13 VGND 0.01585f
C13735 XThC.Tn[9].t30 VGND 0.01732f
C13736 XThC.Tn[9].n6 VGND 0.03865f
C13737 XThC.Tn[9].n7 VGND 0.02648f
C13738 XThC.Tn[9].n8 VGND 0.08716f
C13739 XThC.Tn[9].n9 VGND 0.14365f
C13740 XThC.Tn[9].t15 VGND 0.01585f
C13741 XThC.Tn[9].t34 VGND 0.01732f
C13742 XThC.Tn[9].n10 VGND 0.03865f
C13743 XThC.Tn[9].n11 VGND 0.02648f
C13744 XThC.Tn[9].n12 VGND 0.08716f
C13745 XThC.Tn[9].n13 VGND 0.14365f
C13746 XThC.Tn[9].t17 VGND 0.01585f
C13747 XThC.Tn[9].t35 VGND 0.01732f
C13748 XThC.Tn[9].n14 VGND 0.03865f
C13749 XThC.Tn[9].n15 VGND 0.02648f
C13750 XThC.Tn[9].n16 VGND 0.08716f
C13751 XThC.Tn[9].n17 VGND 0.14365f
C13752 XThC.Tn[9].t39 VGND 0.01585f
C13753 XThC.Tn[9].t24 VGND 0.01732f
C13754 XThC.Tn[9].n18 VGND 0.03865f
C13755 XThC.Tn[9].n19 VGND 0.02648f
C13756 XThC.Tn[9].n20 VGND 0.08716f
C13757 XThC.Tn[9].n21 VGND 0.14365f
C13758 XThC.Tn[9].t40 VGND 0.01585f
C13759 XThC.Tn[9].t25 VGND 0.01732f
C13760 XThC.Tn[9].n22 VGND 0.03865f
C13761 XThC.Tn[9].n23 VGND 0.02648f
C13762 XThC.Tn[9].n24 VGND 0.08716f
C13763 XThC.Tn[9].n25 VGND 0.14365f
C13764 XThC.Tn[9].t22 VGND 0.01585f
C13765 XThC.Tn[9].t38 VGND 0.01732f
C13766 XThC.Tn[9].n26 VGND 0.03865f
C13767 XThC.Tn[9].n27 VGND 0.02648f
C13768 XThC.Tn[9].n28 VGND 0.08716f
C13769 XThC.Tn[9].n29 VGND 0.14365f
C13770 XThC.Tn[9].t28 VGND 0.01585f
C13771 XThC.Tn[9].t14 VGND 0.01732f
C13772 XThC.Tn[9].n30 VGND 0.03865f
C13773 XThC.Tn[9].n31 VGND 0.02648f
C13774 XThC.Tn[9].n32 VGND 0.08716f
C13775 XThC.Tn[9].n33 VGND 0.14365f
C13776 XThC.Tn[9].t31 VGND 0.01585f
C13777 XThC.Tn[9].t16 VGND 0.01732f
C13778 XThC.Tn[9].n34 VGND 0.03865f
C13779 XThC.Tn[9].n35 VGND 0.02648f
C13780 XThC.Tn[9].n36 VGND 0.08716f
C13781 XThC.Tn[9].n37 VGND 0.14365f
C13782 XThC.Tn[9].t19 VGND 0.01585f
C13783 XThC.Tn[9].t36 VGND 0.01732f
C13784 XThC.Tn[9].n38 VGND 0.03865f
C13785 XThC.Tn[9].n39 VGND 0.02648f
C13786 XThC.Tn[9].n40 VGND 0.08716f
C13787 XThC.Tn[9].n41 VGND 0.14365f
C13788 XThC.Tn[9].t21 VGND 0.01585f
C13789 XThC.Tn[9].t37 VGND 0.01732f
C13790 XThC.Tn[9].n42 VGND 0.03865f
C13791 XThC.Tn[9].n43 VGND 0.02648f
C13792 XThC.Tn[9].n44 VGND 0.08716f
C13793 XThC.Tn[9].n45 VGND 0.14365f
C13794 XThC.Tn[9].t32 VGND 0.01585f
C13795 XThC.Tn[9].t18 VGND 0.01732f
C13796 XThC.Tn[9].n46 VGND 0.03865f
C13797 XThC.Tn[9].n47 VGND 0.02648f
C13798 XThC.Tn[9].n48 VGND 0.08716f
C13799 XThC.Tn[9].n49 VGND 0.14365f
C13800 XThC.Tn[9].t42 VGND 0.01585f
C13801 XThC.Tn[9].t27 VGND 0.01732f
C13802 XThC.Tn[9].n50 VGND 0.03865f
C13803 XThC.Tn[9].n51 VGND 0.02648f
C13804 XThC.Tn[9].n52 VGND 0.08716f
C13805 XThC.Tn[9].n53 VGND 0.14365f
C13806 XThC.Tn[9].t43 VGND 0.01585f
C13807 XThC.Tn[9].t29 VGND 0.01732f
C13808 XThC.Tn[9].n54 VGND 0.03865f
C13809 XThC.Tn[9].n55 VGND 0.02648f
C13810 XThC.Tn[9].n56 VGND 0.08716f
C13811 XThC.Tn[9].n57 VGND 0.14365f
C13812 XThC.Tn[9].t23 VGND 0.01585f
C13813 XThC.Tn[9].t41 VGND 0.01732f
C13814 XThC.Tn[9].n58 VGND 0.03865f
C13815 XThC.Tn[9].n59 VGND 0.02648f
C13816 XThC.Tn[9].n60 VGND 0.08716f
C13817 XThC.Tn[9].n61 VGND 0.14365f
C13818 XThC.Tn[9].t33 VGND 0.01585f
C13819 XThC.Tn[9].t20 VGND 0.01732f
C13820 XThC.Tn[9].n62 VGND 0.03865f
C13821 XThC.Tn[9].n63 VGND 0.02648f
C13822 XThC.Tn[9].n64 VGND 0.08716f
C13823 XThC.Tn[9].n65 VGND 0.14365f
C13824 XThC.Tn[9].n66 VGND 0.61747f
C13825 XThC.Tn[9].n67 VGND 0.26115f
C13826 XThC.Tn[9].t4 VGND 0.02f
C13827 XThC.Tn[9].t7 VGND 0.02f
C13828 XThC.Tn[9].n68 VGND 0.04321f
C13829 XThC.Tn[9].t6 VGND 0.02f
C13830 XThC.Tn[9].t5 VGND 0.02f
C13831 XThC.Tn[9].n69 VGND 0.06812f
C13832 XThC.Tn[9].n70 VGND 0.1804f
C13833 XThC.Tn[9].n71 VGND 0.01328f
C13834 XThC.Tn[9].t1 VGND 0.02f
C13835 XThC.Tn[9].t0 VGND 0.02f
C13836 XThC.Tn[9].n72 VGND 0.06073f
C13837 XThC.Tn[9].t3 VGND 0.02f
C13838 XThC.Tn[9].t2 VGND 0.02f
C13839 XThC.Tn[9].n73 VGND 0.04446f
C13840 XThC.Tn[9].n74 VGND 0.19787f
C13841 XThC.Tn[5].t7 VGND 0.01807f
C13842 XThC.Tn[5].t6 VGND 0.01807f
C13843 XThC.Tn[5].n0 VGND 0.03647f
C13844 XThC.Tn[5].t5 VGND 0.01807f
C13845 XThC.Tn[5].t4 VGND 0.01807f
C13846 XThC.Tn[5].n1 VGND 0.04267f
C13847 XThC.Tn[5].n2 VGND 0.12799f
C13848 XThC.Tn[5].t9 VGND 0.01174f
C13849 XThC.Tn[5].t8 VGND 0.01174f
C13850 XThC.Tn[5].n3 VGND 0.02674f
C13851 XThC.Tn[5].t11 VGND 0.01174f
C13852 XThC.Tn[5].t10 VGND 0.01174f
C13853 XThC.Tn[5].n4 VGND 0.02674f
C13854 XThC.Tn[5].t2 VGND 0.01174f
C13855 XThC.Tn[5].t1 VGND 0.01174f
C13856 XThC.Tn[5].n5 VGND 0.02674f
C13857 XThC.Tn[5].t0 VGND 0.01174f
C13858 XThC.Tn[5].t3 VGND 0.01174f
C13859 XThC.Tn[5].n6 VGND 0.04456f
C13860 XThC.Tn[5].n7 VGND 0.12735f
C13861 XThC.Tn[5].n8 VGND 0.07873f
C13862 XThC.Tn[5].n9 VGND 0.08885f
C13863 XThC.Tn[5].t15 VGND 0.01432f
C13864 XThC.Tn[5].t33 VGND 0.01564f
C13865 XThC.Tn[5].n10 VGND 0.03492f
C13866 XThC.Tn[5].n11 VGND 0.02392f
C13867 XThC.Tn[5].n12 VGND 0.07852f
C13868 XThC.Tn[5].t34 VGND 0.01432f
C13869 XThC.Tn[5].t19 VGND 0.01564f
C13870 XThC.Tn[5].n13 VGND 0.03492f
C13871 XThC.Tn[5].n14 VGND 0.02392f
C13872 XThC.Tn[5].n15 VGND 0.07873f
C13873 XThC.Tn[5].n16 VGND 0.12976f
C13874 XThC.Tn[5].t36 VGND 0.01432f
C13875 XThC.Tn[5].t23 VGND 0.01564f
C13876 XThC.Tn[5].n17 VGND 0.03492f
C13877 XThC.Tn[5].n18 VGND 0.02392f
C13878 XThC.Tn[5].n19 VGND 0.07873f
C13879 XThC.Tn[5].n20 VGND 0.12976f
C13880 XThC.Tn[5].t38 VGND 0.01432f
C13881 XThC.Tn[5].t24 VGND 0.01564f
C13882 XThC.Tn[5].n21 VGND 0.03492f
C13883 XThC.Tn[5].n22 VGND 0.02392f
C13884 XThC.Tn[5].n23 VGND 0.07873f
C13885 XThC.Tn[5].n24 VGND 0.12976f
C13886 XThC.Tn[5].t28 VGND 0.01432f
C13887 XThC.Tn[5].t13 VGND 0.01564f
C13888 XThC.Tn[5].n25 VGND 0.03492f
C13889 XThC.Tn[5].n26 VGND 0.02392f
C13890 XThC.Tn[5].n27 VGND 0.07873f
C13891 XThC.Tn[5].n28 VGND 0.12976f
C13892 XThC.Tn[5].t29 VGND 0.01432f
C13893 XThC.Tn[5].t14 VGND 0.01564f
C13894 XThC.Tn[5].n29 VGND 0.03492f
C13895 XThC.Tn[5].n30 VGND 0.02392f
C13896 XThC.Tn[5].n31 VGND 0.07873f
C13897 XThC.Tn[5].n32 VGND 0.12976f
C13898 XThC.Tn[5].t43 VGND 0.01432f
C13899 XThC.Tn[5].t27 VGND 0.01564f
C13900 XThC.Tn[5].n33 VGND 0.03492f
C13901 XThC.Tn[5].n34 VGND 0.02392f
C13902 XThC.Tn[5].n35 VGND 0.07873f
C13903 XThC.Tn[5].n36 VGND 0.12976f
C13904 XThC.Tn[5].t17 VGND 0.01432f
C13905 XThC.Tn[5].t35 VGND 0.01564f
C13906 XThC.Tn[5].n37 VGND 0.03492f
C13907 XThC.Tn[5].n38 VGND 0.02392f
C13908 XThC.Tn[5].n39 VGND 0.07873f
C13909 XThC.Tn[5].n40 VGND 0.12976f
C13910 XThC.Tn[5].t20 VGND 0.01432f
C13911 XThC.Tn[5].t37 VGND 0.01564f
C13912 XThC.Tn[5].n41 VGND 0.03492f
C13913 XThC.Tn[5].n42 VGND 0.02392f
C13914 XThC.Tn[5].n43 VGND 0.07873f
C13915 XThC.Tn[5].n44 VGND 0.12976f
C13916 XThC.Tn[5].t40 VGND 0.01432f
C13917 XThC.Tn[5].t25 VGND 0.01564f
C13918 XThC.Tn[5].n45 VGND 0.03492f
C13919 XThC.Tn[5].n46 VGND 0.02392f
C13920 XThC.Tn[5].n47 VGND 0.07873f
C13921 XThC.Tn[5].n48 VGND 0.12976f
C13922 XThC.Tn[5].t42 VGND 0.01432f
C13923 XThC.Tn[5].t26 VGND 0.01564f
C13924 XThC.Tn[5].n49 VGND 0.03492f
C13925 XThC.Tn[5].n50 VGND 0.02392f
C13926 XThC.Tn[5].n51 VGND 0.07873f
C13927 XThC.Tn[5].n52 VGND 0.12976f
C13928 XThC.Tn[5].t21 VGND 0.01432f
C13929 XThC.Tn[5].t39 VGND 0.01564f
C13930 XThC.Tn[5].n53 VGND 0.03492f
C13931 XThC.Tn[5].n54 VGND 0.02392f
C13932 XThC.Tn[5].n55 VGND 0.07873f
C13933 XThC.Tn[5].n56 VGND 0.12976f
C13934 XThC.Tn[5].t31 VGND 0.01432f
C13935 XThC.Tn[5].t16 VGND 0.01564f
C13936 XThC.Tn[5].n57 VGND 0.03492f
C13937 XThC.Tn[5].n58 VGND 0.02392f
C13938 XThC.Tn[5].n59 VGND 0.07873f
C13939 XThC.Tn[5].n60 VGND 0.12976f
C13940 XThC.Tn[5].t32 VGND 0.01432f
C13941 XThC.Tn[5].t18 VGND 0.01564f
C13942 XThC.Tn[5].n61 VGND 0.03492f
C13943 XThC.Tn[5].n62 VGND 0.02392f
C13944 XThC.Tn[5].n63 VGND 0.07873f
C13945 XThC.Tn[5].n64 VGND 0.12976f
C13946 XThC.Tn[5].t12 VGND 0.01432f
C13947 XThC.Tn[5].t30 VGND 0.01564f
C13948 XThC.Tn[5].n65 VGND 0.03492f
C13949 XThC.Tn[5].n66 VGND 0.02392f
C13950 XThC.Tn[5].n67 VGND 0.07873f
C13951 XThC.Tn[5].n68 VGND 0.12976f
C13952 XThC.Tn[5].t22 VGND 0.01432f
C13953 XThC.Tn[5].t41 VGND 0.01564f
C13954 XThC.Tn[5].n69 VGND 0.03492f
C13955 XThC.Tn[5].n70 VGND 0.02392f
C13956 XThC.Tn[5].n71 VGND 0.07873f
C13957 XThC.Tn[5].n72 VGND 0.12976f
C13958 XThC.Tn[5].n73 VGND 0.14766f
C13959 XThR.Tn[9].t10 VGND 0.02425f
C13960 XThR.Tn[9].t8 VGND 0.02425f
C13961 XThR.Tn[9].n0 VGND 0.07362f
C13962 XThR.Tn[9].t11 VGND 0.02425f
C13963 XThR.Tn[9].t9 VGND 0.02425f
C13964 XThR.Tn[9].n1 VGND 0.0539f
C13965 XThR.Tn[9].n2 VGND 0.24507f
C13966 XThR.Tn[9].t5 VGND 0.01576f
C13967 XThR.Tn[9].t7 VGND 0.01576f
C13968 XThR.Tn[9].n3 VGND 0.03931f
C13969 XThR.Tn[9].t4 VGND 0.01576f
C13970 XThR.Tn[9].t6 VGND 0.01576f
C13971 XThR.Tn[9].n4 VGND 0.03152f
C13972 XThR.Tn[9].n5 VGND 0.07929f
C13973 XThR.Tn[9].t17 VGND 0.01895f
C13974 XThR.Tn[9].t71 VGND 0.02075f
C13975 XThR.Tn[9].n6 VGND 0.05067f
C13976 XThR.Tn[9].n7 VGND 0.09733f
C13977 XThR.Tn[9].t35 VGND 0.01895f
C13978 XThR.Tn[9].t28 VGND 0.02075f
C13979 XThR.Tn[9].n8 VGND 0.05067f
C13980 XThR.Tn[9].t50 VGND 0.01889f
C13981 XThR.Tn[9].t19 VGND 0.02068f
C13982 XThR.Tn[9].n9 VGND 0.05272f
C13983 XThR.Tn[9].n10 VGND 0.03704f
C13984 XThR.Tn[9].n11 VGND 0.00677f
C13985 XThR.Tn[9].n12 VGND 0.11885f
C13986 XThR.Tn[9].t72 VGND 0.01895f
C13987 XThR.Tn[9].t64 VGND 0.02075f
C13988 XThR.Tn[9].n13 VGND 0.05067f
C13989 XThR.Tn[9].t26 VGND 0.01889f
C13990 XThR.Tn[9].t59 VGND 0.02068f
C13991 XThR.Tn[9].n14 VGND 0.05272f
C13992 XThR.Tn[9].n15 VGND 0.03704f
C13993 XThR.Tn[9].n16 VGND 0.00677f
C13994 XThR.Tn[9].n17 VGND 0.11885f
C13995 XThR.Tn[9].t29 VGND 0.01895f
C13996 XThR.Tn[9].t21 VGND 0.02075f
C13997 XThR.Tn[9].n18 VGND 0.05067f
C13998 XThR.Tn[9].t41 VGND 0.01889f
C13999 XThR.Tn[9].t15 VGND 0.02068f
C14000 XThR.Tn[9].n19 VGND 0.05272f
C14001 XThR.Tn[9].n20 VGND 0.03704f
C14002 XThR.Tn[9].n21 VGND 0.00677f
C14003 XThR.Tn[9].n22 VGND 0.11885f
C14004 XThR.Tn[9].t56 VGND 0.01895f
C14005 XThR.Tn[9].t46 VGND 0.02075f
C14006 XThR.Tn[9].n23 VGND 0.05067f
C14007 XThR.Tn[9].t73 VGND 0.01889f
C14008 XThR.Tn[9].t42 VGND 0.02068f
C14009 XThR.Tn[9].n24 VGND 0.05272f
C14010 XThR.Tn[9].n25 VGND 0.03704f
C14011 XThR.Tn[9].n26 VGND 0.00677f
C14012 XThR.Tn[9].n27 VGND 0.11885f
C14013 XThR.Tn[9].t31 VGND 0.01895f
C14014 XThR.Tn[9].t23 VGND 0.02075f
C14015 XThR.Tn[9].n28 VGND 0.05067f
C14016 XThR.Tn[9].t44 VGND 0.01889f
C14017 XThR.Tn[9].t16 VGND 0.02068f
C14018 XThR.Tn[9].n29 VGND 0.05272f
C14019 XThR.Tn[9].n30 VGND 0.03704f
C14020 XThR.Tn[9].n31 VGND 0.00677f
C14021 XThR.Tn[9].n32 VGND 0.11885f
C14022 XThR.Tn[9].t67 VGND 0.01895f
C14023 XThR.Tn[9].t37 VGND 0.02075f
C14024 XThR.Tn[9].n33 VGND 0.05067f
C14025 XThR.Tn[9].t20 VGND 0.01889f
C14026 XThR.Tn[9].t33 VGND 0.02068f
C14027 XThR.Tn[9].n34 VGND 0.05272f
C14028 XThR.Tn[9].n35 VGND 0.03704f
C14029 XThR.Tn[9].n36 VGND 0.00677f
C14030 XThR.Tn[9].n37 VGND 0.11885f
C14031 XThR.Tn[9].t36 VGND 0.01895f
C14032 XThR.Tn[9].t32 VGND 0.02075f
C14033 XThR.Tn[9].n38 VGND 0.05067f
C14034 XThR.Tn[9].t51 VGND 0.01889f
C14035 XThR.Tn[9].t25 VGND 0.02068f
C14036 XThR.Tn[9].n39 VGND 0.05272f
C14037 XThR.Tn[9].n40 VGND 0.03704f
C14038 XThR.Tn[9].n41 VGND 0.00677f
C14039 XThR.Tn[9].n42 VGND 0.11885f
C14040 XThR.Tn[9].t39 VGND 0.01895f
C14041 XThR.Tn[9].t45 VGND 0.02075f
C14042 XThR.Tn[9].n43 VGND 0.05067f
C14043 XThR.Tn[9].t55 VGND 0.01889f
C14044 XThR.Tn[9].t40 VGND 0.02068f
C14045 XThR.Tn[9].n44 VGND 0.05272f
C14046 XThR.Tn[9].n45 VGND 0.03704f
C14047 XThR.Tn[9].n46 VGND 0.00677f
C14048 XThR.Tn[9].n47 VGND 0.11885f
C14049 XThR.Tn[9].t58 VGND 0.01895f
C14050 XThR.Tn[9].t66 VGND 0.02075f
C14051 XThR.Tn[9].n48 VGND 0.05067f
C14052 XThR.Tn[9].t13 VGND 0.01889f
C14053 XThR.Tn[9].t60 VGND 0.02068f
C14054 XThR.Tn[9].n49 VGND 0.05272f
C14055 XThR.Tn[9].n50 VGND 0.03704f
C14056 XThR.Tn[9].n51 VGND 0.00677f
C14057 XThR.Tn[9].n52 VGND 0.11885f
C14058 XThR.Tn[9].t48 VGND 0.01895f
C14059 XThR.Tn[9].t24 VGND 0.02075f
C14060 XThR.Tn[9].n53 VGND 0.05067f
C14061 XThR.Tn[9].t65 VGND 0.01889f
C14062 XThR.Tn[9].t18 VGND 0.02068f
C14063 XThR.Tn[9].n54 VGND 0.05272f
C14064 XThR.Tn[9].n55 VGND 0.03704f
C14065 XThR.Tn[9].n56 VGND 0.00677f
C14066 XThR.Tn[9].n57 VGND 0.11885f
C14067 XThR.Tn[9].t70 VGND 0.01895f
C14068 XThR.Tn[9].t62 VGND 0.02075f
C14069 XThR.Tn[9].n58 VGND 0.05067f
C14070 XThR.Tn[9].t22 VGND 0.01889f
C14071 XThR.Tn[9].t52 VGND 0.02068f
C14072 XThR.Tn[9].n59 VGND 0.05272f
C14073 XThR.Tn[9].n60 VGND 0.03704f
C14074 XThR.Tn[9].n61 VGND 0.00677f
C14075 XThR.Tn[9].n62 VGND 0.11885f
C14076 XThR.Tn[9].t38 VGND 0.01895f
C14077 XThR.Tn[9].t34 VGND 0.02075f
C14078 XThR.Tn[9].n63 VGND 0.05067f
C14079 XThR.Tn[9].t53 VGND 0.01889f
C14080 XThR.Tn[9].t27 VGND 0.02068f
C14081 XThR.Tn[9].n64 VGND 0.05272f
C14082 XThR.Tn[9].n65 VGND 0.03704f
C14083 XThR.Tn[9].n66 VGND 0.00677f
C14084 XThR.Tn[9].n67 VGND 0.11885f
C14085 XThR.Tn[9].t57 VGND 0.01895f
C14086 XThR.Tn[9].t47 VGND 0.02075f
C14087 XThR.Tn[9].n68 VGND 0.05067f
C14088 XThR.Tn[9].t12 VGND 0.01889f
C14089 XThR.Tn[9].t43 VGND 0.02068f
C14090 XThR.Tn[9].n69 VGND 0.05272f
C14091 XThR.Tn[9].n70 VGND 0.03704f
C14092 XThR.Tn[9].n71 VGND 0.00677f
C14093 XThR.Tn[9].n72 VGND 0.11885f
C14094 XThR.Tn[9].t14 VGND 0.01895f
C14095 XThR.Tn[9].t69 VGND 0.02075f
C14096 XThR.Tn[9].n73 VGND 0.05067f
C14097 XThR.Tn[9].t30 VGND 0.01889f
C14098 XThR.Tn[9].t61 VGND 0.02068f
C14099 XThR.Tn[9].n74 VGND 0.05272f
C14100 XThR.Tn[9].n75 VGND 0.03704f
C14101 XThR.Tn[9].n76 VGND 0.00677f
C14102 XThR.Tn[9].n77 VGND 0.11885f
C14103 XThR.Tn[9].t49 VGND 0.01895f
C14104 XThR.Tn[9].t63 VGND 0.02075f
C14105 XThR.Tn[9].n78 VGND 0.05067f
C14106 XThR.Tn[9].t68 VGND 0.01889f
C14107 XThR.Tn[9].t54 VGND 0.02068f
C14108 XThR.Tn[9].n79 VGND 0.05272f
C14109 XThR.Tn[9].n80 VGND 0.03704f
C14110 XThR.Tn[9].n81 VGND 0.00677f
C14111 XThR.Tn[9].n82 VGND 0.11885f
C14112 XThR.Tn[9].n83 VGND 0.10801f
C14113 XThR.Tn[9].n84 VGND 0.35039f
C14114 XThR.Tn[9].t2 VGND 0.02425f
C14115 XThR.Tn[9].t0 VGND 0.02425f
C14116 XThR.Tn[9].n85 VGND 0.05239f
C14117 XThR.Tn[9].t3 VGND 0.02425f
C14118 XThR.Tn[9].t1 VGND 0.02425f
C14119 XThR.Tn[9].n86 VGND 0.07973f
C14120 XThR.Tn[9].n87 VGND 0.22139f
C14121 XThR.Tn[9].n88 VGND 0.02964f
C14122 XThC.Tn[6].t7 VGND 0.0182f
C14123 XThC.Tn[6].t6 VGND 0.0182f
C14124 XThC.Tn[6].n0 VGND 0.03674f
C14125 XThC.Tn[6].t5 VGND 0.0182f
C14126 XThC.Tn[6].t4 VGND 0.0182f
C14127 XThC.Tn[6].n1 VGND 0.04298f
C14128 XThC.Tn[6].n2 VGND 0.12033f
C14129 XThC.Tn[6].t8 VGND 0.01183f
C14130 XThC.Tn[6].t11 VGND 0.01183f
C14131 XThC.Tn[6].n3 VGND 0.02694f
C14132 XThC.Tn[6].t10 VGND 0.01183f
C14133 XThC.Tn[6].t9 VGND 0.01183f
C14134 XThC.Tn[6].n4 VGND 0.02694f
C14135 XThC.Tn[6].t1 VGND 0.01183f
C14136 XThC.Tn[6].t0 VGND 0.01183f
C14137 XThC.Tn[6].n5 VGND 0.02694f
C14138 XThC.Tn[6].t3 VGND 0.01183f
C14139 XThC.Tn[6].t2 VGND 0.01183f
C14140 XThC.Tn[6].n6 VGND 0.04489f
C14141 XThC.Tn[6].n7 VGND 0.12829f
C14142 XThC.Tn[6].n8 VGND 0.07931f
C14143 XThC.Tn[6].n9 VGND 0.0895f
C14144 XThC.Tn[6].t23 VGND 0.01443f
C14145 XThC.Tn[6].t26 VGND 0.01576f
C14146 XThC.Tn[6].n10 VGND 0.03517f
C14147 XThC.Tn[6].n11 VGND 0.0241f
C14148 XThC.Tn[6].n12 VGND 0.0791f
C14149 XThC.Tn[6].t40 VGND 0.01443f
C14150 XThC.Tn[6].t13 VGND 0.01576f
C14151 XThC.Tn[6].n13 VGND 0.03517f
C14152 XThC.Tn[6].n14 VGND 0.0241f
C14153 XThC.Tn[6].n15 VGND 0.07932f
C14154 XThC.Tn[6].n16 VGND 0.13072f
C14155 XThC.Tn[6].t42 VGND 0.01443f
C14156 XThC.Tn[6].t17 VGND 0.01576f
C14157 XThC.Tn[6].n17 VGND 0.03517f
C14158 XThC.Tn[6].n18 VGND 0.0241f
C14159 XThC.Tn[6].n19 VGND 0.07932f
C14160 XThC.Tn[6].n20 VGND 0.13072f
C14161 XThC.Tn[6].t12 VGND 0.01443f
C14162 XThC.Tn[6].t18 VGND 0.01576f
C14163 XThC.Tn[6].n21 VGND 0.03517f
C14164 XThC.Tn[6].n22 VGND 0.0241f
C14165 XThC.Tn[6].n23 VGND 0.07932f
C14166 XThC.Tn[6].n24 VGND 0.13072f
C14167 XThC.Tn[6].t33 VGND 0.01443f
C14168 XThC.Tn[6].t37 VGND 0.01576f
C14169 XThC.Tn[6].n25 VGND 0.03517f
C14170 XThC.Tn[6].n26 VGND 0.0241f
C14171 XThC.Tn[6].n27 VGND 0.07932f
C14172 XThC.Tn[6].n28 VGND 0.13072f
C14173 XThC.Tn[6].t35 VGND 0.01443f
C14174 XThC.Tn[6].t38 VGND 0.01576f
C14175 XThC.Tn[6].n29 VGND 0.03517f
C14176 XThC.Tn[6].n30 VGND 0.0241f
C14177 XThC.Tn[6].n31 VGND 0.07932f
C14178 XThC.Tn[6].n32 VGND 0.13072f
C14179 XThC.Tn[6].t16 VGND 0.01443f
C14180 XThC.Tn[6].t22 VGND 0.01576f
C14181 XThC.Tn[6].n33 VGND 0.03517f
C14182 XThC.Tn[6].n34 VGND 0.0241f
C14183 XThC.Tn[6].n35 VGND 0.07932f
C14184 XThC.Tn[6].n36 VGND 0.13072f
C14185 XThC.Tn[6].t25 VGND 0.01443f
C14186 XThC.Tn[6].t29 VGND 0.01576f
C14187 XThC.Tn[6].n37 VGND 0.03517f
C14188 XThC.Tn[6].n38 VGND 0.0241f
C14189 XThC.Tn[6].n39 VGND 0.07932f
C14190 XThC.Tn[6].n40 VGND 0.13072f
C14191 XThC.Tn[6].t27 VGND 0.01443f
C14192 XThC.Tn[6].t31 VGND 0.01576f
C14193 XThC.Tn[6].n41 VGND 0.03517f
C14194 XThC.Tn[6].n42 VGND 0.0241f
C14195 XThC.Tn[6].n43 VGND 0.07932f
C14196 XThC.Tn[6].n44 VGND 0.13072f
C14197 XThC.Tn[6].t14 VGND 0.01443f
C14198 XThC.Tn[6].t19 VGND 0.01576f
C14199 XThC.Tn[6].n45 VGND 0.03517f
C14200 XThC.Tn[6].n46 VGND 0.0241f
C14201 XThC.Tn[6].n47 VGND 0.07932f
C14202 XThC.Tn[6].n48 VGND 0.13072f
C14203 XThC.Tn[6].t15 VGND 0.01443f
C14204 XThC.Tn[6].t21 VGND 0.01576f
C14205 XThC.Tn[6].n49 VGND 0.03517f
C14206 XThC.Tn[6].n50 VGND 0.0241f
C14207 XThC.Tn[6].n51 VGND 0.07932f
C14208 XThC.Tn[6].n52 VGND 0.13072f
C14209 XThC.Tn[6].t28 VGND 0.01443f
C14210 XThC.Tn[6].t32 VGND 0.01576f
C14211 XThC.Tn[6].n53 VGND 0.03517f
C14212 XThC.Tn[6].n54 VGND 0.0241f
C14213 XThC.Tn[6].n55 VGND 0.07932f
C14214 XThC.Tn[6].n56 VGND 0.13072f
C14215 XThC.Tn[6].t36 VGND 0.01443f
C14216 XThC.Tn[6].t41 VGND 0.01576f
C14217 XThC.Tn[6].n57 VGND 0.03517f
C14218 XThC.Tn[6].n58 VGND 0.0241f
C14219 XThC.Tn[6].n59 VGND 0.07932f
C14220 XThC.Tn[6].n60 VGND 0.13072f
C14221 XThC.Tn[6].t39 VGND 0.01443f
C14222 XThC.Tn[6].t43 VGND 0.01576f
C14223 XThC.Tn[6].n61 VGND 0.03517f
C14224 XThC.Tn[6].n62 VGND 0.0241f
C14225 XThC.Tn[6].n63 VGND 0.07932f
C14226 XThC.Tn[6].n64 VGND 0.13072f
C14227 XThC.Tn[6].t20 VGND 0.01443f
C14228 XThC.Tn[6].t24 VGND 0.01576f
C14229 XThC.Tn[6].n65 VGND 0.03517f
C14230 XThC.Tn[6].n66 VGND 0.0241f
C14231 XThC.Tn[6].n67 VGND 0.07932f
C14232 XThC.Tn[6].n68 VGND 0.13072f
C14233 XThC.Tn[6].t30 VGND 0.01443f
C14234 XThC.Tn[6].t34 VGND 0.01576f
C14235 XThC.Tn[6].n69 VGND 0.03517f
C14236 XThC.Tn[6].n70 VGND 0.0241f
C14237 XThC.Tn[6].n71 VGND 0.07932f
C14238 XThC.Tn[6].n72 VGND 0.13072f
C14239 XThC.Tn[6].n73 VGND 0.14537f
C14240 XThC.Tn[6].n74 VGND 0.03808f
C14241 XThC.XTBN.Y.n0 VGND 0.01531f
C14242 XThC.XTBN.Y.t50 VGND 0.01024f
C14243 XThC.XTBN.Y.t118 VGND 0.00603f
C14244 XThC.XTBN.Y.t18 VGND 0.01024f
C14245 XThC.XTBN.Y.t83 VGND 0.00603f
C14246 XThC.XTBN.Y.n1 VGND 0.01477f
C14247 XThC.XTBN.Y.n2 VGND 0.00524f
C14248 XThC.XTBN.Y.t120 VGND 0.01024f
C14249 XThC.XTBN.Y.t71 VGND 0.00603f
C14250 XThC.XTBN.Y.t114 VGND 0.01024f
C14251 XThC.XTBN.Y.t62 VGND 0.00603f
C14252 XThC.XTBN.Y.n3 VGND 0.0138f
C14253 XThC.XTBN.Y.n4 VGND 0.00676f
C14254 XThC.XTBN.Y.n5 VGND 0.01477f
C14255 XThC.XTBN.Y.n6 VGND 0.00676f
C14256 XThC.XTBN.Y.n7 VGND 0.00548f
C14257 XThC.XTBN.Y.n8 VGND 0.00561f
C14258 XThC.XTBN.Y.n9 VGND 0.00676f
C14259 XThC.XTBN.Y.n10 VGND 0.02164f
C14260 XThC.XTBN.Y.n11 VGND 0.00584f
C14261 XThC.XTBN.Y.n12 VGND 0.00877f
C14262 XThC.XTBN.Y.t121 VGND 0.00603f
C14263 XThC.XTBN.Y.t79 VGND 0.01024f
C14264 XThC.XTBN.Y.t84 VGND 0.00603f
C14265 XThC.XTBN.Y.t36 VGND 0.01024f
C14266 XThC.XTBN.Y.n13 VGND 0.01477f
C14267 XThC.XTBN.Y.n14 VGND 0.00524f
C14268 XThC.XTBN.Y.t73 VGND 0.00603f
C14269 XThC.XTBN.Y.t26 VGND 0.01024f
C14270 XThC.XTBN.Y.t64 VGND 0.00603f
C14271 XThC.XTBN.Y.t21 VGND 0.01024f
C14272 XThC.XTBN.Y.n15 VGND 0.0138f
C14273 XThC.XTBN.Y.n16 VGND 0.00676f
C14274 XThC.XTBN.Y.n17 VGND 0.01477f
C14275 XThC.XTBN.Y.n18 VGND 0.00676f
C14276 XThC.XTBN.Y.n19 VGND 0.00548f
C14277 XThC.XTBN.Y.n20 VGND 0.00561f
C14278 XThC.XTBN.Y.n21 VGND 0.00676f
C14279 XThC.XTBN.Y.n22 VGND 0.02164f
C14280 XThC.XTBN.Y.n23 VGND 0.00584f
C14281 XThC.XTBN.Y.n24 VGND 0.00417f
C14282 XThC.XTBN.Y.n25 VGND 0.11789f
C14283 XThC.XTBN.Y.t106 VGND 0.01024f
C14284 XThC.XTBN.Y.t89 VGND 0.00603f
C14285 XThC.XTBN.Y.t70 VGND 0.01024f
C14286 XThC.XTBN.Y.t41 VGND 0.00603f
C14287 XThC.XTBN.Y.n26 VGND 0.01477f
C14288 XThC.XTBN.Y.n27 VGND 0.00524f
C14289 XThC.XTBN.Y.t56 VGND 0.01024f
C14290 XThC.XTBN.Y.t35 VGND 0.00603f
C14291 XThC.XTBN.Y.t48 VGND 0.01024f
C14292 XThC.XTBN.Y.t32 VGND 0.00603f
C14293 XThC.XTBN.Y.n28 VGND 0.0138f
C14294 XThC.XTBN.Y.n29 VGND 0.00676f
C14295 XThC.XTBN.Y.n30 VGND 0.01477f
C14296 XThC.XTBN.Y.n31 VGND 0.00676f
C14297 XThC.XTBN.Y.n32 VGND 0.00548f
C14298 XThC.XTBN.Y.n33 VGND 0.00561f
C14299 XThC.XTBN.Y.n34 VGND 0.00676f
C14300 XThC.XTBN.Y.n35 VGND 0.02164f
C14301 XThC.XTBN.Y.n36 VGND 0.00584f
C14302 XThC.XTBN.Y.n37 VGND 0.00417f
C14303 XThC.XTBN.Y.n38 VGND 0.07443f
C14304 XThC.XTBN.Y.t43 VGND 0.00603f
C14305 XThC.XTBN.Y.t39 VGND 0.01024f
C14306 XThC.XTBN.Y.t10 VGND 0.00603f
C14307 XThC.XTBN.Y.t122 VGND 0.01024f
C14308 XThC.XTBN.Y.n39 VGND 0.01477f
C14309 XThC.XTBN.Y.n40 VGND 0.00524f
C14310 XThC.XTBN.Y.t112 VGND 0.00603f
C14311 XThC.XTBN.Y.t109 VGND 0.01024f
C14312 XThC.XTBN.Y.t108 VGND 0.00603f
C14313 XThC.XTBN.Y.t102 VGND 0.01024f
C14314 XThC.XTBN.Y.n41 VGND 0.0138f
C14315 XThC.XTBN.Y.n42 VGND 0.00676f
C14316 XThC.XTBN.Y.n43 VGND 0.01477f
C14317 XThC.XTBN.Y.n44 VGND 0.00676f
C14318 XThC.XTBN.Y.n45 VGND 0.00548f
C14319 XThC.XTBN.Y.n46 VGND 0.00561f
C14320 XThC.XTBN.Y.n47 VGND 0.00676f
C14321 XThC.XTBN.Y.n48 VGND 0.02164f
C14322 XThC.XTBN.Y.n49 VGND 0.00584f
C14323 XThC.XTBN.Y.n50 VGND 0.00417f
C14324 XThC.XTBN.Y.n51 VGND 0.07443f
C14325 XThC.XTBN.Y.t47 VGND 0.01024f
C14326 XThC.XTBN.Y.t31 VGND 0.00603f
C14327 XThC.XTBN.Y.t17 VGND 0.01024f
C14328 XThC.XTBN.Y.t104 VGND 0.00603f
C14329 XThC.XTBN.Y.n52 VGND 0.01477f
C14330 XThC.XTBN.Y.n53 VGND 0.00524f
C14331 XThC.XTBN.Y.t116 VGND 0.01024f
C14332 XThC.XTBN.Y.t94 VGND 0.00603f
C14333 XThC.XTBN.Y.t111 VGND 0.01024f
C14334 XThC.XTBN.Y.t92 VGND 0.00603f
C14335 XThC.XTBN.Y.n54 VGND 0.0138f
C14336 XThC.XTBN.Y.n55 VGND 0.00676f
C14337 XThC.XTBN.Y.n56 VGND 0.01477f
C14338 XThC.XTBN.Y.n57 VGND 0.00676f
C14339 XThC.XTBN.Y.n58 VGND 0.00548f
C14340 XThC.XTBN.Y.n59 VGND 0.00561f
C14341 XThC.XTBN.Y.n60 VGND 0.00676f
C14342 XThC.XTBN.Y.n61 VGND 0.02164f
C14343 XThC.XTBN.Y.n62 VGND 0.00584f
C14344 XThC.XTBN.Y.n63 VGND 0.00417f
C14345 XThC.XTBN.Y.n64 VGND 0.07443f
C14346 XThC.XTBN.Y.t107 VGND 0.00603f
C14347 XThC.XTBN.Y.t101 VGND 0.01024f
C14348 XThC.XTBN.Y.t72 VGND 0.00603f
C14349 XThC.XTBN.Y.t63 VGND 0.01024f
C14350 XThC.XTBN.Y.n65 VGND 0.01477f
C14351 XThC.XTBN.Y.n66 VGND 0.00524f
C14352 XThC.XTBN.Y.t57 VGND 0.00603f
C14353 XThC.XTBN.Y.t52 VGND 0.01024f
C14354 XThC.XTBN.Y.t49 VGND 0.00603f
C14355 XThC.XTBN.Y.t44 VGND 0.01024f
C14356 XThC.XTBN.Y.n67 VGND 0.0138f
C14357 XThC.XTBN.Y.n68 VGND 0.00676f
C14358 XThC.XTBN.Y.n69 VGND 0.01477f
C14359 XThC.XTBN.Y.n70 VGND 0.00676f
C14360 XThC.XTBN.Y.n71 VGND 0.00548f
C14361 XThC.XTBN.Y.n72 VGND 0.00561f
C14362 XThC.XTBN.Y.n73 VGND 0.00676f
C14363 XThC.XTBN.Y.n74 VGND 0.02164f
C14364 XThC.XTBN.Y.n75 VGND 0.00584f
C14365 XThC.XTBN.Y.n76 VGND 0.00417f
C14366 XThC.XTBN.Y.n77 VGND 0.07443f
C14367 XThC.XTBN.Y.t25 VGND 0.01024f
C14368 XThC.XTBN.Y.t123 VGND 0.00603f
C14369 XThC.XTBN.Y.t100 VGND 0.01024f
C14370 XThC.XTBN.Y.t85 VGND 0.00603f
C14371 XThC.XTBN.Y.n78 VGND 0.01477f
C14372 XThC.XTBN.Y.n79 VGND 0.00524f
C14373 XThC.XTBN.Y.t93 VGND 0.01024f
C14374 XThC.XTBN.Y.t74 VGND 0.00603f
C14375 XThC.XTBN.Y.t90 VGND 0.01024f
C14376 XThC.XTBN.Y.t65 VGND 0.00603f
C14377 XThC.XTBN.Y.n80 VGND 0.0138f
C14378 XThC.XTBN.Y.n81 VGND 0.00676f
C14379 XThC.XTBN.Y.n82 VGND 0.01477f
C14380 XThC.XTBN.Y.n83 VGND 0.00676f
C14381 XThC.XTBN.Y.n84 VGND 0.00548f
C14382 XThC.XTBN.Y.n85 VGND 0.00561f
C14383 XThC.XTBN.Y.n86 VGND 0.00676f
C14384 XThC.XTBN.Y.n87 VGND 0.02164f
C14385 XThC.XTBN.Y.n88 VGND 0.00584f
C14386 XThC.XTBN.Y.n89 VGND 0.00417f
C14387 XThC.XTBN.Y.n90 VGND 0.06646f
C14388 XThC.XTBN.Y.t46 VGND 0.01024f
C14389 XThC.XTBN.Y.t67 VGND 0.00603f
C14390 XThC.XTBN.Y.n91 VGND 0.00619f
C14391 XThC.XTBN.Y.t6 VGND 0.01024f
C14392 XThC.XTBN.Y.t24 VGND 0.00603f
C14393 XThC.XTBN.Y.n92 VGND 0.01243f
C14394 XThC.XTBN.Y.t12 VGND 0.01024f
C14395 XThC.XTBN.Y.t29 VGND 0.00603f
C14396 XThC.XTBN.Y.n93 VGND 0.01348f
C14397 XThC.XTBN.Y.n94 VGND 0.0076f
C14398 XThC.XTBN.Y.n95 VGND 0.01252f
C14399 XThC.XTBN.Y.n96 VGND 0.00434f
C14400 XThC.XTBN.Y.n97 VGND 0.00603f
C14401 XThC.XTBN.Y.n98 VGND 0.01348f
C14402 XThC.XTBN.Y.t54 VGND 0.01024f
C14403 XThC.XTBN.Y.t76 VGND 0.00603f
C14404 XThC.XTBN.Y.n99 VGND 0.01227f
C14405 XThC.XTBN.Y.n100 VGND 0.00676f
C14406 XThC.XTBN.Y.n101 VGND 0.01009f
C14407 XThC.XTBN.Y.t55 VGND 0.00603f
C14408 XThC.XTBN.Y.t38 VGND 0.01024f
C14409 XThC.XTBN.Y.n102 VGND 0.00619f
C14410 XThC.XTBN.Y.t16 VGND 0.00603f
C14411 XThC.XTBN.Y.t113 VGND 0.01024f
C14412 XThC.XTBN.Y.n103 VGND 0.01243f
C14413 XThC.XTBN.Y.t19 VGND 0.00603f
C14414 XThC.XTBN.Y.t119 VGND 0.01024f
C14415 XThC.XTBN.Y.n104 VGND 0.01348f
C14416 XThC.XTBN.Y.n105 VGND 0.0076f
C14417 XThC.XTBN.Y.n106 VGND 0.01252f
C14418 XThC.XTBN.Y.n107 VGND 0.00434f
C14419 XThC.XTBN.Y.n108 VGND 0.00603f
C14420 XThC.XTBN.Y.n109 VGND 0.01348f
C14421 XThC.XTBN.Y.t59 VGND 0.00603f
C14422 XThC.XTBN.Y.t42 VGND 0.01024f
C14423 XThC.XTBN.Y.n110 VGND 0.01227f
C14424 XThC.XTBN.Y.n111 VGND 0.00676f
C14425 XThC.XTBN.Y.n112 VGND 0.00747f
C14426 XThC.XTBN.Y.n113 VGND 0.11256f
C14427 XThC.XTBN.Y.t30 VGND 0.01024f
C14428 XThC.XTBN.Y.t8 VGND 0.00603f
C14429 XThC.XTBN.Y.n114 VGND 0.00619f
C14430 XThC.XTBN.Y.t98 VGND 0.01024f
C14431 XThC.XTBN.Y.t82 VGND 0.00603f
C14432 XThC.XTBN.Y.n115 VGND 0.01243f
C14433 XThC.XTBN.Y.t103 VGND 0.01024f
C14434 XThC.XTBN.Y.t87 VGND 0.00603f
C14435 XThC.XTBN.Y.n116 VGND 0.01348f
C14436 XThC.XTBN.Y.n117 VGND 0.0076f
C14437 XThC.XTBN.Y.n118 VGND 0.01252f
C14438 XThC.XTBN.Y.n119 VGND 0.00434f
C14439 XThC.XTBN.Y.n120 VGND 0.00603f
C14440 XThC.XTBN.Y.n121 VGND 0.01348f
C14441 XThC.XTBN.Y.t34 VGND 0.01024f
C14442 XThC.XTBN.Y.t15 VGND 0.00603f
C14443 XThC.XTBN.Y.n122 VGND 0.01227f
C14444 XThC.XTBN.Y.n123 VGND 0.00676f
C14445 XThC.XTBN.Y.n124 VGND 0.00747f
C14446 XThC.XTBN.Y.n125 VGND 0.07521f
C14447 XThC.XTBN.Y.t110 VGND 0.00603f
C14448 XThC.XTBN.Y.t96 VGND 0.01024f
C14449 XThC.XTBN.Y.n126 VGND 0.00619f
C14450 XThC.XTBN.Y.t68 VGND 0.00603f
C14451 XThC.XTBN.Y.t51 VGND 0.01024f
C14452 XThC.XTBN.Y.n127 VGND 0.01243f
C14453 XThC.XTBN.Y.t77 VGND 0.00603f
C14454 XThC.XTBN.Y.t58 VGND 0.01024f
C14455 XThC.XTBN.Y.n128 VGND 0.01348f
C14456 XThC.XTBN.Y.n129 VGND 0.0076f
C14457 XThC.XTBN.Y.n130 VGND 0.01252f
C14458 XThC.XTBN.Y.n131 VGND 0.00434f
C14459 XThC.XTBN.Y.n132 VGND 0.00603f
C14460 XThC.XTBN.Y.n133 VGND 0.01348f
C14461 XThC.XTBN.Y.t115 VGND 0.00603f
C14462 XThC.XTBN.Y.t99 VGND 0.01024f
C14463 XThC.XTBN.Y.n134 VGND 0.01227f
C14464 XThC.XTBN.Y.n135 VGND 0.00676f
C14465 XThC.XTBN.Y.n136 VGND 0.00747f
C14466 XThC.XTBN.Y.n137 VGND 0.07521f
C14467 XThC.XTBN.Y.t88 VGND 0.01024f
C14468 XThC.XTBN.Y.t60 VGND 0.00603f
C14469 XThC.XTBN.Y.n138 VGND 0.00619f
C14470 XThC.XTBN.Y.t37 VGND 0.01024f
C14471 XThC.XTBN.Y.t20 VGND 0.00603f
C14472 XThC.XTBN.Y.n139 VGND 0.01243f
C14473 XThC.XTBN.Y.t40 VGND 0.01024f
C14474 XThC.XTBN.Y.t22 VGND 0.00603f
C14475 XThC.XTBN.Y.n140 VGND 0.01348f
C14476 XThC.XTBN.Y.n141 VGND 0.0076f
C14477 XThC.XTBN.Y.n142 VGND 0.01252f
C14478 XThC.XTBN.Y.n143 VGND 0.00434f
C14479 XThC.XTBN.Y.n144 VGND 0.00603f
C14480 XThC.XTBN.Y.n145 VGND 0.01348f
C14481 XThC.XTBN.Y.t91 VGND 0.01024f
C14482 XThC.XTBN.Y.t66 VGND 0.00603f
C14483 XThC.XTBN.Y.n146 VGND 0.01227f
C14484 XThC.XTBN.Y.n147 VGND 0.00676f
C14485 XThC.XTBN.Y.n148 VGND 0.00747f
C14486 XThC.XTBN.Y.n149 VGND 0.07534f
C14487 XThC.XTBN.Y.t45 VGND 0.00603f
C14488 XThC.XTBN.Y.t7 VGND 0.01024f
C14489 XThC.XTBN.Y.n150 VGND 0.00619f
C14490 XThC.XTBN.Y.t5 VGND 0.00603f
C14491 XThC.XTBN.Y.t81 VGND 0.01024f
C14492 XThC.XTBN.Y.n151 VGND 0.01243f
C14493 XThC.XTBN.Y.t11 VGND 0.00603f
C14494 XThC.XTBN.Y.t86 VGND 0.01024f
C14495 XThC.XTBN.Y.n152 VGND 0.01348f
C14496 XThC.XTBN.Y.n153 VGND 0.0076f
C14497 XThC.XTBN.Y.n154 VGND 0.01252f
C14498 XThC.XTBN.Y.n155 VGND 0.00434f
C14499 XThC.XTBN.Y.n156 VGND 0.00603f
C14500 XThC.XTBN.Y.n157 VGND 0.01348f
C14501 XThC.XTBN.Y.t53 VGND 0.00603f
C14502 XThC.XTBN.Y.t13 VGND 0.01024f
C14503 XThC.XTBN.Y.n158 VGND 0.01227f
C14504 XThC.XTBN.Y.n159 VGND 0.00676f
C14505 XThC.XTBN.Y.n160 VGND 0.00747f
C14506 XThC.XTBN.Y.n161 VGND 0.07521f
C14507 XThC.XTBN.Y.t23 VGND 0.01024f
C14508 XThC.XTBN.Y.t117 VGND 0.00603f
C14509 XThC.XTBN.Y.n162 VGND 0.00619f
C14510 XThC.XTBN.Y.t95 VGND 0.01024f
C14511 XThC.XTBN.Y.t78 VGND 0.00603f
C14512 XThC.XTBN.Y.n163 VGND 0.01243f
C14513 XThC.XTBN.Y.t97 VGND 0.01024f
C14514 XThC.XTBN.Y.t80 VGND 0.00603f
C14515 XThC.XTBN.Y.n164 VGND 0.01348f
C14516 XThC.XTBN.Y.n165 VGND 0.0076f
C14517 XThC.XTBN.Y.n166 VGND 0.01252f
C14518 XThC.XTBN.Y.n167 VGND 0.00434f
C14519 XThC.XTBN.Y.n168 VGND 0.00603f
C14520 XThC.XTBN.Y.n169 VGND 0.01348f
C14521 XThC.XTBN.Y.t28 VGND 0.01024f
C14522 XThC.XTBN.Y.t4 VGND 0.00603f
C14523 XThC.XTBN.Y.n170 VGND 0.01227f
C14524 XThC.XTBN.Y.n171 VGND 0.00676f
C14525 XThC.XTBN.Y.n172 VGND 0.00747f
C14526 XThC.XTBN.Y.n173 VGND 0.08751f
C14527 XThC.XTBN.Y.n174 VGND 0.11019f
C14528 XThC.XTBN.Y.t105 VGND 0.00603f
C14529 XThC.XTBN.Y.t75 VGND 0.01024f
C14530 XThC.XTBN.Y.t69 VGND 0.00603f
C14531 XThC.XTBN.Y.t33 VGND 0.01024f
C14532 XThC.XTBN.Y.n175 VGND 0.01477f
C14533 XThC.XTBN.Y.t61 VGND 0.00603f
C14534 XThC.XTBN.Y.t27 VGND 0.01024f
C14535 XThC.XTBN.Y.n176 VGND 0.02293f
C14536 XThC.XTBN.Y.n177 VGND 0.00676f
C14537 XThC.XTBN.Y.n178 VGND 0.00561f
C14538 XThC.XTBN.Y.n179 VGND 0.00561f
C14539 XThC.XTBN.Y.n180 VGND 0.00676f
C14540 XThC.XTBN.Y.n181 VGND 0.01477f
C14541 XThC.XTBN.Y.t14 VGND 0.00603f
C14542 XThC.XTBN.Y.t9 VGND 0.01024f
C14543 XThC.XTBN.Y.n182 VGND 0.0138f
C14544 XThC.XTBN.Y.n183 VGND 0.00676f
C14545 XThC.XTBN.Y.n184 VGND 0.00372f
C14546 XThC.XTBN.Y.n185 VGND 0.00408f
C14547 XThC.XTBN.Y.n186 VGND 0.11129f
C14548 XThC.XTBN.Y.n187 VGND 0.02169f
C14549 XThC.XTBN.Y.t3 VGND 0.00428f
C14550 XThC.XTBN.Y.t2 VGND 0.00428f
C14551 XThC.XTBN.Y.n188 VGND 0.0094f
C14552 XThC.XTBN.Y.n189 VGND 0.00607f
C14553 XThC.XTBN.Y.n190 VGND 0.00526f
C14554 XThC.XTBN.Y.t0 VGND 0.00658f
C14555 XThC.XTBN.Y.t1 VGND 0.00658f
C14556 XThC.XTBN.Y.n191 VGND 0.01513f
C14557 XThC.XTBN.Y.n192 VGND 0.0307f
C14558 XThR.Tn[12].t11 VGND 0.02425f
C14559 XThR.Tn[12].t9 VGND 0.02425f
C14560 XThR.Tn[12].n0 VGND 0.07362f
C14561 XThR.Tn[12].t8 VGND 0.02425f
C14562 XThR.Tn[12].t10 VGND 0.02425f
C14563 XThR.Tn[12].n1 VGND 0.0539f
C14564 XThR.Tn[12].n2 VGND 0.24508f
C14565 XThR.Tn[12].t7 VGND 0.01576f
C14566 XThR.Tn[12].t5 VGND 0.01576f
C14567 XThR.Tn[12].n3 VGND 0.03931f
C14568 XThR.Tn[12].t6 VGND 0.01576f
C14569 XThR.Tn[12].t4 VGND 0.01576f
C14570 XThR.Tn[12].n4 VGND 0.03152f
C14571 XThR.Tn[12].n5 VGND 0.07268f
C14572 XThR.Tn[12].t36 VGND 0.01895f
C14573 XThR.Tn[12].t28 VGND 0.02075f
C14574 XThR.Tn[12].n6 VGND 0.05067f
C14575 XThR.Tn[12].n7 VGND 0.09734f
C14576 XThR.Tn[12].t53 VGND 0.01895f
C14577 XThR.Tn[12].t43 VGND 0.02075f
C14578 XThR.Tn[12].n8 VGND 0.05067f
C14579 XThR.Tn[12].t71 VGND 0.01889f
C14580 XThR.Tn[12].t21 VGND 0.02068f
C14581 XThR.Tn[12].n9 VGND 0.05272f
C14582 XThR.Tn[12].n10 VGND 0.03704f
C14583 XThR.Tn[12].n11 VGND 0.00677f
C14584 XThR.Tn[12].n12 VGND 0.11886f
C14585 XThR.Tn[12].t30 VGND 0.01895f
C14586 XThR.Tn[12].t20 VGND 0.02075f
C14587 XThR.Tn[12].n13 VGND 0.05067f
C14588 XThR.Tn[12].t49 VGND 0.01889f
C14589 XThR.Tn[12].t60 VGND 0.02068f
C14590 XThR.Tn[12].n14 VGND 0.05272f
C14591 XThR.Tn[12].n15 VGND 0.03704f
C14592 XThR.Tn[12].n16 VGND 0.00677f
C14593 XThR.Tn[12].n17 VGND 0.11886f
C14594 XThR.Tn[12].t45 VGND 0.01895f
C14595 XThR.Tn[12].t38 VGND 0.02075f
C14596 XThR.Tn[12].n18 VGND 0.05067f
C14597 XThR.Tn[12].t63 VGND 0.01889f
C14598 XThR.Tn[12].t15 VGND 0.02068f
C14599 XThR.Tn[12].n19 VGND 0.05272f
C14600 XThR.Tn[12].n20 VGND 0.03704f
C14601 XThR.Tn[12].n21 VGND 0.00677f
C14602 XThR.Tn[12].n22 VGND 0.11886f
C14603 XThR.Tn[12].t70 VGND 0.01895f
C14604 XThR.Tn[12].t66 VGND 0.02075f
C14605 XThR.Tn[12].n23 VGND 0.05067f
C14606 XThR.Tn[12].t33 VGND 0.01889f
C14607 XThR.Tn[12].t46 VGND 0.02068f
C14608 XThR.Tn[12].n24 VGND 0.05272f
C14609 XThR.Tn[12].n25 VGND 0.03704f
C14610 XThR.Tn[12].n26 VGND 0.00677f
C14611 XThR.Tn[12].n27 VGND 0.11886f
C14612 XThR.Tn[12].t48 VGND 0.01895f
C14613 XThR.Tn[12].t39 VGND 0.02075f
C14614 XThR.Tn[12].n28 VGND 0.05067f
C14615 XThR.Tn[12].t64 VGND 0.01889f
C14616 XThR.Tn[12].t17 VGND 0.02068f
C14617 XThR.Tn[12].n29 VGND 0.05272f
C14618 XThR.Tn[12].n30 VGND 0.03704f
C14619 XThR.Tn[12].n31 VGND 0.00677f
C14620 XThR.Tn[12].n32 VGND 0.11886f
C14621 XThR.Tn[12].t23 VGND 0.01895f
C14622 XThR.Tn[12].t56 VGND 0.02075f
C14623 XThR.Tn[12].n33 VGND 0.05067f
C14624 XThR.Tn[12].t41 VGND 0.01889f
C14625 XThR.Tn[12].t37 VGND 0.02068f
C14626 XThR.Tn[12].n34 VGND 0.05272f
C14627 XThR.Tn[12].n35 VGND 0.03704f
C14628 XThR.Tn[12].n36 VGND 0.00677f
C14629 XThR.Tn[12].n37 VGND 0.11886f
C14630 XThR.Tn[12].t54 VGND 0.01895f
C14631 XThR.Tn[12].t51 VGND 0.02075f
C14632 XThR.Tn[12].n38 VGND 0.05067f
C14633 XThR.Tn[12].t72 VGND 0.01889f
C14634 XThR.Tn[12].t29 VGND 0.02068f
C14635 XThR.Tn[12].n39 VGND 0.05272f
C14636 XThR.Tn[12].n40 VGND 0.03704f
C14637 XThR.Tn[12].n41 VGND 0.00677f
C14638 XThR.Tn[12].n42 VGND 0.11886f
C14639 XThR.Tn[12].t59 VGND 0.01895f
C14640 XThR.Tn[12].t65 VGND 0.02075f
C14641 XThR.Tn[12].n43 VGND 0.05067f
C14642 XThR.Tn[12].t14 VGND 0.01889f
C14643 XThR.Tn[12].t44 VGND 0.02068f
C14644 XThR.Tn[12].n44 VGND 0.05272f
C14645 XThR.Tn[12].n45 VGND 0.03704f
C14646 XThR.Tn[12].n46 VGND 0.00677f
C14647 XThR.Tn[12].n47 VGND 0.11886f
C14648 XThR.Tn[12].t12 VGND 0.01895f
C14649 XThR.Tn[12].t22 VGND 0.02075f
C14650 XThR.Tn[12].n48 VGND 0.05067f
C14651 XThR.Tn[12].t35 VGND 0.01889f
C14652 XThR.Tn[12].t61 VGND 0.02068f
C14653 XThR.Tn[12].n49 VGND 0.05272f
C14654 XThR.Tn[12].n50 VGND 0.03704f
C14655 XThR.Tn[12].n51 VGND 0.00677f
C14656 XThR.Tn[12].n52 VGND 0.11886f
C14657 XThR.Tn[12].t68 VGND 0.01895f
C14658 XThR.Tn[12].t40 VGND 0.02075f
C14659 XThR.Tn[12].n53 VGND 0.05067f
C14660 XThR.Tn[12].t26 VGND 0.01889f
C14661 XThR.Tn[12].t19 VGND 0.02068f
C14662 XThR.Tn[12].n54 VGND 0.05272f
C14663 XThR.Tn[12].n55 VGND 0.03704f
C14664 XThR.Tn[12].n56 VGND 0.00677f
C14665 XThR.Tn[12].n57 VGND 0.11886f
C14666 XThR.Tn[12].t25 VGND 0.01895f
C14667 XThR.Tn[12].t16 VGND 0.02075f
C14668 XThR.Tn[12].n58 VGND 0.05067f
C14669 XThR.Tn[12].t42 VGND 0.01889f
C14670 XThR.Tn[12].t55 VGND 0.02068f
C14671 XThR.Tn[12].n59 VGND 0.05272f
C14672 XThR.Tn[12].n60 VGND 0.03704f
C14673 XThR.Tn[12].n61 VGND 0.00677f
C14674 XThR.Tn[12].n62 VGND 0.11886f
C14675 XThR.Tn[12].t57 VGND 0.01895f
C14676 XThR.Tn[12].t52 VGND 0.02075f
C14677 XThR.Tn[12].n63 VGND 0.05067f
C14678 XThR.Tn[12].t13 VGND 0.01889f
C14679 XThR.Tn[12].t31 VGND 0.02068f
C14680 XThR.Tn[12].n64 VGND 0.05272f
C14681 XThR.Tn[12].n65 VGND 0.03704f
C14682 XThR.Tn[12].n66 VGND 0.00677f
C14683 XThR.Tn[12].n67 VGND 0.11886f
C14684 XThR.Tn[12].t73 VGND 0.01895f
C14685 XThR.Tn[12].t67 VGND 0.02075f
C14686 XThR.Tn[12].n68 VGND 0.05067f
C14687 XThR.Tn[12].t34 VGND 0.01889f
C14688 XThR.Tn[12].t47 VGND 0.02068f
C14689 XThR.Tn[12].n69 VGND 0.05272f
C14690 XThR.Tn[12].n70 VGND 0.03704f
C14691 XThR.Tn[12].n71 VGND 0.00677f
C14692 XThR.Tn[12].n72 VGND 0.11886f
C14693 XThR.Tn[12].t32 VGND 0.01895f
C14694 XThR.Tn[12].t24 VGND 0.02075f
C14695 XThR.Tn[12].n73 VGND 0.05067f
C14696 XThR.Tn[12].t50 VGND 0.01889f
C14697 XThR.Tn[12].t62 VGND 0.02068f
C14698 XThR.Tn[12].n74 VGND 0.05272f
C14699 XThR.Tn[12].n75 VGND 0.03704f
C14700 XThR.Tn[12].n76 VGND 0.00677f
C14701 XThR.Tn[12].n77 VGND 0.11886f
C14702 XThR.Tn[12].t69 VGND 0.01895f
C14703 XThR.Tn[12].t18 VGND 0.02075f
C14704 XThR.Tn[12].n78 VGND 0.05067f
C14705 XThR.Tn[12].t27 VGND 0.01889f
C14706 XThR.Tn[12].t58 VGND 0.02068f
C14707 XThR.Tn[12].n79 VGND 0.05272f
C14708 XThR.Tn[12].n80 VGND 0.03704f
C14709 XThR.Tn[12].n81 VGND 0.00677f
C14710 XThR.Tn[12].n82 VGND 0.11886f
C14711 XThR.Tn[12].n83 VGND 0.10802f
C14712 XThR.Tn[12].n84 VGND 0.36839f
C14713 XThR.Tn[12].t2 VGND 0.02425f
C14714 XThR.Tn[12].t0 VGND 0.02425f
C14715 XThR.Tn[12].n85 VGND 0.05239f
C14716 XThR.Tn[12].t3 VGND 0.02425f
C14717 XThR.Tn[12].t1 VGND 0.02425f
C14718 XThR.Tn[12].n86 VGND 0.07973f
C14719 XThR.Tn[12].n87 VGND 0.2214f
C14720 XThR.Tn[12].n88 VGND 0.01091f
C14721 XThR.Tn[14].t8 VGND 0.02436f
C14722 XThR.Tn[14].t9 VGND 0.02436f
C14723 XThR.Tn[14].n0 VGND 0.07395f
C14724 XThR.Tn[14].t10 VGND 0.02436f
C14725 XThR.Tn[14].t11 VGND 0.02436f
C14726 XThR.Tn[14].n1 VGND 0.05414f
C14727 XThR.Tn[14].n2 VGND 0.24618f
C14728 XThR.Tn[14].t6 VGND 0.01583f
C14729 XThR.Tn[14].t7 VGND 0.01583f
C14730 XThR.Tn[14].n3 VGND 0.03948f
C14731 XThR.Tn[14].t4 VGND 0.01583f
C14732 XThR.Tn[14].t5 VGND 0.01583f
C14733 XThR.Tn[14].n4 VGND 0.03166f
C14734 XThR.Tn[14].n5 VGND 0.07301f
C14735 XThR.Tn[14].t69 VGND 0.01904f
C14736 XThR.Tn[14].t62 VGND 0.02084f
C14737 XThR.Tn[14].n6 VGND 0.0509f
C14738 XThR.Tn[14].n7 VGND 0.09778f
C14739 XThR.Tn[14].t24 VGND 0.01904f
C14740 XThR.Tn[14].t13 VGND 0.02084f
C14741 XThR.Tn[14].n8 VGND 0.0509f
C14742 XThR.Tn[14].t28 VGND 0.01897f
C14743 XThR.Tn[14].t60 VGND 0.02078f
C14744 XThR.Tn[14].n9 VGND 0.05296f
C14745 XThR.Tn[14].n10 VGND 0.03721f
C14746 XThR.Tn[14].n11 VGND 0.0068f
C14747 XThR.Tn[14].n12 VGND 0.11939f
C14748 XThR.Tn[14].t64 VGND 0.01904f
C14749 XThR.Tn[14].t54 VGND 0.02084f
C14750 XThR.Tn[14].n13 VGND 0.0509f
C14751 XThR.Tn[14].t67 VGND 0.01897f
C14752 XThR.Tn[14].t34 VGND 0.02078f
C14753 XThR.Tn[14].n14 VGND 0.05296f
C14754 XThR.Tn[14].n15 VGND 0.03721f
C14755 XThR.Tn[14].n16 VGND 0.0068f
C14756 XThR.Tn[14].n17 VGND 0.11939f
C14757 XThR.Tn[14].t14 VGND 0.01904f
C14758 XThR.Tn[14].t72 VGND 0.02084f
C14759 XThR.Tn[14].n18 VGND 0.0509f
C14760 XThR.Tn[14].t17 VGND 0.01897f
C14761 XThR.Tn[14].t52 VGND 0.02078f
C14762 XThR.Tn[14].n19 VGND 0.05296f
C14763 XThR.Tn[14].n20 VGND 0.03721f
C14764 XThR.Tn[14].n21 VGND 0.0068f
C14765 XThR.Tn[14].n22 VGND 0.11939f
C14766 XThR.Tn[14].t44 VGND 0.01904f
C14767 XThR.Tn[14].t38 VGND 0.02084f
C14768 XThR.Tn[14].n23 VGND 0.0509f
C14769 XThR.Tn[14].t47 VGND 0.01897f
C14770 XThR.Tn[14].t18 VGND 0.02078f
C14771 XThR.Tn[14].n24 VGND 0.05296f
C14772 XThR.Tn[14].n25 VGND 0.03721f
C14773 XThR.Tn[14].n26 VGND 0.0068f
C14774 XThR.Tn[14].n27 VGND 0.11939f
C14775 XThR.Tn[14].t15 VGND 0.01904f
C14776 XThR.Tn[14].t73 VGND 0.02084f
C14777 XThR.Tn[14].n28 VGND 0.0509f
C14778 XThR.Tn[14].t21 VGND 0.01897f
C14779 XThR.Tn[14].t53 VGND 0.02078f
C14780 XThR.Tn[14].n29 VGND 0.05296f
C14781 XThR.Tn[14].n30 VGND 0.03721f
C14782 XThR.Tn[14].n31 VGND 0.0068f
C14783 XThR.Tn[14].n32 VGND 0.11939f
C14784 XThR.Tn[14].t57 VGND 0.01904f
C14785 XThR.Tn[14].t25 VGND 0.02084f
C14786 XThR.Tn[14].n33 VGND 0.0509f
C14787 XThR.Tn[14].t61 VGND 0.01897f
C14788 XThR.Tn[14].t71 VGND 0.02078f
C14789 XThR.Tn[14].n34 VGND 0.05296f
C14790 XThR.Tn[14].n35 VGND 0.03721f
C14791 XThR.Tn[14].n36 VGND 0.0068f
C14792 XThR.Tn[14].n37 VGND 0.11939f
C14793 XThR.Tn[14].t23 VGND 0.01904f
C14794 XThR.Tn[14].t19 VGND 0.02084f
C14795 XThR.Tn[14].n38 VGND 0.0509f
C14796 XThR.Tn[14].t29 VGND 0.01897f
C14797 XThR.Tn[14].t66 VGND 0.02078f
C14798 XThR.Tn[14].n39 VGND 0.05296f
C14799 XThR.Tn[14].n40 VGND 0.03721f
C14800 XThR.Tn[14].n41 VGND 0.0068f
C14801 XThR.Tn[14].n42 VGND 0.11939f
C14802 XThR.Tn[14].t27 VGND 0.01904f
C14803 XThR.Tn[14].t36 VGND 0.02084f
C14804 XThR.Tn[14].n43 VGND 0.0509f
C14805 XThR.Tn[14].t33 VGND 0.01897f
C14806 XThR.Tn[14].t16 VGND 0.02078f
C14807 XThR.Tn[14].n44 VGND 0.05296f
C14808 XThR.Tn[14].n45 VGND 0.03721f
C14809 XThR.Tn[14].n46 VGND 0.0068f
C14810 XThR.Tn[14].n47 VGND 0.11939f
C14811 XThR.Tn[14].t46 VGND 0.01904f
C14812 XThR.Tn[14].t56 VGND 0.02084f
C14813 XThR.Tn[14].n48 VGND 0.0509f
C14814 XThR.Tn[14].t50 VGND 0.01897f
C14815 XThR.Tn[14].t35 VGND 0.02078f
C14816 XThR.Tn[14].n49 VGND 0.05296f
C14817 XThR.Tn[14].n50 VGND 0.03721f
C14818 XThR.Tn[14].n51 VGND 0.0068f
C14819 XThR.Tn[14].n52 VGND 0.11939f
C14820 XThR.Tn[14].t40 VGND 0.01904f
C14821 XThR.Tn[14].t12 VGND 0.02084f
C14822 XThR.Tn[14].n53 VGND 0.0509f
C14823 XThR.Tn[14].t42 VGND 0.01897f
C14824 XThR.Tn[14].t55 VGND 0.02078f
C14825 XThR.Tn[14].n54 VGND 0.05296f
C14826 XThR.Tn[14].n55 VGND 0.03721f
C14827 XThR.Tn[14].n56 VGND 0.0068f
C14828 XThR.Tn[14].n57 VGND 0.11939f
C14829 XThR.Tn[14].t59 VGND 0.01904f
C14830 XThR.Tn[14].t49 VGND 0.02084f
C14831 XThR.Tn[14].n58 VGND 0.0509f
C14832 XThR.Tn[14].t63 VGND 0.01897f
C14833 XThR.Tn[14].t30 VGND 0.02078f
C14834 XThR.Tn[14].n59 VGND 0.05296f
C14835 XThR.Tn[14].n60 VGND 0.03721f
C14836 XThR.Tn[14].n61 VGND 0.0068f
C14837 XThR.Tn[14].n62 VGND 0.11939f
C14838 XThR.Tn[14].t26 VGND 0.01904f
C14839 XThR.Tn[14].t22 VGND 0.02084f
C14840 XThR.Tn[14].n63 VGND 0.0509f
C14841 XThR.Tn[14].t31 VGND 0.01897f
C14842 XThR.Tn[14].t68 VGND 0.02078f
C14843 XThR.Tn[14].n64 VGND 0.05296f
C14844 XThR.Tn[14].n65 VGND 0.03721f
C14845 XThR.Tn[14].n66 VGND 0.0068f
C14846 XThR.Tn[14].n67 VGND 0.11939f
C14847 XThR.Tn[14].t45 VGND 0.01904f
C14848 XThR.Tn[14].t39 VGND 0.02084f
C14849 XThR.Tn[14].n68 VGND 0.0509f
C14850 XThR.Tn[14].t48 VGND 0.01897f
C14851 XThR.Tn[14].t20 VGND 0.02078f
C14852 XThR.Tn[14].n69 VGND 0.05296f
C14853 XThR.Tn[14].n70 VGND 0.03721f
C14854 XThR.Tn[14].n71 VGND 0.0068f
C14855 XThR.Tn[14].n72 VGND 0.11939f
C14856 XThR.Tn[14].t65 VGND 0.01904f
C14857 XThR.Tn[14].t58 VGND 0.02084f
C14858 XThR.Tn[14].n73 VGND 0.0509f
C14859 XThR.Tn[14].t70 VGND 0.01897f
C14860 XThR.Tn[14].t37 VGND 0.02078f
C14861 XThR.Tn[14].n74 VGND 0.05296f
C14862 XThR.Tn[14].n75 VGND 0.03721f
C14863 XThR.Tn[14].n76 VGND 0.0068f
C14864 XThR.Tn[14].n77 VGND 0.11939f
C14865 XThR.Tn[14].t41 VGND 0.01904f
C14866 XThR.Tn[14].t51 VGND 0.02084f
C14867 XThR.Tn[14].n78 VGND 0.0509f
C14868 XThR.Tn[14].t43 VGND 0.01897f
C14869 XThR.Tn[14].t32 VGND 0.02078f
C14870 XThR.Tn[14].n79 VGND 0.05296f
C14871 XThR.Tn[14].n80 VGND 0.03721f
C14872 XThR.Tn[14].n81 VGND 0.0068f
C14873 XThR.Tn[14].n82 VGND 0.11939f
C14874 XThR.Tn[14].n83 VGND 0.1085f
C14875 XThR.Tn[14].n84 VGND 0.43586f
C14876 XThR.Tn[14].t2 VGND 0.02436f
C14877 XThR.Tn[14].t3 VGND 0.02436f
C14878 XThR.Tn[14].n85 VGND 0.05262f
C14879 XThR.Tn[14].t0 VGND 0.02436f
C14880 XThR.Tn[14].t1 VGND 0.02436f
C14881 XThR.Tn[14].n86 VGND 0.08009f
C14882 XThR.Tn[14].n87 VGND 0.22239f
C14883 XThR.Tn[14].n88 VGND 0.01096f
C14884 XThR.Tn[6].t7 VGND 0.02335f
C14885 XThR.Tn[6].t4 VGND 0.02335f
C14886 XThR.Tn[6].n0 VGND 0.04712f
C14887 XThR.Tn[6].t6 VGND 0.02335f
C14888 XThR.Tn[6].t5 VGND 0.02335f
C14889 XThR.Tn[6].n1 VGND 0.05514f
C14890 XThR.Tn[6].n2 VGND 0.16538f
C14891 XThR.Tn[6].t8 VGND 0.01517f
C14892 XThR.Tn[6].t9 VGND 0.01517f
C14893 XThR.Tn[6].n3 VGND 0.03456f
C14894 XThR.Tn[6].t11 VGND 0.01517f
C14895 XThR.Tn[6].t10 VGND 0.01517f
C14896 XThR.Tn[6].n4 VGND 0.03456f
C14897 XThR.Tn[6].t0 VGND 0.01517f
C14898 XThR.Tn[6].t1 VGND 0.01517f
C14899 XThR.Tn[6].n5 VGND 0.05758f
C14900 XThR.Tn[6].t3 VGND 0.01517f
C14901 XThR.Tn[6].t2 VGND 0.01517f
C14902 XThR.Tn[6].n6 VGND 0.03456f
C14903 XThR.Tn[6].n7 VGND 0.16456f
C14904 XThR.Tn[6].n8 VGND 0.10173f
C14905 XThR.Tn[6].n9 VGND 0.11481f
C14906 XThR.Tn[6].t62 VGND 0.01825f
C14907 XThR.Tn[6].t56 VGND 0.01998f
C14908 XThR.Tn[6].n10 VGND 0.04879f
C14909 XThR.Tn[6].n11 VGND 0.09372f
C14910 XThR.Tn[6].t20 VGND 0.01825f
C14911 XThR.Tn[6].t72 VGND 0.01998f
C14912 XThR.Tn[6].n12 VGND 0.04879f
C14913 XThR.Tn[6].t36 VGND 0.01819f
C14914 XThR.Tn[6].t68 VGND 0.01991f
C14915 XThR.Tn[6].n13 VGND 0.05076f
C14916 XThR.Tn[6].n14 VGND 0.03566f
C14917 XThR.Tn[6].n15 VGND 0.00652f
C14918 XThR.Tn[6].n16 VGND 0.11444f
C14919 XThR.Tn[6].t57 VGND 0.01825f
C14920 XThR.Tn[6].t49 VGND 0.01998f
C14921 XThR.Tn[6].n17 VGND 0.04879f
C14922 XThR.Tn[6].t14 VGND 0.01819f
C14923 XThR.Tn[6].t45 VGND 0.01991f
C14924 XThR.Tn[6].n18 VGND 0.05076f
C14925 XThR.Tn[6].n19 VGND 0.03566f
C14926 XThR.Tn[6].n20 VGND 0.00652f
C14927 XThR.Tn[6].n21 VGND 0.11444f
C14928 XThR.Tn[6].t73 VGND 0.01825f
C14929 XThR.Tn[6].t66 VGND 0.01998f
C14930 XThR.Tn[6].n22 VGND 0.04879f
C14931 XThR.Tn[6].t26 VGND 0.01819f
C14932 XThR.Tn[6].t63 VGND 0.01991f
C14933 XThR.Tn[6].n23 VGND 0.05076f
C14934 XThR.Tn[6].n24 VGND 0.03566f
C14935 XThR.Tn[6].n25 VGND 0.00652f
C14936 XThR.Tn[6].n26 VGND 0.11444f
C14937 XThR.Tn[6].t35 VGND 0.01825f
C14938 XThR.Tn[6].t31 VGND 0.01998f
C14939 XThR.Tn[6].n27 VGND 0.04879f
C14940 XThR.Tn[6].t59 VGND 0.01819f
C14941 XThR.Tn[6].t27 VGND 0.01991f
C14942 XThR.Tn[6].n28 VGND 0.05076f
C14943 XThR.Tn[6].n29 VGND 0.03566f
C14944 XThR.Tn[6].n30 VGND 0.00652f
C14945 XThR.Tn[6].n31 VGND 0.11444f
C14946 XThR.Tn[6].t13 VGND 0.01825f
C14947 XThR.Tn[6].t67 VGND 0.01998f
C14948 XThR.Tn[6].n32 VGND 0.04879f
C14949 XThR.Tn[6].t29 VGND 0.01819f
C14950 XThR.Tn[6].t64 VGND 0.01991f
C14951 XThR.Tn[6].n33 VGND 0.05076f
C14952 XThR.Tn[6].n34 VGND 0.03566f
C14953 XThR.Tn[6].n35 VGND 0.00652f
C14954 XThR.Tn[6].n36 VGND 0.11444f
C14955 XThR.Tn[6].t51 VGND 0.01825f
C14956 XThR.Tn[6].t22 VGND 0.01998f
C14957 XThR.Tn[6].n37 VGND 0.04879f
C14958 XThR.Tn[6].t70 VGND 0.01819f
C14959 XThR.Tn[6].t19 VGND 0.01991f
C14960 XThR.Tn[6].n38 VGND 0.05076f
C14961 XThR.Tn[6].n39 VGND 0.03566f
C14962 XThR.Tn[6].n40 VGND 0.00652f
C14963 XThR.Tn[6].n41 VGND 0.11444f
C14964 XThR.Tn[6].t21 VGND 0.01825f
C14965 XThR.Tn[6].t17 VGND 0.01998f
C14966 XThR.Tn[6].n42 VGND 0.04879f
C14967 XThR.Tn[6].t37 VGND 0.01819f
C14968 XThR.Tn[6].t12 VGND 0.01991f
C14969 XThR.Tn[6].n43 VGND 0.05076f
C14970 XThR.Tn[6].n44 VGND 0.03566f
C14971 XThR.Tn[6].n45 VGND 0.00652f
C14972 XThR.Tn[6].n46 VGND 0.11444f
C14973 XThR.Tn[6].t24 VGND 0.01825f
C14974 XThR.Tn[6].t30 VGND 0.01998f
C14975 XThR.Tn[6].n47 VGND 0.04879f
C14976 XThR.Tn[6].t43 VGND 0.01819f
C14977 XThR.Tn[6].t25 VGND 0.01991f
C14978 XThR.Tn[6].n48 VGND 0.05076f
C14979 XThR.Tn[6].n49 VGND 0.03566f
C14980 XThR.Tn[6].n50 VGND 0.00652f
C14981 XThR.Tn[6].n51 VGND 0.11444f
C14982 XThR.Tn[6].t40 VGND 0.01825f
C14983 XThR.Tn[6].t50 VGND 0.01998f
C14984 XThR.Tn[6].n52 VGND 0.04879f
C14985 XThR.Tn[6].t61 VGND 0.01819f
C14986 XThR.Tn[6].t47 VGND 0.01991f
C14987 XThR.Tn[6].n53 VGND 0.05076f
C14988 XThR.Tn[6].n54 VGND 0.03566f
C14989 XThR.Tn[6].n55 VGND 0.00652f
C14990 XThR.Tn[6].n56 VGND 0.11444f
C14991 XThR.Tn[6].t33 VGND 0.01825f
C14992 XThR.Tn[6].t69 VGND 0.01998f
C14993 XThR.Tn[6].n57 VGND 0.04879f
C14994 XThR.Tn[6].t54 VGND 0.01819f
C14995 XThR.Tn[6].t65 VGND 0.01991f
C14996 XThR.Tn[6].n58 VGND 0.05076f
C14997 XThR.Tn[6].n59 VGND 0.03566f
C14998 XThR.Tn[6].n60 VGND 0.00652f
C14999 XThR.Tn[6].n61 VGND 0.11444f
C15000 XThR.Tn[6].t53 VGND 0.01825f
C15001 XThR.Tn[6].t44 VGND 0.01998f
C15002 XThR.Tn[6].n62 VGND 0.04879f
C15003 XThR.Tn[6].t71 VGND 0.01819f
C15004 XThR.Tn[6].t39 VGND 0.01991f
C15005 XThR.Tn[6].n63 VGND 0.05076f
C15006 XThR.Tn[6].n64 VGND 0.03566f
C15007 XThR.Tn[6].n65 VGND 0.00652f
C15008 XThR.Tn[6].n66 VGND 0.11444f
C15009 XThR.Tn[6].t23 VGND 0.01825f
C15010 XThR.Tn[6].t18 VGND 0.01998f
C15011 XThR.Tn[6].n67 VGND 0.04879f
C15012 XThR.Tn[6].t41 VGND 0.01819f
C15013 XThR.Tn[6].t15 VGND 0.01991f
C15014 XThR.Tn[6].n68 VGND 0.05076f
C15015 XThR.Tn[6].n69 VGND 0.03566f
C15016 XThR.Tn[6].n70 VGND 0.00652f
C15017 XThR.Tn[6].n71 VGND 0.11444f
C15018 XThR.Tn[6].t38 VGND 0.01825f
C15019 XThR.Tn[6].t32 VGND 0.01998f
C15020 XThR.Tn[6].n72 VGND 0.04879f
C15021 XThR.Tn[6].t60 VGND 0.01819f
C15022 XThR.Tn[6].t28 VGND 0.01991f
C15023 XThR.Tn[6].n73 VGND 0.05076f
C15024 XThR.Tn[6].n74 VGND 0.03566f
C15025 XThR.Tn[6].n75 VGND 0.00652f
C15026 XThR.Tn[6].n76 VGND 0.11444f
C15027 XThR.Tn[6].t58 VGND 0.01825f
C15028 XThR.Tn[6].t52 VGND 0.01998f
C15029 XThR.Tn[6].n77 VGND 0.04879f
C15030 XThR.Tn[6].t16 VGND 0.01819f
C15031 XThR.Tn[6].t48 VGND 0.01991f
C15032 XThR.Tn[6].n78 VGND 0.05076f
C15033 XThR.Tn[6].n79 VGND 0.03566f
C15034 XThR.Tn[6].n80 VGND 0.00652f
C15035 XThR.Tn[6].n81 VGND 0.11444f
C15036 XThR.Tn[6].t34 VGND 0.01825f
C15037 XThR.Tn[6].t46 VGND 0.01998f
C15038 XThR.Tn[6].n82 VGND 0.04879f
C15039 XThR.Tn[6].t55 VGND 0.01819f
C15040 XThR.Tn[6].t42 VGND 0.01991f
C15041 XThR.Tn[6].n83 VGND 0.05076f
C15042 XThR.Tn[6].n84 VGND 0.03566f
C15043 XThR.Tn[6].n85 VGND 0.00652f
C15044 XThR.Tn[6].n86 VGND 0.11444f
C15045 XThR.Tn[6].n87 VGND 0.104f
C15046 XThR.Tn[6].n88 VGND 0.17311f
C15047 XThC.Tn[10].t4 VGND 0.01306f
C15048 XThC.Tn[10].t1 VGND 0.01306f
C15049 XThC.Tn[10].n0 VGND 0.03258f
C15050 XThC.Tn[10].t3 VGND 0.01306f
C15051 XThC.Tn[10].t5 VGND 0.01306f
C15052 XThC.Tn[10].n1 VGND 0.02613f
C15053 XThC.Tn[10].n2 VGND 0.06572f
C15054 XThC.Tn[10].n3 VGND 0.02851f
C15055 XThC.Tn[10].t38 VGND 0.01593f
C15056 XThC.Tn[10].t36 VGND 0.0174f
C15057 XThC.Tn[10].n4 VGND 0.03884f
C15058 XThC.Tn[10].n5 VGND 0.02661f
C15059 XThC.Tn[10].n6 VGND 0.08734f
C15060 XThC.Tn[10].t24 VGND 0.01593f
C15061 XThC.Tn[10].t21 VGND 0.0174f
C15062 XThC.Tn[10].n7 VGND 0.03884f
C15063 XThC.Tn[10].n8 VGND 0.02661f
C15064 XThC.Tn[10].n9 VGND 0.08758f
C15065 XThC.Tn[10].n10 VGND 0.14434f
C15066 XThC.Tn[10].t29 VGND 0.01593f
C15067 XThC.Tn[10].t23 VGND 0.0174f
C15068 XThC.Tn[10].n11 VGND 0.03884f
C15069 XThC.Tn[10].n12 VGND 0.02661f
C15070 XThC.Tn[10].n13 VGND 0.08758f
C15071 XThC.Tn[10].n14 VGND 0.14434f
C15072 XThC.Tn[10].t30 VGND 0.01593f
C15073 XThC.Tn[10].t25 VGND 0.0174f
C15074 XThC.Tn[10].n15 VGND 0.03884f
C15075 XThC.Tn[10].n16 VGND 0.02661f
C15076 XThC.Tn[10].n17 VGND 0.08758f
C15077 XThC.Tn[10].n18 VGND 0.14434f
C15078 XThC.Tn[10].t17 VGND 0.01593f
C15079 XThC.Tn[10].t14 VGND 0.0174f
C15080 XThC.Tn[10].n19 VGND 0.03884f
C15081 XThC.Tn[10].n20 VGND 0.02661f
C15082 XThC.Tn[10].n21 VGND 0.08758f
C15083 XThC.Tn[10].n22 VGND 0.14434f
C15084 XThC.Tn[10].t18 VGND 0.01593f
C15085 XThC.Tn[10].t15 VGND 0.0174f
C15086 XThC.Tn[10].n23 VGND 0.03884f
C15087 XThC.Tn[10].n24 VGND 0.02661f
C15088 XThC.Tn[10].n25 VGND 0.08758f
C15089 XThC.Tn[10].n26 VGND 0.14434f
C15090 XThC.Tn[10].t34 VGND 0.01593f
C15091 XThC.Tn[10].t28 VGND 0.0174f
C15092 XThC.Tn[10].n27 VGND 0.03884f
C15093 XThC.Tn[10].n28 VGND 0.02661f
C15094 XThC.Tn[10].n29 VGND 0.08758f
C15095 XThC.Tn[10].n30 VGND 0.14434f
C15096 XThC.Tn[10].t41 VGND 0.01593f
C15097 XThC.Tn[10].t37 VGND 0.0174f
C15098 XThC.Tn[10].n31 VGND 0.03884f
C15099 XThC.Tn[10].n32 VGND 0.02661f
C15100 XThC.Tn[10].n33 VGND 0.08758f
C15101 XThC.Tn[10].n34 VGND 0.14434f
C15102 XThC.Tn[10].t43 VGND 0.01593f
C15103 XThC.Tn[10].t39 VGND 0.0174f
C15104 XThC.Tn[10].n35 VGND 0.03884f
C15105 XThC.Tn[10].n36 VGND 0.02661f
C15106 XThC.Tn[10].n37 VGND 0.08758f
C15107 XThC.Tn[10].n38 VGND 0.14434f
C15108 XThC.Tn[10].t31 VGND 0.01593f
C15109 XThC.Tn[10].t26 VGND 0.0174f
C15110 XThC.Tn[10].n39 VGND 0.03884f
C15111 XThC.Tn[10].n40 VGND 0.02661f
C15112 XThC.Tn[10].n41 VGND 0.08758f
C15113 XThC.Tn[10].n42 VGND 0.14434f
C15114 XThC.Tn[10].t33 VGND 0.01593f
C15115 XThC.Tn[10].t27 VGND 0.0174f
C15116 XThC.Tn[10].n43 VGND 0.03884f
C15117 XThC.Tn[10].n44 VGND 0.02661f
C15118 XThC.Tn[10].n45 VGND 0.08758f
C15119 XThC.Tn[10].n46 VGND 0.14434f
C15120 XThC.Tn[10].t12 VGND 0.01593f
C15121 XThC.Tn[10].t40 VGND 0.0174f
C15122 XThC.Tn[10].n47 VGND 0.03884f
C15123 XThC.Tn[10].n48 VGND 0.02661f
C15124 XThC.Tn[10].n49 VGND 0.08758f
C15125 XThC.Tn[10].n50 VGND 0.14434f
C15126 XThC.Tn[10].t20 VGND 0.01593f
C15127 XThC.Tn[10].t16 VGND 0.0174f
C15128 XThC.Tn[10].n51 VGND 0.03884f
C15129 XThC.Tn[10].n52 VGND 0.02661f
C15130 XThC.Tn[10].n53 VGND 0.08758f
C15131 XThC.Tn[10].n54 VGND 0.14434f
C15132 XThC.Tn[10].t22 VGND 0.01593f
C15133 XThC.Tn[10].t19 VGND 0.0174f
C15134 XThC.Tn[10].n55 VGND 0.03884f
C15135 XThC.Tn[10].n56 VGND 0.02661f
C15136 XThC.Tn[10].n57 VGND 0.08758f
C15137 XThC.Tn[10].n58 VGND 0.14434f
C15138 XThC.Tn[10].t35 VGND 0.01593f
C15139 XThC.Tn[10].t32 VGND 0.0174f
C15140 XThC.Tn[10].n59 VGND 0.03884f
C15141 XThC.Tn[10].n60 VGND 0.02661f
C15142 XThC.Tn[10].n61 VGND 0.08758f
C15143 XThC.Tn[10].n62 VGND 0.14434f
C15144 XThC.Tn[10].t13 VGND 0.01593f
C15145 XThC.Tn[10].t42 VGND 0.0174f
C15146 XThC.Tn[10].n63 VGND 0.03884f
C15147 XThC.Tn[10].n64 VGND 0.02661f
C15148 XThC.Tn[10].n65 VGND 0.08758f
C15149 XThC.Tn[10].n66 VGND 0.14434f
C15150 XThC.Tn[10].n67 VGND 0.61921f
C15151 XThC.Tn[10].n68 VGND 0.2357f
C15152 XThC.Tn[10].t7 VGND 0.0201f
C15153 XThC.Tn[10].t6 VGND 0.0201f
C15154 XThC.Tn[10].n69 VGND 0.04342f
C15155 XThC.Tn[10].t2 VGND 0.0201f
C15156 XThC.Tn[10].t10 VGND 0.0201f
C15157 XThC.Tn[10].n70 VGND 0.06609f
C15158 XThC.Tn[10].n71 VGND 0.18363f
C15159 XThC.Tn[10].n72 VGND 0.02887f
C15160 XThC.Tn[10].t8 VGND 0.0201f
C15161 XThC.Tn[10].t9 VGND 0.0201f
C15162 XThC.Tn[10].n73 VGND 0.04468f
C15163 XThC.Tn[10].t0 VGND 0.0201f
C15164 XThC.Tn[10].t11 VGND 0.0201f
C15165 XThC.Tn[10].n74 VGND 0.06102f
C15166 XThC.Tn[10].n75 VGND 0.19884f
C15167 Iout.n0 VGND 0.23929f
C15168 Iout.n1 VGND 1.25122f
C15169 Iout.n2 VGND 0.23929f
C15170 Iout.n3 VGND 0.23929f
C15171 Iout.t96 VGND 0.02304f
C15172 Iout.n4 VGND 0.05124f
C15173 Iout.n5 VGND 0.20242f
C15174 Iout.n6 VGND 0.23929f
C15175 Iout.n7 VGND 1.25122f
C15176 Iout.n8 VGND 0.23929f
C15177 Iout.t196 VGND 0.02304f
C15178 Iout.n9 VGND 0.05124f
C15179 Iout.n10 VGND 0.20242f
C15180 Iout.n11 VGND 0.23929f
C15181 Iout.n12 VGND 1.25122f
C15182 Iout.n13 VGND 0.23929f
C15183 Iout.t132 VGND 0.02304f
C15184 Iout.n14 VGND 0.05124f
C15185 Iout.n15 VGND 0.20242f
C15186 Iout.n16 VGND 0.23929f
C15187 Iout.n17 VGND 1.25122f
C15188 Iout.n18 VGND 0.23929f
C15189 Iout.t116 VGND 0.02304f
C15190 Iout.n19 VGND 0.05124f
C15191 Iout.n20 VGND 0.20242f
C15192 Iout.n21 VGND 0.49611f
C15193 Iout.t224 VGND 0.02304f
C15194 Iout.n22 VGND 0.05124f
C15195 Iout.n23 VGND 0.29851f
C15196 Iout.n24 VGND 0.23929f
C15197 Iout.n25 VGND 0.23929f
C15198 Iout.n26 VGND 0.23929f
C15199 Iout.n27 VGND 0.23929f
C15200 Iout.n28 VGND 0.23929f
C15201 Iout.n29 VGND 0.23929f
C15202 Iout.n30 VGND 0.23929f
C15203 Iout.n31 VGND 0.23929f
C15204 Iout.n32 VGND 0.23929f
C15205 Iout.n33 VGND 0.23929f
C15206 Iout.n34 VGND 0.23929f
C15207 Iout.n35 VGND 0.23929f
C15208 Iout.n36 VGND 0.23929f
C15209 Iout.n37 VGND 0.23929f
C15210 Iout.t46 VGND 0.02304f
C15211 Iout.n38 VGND 0.05124f
C15212 Iout.n39 VGND 0.02606f
C15213 Iout.n40 VGND 0.23929f
C15214 Iout.n41 VGND 0.04775f
C15215 Iout.t205 VGND 0.02304f
C15216 Iout.n42 VGND 0.05124f
C15217 Iout.n43 VGND 0.02606f
C15218 Iout.t201 VGND 0.02304f
C15219 Iout.n44 VGND 0.05124f
C15220 Iout.n45 VGND 0.02606f
C15221 Iout.n46 VGND 0.23929f
C15222 Iout.t189 VGND 0.02304f
C15223 Iout.n47 VGND 0.05124f
C15224 Iout.n48 VGND 0.02606f
C15225 Iout.n49 VGND 0.23929f
C15226 Iout.t206 VGND 0.02304f
C15227 Iout.n50 VGND 0.05124f
C15228 Iout.n51 VGND 0.02606f
C15229 Iout.n52 VGND 0.23929f
C15230 Iout.t188 VGND 0.02304f
C15231 Iout.n53 VGND 0.05124f
C15232 Iout.n54 VGND 0.02606f
C15233 Iout.n55 VGND 0.23929f
C15234 Iout.t53 VGND 0.02304f
C15235 Iout.n56 VGND 0.05124f
C15236 Iout.n57 VGND 0.02606f
C15237 Iout.n58 VGND 0.23929f
C15238 Iout.t249 VGND 0.02304f
C15239 Iout.n59 VGND 0.05124f
C15240 Iout.n60 VGND 0.02606f
C15241 Iout.n61 VGND 0.23929f
C15242 Iout.t108 VGND 0.02304f
C15243 Iout.n62 VGND 0.05124f
C15244 Iout.n63 VGND 0.02606f
C15245 Iout.n64 VGND 0.23929f
C15246 Iout.t212 VGND 0.02304f
C15247 Iout.n65 VGND 0.05124f
C15248 Iout.n66 VGND 0.02606f
C15249 Iout.n67 VGND 0.23929f
C15250 Iout.t210 VGND 0.02304f
C15251 Iout.n68 VGND 0.05124f
C15252 Iout.n69 VGND 0.02606f
C15253 Iout.n70 VGND 0.23929f
C15254 Iout.t144 VGND 0.02304f
C15255 Iout.n71 VGND 0.05124f
C15256 Iout.n72 VGND 0.02606f
C15257 Iout.n73 VGND 0.23929f
C15258 Iout.t166 VGND 0.02304f
C15259 Iout.n74 VGND 0.05124f
C15260 Iout.n75 VGND 0.02606f
C15261 Iout.n76 VGND 0.23929f
C15262 Iout.t184 VGND 0.02304f
C15263 Iout.n77 VGND 0.05124f
C15264 Iout.n78 VGND 0.02606f
C15265 Iout.n79 VGND 0.23929f
C15266 Iout.n80 VGND 0.23929f
C15267 Iout.t51 VGND 0.02304f
C15268 Iout.n81 VGND 0.05124f
C15269 Iout.n82 VGND 0.02606f
C15270 Iout.n83 VGND 0.23929f
C15271 Iout.n84 VGND 0.04775f
C15272 Iout.t58 VGND 0.02304f
C15273 Iout.n85 VGND 0.05124f
C15274 Iout.n86 VGND 0.02606f
C15275 Iout.t13 VGND 0.02304f
C15276 Iout.n87 VGND 0.05124f
C15277 Iout.n88 VGND 0.02606f
C15278 Iout.n89 VGND 0.23929f
C15279 Iout.t199 VGND 0.02304f
C15280 Iout.n90 VGND 0.05124f
C15281 Iout.n91 VGND 0.02606f
C15282 Iout.n92 VGND 0.23929f
C15283 Iout.t71 VGND 0.02304f
C15284 Iout.n93 VGND 0.05124f
C15285 Iout.n94 VGND 0.02606f
C15286 Iout.n95 VGND 0.23929f
C15287 Iout.t43 VGND 0.02304f
C15288 Iout.n96 VGND 0.05124f
C15289 Iout.n97 VGND 0.02606f
C15290 Iout.n98 VGND 0.23929f
C15291 Iout.t164 VGND 0.02304f
C15292 Iout.n99 VGND 0.05124f
C15293 Iout.n100 VGND 0.02606f
C15294 Iout.n101 VGND 0.23929f
C15295 Iout.t40 VGND 0.02304f
C15296 Iout.n102 VGND 0.05124f
C15297 Iout.n103 VGND 0.02606f
C15298 Iout.n104 VGND 0.23929f
C15299 Iout.t111 VGND 0.02304f
C15300 Iout.n105 VGND 0.05124f
C15301 Iout.n106 VGND 0.02606f
C15302 Iout.n107 VGND 0.23929f
C15303 Iout.t158 VGND 0.02304f
C15304 Iout.n108 VGND 0.05124f
C15305 Iout.n109 VGND 0.02606f
C15306 Iout.n110 VGND 0.23929f
C15307 Iout.t70 VGND 0.02304f
C15308 Iout.n111 VGND 0.05124f
C15309 Iout.n112 VGND 0.02606f
C15310 Iout.n113 VGND 0.23929f
C15311 Iout.t163 VGND 0.02304f
C15312 Iout.n114 VGND 0.05124f
C15313 Iout.n115 VGND 0.02606f
C15314 Iout.n116 VGND 0.23929f
C15315 Iout.t128 VGND 0.02304f
C15316 Iout.n117 VGND 0.05124f
C15317 Iout.n118 VGND 0.02606f
C15318 Iout.n119 VGND 0.23929f
C15319 Iout.t48 VGND 0.02304f
C15320 Iout.n120 VGND 0.05124f
C15321 Iout.n121 VGND 0.02606f
C15322 Iout.n122 VGND 0.04775f
C15323 Iout.t148 VGND 0.02304f
C15324 Iout.n123 VGND 0.05124f
C15325 Iout.n124 VGND 0.02606f
C15326 Iout.n125 VGND 0.23929f
C15327 Iout.n126 VGND 0.23929f
C15328 Iout.t207 VGND 0.02304f
C15329 Iout.n127 VGND 0.05124f
C15330 Iout.n128 VGND 0.02606f
C15331 Iout.n129 VGND 0.04775f
C15332 Iout.t194 VGND 0.02304f
C15333 Iout.n130 VGND 0.05124f
C15334 Iout.n131 VGND 0.02606f
C15335 Iout.n132 VGND 0.23929f
C15336 Iout.t145 VGND 0.02304f
C15337 Iout.n133 VGND 0.05124f
C15338 Iout.n134 VGND 0.02606f
C15339 Iout.n135 VGND 0.04775f
C15340 Iout.t47 VGND 0.02304f
C15341 Iout.n136 VGND 0.05124f
C15342 Iout.n137 VGND 0.02606f
C15343 Iout.n138 VGND 0.23929f
C15344 Iout.n139 VGND 0.23929f
C15345 Iout.t63 VGND 0.02304f
C15346 Iout.n140 VGND 0.05124f
C15347 Iout.n141 VGND 0.02606f
C15348 Iout.n142 VGND 0.04775f
C15349 Iout.t181 VGND 0.02304f
C15350 Iout.n143 VGND 0.05124f
C15351 Iout.n144 VGND 0.02606f
C15352 Iout.n145 VGND 0.14126f
C15353 Iout.t105 VGND 0.02304f
C15354 Iout.n146 VGND 0.05124f
C15355 Iout.n147 VGND 0.02606f
C15356 Iout.n148 VGND 0.04775f
C15357 Iout.t61 VGND 0.02304f
C15358 Iout.n149 VGND 0.05124f
C15359 Iout.n150 VGND 0.02606f
C15360 Iout.n151 VGND 0.23929f
C15361 Iout.n152 VGND 0.14126f
C15362 Iout.n153 VGND 0.23929f
C15363 Iout.n154 VGND 0.23929f
C15364 Iout.n155 VGND 0.23929f
C15365 Iout.t253 VGND 0.02304f
C15366 Iout.n156 VGND 0.05124f
C15367 Iout.n157 VGND 0.02606f
C15368 Iout.n158 VGND 0.23929f
C15369 Iout.n159 VGND 0.23929f
C15370 Iout.n160 VGND 0.23929f
C15371 Iout.n161 VGND 0.23929f
C15372 Iout.n162 VGND 0.23929f
C15373 Iout.n163 VGND 0.23929f
C15374 Iout.n164 VGND 0.23929f
C15375 Iout.n165 VGND 0.23929f
C15376 Iout.n166 VGND 0.23929f
C15377 Iout.n167 VGND 0.23929f
C15378 Iout.t6 VGND 0.02304f
C15379 Iout.n168 VGND 0.05124f
C15380 Iout.n169 VGND 0.02606f
C15381 Iout.n170 VGND 0.23929f
C15382 Iout.n171 VGND 0.04775f
C15383 Iout.t225 VGND 0.02304f
C15384 Iout.n172 VGND 0.05124f
C15385 Iout.n173 VGND 0.02606f
C15386 Iout.t29 VGND 0.02304f
C15387 Iout.n174 VGND 0.05124f
C15388 Iout.n175 VGND 0.02606f
C15389 Iout.n176 VGND 0.23929f
C15390 Iout.t98 VGND 0.02304f
C15391 Iout.n177 VGND 0.05124f
C15392 Iout.n178 VGND 0.02606f
C15393 Iout.n179 VGND 0.23929f
C15394 Iout.t7 VGND 0.02304f
C15395 Iout.n180 VGND 0.05124f
C15396 Iout.n181 VGND 0.02606f
C15397 Iout.n182 VGND 0.23929f
C15398 Iout.t177 VGND 0.02304f
C15399 Iout.n183 VGND 0.05124f
C15400 Iout.n184 VGND 0.02606f
C15401 Iout.n185 VGND 0.23929f
C15402 Iout.t255 VGND 0.02304f
C15403 Iout.n186 VGND 0.05124f
C15404 Iout.n187 VGND 0.02606f
C15405 Iout.n188 VGND 0.23929f
C15406 Iout.t123 VGND 0.02304f
C15407 Iout.n189 VGND 0.05124f
C15408 Iout.n190 VGND 0.02606f
C15409 Iout.n191 VGND 0.14126f
C15410 Iout.t236 VGND 0.02304f
C15411 Iout.n192 VGND 0.05124f
C15412 Iout.n193 VGND 0.02606f
C15413 Iout.n194 VGND 0.04775f
C15414 Iout.t242 VGND 0.02304f
C15415 Iout.n195 VGND 0.05124f
C15416 Iout.n196 VGND 0.02606f
C15417 Iout.n197 VGND 0.14126f
C15418 Iout.n198 VGND 0.04775f
C15419 Iout.t95 VGND 0.02304f
C15420 Iout.n199 VGND 0.05124f
C15421 Iout.n200 VGND 0.02606f
C15422 Iout.n201 VGND 0.04775f
C15423 Iout.t14 VGND 0.02304f
C15424 Iout.n202 VGND 0.05124f
C15425 Iout.n203 VGND 0.02606f
C15426 Iout.n204 VGND 0.14126f
C15427 Iout.n205 VGND 0.04775f
C15428 Iout.t99 VGND 0.02304f
C15429 Iout.n206 VGND 0.05124f
C15430 Iout.n207 VGND 0.02606f
C15431 Iout.n208 VGND 0.14126f
C15432 Iout.n209 VGND 0.04775f
C15433 Iout.t37 VGND 0.02304f
C15434 Iout.n210 VGND 0.05124f
C15435 Iout.n211 VGND 0.02606f
C15436 Iout.n212 VGND 0.14126f
C15437 Iout.n213 VGND 0.04775f
C15438 Iout.t34 VGND 0.02304f
C15439 Iout.n214 VGND 0.05124f
C15440 Iout.n215 VGND 0.02606f
C15441 Iout.n216 VGND 0.14126f
C15442 Iout.n217 VGND 0.04775f
C15443 Iout.t134 VGND 0.02304f
C15444 Iout.n218 VGND 0.05124f
C15445 Iout.n219 VGND 0.02606f
C15446 Iout.n220 VGND 0.14126f
C15447 Iout.n221 VGND 0.04775f
C15448 Iout.t127 VGND 0.02304f
C15449 Iout.n222 VGND 0.05124f
C15450 Iout.n223 VGND 0.02606f
C15451 Iout.n224 VGND 0.14126f
C15452 Iout.n225 VGND 0.04775f
C15453 Iout.t28 VGND 0.02304f
C15454 Iout.n226 VGND 0.05124f
C15455 Iout.n227 VGND 0.02606f
C15456 Iout.n228 VGND 0.04775f
C15457 Iout.n229 VGND 0.14126f
C15458 Iout.n230 VGND 0.23929f
C15459 Iout.n231 VGND 0.04775f
C15460 Iout.t84 VGND 0.02304f
C15461 Iout.n232 VGND 0.05124f
C15462 Iout.n233 VGND 0.02606f
C15463 Iout.n234 VGND 0.04775f
C15464 Iout.t82 VGND 0.02304f
C15465 Iout.n235 VGND 0.05124f
C15466 Iout.n236 VGND 0.02606f
C15467 Iout.n237 VGND 0.04775f
C15468 Iout.t220 VGND 0.02304f
C15469 Iout.n238 VGND 0.05124f
C15470 Iout.n239 VGND 0.02606f
C15471 Iout.n240 VGND 0.04775f
C15472 Iout.t213 VGND 0.02304f
C15473 Iout.n241 VGND 0.05124f
C15474 Iout.n242 VGND 0.02606f
C15475 Iout.n243 VGND 0.04775f
C15476 Iout.t216 VGND 0.02304f
C15477 Iout.n244 VGND 0.05124f
C15478 Iout.n245 VGND 0.02606f
C15479 Iout.n246 VGND 0.04775f
C15480 Iout.t86 VGND 0.02304f
C15481 Iout.n247 VGND 0.05124f
C15482 Iout.n248 VGND 0.02606f
C15483 Iout.n249 VGND 0.04775f
C15484 Iout.t238 VGND 0.02304f
C15485 Iout.n250 VGND 0.05124f
C15486 Iout.n251 VGND 0.02606f
C15487 Iout.t45 VGND 0.02304f
C15488 Iout.n252 VGND 0.05124f
C15489 Iout.n253 VGND 0.02606f
C15490 Iout.n254 VGND 0.04775f
C15491 Iout.t161 VGND 0.02304f
C15492 Iout.n255 VGND 0.05124f
C15493 Iout.n256 VGND 0.02606f
C15494 Iout.n257 VGND 0.04775f
C15495 Iout.n258 VGND 0.23929f
C15496 Iout.t203 VGND 0.02304f
C15497 Iout.n259 VGND 0.05124f
C15498 Iout.n260 VGND 0.02606f
C15499 Iout.n261 VGND 0.04775f
C15500 Iout.n262 VGND 0.23929f
C15501 Iout.n263 VGND 0.23929f
C15502 Iout.n264 VGND 0.04775f
C15503 Iout.t41 VGND 0.02304f
C15504 Iout.n265 VGND 0.05124f
C15505 Iout.n266 VGND 0.02606f
C15506 Iout.n267 VGND 0.04775f
C15507 Iout.n268 VGND 0.23929f
C15508 Iout.n269 VGND 0.23929f
C15509 Iout.n270 VGND 0.04775f
C15510 Iout.t130 VGND 0.02304f
C15511 Iout.n271 VGND 0.05124f
C15512 Iout.n272 VGND 0.02606f
C15513 Iout.n273 VGND 0.04775f
C15514 Iout.n274 VGND 0.23929f
C15515 Iout.n275 VGND 0.23929f
C15516 Iout.n276 VGND 0.04775f
C15517 Iout.t19 VGND 0.02304f
C15518 Iout.n277 VGND 0.05124f
C15519 Iout.n278 VGND 0.02606f
C15520 Iout.n279 VGND 0.04775f
C15521 Iout.n280 VGND 0.23929f
C15522 Iout.n281 VGND 0.23929f
C15523 Iout.n282 VGND 0.04775f
C15524 Iout.t42 VGND 0.02304f
C15525 Iout.n283 VGND 0.05124f
C15526 Iout.n284 VGND 0.02606f
C15527 Iout.n285 VGND 0.04775f
C15528 Iout.n286 VGND 0.23929f
C15529 Iout.n287 VGND 0.23929f
C15530 Iout.n288 VGND 0.04775f
C15531 Iout.t102 VGND 0.02304f
C15532 Iout.n289 VGND 0.05124f
C15533 Iout.n290 VGND 0.02606f
C15534 Iout.n291 VGND 0.04775f
C15535 Iout.n292 VGND 0.23929f
C15536 Iout.n293 VGND 0.23929f
C15537 Iout.n294 VGND 0.04775f
C15538 Iout.t214 VGND 0.02304f
C15539 Iout.n295 VGND 0.05124f
C15540 Iout.n296 VGND 0.02606f
C15541 Iout.n297 VGND 0.04775f
C15542 Iout.n298 VGND 0.23929f
C15543 Iout.n299 VGND 0.23929f
C15544 Iout.n300 VGND 0.04775f
C15545 Iout.t2 VGND 0.02304f
C15546 Iout.n301 VGND 0.05124f
C15547 Iout.n302 VGND 0.02606f
C15548 Iout.n303 VGND 0.04775f
C15549 Iout.n304 VGND 0.23929f
C15550 Iout.t136 VGND 0.02304f
C15551 Iout.n305 VGND 0.05124f
C15552 Iout.n306 VGND 0.02606f
C15553 Iout.n307 VGND 0.04775f
C15554 Iout.t221 VGND 0.02304f
C15555 Iout.n308 VGND 0.05124f
C15556 Iout.n309 VGND 0.02606f
C15557 Iout.n310 VGND 0.04775f
C15558 Iout.t81 VGND 0.02304f
C15559 Iout.n311 VGND 0.05124f
C15560 Iout.n312 VGND 0.02606f
C15561 Iout.n313 VGND 0.04775f
C15562 Iout.t173 VGND 0.02304f
C15563 Iout.n314 VGND 0.05124f
C15564 Iout.n315 VGND 0.02606f
C15565 Iout.n316 VGND 0.04775f
C15566 Iout.t77 VGND 0.02304f
C15567 Iout.n317 VGND 0.05124f
C15568 Iout.n318 VGND 0.02606f
C15569 Iout.n319 VGND 0.04775f
C15570 Iout.t183 VGND 0.02304f
C15571 Iout.n320 VGND 0.05124f
C15572 Iout.n321 VGND 0.02606f
C15573 Iout.n322 VGND 0.04775f
C15574 Iout.t209 VGND 0.02304f
C15575 Iout.n323 VGND 0.05124f
C15576 Iout.n324 VGND 0.02606f
C15577 Iout.n325 VGND 0.04775f
C15578 Iout.t93 VGND 0.02304f
C15579 Iout.n326 VGND 0.05124f
C15580 Iout.n327 VGND 0.02606f
C15581 Iout.n328 VGND 0.04775f
C15582 Iout.t74 VGND 0.02304f
C15583 Iout.n329 VGND 0.05124f
C15584 Iout.n330 VGND 0.02606f
C15585 Iout.n331 VGND 0.04775f
C15586 Iout.n332 VGND 0.23929f
C15587 Iout.t180 VGND 0.02304f
C15588 Iout.n333 VGND 0.05124f
C15589 Iout.n334 VGND 0.02606f
C15590 Iout.n335 VGND 0.04775f
C15591 Iout.t73 VGND 0.02304f
C15592 Iout.n336 VGND 0.05124f
C15593 Iout.n337 VGND 0.02606f
C15594 Iout.n338 VGND 0.04775f
C15595 Iout.t115 VGND 0.02304f
C15596 Iout.n339 VGND 0.05124f
C15597 Iout.n340 VGND 0.02606f
C15598 Iout.n341 VGND 0.04775f
C15599 Iout.t185 VGND 0.02304f
C15600 Iout.n342 VGND 0.05124f
C15601 Iout.n343 VGND 0.02606f
C15602 Iout.n344 VGND 0.04775f
C15603 Iout.t33 VGND 0.02304f
C15604 Iout.n345 VGND 0.05124f
C15605 Iout.n346 VGND 0.02606f
C15606 Iout.n347 VGND 0.04775f
C15607 Iout.t179 VGND 0.02304f
C15608 Iout.n348 VGND 0.05124f
C15609 Iout.n349 VGND 0.02606f
C15610 Iout.n350 VGND 0.04775f
C15611 Iout.t143 VGND 0.02304f
C15612 Iout.n351 VGND 0.05124f
C15613 Iout.n352 VGND 0.02606f
C15614 Iout.n353 VGND 0.04775f
C15615 Iout.t248 VGND 0.02304f
C15616 Iout.n354 VGND 0.05124f
C15617 Iout.n355 VGND 0.02606f
C15618 Iout.n356 VGND 0.04775f
C15619 Iout.t57 VGND 0.02304f
C15620 Iout.n357 VGND 0.05124f
C15621 Iout.n358 VGND 0.02606f
C15622 Iout.n359 VGND 0.04775f
C15623 Iout.t160 VGND 0.02304f
C15624 Iout.n360 VGND 0.05124f
C15625 Iout.n361 VGND 0.02606f
C15626 Iout.n362 VGND 0.04775f
C15627 Iout.t165 VGND 0.02304f
C15628 Iout.n363 VGND 0.05124f
C15629 Iout.n364 VGND 0.02606f
C15630 Iout.n365 VGND 0.04775f
C15631 Iout.t245 VGND 0.02304f
C15632 Iout.n366 VGND 0.05124f
C15633 Iout.n367 VGND 0.02606f
C15634 Iout.n368 VGND 0.04775f
C15635 Iout.n369 VGND 0.23929f
C15636 Iout.t240 VGND 0.02304f
C15637 Iout.n370 VGND 0.05124f
C15638 Iout.n371 VGND 0.02606f
C15639 Iout.n372 VGND 0.04775f
C15640 Iout.n373 VGND 0.23929f
C15641 Iout.n374 VGND 0.23929f
C15642 Iout.n375 VGND 0.04775f
C15643 Iout.t153 VGND 0.02304f
C15644 Iout.n376 VGND 0.05124f
C15645 Iout.n377 VGND 0.02606f
C15646 Iout.t120 VGND 0.02304f
C15647 Iout.n378 VGND 0.05124f
C15648 Iout.n379 VGND 0.02606f
C15649 Iout.n380 VGND 0.04775f
C15650 Iout.n381 VGND 0.23929f
C15651 Iout.n382 VGND 0.23929f
C15652 Iout.n383 VGND 0.04775f
C15653 Iout.t250 VGND 0.02304f
C15654 Iout.n384 VGND 0.05124f
C15655 Iout.n385 VGND 0.02606f
C15656 Iout.t155 VGND 0.02304f
C15657 Iout.n386 VGND 0.05124f
C15658 Iout.n387 VGND 0.02606f
C15659 Iout.n388 VGND 0.04775f
C15660 Iout.n389 VGND 0.23929f
C15661 Iout.n390 VGND 0.23929f
C15662 Iout.n391 VGND 0.04775f
C15663 Iout.t23 VGND 0.02304f
C15664 Iout.n392 VGND 0.05124f
C15665 Iout.n393 VGND 0.02606f
C15666 Iout.t67 VGND 0.02304f
C15667 Iout.n394 VGND 0.05124f
C15668 Iout.n395 VGND 0.02606f
C15669 Iout.n396 VGND 0.04775f
C15670 Iout.n397 VGND 0.23929f
C15671 Iout.n398 VGND 0.23929f
C15672 Iout.n399 VGND 0.04775f
C15673 Iout.t133 VGND 0.02304f
C15674 Iout.n400 VGND 0.05124f
C15675 Iout.n401 VGND 0.02606f
C15676 Iout.t68 VGND 0.02304f
C15677 Iout.n402 VGND 0.05124f
C15678 Iout.n403 VGND 0.02606f
C15679 Iout.n404 VGND 0.04775f
C15680 Iout.n405 VGND 0.23929f
C15681 Iout.n406 VGND 0.23929f
C15682 Iout.n407 VGND 0.04775f
C15683 Iout.t150 VGND 0.02304f
C15684 Iout.n408 VGND 0.05124f
C15685 Iout.n409 VGND 0.02606f
C15686 Iout.t222 VGND 0.02304f
C15687 Iout.n410 VGND 0.05124f
C15688 Iout.n411 VGND 0.02606f
C15689 Iout.n412 VGND 0.04775f
C15690 Iout.n413 VGND 0.23929f
C15691 Iout.n414 VGND 0.23929f
C15692 Iout.n415 VGND 0.04775f
C15693 Iout.t38 VGND 0.02304f
C15694 Iout.n416 VGND 0.05124f
C15695 Iout.n417 VGND 0.02606f
C15696 Iout.t109 VGND 0.02304f
C15697 Iout.n418 VGND 0.05124f
C15698 Iout.n419 VGND 0.02606f
C15699 Iout.n420 VGND 0.04775f
C15700 Iout.n421 VGND 0.23929f
C15701 Iout.n422 VGND 0.23929f
C15702 Iout.n423 VGND 0.04775f
C15703 Iout.t191 VGND 0.02304f
C15704 Iout.n424 VGND 0.05124f
C15705 Iout.n425 VGND 0.02606f
C15706 Iout.t157 VGND 0.02304f
C15707 Iout.n426 VGND 0.05124f
C15708 Iout.n427 VGND 0.02606f
C15709 Iout.n428 VGND 0.04775f
C15710 Iout.n429 VGND 0.23929f
C15711 Iout.n430 VGND 0.23929f
C15712 Iout.n431 VGND 0.04775f
C15713 Iout.t20 VGND 0.02304f
C15714 Iout.n432 VGND 0.05124f
C15715 Iout.n433 VGND 0.02606f
C15716 Iout.t187 VGND 0.02304f
C15717 Iout.n434 VGND 0.05124f
C15718 Iout.n435 VGND 0.02606f
C15719 Iout.n436 VGND 0.23929f
C15720 Iout.n437 VGND 0.04775f
C15721 Iout.t208 VGND 0.02304f
C15722 Iout.n438 VGND 0.05124f
C15723 Iout.n439 VGND 0.02606f
C15724 Iout.n440 VGND 0.04775f
C15725 Iout.t162 VGND 0.02304f
C15726 Iout.n441 VGND 0.05124f
C15727 Iout.n442 VGND 0.02606f
C15728 Iout.n443 VGND 0.04775f
C15729 Iout.n444 VGND 0.23929f
C15730 Iout.n445 VGND 0.23929f
C15731 Iout.n446 VGND 0.04775f
C15732 Iout.t169 VGND 0.02304f
C15733 Iout.n447 VGND 0.05124f
C15734 Iout.n448 VGND 0.02606f
C15735 Iout.t251 VGND 0.02304f
C15736 Iout.n449 VGND 0.05124f
C15737 Iout.n450 VGND 0.02606f
C15738 Iout.n451 VGND 0.04775f
C15739 Iout.t66 VGND 0.02304f
C15740 Iout.n452 VGND 0.05124f
C15741 Iout.n453 VGND 0.02606f
C15742 Iout.n454 VGND 0.04775f
C15743 Iout.n455 VGND 0.23929f
C15744 Iout.n456 VGND 0.23929f
C15745 Iout.n457 VGND 0.04775f
C15746 Iout.t149 VGND 0.02304f
C15747 Iout.n458 VGND 0.05124f
C15748 Iout.n459 VGND 0.02606f
C15749 Iout.t65 VGND 0.02304f
C15750 Iout.n460 VGND 0.05124f
C15751 Iout.n461 VGND 0.02606f
C15752 Iout.n462 VGND 0.04775f
C15753 Iout.t16 VGND 0.02304f
C15754 Iout.n463 VGND 0.05124f
C15755 Iout.n464 VGND 0.02606f
C15756 Iout.n465 VGND 0.04775f
C15757 Iout.n466 VGND 0.23929f
C15758 Iout.n467 VGND 0.23929f
C15759 Iout.n468 VGND 0.04775f
C15760 Iout.t151 VGND 0.02304f
C15761 Iout.n469 VGND 0.05124f
C15762 Iout.n470 VGND 0.02606f
C15763 Iout.n471 VGND 0.04775f
C15764 Iout.t219 VGND 0.02304f
C15765 Iout.n472 VGND 0.05124f
C15766 Iout.n473 VGND 0.02606f
C15767 Iout.n474 VGND 0.04775f
C15768 Iout.n475 VGND 0.23929f
C15769 Iout.n476 VGND 0.23929f
C15770 Iout.n477 VGND 0.04775f
C15771 Iout.t4 VGND 0.02304f
C15772 Iout.n478 VGND 0.05124f
C15773 Iout.n479 VGND 0.02606f
C15774 Iout.t80 VGND 0.02304f
C15775 Iout.n480 VGND 0.05124f
C15776 Iout.n481 VGND 0.02606f
C15777 Iout.n482 VGND 0.04775f
C15778 Iout.t55 VGND 0.02304f
C15779 Iout.n483 VGND 0.05124f
C15780 Iout.n484 VGND 0.02606f
C15781 Iout.n485 VGND 0.04775f
C15782 Iout.n486 VGND 0.23929f
C15783 Iout.n487 VGND 0.23929f
C15784 Iout.n488 VGND 0.04775f
C15785 Iout.t69 VGND 0.02304f
C15786 Iout.n489 VGND 0.05124f
C15787 Iout.n490 VGND 0.02606f
C15788 Iout.t91 VGND 0.02304f
C15789 Iout.n491 VGND 0.05124f
C15790 Iout.n492 VGND 0.02606f
C15791 Iout.n493 VGND 0.04775f
C15792 Iout.t192 VGND 0.02304f
C15793 Iout.n494 VGND 0.05124f
C15794 Iout.n495 VGND 0.02606f
C15795 Iout.n496 VGND 0.04775f
C15796 Iout.n497 VGND 0.23929f
C15797 Iout.n498 VGND 0.14126f
C15798 Iout.n499 VGND 0.04775f
C15799 Iout.t147 VGND 0.02304f
C15800 Iout.n500 VGND 0.05124f
C15801 Iout.n501 VGND 0.02606f
C15802 Iout.n502 VGND 0.14126f
C15803 Iout.n503 VGND 0.04775f
C15804 Iout.t126 VGND 0.02304f
C15805 Iout.n504 VGND 0.05124f
C15806 Iout.n505 VGND 0.02606f
C15807 Iout.n506 VGND 0.04775f
C15808 Iout.t131 VGND 0.02304f
C15809 Iout.n507 VGND 0.05124f
C15810 Iout.n508 VGND 0.02606f
C15811 Iout.t124 VGND 0.02304f
C15812 Iout.n509 VGND 0.05124f
C15813 Iout.n510 VGND 0.02606f
C15814 Iout.n511 VGND 0.14126f
C15815 Iout.n512 VGND 0.04775f
C15816 Iout.t11 VGND 0.02304f
C15817 Iout.n513 VGND 0.05124f
C15818 Iout.n514 VGND 0.02606f
C15819 Iout.n515 VGND 0.04775f
C15820 Iout.n516 VGND 0.14126f
C15821 Iout.n517 VGND 0.23929f
C15822 Iout.n518 VGND 0.04775f
C15823 Iout.t83 VGND 0.02304f
C15824 Iout.n519 VGND 0.05124f
C15825 Iout.n520 VGND 0.02606f
C15826 Iout.n521 VGND 0.04775f
C15827 Iout.n522 VGND 0.23929f
C15828 Iout.n523 VGND 0.23929f
C15829 Iout.n524 VGND 0.04775f
C15830 Iout.t146 VGND 0.02304f
C15831 Iout.n525 VGND 0.05124f
C15832 Iout.n526 VGND 0.02606f
C15833 Iout.n527 VGND 0.04775f
C15834 Iout.n528 VGND 0.23929f
C15835 Iout.n529 VGND 0.23929f
C15836 Iout.n530 VGND 0.04775f
C15837 Iout.t79 VGND 0.02304f
C15838 Iout.n531 VGND 0.05124f
C15839 Iout.n532 VGND 0.02606f
C15840 Iout.n533 VGND 0.04775f
C15841 Iout.t113 VGND 0.02304f
C15842 Iout.n534 VGND 0.05124f
C15843 Iout.n535 VGND 0.02606f
C15844 Iout.t172 VGND 0.02304f
C15845 Iout.n536 VGND 0.05124f
C15846 Iout.n537 VGND 0.02606f
C15847 Iout.n538 VGND 0.04775f
C15848 Iout.n539 VGND 0.23929f
C15849 Iout.n540 VGND 0.23929f
C15850 Iout.n541 VGND 0.04775f
C15851 Iout.t233 VGND 0.02304f
C15852 Iout.n542 VGND 0.05124f
C15853 Iout.n543 VGND 0.02606f
C15854 Iout.n544 VGND 0.04775f
C15855 Iout.n545 VGND 0.23929f
C15856 Iout.n546 VGND 0.23929f
C15857 Iout.n547 VGND 0.04775f
C15858 Iout.t25 VGND 0.02304f
C15859 Iout.n548 VGND 0.05124f
C15860 Iout.n549 VGND 0.02606f
C15861 Iout.n550 VGND 0.04775f
C15862 Iout.n551 VGND 0.23929f
C15863 Iout.n552 VGND 0.23929f
C15864 Iout.n553 VGND 0.04775f
C15865 Iout.t72 VGND 0.02304f
C15866 Iout.n554 VGND 0.05124f
C15867 Iout.n555 VGND 0.02606f
C15868 Iout.n556 VGND 0.04775f
C15869 Iout.t223 VGND 0.02304f
C15870 Iout.n557 VGND 0.05124f
C15871 Iout.n558 VGND 0.02606f
C15872 Iout.t121 VGND 0.02304f
C15873 Iout.n559 VGND 0.05124f
C15874 Iout.n560 VGND 0.02606f
C15875 Iout.n561 VGND 0.04775f
C15876 Iout.n562 VGND 0.23929f
C15877 Iout.t106 VGND 0.02304f
C15878 Iout.n563 VGND 0.05124f
C15879 Iout.n564 VGND 0.02606f
C15880 Iout.n565 VGND 0.04775f
C15881 Iout.n566 VGND 0.23929f
C15882 Iout.n567 VGND 0.23929f
C15883 Iout.n568 VGND 0.04775f
C15884 Iout.t12 VGND 0.02304f
C15885 Iout.n569 VGND 0.05124f
C15886 Iout.n570 VGND 0.02606f
C15887 Iout.n571 VGND 0.04775f
C15888 Iout.n572 VGND 0.23929f
C15889 Iout.t88 VGND 0.02304f
C15890 Iout.n573 VGND 0.05124f
C15891 Iout.n574 VGND 0.02606f
C15892 Iout.n575 VGND 0.04775f
C15893 Iout.t90 VGND 0.02304f
C15894 Iout.n576 VGND 0.05124f
C15895 Iout.n577 VGND 0.02606f
C15896 Iout.n578 VGND 0.04775f
C15897 Iout.n579 VGND 0.23929f
C15898 Iout.n580 VGND 0.23929f
C15899 Iout.n581 VGND 0.04775f
C15900 Iout.t50 VGND 0.02304f
C15901 Iout.n582 VGND 0.05124f
C15902 Iout.n583 VGND 0.02606f
C15903 Iout.n584 VGND 0.04775f
C15904 Iout.n585 VGND 0.23929f
C15905 Iout.n586 VGND 0.23929f
C15906 Iout.n587 VGND 0.04775f
C15907 Iout.t239 VGND 0.02304f
C15908 Iout.n588 VGND 0.05124f
C15909 Iout.n589 VGND 0.02606f
C15910 Iout.n590 VGND 0.04775f
C15911 Iout.n591 VGND 0.23929f
C15912 Iout.n592 VGND 0.23929f
C15913 Iout.n593 VGND 0.04775f
C15914 Iout.t218 VGND 0.02304f
C15915 Iout.n594 VGND 0.05124f
C15916 Iout.n595 VGND 0.02606f
C15917 Iout.n596 VGND 0.04775f
C15918 Iout.n597 VGND 0.23929f
C15919 Iout.n598 VGND 0.23929f
C15920 Iout.n599 VGND 0.04775f
C15921 Iout.t171 VGND 0.02304f
C15922 Iout.n600 VGND 0.05124f
C15923 Iout.n601 VGND 0.02606f
C15924 Iout.n602 VGND 0.04775f
C15925 Iout.n603 VGND 0.23929f
C15926 Iout.n604 VGND 0.23929f
C15927 Iout.n605 VGND 0.04775f
C15928 Iout.t85 VGND 0.02304f
C15929 Iout.n606 VGND 0.05124f
C15930 Iout.n607 VGND 0.02606f
C15931 Iout.n608 VGND 0.04775f
C15932 Iout.n609 VGND 0.23929f
C15933 Iout.n610 VGND 0.23929f
C15934 Iout.n611 VGND 0.04775f
C15935 Iout.t10 VGND 0.02304f
C15936 Iout.n612 VGND 0.05124f
C15937 Iout.n613 VGND 0.02606f
C15938 Iout.n614 VGND 0.04775f
C15939 Iout.n615 VGND 0.23929f
C15940 Iout.n616 VGND 0.23929f
C15941 Iout.n617 VGND 0.04775f
C15942 Iout.t119 VGND 0.02304f
C15943 Iout.n618 VGND 0.05124f
C15944 Iout.n619 VGND 0.02606f
C15945 Iout.n620 VGND 0.04775f
C15946 Iout.n621 VGND 0.23929f
C15947 Iout.n622 VGND 0.23929f
C15948 Iout.n623 VGND 0.04775f
C15949 Iout.t27 VGND 0.02304f
C15950 Iout.n624 VGND 0.05124f
C15951 Iout.n625 VGND 0.02606f
C15952 Iout.n626 VGND 0.04775f
C15953 Iout.n627 VGND 0.23929f
C15954 Iout.n628 VGND 0.23929f
C15955 Iout.n629 VGND 0.04775f
C15956 Iout.t36 VGND 0.02304f
C15957 Iout.n630 VGND 0.05124f
C15958 Iout.n631 VGND 0.02606f
C15959 Iout.n632 VGND 0.04775f
C15960 Iout.n633 VGND 0.23929f
C15961 Iout.n634 VGND 0.23929f
C15962 Iout.n635 VGND 0.04775f
C15963 Iout.t103 VGND 0.02304f
C15964 Iout.n636 VGND 0.05124f
C15965 Iout.n637 VGND 0.02606f
C15966 Iout.n638 VGND 0.04775f
C15967 Iout.n639 VGND 0.23929f
C15968 Iout.n640 VGND 0.23929f
C15969 Iout.n641 VGND 0.04775f
C15970 Iout.t122 VGND 0.02304f
C15971 Iout.n642 VGND 0.05124f
C15972 Iout.n643 VGND 0.02606f
C15973 Iout.n644 VGND 0.04775f
C15974 Iout.n645 VGND 0.23929f
C15975 Iout.n646 VGND 0.23929f
C15976 Iout.n647 VGND 0.04775f
C15977 Iout.t125 VGND 0.02304f
C15978 Iout.n648 VGND 0.05124f
C15979 Iout.n649 VGND 0.02606f
C15980 Iout.n650 VGND 0.04775f
C15981 Iout.n651 VGND 0.23929f
C15982 Iout.n652 VGND 0.23929f
C15983 Iout.n653 VGND 0.04775f
C15984 Iout.t1 VGND 0.02304f
C15985 Iout.n654 VGND 0.05124f
C15986 Iout.n655 VGND 0.02606f
C15987 Iout.n656 VGND 0.04775f
C15988 Iout.t241 VGND 0.02304f
C15989 Iout.n657 VGND 0.05124f
C15990 Iout.n658 VGND 0.02606f
C15991 Iout.n659 VGND 0.04775f
C15992 Iout.t254 VGND 0.02304f
C15993 Iout.n660 VGND 0.05124f
C15994 Iout.n661 VGND 0.02606f
C15995 Iout.n662 VGND 0.04775f
C15996 Iout.t35 VGND 0.02304f
C15997 Iout.n663 VGND 0.05124f
C15998 Iout.n664 VGND 0.02606f
C15999 Iout.n665 VGND 0.04775f
C16000 Iout.t59 VGND 0.02304f
C16001 Iout.n666 VGND 0.05124f
C16002 Iout.n667 VGND 0.02606f
C16003 Iout.n668 VGND 0.04775f
C16004 Iout.t138 VGND 0.02304f
C16005 Iout.n669 VGND 0.05124f
C16006 Iout.n670 VGND 0.02606f
C16007 Iout.n671 VGND 0.04775f
C16008 Iout.t229 VGND 0.02304f
C16009 Iout.n672 VGND 0.05124f
C16010 Iout.n673 VGND 0.02606f
C16011 Iout.n674 VGND 0.04775f
C16012 Iout.t226 VGND 0.02304f
C16013 Iout.n675 VGND 0.05124f
C16014 Iout.n676 VGND 0.02606f
C16015 Iout.n677 VGND 0.04775f
C16016 Iout.t22 VGND 0.02304f
C16017 Iout.n678 VGND 0.05124f
C16018 Iout.n679 VGND 0.02606f
C16019 Iout.n680 VGND 0.04775f
C16020 Iout.t64 VGND 0.02304f
C16021 Iout.n681 VGND 0.05124f
C16022 Iout.n682 VGND 0.02606f
C16023 Iout.n683 VGND 0.04775f
C16024 Iout.t156 VGND 0.02304f
C16025 Iout.n684 VGND 0.05124f
C16026 Iout.n685 VGND 0.02606f
C16027 Iout.n686 VGND 0.04775f
C16028 Iout.t237 VGND 0.02304f
C16029 Iout.n687 VGND 0.05124f
C16030 Iout.n688 VGND 0.02606f
C16031 Iout.n689 VGND 0.04775f
C16032 Iout.t75 VGND 0.02304f
C16033 Iout.n690 VGND 0.05124f
C16034 Iout.n691 VGND 0.02606f
C16035 Iout.t193 VGND 0.02304f
C16036 Iout.n692 VGND 0.05124f
C16037 Iout.n693 VGND 0.02606f
C16038 Iout.n694 VGND 0.04775f
C16039 Iout.t107 VGND 0.02304f
C16040 Iout.n695 VGND 0.05124f
C16041 Iout.n696 VGND 0.02606f
C16042 Iout.n697 VGND 0.04775f
C16043 Iout.n698 VGND 0.23929f
C16044 Iout.t101 VGND 0.02304f
C16045 Iout.n699 VGND 0.05124f
C16046 Iout.n700 VGND 0.02606f
C16047 Iout.n701 VGND 0.04775f
C16048 Iout.n702 VGND 0.23929f
C16049 Iout.n703 VGND 0.23929f
C16050 Iout.n704 VGND 0.04775f
C16051 Iout.t152 VGND 0.02304f
C16052 Iout.n705 VGND 0.05124f
C16053 Iout.n706 VGND 0.02606f
C16054 Iout.n707 VGND 0.04775f
C16055 Iout.n708 VGND 0.23929f
C16056 Iout.n709 VGND 0.23929f
C16057 Iout.n710 VGND 0.04775f
C16058 Iout.t175 VGND 0.02304f
C16059 Iout.n711 VGND 0.05124f
C16060 Iout.n712 VGND 0.02606f
C16061 Iout.n713 VGND 0.04775f
C16062 Iout.n714 VGND 0.23929f
C16063 Iout.n715 VGND 0.23929f
C16064 Iout.n716 VGND 0.04775f
C16065 Iout.t231 VGND 0.02304f
C16066 Iout.n717 VGND 0.05124f
C16067 Iout.n718 VGND 0.02606f
C16068 Iout.n719 VGND 0.04775f
C16069 Iout.n720 VGND 0.23929f
C16070 Iout.n721 VGND 0.23929f
C16071 Iout.n722 VGND 0.04775f
C16072 Iout.t247 VGND 0.02304f
C16073 Iout.n723 VGND 0.05124f
C16074 Iout.n724 VGND 0.02606f
C16075 Iout.n725 VGND 0.04775f
C16076 Iout.n726 VGND 0.23929f
C16077 Iout.n727 VGND 0.23929f
C16078 Iout.n728 VGND 0.04775f
C16079 Iout.t243 VGND 0.02304f
C16080 Iout.n729 VGND 0.05124f
C16081 Iout.n730 VGND 0.02606f
C16082 Iout.n731 VGND 0.04775f
C16083 Iout.n732 VGND 0.23929f
C16084 Iout.n733 VGND 0.23929f
C16085 Iout.n734 VGND 0.04775f
C16086 Iout.t17 VGND 0.02304f
C16087 Iout.n735 VGND 0.05124f
C16088 Iout.n736 VGND 0.02606f
C16089 Iout.n737 VGND 0.04775f
C16090 Iout.n738 VGND 0.23929f
C16091 Iout.n739 VGND 0.23929f
C16092 Iout.n740 VGND 0.04775f
C16093 Iout.t94 VGND 0.02304f
C16094 Iout.n741 VGND 0.05124f
C16095 Iout.n742 VGND 0.02606f
C16096 Iout.n743 VGND 0.04775f
C16097 Iout.n744 VGND 0.23929f
C16098 Iout.n745 VGND 0.23929f
C16099 Iout.n746 VGND 0.04775f
C16100 Iout.t230 VGND 0.02304f
C16101 Iout.n747 VGND 0.05124f
C16102 Iout.n748 VGND 0.02606f
C16103 Iout.n749 VGND 0.04775f
C16104 Iout.n750 VGND 0.23929f
C16105 Iout.n751 VGND 0.23929f
C16106 Iout.n752 VGND 0.04775f
C16107 Iout.t31 VGND 0.02304f
C16108 Iout.n753 VGND 0.05124f
C16109 Iout.n754 VGND 0.02606f
C16110 Iout.n755 VGND 0.04775f
C16111 Iout.n756 VGND 0.23929f
C16112 Iout.n757 VGND 0.23929f
C16113 Iout.n758 VGND 0.04775f
C16114 Iout.t167 VGND 0.02304f
C16115 Iout.n759 VGND 0.05124f
C16116 Iout.n760 VGND 0.02606f
C16117 Iout.n761 VGND 0.04775f
C16118 Iout.n762 VGND 0.23929f
C16119 Iout.n763 VGND 0.23929f
C16120 Iout.n764 VGND 0.04775f
C16121 Iout.t62 VGND 0.02304f
C16122 Iout.n765 VGND 0.05124f
C16123 Iout.n766 VGND 0.02606f
C16124 Iout.n767 VGND 0.04775f
C16125 Iout.n768 VGND 0.23929f
C16126 Iout.n769 VGND 0.23929f
C16127 Iout.n770 VGND 0.04775f
C16128 Iout.t89 VGND 0.02304f
C16129 Iout.n771 VGND 0.05124f
C16130 Iout.n772 VGND 0.02606f
C16131 Iout.n773 VGND 0.04775f
C16132 Iout.n774 VGND 0.23929f
C16133 Iout.n775 VGND 0.23929f
C16134 Iout.n776 VGND 0.04775f
C16135 Iout.t129 VGND 0.02304f
C16136 Iout.n777 VGND 0.05124f
C16137 Iout.n778 VGND 0.02606f
C16138 Iout.n779 VGND 0.04775f
C16139 Iout.n780 VGND 0.23929f
C16140 Iout.t215 VGND 0.02304f
C16141 Iout.n781 VGND 0.05124f
C16142 Iout.n782 VGND 0.02606f
C16143 Iout.n783 VGND 0.04775f
C16144 Iout.t26 VGND 0.02304f
C16145 Iout.n784 VGND 0.05124f
C16146 Iout.n785 VGND 0.02606f
C16147 Iout.n786 VGND 0.04775f
C16148 Iout.t39 VGND 0.02304f
C16149 Iout.n787 VGND 0.05124f
C16150 Iout.n788 VGND 0.02606f
C16151 Iout.n789 VGND 0.04775f
C16152 Iout.t186 VGND 0.02304f
C16153 Iout.n790 VGND 0.05124f
C16154 Iout.n791 VGND 0.02606f
C16155 Iout.n792 VGND 0.04775f
C16156 Iout.t195 VGND 0.02304f
C16157 Iout.n793 VGND 0.05124f
C16158 Iout.n794 VGND 0.02606f
C16159 Iout.n795 VGND 0.04775f
C16160 Iout.t49 VGND 0.02304f
C16161 Iout.n796 VGND 0.05124f
C16162 Iout.n797 VGND 0.02606f
C16163 Iout.n798 VGND 0.04775f
C16164 Iout.t100 VGND 0.02304f
C16165 Iout.n799 VGND 0.05124f
C16166 Iout.n800 VGND 0.02606f
C16167 Iout.n801 VGND 0.04775f
C16168 Iout.t76 VGND 0.02304f
C16169 Iout.n802 VGND 0.05124f
C16170 Iout.n803 VGND 0.02606f
C16171 Iout.n804 VGND 0.04775f
C16172 Iout.t154 VGND 0.02304f
C16173 Iout.n805 VGND 0.05124f
C16174 Iout.n806 VGND 0.02606f
C16175 Iout.n807 VGND 0.04775f
C16176 Iout.t114 VGND 0.02304f
C16177 Iout.n808 VGND 0.05124f
C16178 Iout.n809 VGND 0.02606f
C16179 Iout.n810 VGND 0.04775f
C16180 Iout.t202 VGND 0.02304f
C16181 Iout.n811 VGND 0.05124f
C16182 Iout.n812 VGND 0.02606f
C16183 Iout.n813 VGND 0.04775f
C16184 Iout.t141 VGND 0.02304f
C16185 Iout.n814 VGND 0.05124f
C16186 Iout.n815 VGND 0.02606f
C16187 Iout.n816 VGND 0.04775f
C16188 Iout.t15 VGND 0.02304f
C16189 Iout.n817 VGND 0.05124f
C16190 Iout.n818 VGND 0.02606f
C16191 Iout.n819 VGND 0.04775f
C16192 Iout.t228 VGND 0.02304f
C16193 Iout.n820 VGND 0.05124f
C16194 Iout.n821 VGND 0.02606f
C16195 Iout.n822 VGND 0.04775f
C16196 Iout.t235 VGND 0.02304f
C16197 Iout.n823 VGND 0.05124f
C16198 Iout.n824 VGND 0.02606f
C16199 Iout.n825 VGND 0.04775f
C16200 Iout.n826 VGND 0.23929f
C16201 Iout.t182 VGND 0.02304f
C16202 Iout.n827 VGND 0.05124f
C16203 Iout.n828 VGND 0.02606f
C16204 Iout.n829 VGND 0.08168f
C16205 Iout.n830 VGND 0.49611f
C16206 Iout.n831 VGND 0.04775f
C16207 Iout.t244 VGND 0.02304f
C16208 Iout.n832 VGND 0.05124f
C16209 Iout.n833 VGND 0.02606f
C16210 Iout.t110 VGND 0.02304f
C16211 Iout.n834 VGND 0.05124f
C16212 Iout.n835 VGND 0.02606f
C16213 Iout.n836 VGND 0.04775f
C16214 Iout.n837 VGND 0.49611f
C16215 Iout.n838 VGND 0.08168f
C16216 Iout.t97 VGND 0.02304f
C16217 Iout.n839 VGND 0.05124f
C16218 Iout.n840 VGND 0.02606f
C16219 Iout.t174 VGND 0.02304f
C16220 Iout.n841 VGND 0.05124f
C16221 Iout.n842 VGND 0.02606f
C16222 Iout.n843 VGND 0.08168f
C16223 Iout.n844 VGND 0.49611f
C16224 Iout.n845 VGND 0.04775f
C16225 Iout.t232 VGND 0.02304f
C16226 Iout.n846 VGND 0.05124f
C16227 Iout.n847 VGND 0.02606f
C16228 Iout.t217 VGND 0.02304f
C16229 Iout.n848 VGND 0.05124f
C16230 Iout.n849 VGND 0.02606f
C16231 Iout.n850 VGND 0.04775f
C16232 Iout.n851 VGND 0.49611f
C16233 Iout.n852 VGND 0.08168f
C16234 Iout.t142 VGND 0.02304f
C16235 Iout.n853 VGND 0.05124f
C16236 Iout.n854 VGND 0.02606f
C16237 Iout.t178 VGND 0.02304f
C16238 Iout.n855 VGND 0.05124f
C16239 Iout.n856 VGND 0.02606f
C16240 Iout.n857 VGND 0.08168f
C16241 Iout.n858 VGND 0.49611f
C16242 Iout.n859 VGND 0.04775f
C16243 Iout.t54 VGND 0.02304f
C16244 Iout.n860 VGND 0.05124f
C16245 Iout.n861 VGND 0.02606f
C16246 Iout.t197 VGND 0.02304f
C16247 Iout.n862 VGND 0.05124f
C16248 Iout.n863 VGND 0.02606f
C16249 Iout.n864 VGND 0.04775f
C16250 Iout.n865 VGND 0.49611f
C16251 Iout.n866 VGND 0.08168f
C16252 Iout.t32 VGND 0.02304f
C16253 Iout.n867 VGND 0.05124f
C16254 Iout.n868 VGND 0.02606f
C16255 Iout.t52 VGND 0.02304f
C16256 Iout.n869 VGND 0.05124f
C16257 Iout.n870 VGND 0.02606f
C16258 Iout.n871 VGND 0.08168f
C16259 Iout.n872 VGND 0.49611f
C16260 Iout.n873 VGND 0.04775f
C16261 Iout.t200 VGND 0.02304f
C16262 Iout.n874 VGND 0.05124f
C16263 Iout.n875 VGND 0.02606f
C16264 Iout.t159 VGND 0.02304f
C16265 Iout.n876 VGND 0.05124f
C16266 Iout.n877 VGND 0.02606f
C16267 Iout.n878 VGND 0.04775f
C16268 Iout.n879 VGND 0.49611f
C16269 Iout.n880 VGND 0.08168f
C16270 Iout.t168 VGND 0.02304f
C16271 Iout.n881 VGND 0.05124f
C16272 Iout.n882 VGND 0.02606f
C16273 Iout.t92 VGND 0.02304f
C16274 Iout.n883 VGND 0.05124f
C16275 Iout.n884 VGND 0.02606f
C16276 Iout.n885 VGND 0.08168f
C16277 Iout.n886 VGND 0.49611f
C16278 Iout.n887 VGND 0.04775f
C16279 Iout.t112 VGND 0.02304f
C16280 Iout.n888 VGND 0.05124f
C16281 Iout.n889 VGND 0.02606f
C16282 Iout.t117 VGND 0.02304f
C16283 Iout.n890 VGND 0.05124f
C16284 Iout.n891 VGND 0.02606f
C16285 Iout.n892 VGND 0.04775f
C16286 Iout.n893 VGND 0.49611f
C16287 Iout.n894 VGND 0.08168f
C16288 Iout.t204 VGND 0.02304f
C16289 Iout.n895 VGND 0.05124f
C16290 Iout.n896 VGND 0.02606f
C16291 Iout.t8 VGND 0.02304f
C16292 Iout.n897 VGND 0.05124f
C16293 Iout.n898 VGND 0.02606f
C16294 Iout.n899 VGND 0.08168f
C16295 Iout.n900 VGND 0.49611f
C16296 Iout.n901 VGND 0.04775f
C16297 Iout.t24 VGND 0.02304f
C16298 Iout.n902 VGND 0.05124f
C16299 Iout.n903 VGND 0.02606f
C16300 Iout.t198 VGND 0.02304f
C16301 Iout.n904 VGND 0.05124f
C16302 Iout.n905 VGND 0.02606f
C16303 Iout.n906 VGND 0.04775f
C16304 Iout.n907 VGND 0.49611f
C16305 Iout.n908 VGND 0.08168f
C16306 Iout.t170 VGND 0.02304f
C16307 Iout.n909 VGND 0.05124f
C16308 Iout.n910 VGND 0.02606f
C16309 Iout.t227 VGND 0.02304f
C16310 Iout.n911 VGND 0.05124f
C16311 Iout.n912 VGND 0.02606f
C16312 Iout.n913 VGND 0.08168f
C16313 Iout.n914 VGND 0.49611f
C16314 Iout.n915 VGND 0.04775f
C16315 Iout.t135 VGND 0.02304f
C16316 Iout.n916 VGND 0.05124f
C16317 Iout.n917 VGND 0.02606f
C16318 Iout.t246 VGND 0.02304f
C16319 Iout.n918 VGND 0.05124f
C16320 Iout.n919 VGND 0.02606f
C16321 Iout.n920 VGND 0.04775f
C16322 Iout.n921 VGND 0.49611f
C16323 Iout.n922 VGND 0.08168f
C16324 Iout.t0 VGND 0.02304f
C16325 Iout.n923 VGND 0.05124f
C16326 Iout.n924 VGND 0.02606f
C16327 Iout.n925 VGND 0.08168f
C16328 Iout.t118 VGND 0.02304f
C16329 Iout.n926 VGND 0.05124f
C16330 Iout.n927 VGND 0.02606f
C16331 Iout.n928 VGND 0.08168f
C16332 Iout.n929 VGND 0.49611f
C16333 Iout.n930 VGND 0.04775f
C16334 Iout.t211 VGND 0.02304f
C16335 Iout.n931 VGND 0.05124f
C16336 Iout.n932 VGND 0.02606f
C16337 Iout.n933 VGND 0.04775f
C16338 Iout.t78 VGND 0.02304f
C16339 Iout.n934 VGND 0.05124f
C16340 Iout.n935 VGND 0.20242f
C16341 Iout.n936 VGND 2.65139f
C16342 Iout.n937 VGND 1.25122f
C16343 Iout.t9 VGND 0.02304f
C16344 Iout.n938 VGND 0.05124f
C16345 Iout.n939 VGND 0.20242f
C16346 Iout.n940 VGND 0.04775f
C16347 Iout.n941 VGND 0.23929f
C16348 Iout.n942 VGND 0.23929f
C16349 Iout.n943 VGND 0.04775f
C16350 Iout.t3 VGND 0.02304f
C16351 Iout.n944 VGND 0.05124f
C16352 Iout.n945 VGND 0.02606f
C16353 Iout.n946 VGND 0.04775f
C16354 Iout.n947 VGND 0.23929f
C16355 Iout.n948 VGND 0.23929f
C16356 Iout.n949 VGND 0.04775f
C16357 Iout.t104 VGND 0.02304f
C16358 Iout.n950 VGND 0.05124f
C16359 Iout.n951 VGND 0.02606f
C16360 Iout.n952 VGND 0.04775f
C16361 Iout.t252 VGND 0.02304f
C16362 Iout.n953 VGND 0.05124f
C16363 Iout.n954 VGND 0.20242f
C16364 Iout.n955 VGND 1.25122f
C16365 Iout.n956 VGND 1.25122f
C16366 Iout.t44 VGND 0.02304f
C16367 Iout.n957 VGND 0.05124f
C16368 Iout.n958 VGND 0.20242f
C16369 Iout.n959 VGND 0.04775f
C16370 Iout.n960 VGND 0.23929f
C16371 Iout.n961 VGND 0.23929f
C16372 Iout.n962 VGND 0.04775f
C16373 Iout.t176 VGND 0.02304f
C16374 Iout.n963 VGND 0.05124f
C16375 Iout.n964 VGND 0.02606f
C16376 Iout.n965 VGND 0.04775f
C16377 Iout.n966 VGND 0.23929f
C16378 Iout.n967 VGND 0.23929f
C16379 Iout.n968 VGND 0.04775f
C16380 Iout.t18 VGND 0.02304f
C16381 Iout.n969 VGND 0.05124f
C16382 Iout.n970 VGND 0.02606f
C16383 Iout.n971 VGND 0.04775f
C16384 Iout.t5 VGND 0.02304f
C16385 Iout.n972 VGND 0.05124f
C16386 Iout.n973 VGND 0.20242f
C16387 Iout.n974 VGND 1.25122f
C16388 Iout.n975 VGND 1.25122f
C16389 Iout.t140 VGND 0.02304f
C16390 Iout.n976 VGND 0.05124f
C16391 Iout.n977 VGND 0.20242f
C16392 Iout.n978 VGND 0.04775f
C16393 Iout.n979 VGND 0.23929f
C16394 Iout.n980 VGND 0.23929f
C16395 Iout.n981 VGND 0.04775f
C16396 Iout.t190 VGND 0.02304f
C16397 Iout.n982 VGND 0.05124f
C16398 Iout.n983 VGND 0.02606f
C16399 Iout.n984 VGND 0.04775f
C16400 Iout.n985 VGND 0.23929f
C16401 Iout.n986 VGND 0.23929f
C16402 Iout.n987 VGND 0.04775f
C16403 Iout.t30 VGND 0.02304f
C16404 Iout.n988 VGND 0.05124f
C16405 Iout.n989 VGND 0.02606f
C16406 Iout.n990 VGND 0.04775f
C16407 Iout.t137 VGND 0.02304f
C16408 Iout.n991 VGND 0.05124f
C16409 Iout.n992 VGND 0.20242f
C16410 Iout.n993 VGND 1.25122f
C16411 Iout.n994 VGND 1.25122f
C16412 Iout.t234 VGND 0.02304f
C16413 Iout.n995 VGND 0.05124f
C16414 Iout.n996 VGND 0.20242f
C16415 Iout.n997 VGND 0.04775f
C16416 Iout.n998 VGND 0.23929f
C16417 Iout.n999 VGND 0.23929f
C16418 Iout.n1000 VGND 0.04775f
C16419 Iout.t60 VGND 0.02304f
C16420 Iout.n1001 VGND 0.05124f
C16421 Iout.n1002 VGND 0.02606f
C16422 Iout.n1003 VGND 0.04775f
C16423 Iout.n1004 VGND 0.23929f
C16424 Iout.n1005 VGND 0.23929f
C16425 Iout.n1006 VGND 0.04775f
C16426 Iout.t56 VGND 0.02304f
C16427 Iout.n1007 VGND 0.05124f
C16428 Iout.n1008 VGND 0.02606f
C16429 Iout.n1009 VGND 0.04775f
C16430 Iout.t139 VGND 0.02304f
C16431 Iout.n1010 VGND 0.05124f
C16432 Iout.n1011 VGND 0.20242f
C16433 Iout.n1012 VGND 1.25122f
C16434 Iout.n1013 VGND 1.1235f
C16435 Iout.t87 VGND 0.02304f
C16436 Iout.n1014 VGND 0.05124f
C16437 Iout.n1015 VGND 0.20242f
C16438 Iout.n1016 VGND 0.04775f
C16439 Iout.n1017 VGND 0.23929f
C16440 Iout.n1018 VGND 0.14126f
C16441 Iout.n1019 VGND 0.04775f
C16442 Iout.t21 VGND 0.02304f
C16443 Iout.n1020 VGND 0.05124f
C16444 Iout.n1021 VGND 0.20242f
C16445 Iout.n1022 VGND 0.23244f
C16446 VPWR.n0 VGND 0.04687f
C16447 VPWR.t1722 VGND 0.29639f
C16448 VPWR.t502 VGND 0.13116f
C16449 VPWR.t1873 VGND 0.37815f
C16450 VPWR.t448 VGND 0.14308f
C16451 VPWR.t416 VGND 0.14308f
C16452 VPWR.t412 VGND 0.14308f
C16453 VPWR.t988 VGND 0.14308f
C16454 VPWR.t1501 VGND 0.14308f
C16455 VPWR.t1497 VGND 0.14308f
C16456 VPWR.t992 VGND 0.1005f
C16457 VPWR.n1 VGND 0.1826f
C16458 VPWR.n2 VGND 0.09661f
C16459 VPWR.t503 VGND 0.05716f
C16460 VPWR.n3 VGND 0.0092f
C16461 VPWR.t993 VGND 0.01433f
C16462 VPWR.t1498 VGND 0.01433f
C16463 VPWR.n4 VGND 0.03146f
C16464 VPWR.t1502 VGND 0.01433f
C16465 VPWR.t989 VGND 0.01433f
C16466 VPWR.n5 VGND 0.03141f
C16467 VPWR.n6 VGND 0.0645f
C16468 VPWR.n7 VGND 0.18182f
C16469 VPWR.n8 VGND 0.05756f
C16470 VPWR.n9 VGND 0.04228f
C16471 VPWR.n10 VGND 0.07578f
C16472 VPWR.n11 VGND 0.01119f
C16473 VPWR.n12 VGND 0.0163f
C16474 VPWR.n13 VGND 0.0191f
C16475 VPWR.n14 VGND 0.02802f
C16476 VPWR.n15 VGND 0.08481f
C16477 VPWR.n16 VGND 0.01209f
C16478 VPWR.t1723 VGND 0.05714f
C16479 VPWR.n17 VGND 0.0735f
C16480 VPWR.n18 VGND 0.33563f
C16481 VPWR.n19 VGND 0.97868f
C16482 VPWR.n20 VGND 0.31857f
C16483 VPWR.n21 VGND 1.01577f
C16484 VPWR.n22 VGND 0.13887f
C16485 VPWR.t1970 VGND 0.0112f
C16486 VPWR.t298 VGND 0.01226f
C16487 VPWR.n23 VGND 0.02994f
C16488 VPWR.n24 VGND 0.07953f
C16489 VPWR.t2021 VGND 0.0112f
C16490 VPWR.t187 VGND 0.01226f
C16491 VPWR.n25 VGND 0.02994f
C16492 VPWR.n26 VGND 0.16006f
C16493 VPWR.t1956 VGND 0.0112f
C16494 VPWR.t335 VGND 0.01226f
C16495 VPWR.n27 VGND 0.02994f
C16496 VPWR.n28 VGND 0.12753f
C16497 VPWR.t1995 VGND 0.0112f
C16498 VPWR.t227 VGND 0.01226f
C16499 VPWR.n29 VGND 0.02994f
C16500 VPWR.n30 VGND 0.12753f
C16501 VPWR.t2064 VGND 0.0112f
C16502 VPWR.t40 VGND 0.01226f
C16503 VPWR.n31 VGND 0.02994f
C16504 VPWR.n32 VGND 0.12753f
C16505 VPWR.t1997 VGND 0.0112f
C16506 VPWR.t220 VGND 0.01226f
C16507 VPWR.n33 VGND 0.02994f
C16508 VPWR.n34 VGND 0.12753f
C16509 VPWR.t1943 VGND 0.0112f
C16510 VPWR.t115 VGND 0.01226f
C16511 VPWR.n35 VGND 0.02994f
C16512 VPWR.n36 VGND 0.12753f
C16513 VPWR.t2022 VGND 0.0112f
C16514 VPWR.t155 VGND 0.01226f
C16515 VPWR.n37 VGND 0.02994f
C16516 VPWR.n38 VGND 0.12753f
C16517 VPWR.t2028 VGND 0.0112f
C16518 VPWR.t48 VGND 0.01226f
C16519 VPWR.n39 VGND 0.02994f
C16520 VPWR.n40 VGND 0.12753f
C16521 VPWR.t2069 VGND 0.0112f
C16522 VPWR.t322 VGND 0.01226f
C16523 VPWR.n41 VGND 0.02994f
C16524 VPWR.n42 VGND 0.12753f
C16525 VPWR.t2051 VGND 0.0112f
C16526 VPWR.t214 VGND 0.01226f
C16527 VPWR.n43 VGND 0.02994f
C16528 VPWR.n44 VGND 0.12753f
C16529 VPWR.t1946 VGND 0.0112f
C16530 VPWR.t365 VGND 0.01226f
C16531 VPWR.n45 VGND 0.02994f
C16532 VPWR.n46 VGND 0.12753f
C16533 VPWR.t2026 VGND 0.0112f
C16534 VPWR.t147 VGND 0.01226f
C16535 VPWR.n47 VGND 0.02994f
C16536 VPWR.n48 VGND 0.12753f
C16537 VPWR.t2066 VGND 0.0112f
C16538 VPWR.t32 VGND 0.01226f
C16539 VPWR.n49 VGND 0.02994f
C16540 VPWR.n50 VGND 0.12753f
C16541 VPWR.t1963 VGND 0.0112f
C16542 VPWR.t317 VGND 0.01226f
C16543 VPWR.n51 VGND 0.02994f
C16544 VPWR.n52 VGND 0.12753f
C16545 VPWR.t2053 VGND 0.0112f
C16546 VPWR.t357 VGND 0.01226f
C16547 VPWR.n53 VGND 0.02994f
C16548 VPWR.n54 VGND 0.13808f
C16549 VPWR.n55 VGND 0.11528f
C16550 VPWR.t146 VGND 0.03331f
C16551 VPWR.t251 VGND 0.02961f
C16552 VPWR.n56 VGND 0.09152f
C16553 VPWR.t14 VGND 0.09218f
C16554 VPWR.t21 VGND 0.03331f
C16555 VPWR.t15 VGND 0.02961f
C16556 VPWR.n57 VGND 0.09152f
C16557 VPWR.n58 VGND 0.03437f
C16558 VPWR.n59 VGND 0.13913f
C16559 VPWR.n60 VGND 0.13913f
C16560 VPWR.n61 VGND 0.03437f
C16561 VPWR.t2 VGND 0.03331f
C16562 VPWR.t375 VGND 0.02961f
C16563 VPWR.n62 VGND 0.09152f
C16564 VPWR.t241 VGND 0.09218f
C16565 VPWR.t152 VGND 0.03331f
C16566 VPWR.t242 VGND 0.02961f
C16567 VPWR.n63 VGND 0.09152f
C16568 VPWR.n64 VGND 0.03437f
C16569 VPWR.n65 VGND 0.13913f
C16570 VPWR.n66 VGND 0.13913f
C16571 VPWR.n67 VGND 0.03437f
C16572 VPWR.t122 VGND 0.03331f
C16573 VPWR.t114 VGND 0.02961f
C16574 VPWR.n68 VGND 0.09152f
C16575 VPWR.t95 VGND 0.09218f
C16576 VPWR.t378 VGND 0.03331f
C16577 VPWR.t96 VGND 0.02961f
C16578 VPWR.n69 VGND 0.09152f
C16579 VPWR.n70 VGND 0.03437f
C16580 VPWR.n71 VGND 0.13913f
C16581 VPWR.n72 VGND 0.13913f
C16582 VPWR.n73 VGND 0.03437f
C16583 VPWR.t248 VGND 0.03331f
C16584 VPWR.t329 VGND 0.02961f
C16585 VPWR.n74 VGND 0.09152f
C16586 VPWR.t218 VGND 0.09218f
C16587 VPWR.t232 VGND 0.03331f
C16588 VPWR.t219 VGND 0.02961f
C16589 VPWR.n75 VGND 0.09152f
C16590 VPWR.n76 VGND 0.03437f
C16591 VPWR.n77 VGND 0.13913f
C16592 VPWR.n78 VGND 0.13913f
C16593 VPWR.n79 VGND 0.03437f
C16594 VPWR.t72 VGND 0.03331f
C16595 VPWR.t91 VGND 0.02961f
C16596 VPWR.n80 VGND 0.09152f
C16597 VPWR.t55 VGND 0.09218f
C16598 VPWR.t351 VGND 0.03331f
C16599 VPWR.t56 VGND 0.02961f
C16600 VPWR.n81 VGND 0.09152f
C16601 VPWR.n82 VGND 0.03437f
C16602 VPWR.n83 VGND 0.13913f
C16603 VPWR.n84 VGND 0.13913f
C16604 VPWR.n85 VGND 0.03437f
C16605 VPWR.t195 VGND 0.03331f
C16606 VPWR.t332 VGND 0.02961f
C16607 VPWR.n86 VGND 0.09152f
C16608 VPWR.t176 VGND 0.09218f
C16609 VPWR.t183 VGND 0.03331f
C16610 VPWR.t177 VGND 0.02961f
C16611 VPWR.n87 VGND 0.09152f
C16612 VPWR.n88 VGND 0.03437f
C16613 VPWR.n89 VGND 0.13913f
C16614 VPWR.n90 VGND 0.13913f
C16615 VPWR.n91 VGND 0.03437f
C16616 VPWR.t75 VGND 0.03331f
C16617 VPWR.t69 VGND 0.02961f
C16618 VPWR.n92 VGND 0.09152f
C16619 VPWR.t306 VGND 0.09218f
C16620 VPWR.t310 VGND 0.03331f
C16621 VPWR.t307 VGND 0.02961f
C16622 VPWR.n93 VGND 0.09152f
C16623 VPWR.n94 VGND 0.03437f
C16624 VPWR.n95 VGND 0.13913f
C16625 VPWR.n96 VGND 0.13913f
C16626 VPWR.n97 VGND 0.03437f
C16627 VPWR.t198 VGND 0.03331f
C16628 VPWR.t289 VGND 0.02961f
C16629 VPWR.n98 VGND 0.09152f
C16630 VPWR.t52 VGND 0.14512f
C16631 VPWR.t28 VGND 0.07849f
C16632 VPWR.t159 VGND 0.09218f
C16633 VPWR.t53 VGND 0.03331f
C16634 VPWR.t160 VGND 0.02961f
C16635 VPWR.n99 VGND 0.09152f
C16636 VPWR.t1987 VGND 0.0112f
C16637 VPWR.t287 VGND 0.01226f
C16638 VPWR.n100 VGND 0.02993f
C16639 VPWR.n101 VGND 0.03284f
C16640 VPWR.n102 VGND 0.00697f
C16641 VPWR.n103 VGND 0.01822f
C16642 VPWR.t2032 VGND 0.0112f
C16643 VPWR.t158 VGND 0.01226f
C16644 VPWR.n104 VGND 0.02993f
C16645 VPWR.n105 VGND 0.03284f
C16646 VPWR.t1981 VGND 0.01116f
C16647 VPWR.t51 VGND 0.01222f
C16648 VPWR.n106 VGND 0.03115f
C16649 VPWR.n107 VGND 0.01969f
C16650 VPWR.t1934 VGND 0.01136f
C16651 VPWR.t27 VGND 0.0124f
C16652 VPWR.n108 VGND 0.02768f
C16653 VPWR.n109 VGND 0.02818f
C16654 VPWR.n110 VGND 0.01776f
C16655 VPWR.n111 VGND 0.00697f
C16656 VPWR.n112 VGND 0.01822f
C16657 VPWR.n113 VGND 0.02654f
C16658 VPWR.t2001 VGND 0.0112f
C16659 VPWR.t249 VGND 0.01226f
C16660 VPWR.n114 VGND 0.02993f
C16661 VPWR.n115 VGND 0.03284f
C16662 VPWR.t1951 VGND 0.01116f
C16663 VPWR.t144 VGND 0.01222f
C16664 VPWR.n116 VGND 0.03115f
C16665 VPWR.n117 VGND 0.03694f
C16666 VPWR.n118 VGND 0.00833f
C16667 VPWR.t2048 VGND 0.01136f
C16668 VPWR.t128 VGND 0.0124f
C16669 VPWR.n119 VGND 0.02768f
C16670 VPWR.n120 VGND 0.02818f
C16671 VPWR.n121 VGND 0.01776f
C16672 VPWR.n122 VGND 0.00697f
C16673 VPWR.n123 VGND 0.01822f
C16674 VPWR.n124 VGND 0.02541f
C16675 VPWR.t1940 VGND 0.0112f
C16676 VPWR.t13 VGND 0.01226f
C16677 VPWR.n125 VGND 0.02993f
C16678 VPWR.n126 VGND 0.03284f
C16679 VPWR.t1991 VGND 0.01116f
C16680 VPWR.t19 VGND 0.01222f
C16681 VPWR.n127 VGND 0.03115f
C16682 VPWR.n128 VGND 0.03694f
C16683 VPWR.n129 VGND 0.00833f
C16684 VPWR.t1990 VGND 0.01136f
C16685 VPWR.t277 VGND 0.0124f
C16686 VPWR.n130 VGND 0.02768f
C16687 VPWR.n131 VGND 0.02818f
C16688 VPWR.n132 VGND 0.01776f
C16689 VPWR.n133 VGND 0.00697f
C16690 VPWR.n134 VGND 0.01822f
C16691 VPWR.n135 VGND 0.02384f
C16692 VPWR.n136 VGND 0.21163f
C16693 VPWR.t1954 VGND 0.0112f
C16694 VPWR.t373 VGND 0.01226f
C16695 VPWR.n137 VGND 0.02993f
C16696 VPWR.n138 VGND 0.03284f
C16697 VPWR.t2046 VGND 0.01116f
C16698 VPWR.t0 VGND 0.01222f
C16699 VPWR.n139 VGND 0.03115f
C16700 VPWR.n140 VGND 0.03694f
C16701 VPWR.n141 VGND 0.00833f
C16702 VPWR.t1999 VGND 0.01136f
C16703 VPWR.t252 VGND 0.0124f
C16704 VPWR.n142 VGND 0.02768f
C16705 VPWR.n143 VGND 0.02818f
C16706 VPWR.n144 VGND 0.01776f
C16707 VPWR.n145 VGND 0.00697f
C16708 VPWR.n146 VGND 0.01822f
C16709 VPWR.n147 VGND 0.02384f
C16710 VPWR.n148 VGND 0.17585f
C16711 VPWR.t2004 VGND 0.0112f
C16712 VPWR.t240 VGND 0.01226f
C16713 VPWR.n149 VGND 0.02993f
C16714 VPWR.n150 VGND 0.03284f
C16715 VPWR.t1942 VGND 0.01116f
C16716 VPWR.t150 VGND 0.01222f
C16717 VPWR.n151 VGND 0.03115f
C16718 VPWR.n152 VGND 0.03694f
C16719 VPWR.n153 VGND 0.00833f
C16720 VPWR.t2007 VGND 0.01136f
C16721 VPWR.t233 VGND 0.0124f
C16722 VPWR.n154 VGND 0.02768f
C16723 VPWR.n155 VGND 0.02818f
C16724 VPWR.n156 VGND 0.01776f
C16725 VPWR.n157 VGND 0.00697f
C16726 VPWR.n158 VGND 0.01822f
C16727 VPWR.n159 VGND 0.02384f
C16728 VPWR.n160 VGND 0.17585f
C16729 VPWR.t2052 VGND 0.0112f
C16730 VPWR.t112 VGND 0.01226f
C16731 VPWR.n161 VGND 0.02993f
C16732 VPWR.n162 VGND 0.03284f
C16733 VPWR.t1998 VGND 0.01116f
C16734 VPWR.t120 VGND 0.01222f
C16735 VPWR.n163 VGND 0.03115f
C16736 VPWR.n164 VGND 0.03694f
C16737 VPWR.n165 VGND 0.00833f
C16738 VPWR.t1952 VGND 0.01136f
C16739 VPWR.t379 VGND 0.0124f
C16740 VPWR.n166 VGND 0.02768f
C16741 VPWR.n167 VGND 0.02818f
C16742 VPWR.n168 VGND 0.01776f
C16743 VPWR.n169 VGND 0.00697f
C16744 VPWR.n170 VGND 0.01822f
C16745 VPWR.n171 VGND 0.02384f
C16746 VPWR.n172 VGND 0.17585f
C16747 VPWR.t2058 VGND 0.0112f
C16748 VPWR.t94 VGND 0.01226f
C16749 VPWR.n173 VGND 0.02993f
C16750 VPWR.n174 VGND 0.03284f
C16751 VPWR.t2006 VGND 0.01116f
C16752 VPWR.t376 VGND 0.01222f
C16753 VPWR.n175 VGND 0.03115f
C16754 VPWR.n176 VGND 0.03694f
C16755 VPWR.n177 VGND 0.00833f
C16756 VPWR.t1961 VGND 0.01136f
C16757 VPWR.t360 VGND 0.0124f
C16758 VPWR.n178 VGND 0.02768f
C16759 VPWR.n179 VGND 0.02818f
C16760 VPWR.n180 VGND 0.01776f
C16761 VPWR.n181 VGND 0.00697f
C16762 VPWR.n182 VGND 0.01822f
C16763 VPWR.n183 VGND 0.02384f
C16764 VPWR.n184 VGND 0.17585f
C16765 VPWR.t1973 VGND 0.0112f
C16766 VPWR.t327 VGND 0.01226f
C16767 VPWR.n185 VGND 0.02993f
C16768 VPWR.n186 VGND 0.03284f
C16769 VPWR.t2054 VGND 0.01116f
C16770 VPWR.t246 VGND 0.01222f
C16771 VPWR.n187 VGND 0.03115f
C16772 VPWR.n188 VGND 0.03694f
C16773 VPWR.n189 VGND 0.00833f
C16774 VPWR.t2017 VGND 0.01136f
C16775 VPWR.t199 VGND 0.0124f
C16776 VPWR.n190 VGND 0.02768f
C16777 VPWR.n191 VGND 0.02818f
C16778 VPWR.n192 VGND 0.01776f
C16779 VPWR.n193 VGND 0.00697f
C16780 VPWR.n194 VGND 0.01822f
C16781 VPWR.n195 VGND 0.02384f
C16782 VPWR.n196 VGND 0.17585f
C16783 VPWR.t2009 VGND 0.0112f
C16784 VPWR.t217 VGND 0.01226f
C16785 VPWR.n197 VGND 0.02993f
C16786 VPWR.n198 VGND 0.03284f
C16787 VPWR.t1960 VGND 0.01116f
C16788 VPWR.t230 VGND 0.01222f
C16789 VPWR.n199 VGND 0.03115f
C16790 VPWR.n200 VGND 0.03694f
C16791 VPWR.n201 VGND 0.00833f
C16792 VPWR.t2057 VGND 0.01136f
C16793 VPWR.t97 VGND 0.0124f
C16794 VPWR.n202 VGND 0.02768f
C16795 VPWR.n203 VGND 0.02818f
C16796 VPWR.n204 VGND 0.01776f
C16797 VPWR.n205 VGND 0.00697f
C16798 VPWR.n206 VGND 0.01822f
C16799 VPWR.n207 VGND 0.02384f
C16800 VPWR.n208 VGND 0.17585f
C16801 VPWR.t2060 VGND 0.0112f
C16802 VPWR.t89 VGND 0.01226f
C16803 VPWR.n209 VGND 0.02993f
C16804 VPWR.n210 VGND 0.03284f
C16805 VPWR.t1974 VGND 0.01116f
C16806 VPWR.t70 VGND 0.01222f
C16807 VPWR.n211 VGND 0.03115f
C16808 VPWR.n212 VGND 0.03694f
C16809 VPWR.n213 VGND 0.00833f
C16810 VPWR.t1928 VGND 0.01136f
C16811 VPWR.t62 VGND 0.0124f
C16812 VPWR.n214 VGND 0.02768f
C16813 VPWR.n215 VGND 0.02818f
C16814 VPWR.n216 VGND 0.01776f
C16815 VPWR.n217 VGND 0.00697f
C16816 VPWR.n218 VGND 0.01822f
C16817 VPWR.n219 VGND 0.02384f
C16818 VPWR.n220 VGND 0.17585f
C16819 VPWR.t1931 VGND 0.0112f
C16820 VPWR.t54 VGND 0.01226f
C16821 VPWR.n221 VGND 0.02993f
C16822 VPWR.n222 VGND 0.03284f
C16823 VPWR.t2056 VGND 0.01116f
C16824 VPWR.t349 VGND 0.01222f
C16825 VPWR.n223 VGND 0.03115f
C16826 VPWR.n224 VGND 0.03694f
C16827 VPWR.n225 VGND 0.00833f
C16828 VPWR.t2008 VGND 0.01136f
C16829 VPWR.t225 VGND 0.0124f
C16830 VPWR.n226 VGND 0.02768f
C16831 VPWR.n227 VGND 0.02818f
C16832 VPWR.n228 VGND 0.01776f
C16833 VPWR.n229 VGND 0.00697f
C16834 VPWR.n230 VGND 0.01822f
C16835 VPWR.n231 VGND 0.02384f
C16836 VPWR.n232 VGND 0.17585f
C16837 VPWR.t1972 VGND 0.0112f
C16838 VPWR.t330 VGND 0.01226f
C16839 VPWR.n233 VGND 0.02993f
C16840 VPWR.n234 VGND 0.03284f
C16841 VPWR.t1926 VGND 0.01116f
C16842 VPWR.t193 VGND 0.01222f
C16843 VPWR.n235 VGND 0.03115f
C16844 VPWR.n236 VGND 0.03694f
C16845 VPWR.n237 VGND 0.00833f
C16846 VPWR.t2016 VGND 0.01136f
C16847 VPWR.t201 VGND 0.0124f
C16848 VPWR.n238 VGND 0.02768f
C16849 VPWR.n239 VGND 0.02818f
C16850 VPWR.n240 VGND 0.01776f
C16851 VPWR.n241 VGND 0.00697f
C16852 VPWR.n242 VGND 0.01822f
C16853 VPWR.n243 VGND 0.02384f
C16854 VPWR.n244 VGND 0.17585f
C16855 VPWR.t2027 VGND 0.0112f
C16856 VPWR.t175 VGND 0.01226f
C16857 VPWR.n245 VGND 0.02993f
C16858 VPWR.n246 VGND 0.03284f
C16859 VPWR.t1932 VGND 0.01116f
C16860 VPWR.t181 VGND 0.01222f
C16861 VPWR.n247 VGND 0.03115f
C16862 VPWR.n248 VGND 0.03694f
C16863 VPWR.n249 VGND 0.00833f
C16864 VPWR.t1930 VGND 0.01136f
C16865 VPWR.t57 VGND 0.0124f
C16866 VPWR.n250 VGND 0.02768f
C16867 VPWR.n251 VGND 0.02818f
C16868 VPWR.n252 VGND 0.01776f
C16869 VPWR.n253 VGND 0.00697f
C16870 VPWR.n254 VGND 0.01822f
C16871 VPWR.n255 VGND 0.02384f
C16872 VPWR.n256 VGND 0.17585f
C16873 VPWR.t2068 VGND 0.0112f
C16874 VPWR.t67 VGND 0.01226f
C16875 VPWR.n257 VGND 0.02993f
C16876 VPWR.n258 VGND 0.03284f
C16877 VPWR.t2015 VGND 0.01116f
C16878 VPWR.t73 VGND 0.01222f
C16879 VPWR.n259 VGND 0.03115f
C16880 VPWR.n260 VGND 0.03694f
C16881 VPWR.n261 VGND 0.00833f
C16882 VPWR.t1971 VGND 0.01136f
C16883 VPWR.t333 VGND 0.0124f
C16884 VPWR.n262 VGND 0.02768f
C16885 VPWR.n263 VGND 0.02818f
C16886 VPWR.n264 VGND 0.01776f
C16887 VPWR.n265 VGND 0.00697f
C16888 VPWR.n266 VGND 0.01822f
C16889 VPWR.n267 VGND 0.02384f
C16890 VPWR.n268 VGND 0.17585f
C16891 VPWR.t1980 VGND 0.0112f
C16892 VPWR.t305 VGND 0.01226f
C16893 VPWR.n269 VGND 0.02993f
C16894 VPWR.n270 VGND 0.03284f
C16895 VPWR.t2029 VGND 0.01116f
C16896 VPWR.t308 VGND 0.01222f
C16897 VPWR.n271 VGND 0.03115f
C16898 VPWR.n272 VGND 0.03694f
C16899 VPWR.n273 VGND 0.00833f
C16900 VPWR.t1983 VGND 0.01136f
C16901 VPWR.t293 VGND 0.0124f
C16902 VPWR.n274 VGND 0.02768f
C16903 VPWR.n275 VGND 0.02818f
C16904 VPWR.n276 VGND 0.01776f
C16905 VPWR.n277 VGND 0.00697f
C16906 VPWR.n278 VGND 0.01822f
C16907 VPWR.n279 VGND 0.02384f
C16908 VPWR.n280 VGND 0.17585f
C16909 VPWR.n281 VGND 0.23724f
C16910 VPWR.n282 VGND 0.02384f
C16911 VPWR.n283 VGND 0.01776f
C16912 VPWR.t2030 VGND 0.01136f
C16913 VPWR.t163 VGND 0.0124f
C16914 VPWR.n284 VGND 0.02768f
C16915 VPWR.n285 VGND 0.02818f
C16916 VPWR.n286 VGND 0.00833f
C16917 VPWR.t1933 VGND 0.01116f
C16918 VPWR.t196 VGND 0.01222f
C16919 VPWR.n287 VGND 0.03115f
C16920 VPWR.n288 VGND 0.03694f
C16921 VPWR.n289 VGND 0.03437f
C16922 VPWR.t1426 VGND 0.03331f
C16923 VPWR.t1159 VGND 0.02961f
C16924 VPWR.n290 VGND 0.09152f
C16925 VPWR.t1425 VGND 0.14512f
C16926 VPWR.t1877 VGND 0.07849f
C16927 VPWR.t1158 VGND 0.09218f
C16928 VPWR.t625 VGND 0.03331f
C16929 VPWR.t359 VGND 0.02961f
C16930 VPWR.n291 VGND 0.09152f
C16931 VPWR.n292 VGND 0.01797f
C16932 VPWR.n293 VGND 0.07618f
C16933 VPWR.t358 VGND 0.13333f
C16934 VPWR.t1657 VGND 0.07849f
C16935 VPWR.t624 VGND 0.11957f
C16936 VPWR.t1469 VGND 0.03331f
C16937 VPWR.t749 VGND 0.02961f
C16938 VPWR.n294 VGND 0.09152f
C16939 VPWR.n295 VGND 0.01797f
C16940 VPWR.n296 VGND 0.00728f
C16941 VPWR.n297 VGND 0.10822f
C16942 VPWR.t748 VGND 0.09218f
C16943 VPWR.t804 VGND 0.07849f
C16944 VPWR.t1468 VGND 0.11957f
C16945 VPWR.t820 VGND 0.03331f
C16946 VPWR.t485 VGND 0.02961f
C16947 VPWR.n298 VGND 0.09152f
C16948 VPWR.n299 VGND 0.01797f
C16949 VPWR.n300 VGND 0.00728f
C16950 VPWR.n301 VGND 0.10822f
C16951 VPWR.t484 VGND 0.09218f
C16952 VPWR.t1193 VGND 0.07849f
C16953 VPWR.t819 VGND 0.11957f
C16954 VPWR.t1198 VGND 0.03331f
C16955 VPWR.t1699 VGND 0.02961f
C16956 VPWR.n302 VGND 0.09152f
C16957 VPWR.n303 VGND 0.01797f
C16958 VPWR.n304 VGND 0.00728f
C16959 VPWR.n305 VGND 0.10822f
C16960 VPWR.t1698 VGND 0.09218f
C16961 VPWR.t1194 VGND 0.07849f
C16962 VPWR.t1197 VGND 0.11957f
C16963 VPWR.t1048 VGND 0.03331f
C16964 VPWR.t1188 VGND 0.02961f
C16965 VPWR.n306 VGND 0.09152f
C16966 VPWR.n307 VGND 0.01797f
C16967 VPWR.n308 VGND 0.00728f
C16968 VPWR.n309 VGND 0.10822f
C16969 VPWR.t1187 VGND 0.09218f
C16970 VPWR.t1878 VGND 0.07849f
C16971 VPWR.t1047 VGND 0.11957f
C16972 VPWR.t1835 VGND 0.03331f
C16973 VPWR.t1054 VGND 0.02961f
C16974 VPWR.n310 VGND 0.09152f
C16975 VPWR.n311 VGND 0.01797f
C16976 VPWR.n312 VGND 0.00728f
C16977 VPWR.n313 VGND 0.10822f
C16978 VPWR.t1053 VGND 0.09218f
C16979 VPWR.t1879 VGND 0.07849f
C16980 VPWR.t1834 VGND 0.11957f
C16981 VPWR.t1015 VGND 0.03331f
C16982 VPWR.t647 VGND 0.02961f
C16983 VPWR.n314 VGND 0.09152f
C16984 VPWR.n315 VGND 0.01797f
C16985 VPWR.n316 VGND 0.00728f
C16986 VPWR.n317 VGND 0.10822f
C16987 VPWR.t646 VGND 0.09218f
C16988 VPWR.t1655 VGND 0.07849f
C16989 VPWR.t1014 VGND 0.11957f
C16990 VPWR.t1113 VGND 0.03331f
C16991 VPWR.t1917 VGND 0.02961f
C16992 VPWR.n318 VGND 0.09152f
C16993 VPWR.n319 VGND 0.01797f
C16994 VPWR.n320 VGND 0.00728f
C16995 VPWR.n321 VGND 0.10822f
C16996 VPWR.t1916 VGND 0.09218f
C16997 VPWR.t1658 VGND 0.07849f
C16998 VPWR.t1112 VGND 0.11957f
C16999 VPWR.t719 VGND 0.03331f
C17000 VPWR.t904 VGND 0.02961f
C17001 VPWR.n322 VGND 0.09152f
C17002 VPWR.n323 VGND 0.01797f
C17003 VPWR.n324 VGND 0.00728f
C17004 VPWR.n325 VGND 0.10822f
C17005 VPWR.t903 VGND 0.09218f
C17006 VPWR.t1659 VGND 0.07849f
C17007 VPWR.t718 VGND 0.11957f
C17008 VPWR.t536 VGND 0.03331f
C17009 VPWR.t725 VGND 0.02961f
C17010 VPWR.n326 VGND 0.09152f
C17011 VPWR.n327 VGND 0.01797f
C17012 VPWR.n328 VGND 0.00728f
C17013 VPWR.n329 VGND 0.10822f
C17014 VPWR.t724 VGND 0.09218f
C17015 VPWR.t1653 VGND 0.07849f
C17016 VPWR.t535 VGND 0.11957f
C17017 VPWR.t1714 VGND 0.03331f
C17018 VPWR.t542 VGND 0.02961f
C17019 VPWR.n330 VGND 0.09152f
C17020 VPWR.n331 VGND 0.01797f
C17021 VPWR.n332 VGND 0.00728f
C17022 VPWR.n333 VGND 0.10822f
C17023 VPWR.t541 VGND 0.09218f
C17024 VPWR.t1654 VGND 0.07849f
C17025 VPWR.t1713 VGND 0.11957f
C17026 VPWR.t1060 VGND 0.03331f
C17027 VPWR.t1720 VGND 0.02961f
C17028 VPWR.n334 VGND 0.09152f
C17029 VPWR.n335 VGND 0.01797f
C17030 VPWR.n336 VGND 0.00728f
C17031 VPWR.n337 VGND 0.10822f
C17032 VPWR.t1719 VGND 0.09218f
C17033 VPWR.t1876 VGND 0.07849f
C17034 VPWR.t1059 VGND 0.11957f
C17035 VPWR.t1381 VGND 0.03331f
C17036 VPWR.t1192 VGND 0.02961f
C17037 VPWR.n338 VGND 0.09152f
C17038 VPWR.n339 VGND 0.01797f
C17039 VPWR.n340 VGND 0.00728f
C17040 VPWR.n341 VGND 0.10822f
C17041 VPWR.t1191 VGND 0.09218f
C17042 VPWR.t1880 VGND 0.07849f
C17043 VPWR.t1380 VGND 0.11957f
C17044 VPWR.t422 VGND 0.03331f
C17045 VPWR.t1357 VGND 0.02961f
C17046 VPWR.n342 VGND 0.09152f
C17047 VPWR.n343 VGND 0.01797f
C17048 VPWR.n344 VGND 0.00728f
C17049 VPWR.n345 VGND 0.10822f
C17050 VPWR.t1356 VGND 0.09218f
C17051 VPWR.t1881 VGND 0.07849f
C17052 VPWR.t421 VGND 0.11957f
C17053 VPWR.t1129 VGND 0.03331f
C17054 VPWR.t1608 VGND 0.02961f
C17055 VPWR.n346 VGND 0.09152f
C17056 VPWR.n347 VGND 0.01797f
C17057 VPWR.n348 VGND 0.00728f
C17058 VPWR.n349 VGND 0.10822f
C17059 VPWR.t1607 VGND 0.09218f
C17060 VPWR.t1656 VGND 0.07849f
C17061 VPWR.t1128 VGND 0.11957f
C17062 VPWR.n350 VGND 0.10822f
C17063 VPWR.n351 VGND 0.00728f
C17064 VPWR.n352 VGND 0.01797f
C17065 VPWR.n353 VGND 0.13913f
C17066 VPWR.n354 VGND 1.0094f
C17067 VPWR.n355 VGND 0.13913f
C17068 VPWR.t1419 VGND 0.03331f
C17069 VPWR.t973 VGND 0.02961f
C17070 VPWR.n356 VGND 0.09152f
C17071 VPWR.t1418 VGND 0.14512f
C17072 VPWR.t1279 VGND 0.07849f
C17073 VPWR.t972 VGND 0.09218f
C17074 VPWR.t1611 VGND 0.11957f
C17075 VPWR.t1155 VGND 0.03331f
C17076 VPWR.t836 VGND 0.02961f
C17077 VPWR.n357 VGND 0.09152f
C17078 VPWR.n358 VGND 0.13913f
C17079 VPWR.n359 VGND 0.13913f
C17080 VPWR.t1612 VGND 0.03331f
C17081 VPWR.t1349 VGND 0.02961f
C17082 VPWR.n360 VGND 0.09152f
C17083 VPWR.t498 VGND 0.07849f
C17084 VPWR.t1348 VGND 0.09218f
C17085 VPWR.t1067 VGND 0.11957f
C17086 VPWR.t1373 VGND 0.03331f
C17087 VPWR.t1637 VGND 0.02961f
C17088 VPWR.n361 VGND 0.09152f
C17089 VPWR.n362 VGND 0.13913f
C17090 VPWR.n363 VGND 0.13913f
C17091 VPWR.t1068 VGND 0.03331f
C17092 VPWR.t1553 VGND 0.02961f
C17093 VPWR.n364 VGND 0.09152f
C17094 VPWR.t1278 VGND 0.07849f
C17095 VPWR.t1552 VGND 0.09218f
C17096 VPWR.t545 VGND 0.11957f
C17097 VPWR.t1547 VGND 0.03331f
C17098 VPWR.t689 VGND 0.02961f
C17099 VPWR.n365 VGND 0.09152f
C17100 VPWR.n366 VGND 0.13913f
C17101 VPWR.n367 VGND 0.13913f
C17102 VPWR.t546 VGND 0.03331f
C17103 VPWR.t1793 VGND 0.02961f
C17104 VPWR.n368 VGND 0.09152f
C17105 VPWR.t1660 VGND 0.07849f
C17106 VPWR.t1792 VGND 0.09218f
C17107 VPWR.t1020 VGND 0.11957f
C17108 VPWR.t729 VGND 0.03331f
C17109 VPWR.t914 VGND 0.02961f
C17110 VPWR.n369 VGND 0.09152f
C17111 VPWR.n370 VGND 0.13913f
C17112 VPWR.n371 VGND 0.13913f
C17113 VPWR.t1021 VGND 0.03331f
C17114 VPWR.t1482 VGND 0.02961f
C17115 VPWR.n372 VGND 0.09152f
C17116 VPWR.t1276 VGND 0.07849f
C17117 VPWR.t1481 VGND 0.09218f
C17118 VPWR.t642 VGND 0.11957f
C17119 VPWR.t1921 VGND 0.03331f
C17120 VPWR.t653 VGND 0.02961f
C17121 VPWR.n373 VGND 0.09152f
C17122 VPWR.n374 VGND 0.13913f
C17123 VPWR.n375 VGND 0.13913f
C17124 VPWR.t643 VGND 0.03331f
C17125 VPWR.t1105 VGND 0.02961f
C17126 VPWR.n376 VGND 0.09152f
C17127 VPWR.t1532 VGND 0.07849f
C17128 VPWR.t1104 VGND 0.09218f
C17129 VPWR.t1183 VGND 0.11957f
C17130 VPWR.t1099 VGND 0.03331f
C17131 VPWR.t1462 VGND 0.02961f
C17132 VPWR.n377 VGND 0.09152f
C17133 VPWR.n378 VGND 0.13913f
C17134 VPWR.n379 VGND 0.13913f
C17135 VPWR.t1184 VGND 0.03331f
C17136 VPWR.t1709 VGND 0.02961f
C17137 VPWR.n380 VGND 0.09152f
C17138 VPWR.t501 VGND 0.07849f
C17139 VPWR.t1708 VGND 0.09218f
C17140 VPWR.t682 VGND 0.11957f
C17141 VPWR.t925 VGND 0.03331f
C17142 VPWR.t861 VGND 0.02961f
C17143 VPWR.n381 VGND 0.09152f
C17144 VPWR.n382 VGND 0.13913f
C17145 VPWR.n383 VGND 0.13913f
C17146 VPWR.t683 VGND 0.03331f
C17147 VPWR.t761 VGND 0.02961f
C17148 VPWR.n384 VGND 0.09152f
C17149 VPWR.t499 VGND 0.07849f
C17150 VPWR.t760 VGND 0.09218f
C17151 VPWR.t633 VGND 0.03331f
C17152 VPWR.t319 VGND 0.02961f
C17153 VPWR.n385 VGND 0.09152f
C17154 VPWR.t1815 VGND 0.03331f
C17155 VPWR.t34 VGND 0.02961f
C17156 VPWR.n386 VGND 0.09152f
C17157 VPWR.t1429 VGND 0.14512f
C17158 VPWR.t1673 VGND 0.07849f
C17159 VPWR.t1124 VGND 0.09218f
C17160 VPWR.t1430 VGND 0.03331f
C17161 VPWR.t1125 VGND 0.02961f
C17162 VPWR.n387 VGND 0.09152f
C17163 VPWR.n388 VGND 0.01797f
C17164 VPWR.n389 VGND 0.00728f
C17165 VPWR.n390 VGND 0.10822f
C17166 VPWR.t1728 VGND 0.11957f
C17167 VPWR.t1225 VGND 0.07849f
C17168 VPWR.t1006 VGND 0.09218f
C17169 VPWR.t1729 VGND 0.03331f
C17170 VPWR.t1007 VGND 0.02961f
C17171 VPWR.n391 VGND 0.09152f
C17172 VPWR.n392 VGND 0.01797f
C17173 VPWR.n393 VGND 0.00728f
C17174 VPWR.n394 VGND 0.10822f
C17175 VPWR.t1587 VGND 0.11957f
C17176 VPWR.t1230 VGND 0.07849f
C17177 VPWR.t1366 VGND 0.09218f
C17178 VPWR.t1588 VGND 0.03331f
C17179 VPWR.t1367 VGND 0.02961f
C17180 VPWR.n395 VGND 0.09152f
C17181 VPWR.n396 VGND 0.01797f
C17182 VPWR.n397 VGND 0.00728f
C17183 VPWR.n398 VGND 0.10822f
C17184 VPWR.t1390 VGND 0.11957f
C17185 VPWR.t1229 VGND 0.07849f
C17186 VPWR.t1071 VGND 0.09218f
C17187 VPWR.t1391 VGND 0.03331f
C17188 VPWR.t1072 VGND 0.02961f
C17189 VPWR.n399 VGND 0.09152f
C17190 VPWR.n400 VGND 0.01797f
C17191 VPWR.n401 VGND 0.00728f
C17192 VPWR.n402 VGND 0.10822f
C17193 VPWR.t1855 VGND 0.11957f
C17194 VPWR.t1672 VGND 0.07849f
C17195 VPWR.t1563 VGND 0.09218f
C17196 VPWR.t1856 VGND 0.03331f
C17197 VPWR.t1564 VGND 0.02961f
C17198 VPWR.n403 VGND 0.09152f
C17199 VPWR.n404 VGND 0.01797f
C17200 VPWR.n405 VGND 0.00728f
C17201 VPWR.n406 VGND 0.10822f
C17202 VPWR.t1536 VGND 0.11957f
C17203 VPWR.t1677 VGND 0.07849f
C17204 VPWR.t706 VGND 0.09218f
C17205 VPWR.t1537 VGND 0.03331f
C17206 VPWR.t707 VGND 0.02961f
C17207 VPWR.n407 VGND 0.09152f
C17208 VPWR.n408 VGND 0.01797f
C17209 VPWR.n409 VGND 0.00728f
C17210 VPWR.n410 VGND 0.10822f
C17211 VPWR.t595 VGND 0.11957f
C17212 VPWR.t1676 VGND 0.07849f
C17213 VPWR.t1908 VGND 0.09218f
C17214 VPWR.t596 VGND 0.03331f
C17215 VPWR.t1909 VGND 0.02961f
C17216 VPWR.n411 VGND 0.09152f
C17217 VPWR.n412 VGND 0.01797f
C17218 VPWR.n413 VGND 0.00728f
C17219 VPWR.n414 VGND 0.10822f
C17220 VPWR.t1902 VGND 0.11957f
C17221 VPWR.t1671 VGND 0.07849f
C17222 VPWR.t386 VGND 0.09218f
C17223 VPWR.t1903 VGND 0.03331f
C17224 VPWR.t387 VGND 0.02961f
C17225 VPWR.n415 VGND 0.09152f
C17226 VPWR.n416 VGND 0.01797f
C17227 VPWR.n417 VGND 0.00728f
C17228 VPWR.n418 VGND 0.10822f
C17229 VPWR.t866 VGND 0.11957f
C17230 VPWR.t1227 VGND 0.07849f
C17231 VPWR.t1010 VGND 0.09218f
C17232 VPWR.t867 VGND 0.03331f
C17233 VPWR.t1011 VGND 0.02961f
C17234 VPWR.n419 VGND 0.09152f
C17235 VPWR.n420 VGND 0.01797f
C17236 VPWR.n421 VGND 0.00728f
C17237 VPWR.n422 VGND 0.10822f
C17238 VPWR.t1603 VGND 0.11957f
C17239 VPWR.t1678 VGND 0.07849f
C17240 VPWR.t1830 VGND 0.09218f
C17241 VPWR.t1604 VGND 0.03331f
C17242 VPWR.t1831 VGND 0.02961f
C17243 VPWR.n423 VGND 0.09152f
C17244 VPWR.n424 VGND 0.01797f
C17245 VPWR.n425 VGND 0.00728f
C17246 VPWR.n426 VGND 0.10822f
C17247 VPWR.t1824 VGND 0.11957f
C17248 VPWR.t1228 VGND 0.07849f
C17249 VPWR.t1479 VGND 0.09218f
C17250 VPWR.t1825 VGND 0.03331f
C17251 VPWR.t1480 VGND 0.02961f
C17252 VPWR.n427 VGND 0.09152f
C17253 VPWR.n428 VGND 0.01797f
C17254 VPWR.n429 VGND 0.00728f
C17255 VPWR.n430 VGND 0.10822f
C17256 VPWR.t1473 VGND 0.11957f
C17257 VPWR.t1674 VGND 0.07849f
C17258 VPWR.t1245 VGND 0.09218f
C17259 VPWR.t1474 VGND 0.03331f
C17260 VPWR.t1246 VGND 0.02961f
C17261 VPWR.n431 VGND 0.09152f
C17262 VPWR.n432 VGND 0.01797f
C17263 VPWR.n433 VGND 0.00728f
C17264 VPWR.n434 VGND 0.10822f
C17265 VPWR.t1239 VGND 0.11957f
C17266 VPWR.t1675 VGND 0.07849f
C17267 VPWR.t930 VGND 0.09218f
C17268 VPWR.t1240 VGND 0.03331f
C17269 VPWR.t931 VGND 0.02961f
C17270 VPWR.n435 VGND 0.09152f
C17271 VPWR.n436 VGND 0.01797f
C17272 VPWR.n437 VGND 0.00728f
C17273 VPWR.n438 VGND 0.10822f
C17274 VPWR.t809 VGND 0.11957f
C17275 VPWR.t1232 VGND 0.07849f
C17276 VPWR.t513 VGND 0.09218f
C17277 VPWR.t810 VGND 0.03331f
C17278 VPWR.t514 VGND 0.02961f
C17279 VPWR.n439 VGND 0.09152f
C17280 VPWR.n440 VGND 0.01797f
C17281 VPWR.n441 VGND 0.00728f
C17282 VPWR.n442 VGND 0.10822f
C17283 VPWR.t1001 VGND 0.11957f
C17284 VPWR.t1231 VGND 0.07849f
C17285 VPWR.t636 VGND 0.09218f
C17286 VPWR.t1002 VGND 0.03331f
C17287 VPWR.t637 VGND 0.02961f
C17288 VPWR.n443 VGND 0.09152f
C17289 VPWR.n444 VGND 0.01797f
C17290 VPWR.n445 VGND 0.00728f
C17291 VPWR.n446 VGND 0.10822f
C17292 VPWR.t1814 VGND 0.11957f
C17293 VPWR.t1226 VGND 0.07849f
C17294 VPWR.t33 VGND 0.13333f
C17295 VPWR.n447 VGND 0.07618f
C17296 VPWR.n448 VGND 0.01797f
C17297 VPWR.n449 VGND 0.13913f
C17298 VPWR.n450 VGND 1.01577f
C17299 VPWR.n451 VGND 0.13913f
C17300 VPWR.t695 VGND 0.03331f
C17301 VPWR.t149 VGND 0.02961f
C17302 VPWR.n452 VGND 0.09152f
C17303 VPWR.t1816 VGND 0.09218f
C17304 VPWR.t1492 VGND 0.03331f
C17305 VPWR.t1817 VGND 0.02961f
C17306 VPWR.n453 VGND 0.09152f
C17307 VPWR.n454 VGND 0.13913f
C17308 VPWR.n455 VGND 0.13913f
C17309 VPWR.t454 VGND 0.03331f
C17310 VPWR.t1618 VGND 0.02961f
C17311 VPWR.n456 VGND 0.09152f
C17312 VPWR.t813 VGND 0.09218f
C17313 VPWR.t472 VGND 0.03331f
C17314 VPWR.t814 VGND 0.02961f
C17315 VPWR.n457 VGND 0.09152f
C17316 VPWR.n458 VGND 0.13913f
C17317 VPWR.n459 VGND 0.13913f
C17318 VPWR.t1578 VGND 0.03331f
C17319 VPWR.t1759 VGND 0.02961f
C17320 VPWR.n460 VGND 0.09152f
C17321 VPWR.t1581 VGND 0.09218f
C17322 VPWR.t665 VGND 0.03331f
C17323 VPWR.t1582 VGND 0.02961f
C17324 VPWR.n461 VGND 0.09152f
C17325 VPWR.n462 VGND 0.13913f
C17326 VPWR.n463 VGND 0.13913f
C17327 VPWR.t480 VGND 0.03331f
C17328 VPWR.t673 VGND 0.02961f
C17329 VPWR.n464 VGND 0.09152f
C17330 VPWR.t1116 VGND 0.09218f
C17331 VPWR.t859 VGND 0.03331f
C17332 VPWR.t1117 VGND 0.02961f
C17333 VPWR.n465 VGND 0.09152f
C17334 VPWR.n466 VGND 0.13913f
C17335 VPWR.n467 VGND 0.13913f
C17336 VPWR.t737 VGND 0.03331f
C17337 VPWR.t871 VGND 0.02961f
C17338 VPWR.n468 VGND 0.09152f
C17339 VPWR.t1892 VGND 0.09218f
C17340 VPWR.t964 VGND 0.03331f
C17341 VPWR.t1893 VGND 0.02961f
C17342 VPWR.n469 VGND 0.09152f
C17343 VPWR.n470 VGND 0.13913f
C17344 VPWR.n471 VGND 0.13913f
C17345 VPWR.t1568 VGND 0.03331f
C17346 VPWR.t968 VGND 0.02961f
C17347 VPWR.n472 VGND 0.09152f
C17348 VPWR.t1571 VGND 0.09218f
C17349 VPWR.t1028 VGND 0.03331f
C17350 VPWR.t1572 VGND 0.02961f
C17351 VPWR.n473 VGND 0.09152f
C17352 VPWR.n474 VGND 0.13913f
C17353 VPWR.n475 VGND 0.13913f
C17354 VPWR.t1407 VGND 0.03331f
C17355 VPWR.t1858 VGND 0.02961f
C17356 VPWR.n476 VGND 0.09152f
C17357 VPWR.t1384 VGND 0.09218f
C17358 VPWR.t842 VGND 0.03331f
C17359 VPWR.t1385 VGND 0.02961f
C17360 VPWR.n477 VGND 0.09152f
C17361 VPWR.n478 VGND 0.13913f
C17362 VPWR.n479 VGND 0.13913f
C17363 VPWR.t711 VGND 0.03331f
C17364 VPWR.t1520 VGND 0.02961f
C17365 VPWR.n480 VGND 0.09152f
C17366 VPWR.t1437 VGND 0.14512f
C17367 VPWR.t1097 VGND 0.07849f
C17368 VPWR.t831 VGND 0.09218f
C17369 VPWR.t1438 VGND 0.03331f
C17370 VPWR.t832 VGND 0.02961f
C17371 VPWR.n481 VGND 0.09152f
C17372 VPWR.t1428 VGND 0.03331f
C17373 VPWR.t1157 VGND 0.02961f
C17374 VPWR.n482 VGND 0.09152f
C17375 VPWR.t1427 VGND 0.14512f
C17376 VPWR.t1233 VGND 0.07849f
C17377 VPWR.t1156 VGND 0.09218f
C17378 VPWR.t623 VGND 0.03331f
C17379 VPWR.t367 VGND 0.02961f
C17380 VPWR.n483 VGND 0.09152f
C17381 VPWR.n484 VGND 0.01797f
C17382 VPWR.n485 VGND 0.07618f
C17383 VPWR.t366 VGND 0.13333f
C17384 VPWR.t1555 VGND 0.07849f
C17385 VPWR.t622 VGND 0.11957f
C17386 VPWR.t1467 VGND 0.03331f
C17387 VPWR.t747 VGND 0.02961f
C17388 VPWR.n486 VGND 0.09152f
C17389 VPWR.n487 VGND 0.01797f
C17390 VPWR.n488 VGND 0.00728f
C17391 VPWR.n489 VGND 0.10822f
C17392 VPWR.t746 VGND 0.09218f
C17393 VPWR.t1238 VGND 0.07849f
C17394 VPWR.t1466 VGND 0.11957f
C17395 VPWR.t816 VGND 0.03331f
C17396 VPWR.t685 VGND 0.02961f
C17397 VPWR.n490 VGND 0.09152f
C17398 VPWR.n491 VGND 0.01797f
C17399 VPWR.n492 VGND 0.00728f
C17400 VPWR.n493 VGND 0.10822f
C17401 VPWR.t684 VGND 0.09218f
C17402 VPWR.t1449 VGND 0.07849f
C17403 VPWR.t815 VGND 0.11957f
C17404 VPWR.t1196 VGND 0.03331f
C17405 VPWR.t1695 VGND 0.02961f
C17406 VPWR.n494 VGND 0.09152f
C17407 VPWR.n495 VGND 0.01797f
C17408 VPWR.n496 VGND 0.00728f
C17409 VPWR.n497 VGND 0.10822f
C17410 VPWR.t1694 VGND 0.09218f
C17411 VPWR.t1450 VGND 0.07849f
C17412 VPWR.t1195 VGND 0.11957f
C17413 VPWR.t1046 VGND 0.03331f
C17414 VPWR.t1186 VGND 0.02961f
C17415 VPWR.n498 VGND 0.09152f
C17416 VPWR.n499 VGND 0.01797f
C17417 VPWR.n500 VGND 0.00728f
C17418 VPWR.n501 VGND 0.10822f
C17419 VPWR.t1185 VGND 0.09218f
C17420 VPWR.t1234 VGND 0.07849f
C17421 VPWR.t1045 VGND 0.11957f
C17422 VPWR.t1833 VGND 0.03331f
C17423 VPWR.t1050 VGND 0.02961f
C17424 VPWR.n502 VGND 0.09152f
C17425 VPWR.n503 VGND 0.01797f
C17426 VPWR.n504 VGND 0.00728f
C17427 VPWR.n505 VGND 0.10822f
C17428 VPWR.t1049 VGND 0.09218f
C17429 VPWR.t1235 VGND 0.07849f
C17430 VPWR.t1832 VGND 0.11957f
C17431 VPWR.t1013 VGND 0.03331f
C17432 VPWR.t645 VGND 0.02961f
C17433 VPWR.n506 VGND 0.09152f
C17434 VPWR.n507 VGND 0.01797f
C17435 VPWR.n508 VGND 0.00728f
C17436 VPWR.n509 VGND 0.10822f
C17437 VPWR.t644 VGND 0.09218f
C17438 VPWR.t1453 VGND 0.07849f
C17439 VPWR.t1012 VGND 0.11957f
C17440 VPWR.t1109 VGND 0.03331f
C17441 VPWR.t1913 VGND 0.02961f
C17442 VPWR.n510 VGND 0.09152f
C17443 VPWR.n511 VGND 0.01797f
C17444 VPWR.n512 VGND 0.00728f
C17445 VPWR.n513 VGND 0.10822f
C17446 VPWR.t1912 VGND 0.09218f
C17447 VPWR.t1556 VGND 0.07849f
C17448 VPWR.t1108 VGND 0.11957f
C17449 VPWR.t717 VGND 0.03331f
C17450 VPWR.t918 VGND 0.02961f
C17451 VPWR.n514 VGND 0.09152f
C17452 VPWR.n515 VGND 0.01797f
C17453 VPWR.n516 VGND 0.00728f
C17454 VPWR.n517 VGND 0.10822f
C17455 VPWR.t917 VGND 0.09218f
C17456 VPWR.t1557 VGND 0.07849f
C17457 VPWR.t716 VGND 0.11957f
C17458 VPWR.t709 VGND 0.03331f
C17459 VPWR.t721 VGND 0.02961f
C17460 VPWR.n518 VGND 0.09152f
C17461 VPWR.n519 VGND 0.01797f
C17462 VPWR.n520 VGND 0.00728f
C17463 VPWR.n521 VGND 0.10822f
C17464 VPWR.t720 VGND 0.09218f
C17465 VPWR.t1451 VGND 0.07849f
C17466 VPWR.t708 VGND 0.11957f
C17467 VPWR.t828 VGND 0.03331f
C17468 VPWR.t538 VGND 0.02961f
C17469 VPWR.n522 VGND 0.09152f
C17470 VPWR.n523 VGND 0.01797f
C17471 VPWR.n524 VGND 0.00728f
C17472 VPWR.n525 VGND 0.10822f
C17473 VPWR.t537 VGND 0.09218f
C17474 VPWR.t1452 VGND 0.07849f
C17475 VPWR.t827 VGND 0.11957f
C17476 VPWR.t1058 VGND 0.03331f
C17477 VPWR.t1716 VGND 0.02961f
C17478 VPWR.n526 VGND 0.09152f
C17479 VPWR.n527 VGND 0.01797f
C17480 VPWR.n528 VGND 0.00728f
C17481 VPWR.n529 VGND 0.10822f
C17482 VPWR.t1715 VGND 0.09218f
C17483 VPWR.t1558 VGND 0.07849f
C17484 VPWR.t1057 VGND 0.11957f
C17485 VPWR.t1383 VGND 0.03331f
C17486 VPWR.t1190 VGND 0.02961f
C17487 VPWR.n530 VGND 0.09152f
C17488 VPWR.n531 VGND 0.01797f
C17489 VPWR.n532 VGND 0.00728f
C17490 VPWR.n533 VGND 0.10822f
C17491 VPWR.t1189 VGND 0.09218f
C17492 VPWR.t1236 VGND 0.07849f
C17493 VPWR.t1382 VGND 0.11957f
C17494 VPWR.t420 VGND 0.03331f
C17495 VPWR.t1359 VGND 0.02961f
C17496 VPWR.n534 VGND 0.09152f
C17497 VPWR.n535 VGND 0.01797f
C17498 VPWR.n536 VGND 0.00728f
C17499 VPWR.n537 VGND 0.10822f
C17500 VPWR.t1358 VGND 0.09218f
C17501 VPWR.t1237 VGND 0.07849f
C17502 VPWR.t419 VGND 0.11957f
C17503 VPWR.t1127 VGND 0.03331f
C17504 VPWR.t424 VGND 0.02961f
C17505 VPWR.n538 VGND 0.09152f
C17506 VPWR.n539 VGND 0.01797f
C17507 VPWR.n540 VGND 0.00728f
C17508 VPWR.n541 VGND 0.10822f
C17509 VPWR.t423 VGND 0.09218f
C17510 VPWR.t1554 VGND 0.07849f
C17511 VPWR.t1126 VGND 0.11957f
C17512 VPWR.n542 VGND 0.10822f
C17513 VPWR.n543 VGND 0.00728f
C17514 VPWR.n544 VGND 0.01797f
C17515 VPWR.n545 VGND 0.13913f
C17516 VPWR.n546 VGND 1.0094f
C17517 VPWR.n547 VGND 0.13913f
C17518 VPWR.t1413 VGND 0.03331f
C17519 VPWR.t900 VGND 0.02961f
C17520 VPWR.n548 VGND 0.09152f
C17521 VPWR.t1412 VGND 0.14512f
C17522 VPWR.t1274 VGND 0.07849f
C17523 VPWR.t899 VGND 0.09218f
C17524 VPWR.t1597 VGND 0.11957f
C17525 VPWR.t534 VGND 0.03331f
C17526 VPWR.t1087 VGND 0.02961f
C17527 VPWR.n549 VGND 0.09152f
C17528 VPWR.n550 VGND 0.13913f
C17529 VPWR.n551 VGND 0.13913f
C17530 VPWR.t1598 VGND 0.03331f
C17531 VPWR.t1397 VGND 0.02961f
C17532 VPWR.n552 VGND 0.09152f
C17533 VPWR.t430 VGND 0.07849f
C17534 VPWR.t1396 VGND 0.09218f
C17535 VPWR.t1632 VGND 0.11957f
C17536 VPWR.t1361 VGND 0.03331f
C17537 VPWR.t1036 VGND 0.02961f
C17538 VPWR.n553 VGND 0.09152f
C17539 VPWR.n554 VGND 0.13913f
C17540 VPWR.n555 VGND 0.13913f
C17541 VPWR.t1633 VGND 0.03331f
C17542 VPWR.t518 VGND 0.02961f
C17543 VPWR.n556 VGND 0.09152f
C17544 VPWR.t1273 VGND 0.07849f
C17545 VPWR.t517 VGND 0.09218f
C17546 VPWR.t559 VGND 0.11957f
C17547 VPWR.t1514 VGND 0.03331f
C17548 VPWR.t568 VGND 0.02961f
C17549 VPWR.n557 VGND 0.09152f
C17550 VPWR.n558 VGND 0.13913f
C17551 VPWR.n559 VGND 0.13913f
C17552 VPWR.t560 VGND 0.03331f
C17553 VPWR.t743 VGND 0.02961f
C17554 VPWR.n560 VGND 0.09152f
C17555 VPWR.t1218 VGND 0.07849f
C17556 VPWR.t742 VGND 0.09218f
C17557 VPWR.t905 VGND 0.11957f
C17558 VPWR.t1801 VGND 0.03331f
C17559 VPWR.t574 VGND 0.02961f
C17560 VPWR.n561 VGND 0.09152f
C17561 VPWR.n562 VGND 0.13913f
C17562 VPWR.n563 VGND 0.13913f
C17563 VPWR.t906 VGND 0.03331f
C17564 VPWR.t960 VGND 0.02961f
C17565 VPWR.n564 VGND 0.09152f
C17566 VPWR.t1271 VGND 0.07849f
C17567 VPWR.t959 VGND 0.09218f
C17568 VPWR.t612 VGND 0.11957f
C17569 VPWR.t952 VGND 0.03331f
C17570 VPWR.t621 VGND 0.02961f
C17571 VPWR.n565 VGND 0.09152f
C17572 VPWR.n566 VGND 0.13913f
C17573 VPWR.n567 VGND 0.13913f
C17574 VPWR.t613 VGND 0.03331f
C17575 VPWR.t1689 VGND 0.02961f
C17576 VPWR.n568 VGND 0.09152f
C17577 VPWR.t428 VGND 0.07849f
C17578 VPWR.t1688 VGND 0.09218f
C17579 VPWR.t1762 VGND 0.11957f
C17580 VPWR.t1681 VGND 0.03331f
C17581 VPWR.t468 VGND 0.02961f
C17582 VPWR.n569 VGND 0.09152f
C17583 VPWR.n570 VGND 0.13913f
C17584 VPWR.n571 VGND 0.13913f
C17585 VPWR.t1763 VGND 0.03331f
C17586 VPWR.t462 VGND 0.02961f
C17587 VPWR.n572 VGND 0.09152f
C17588 VPWR.t1217 VGND 0.07849f
C17589 VPWR.t461 VGND 0.09218f
C17590 VPWR.t939 VGND 0.11957f
C17591 VPWR.t1701 VGND 0.03331f
C17592 VPWR.t1783 VGND 0.02961f
C17593 VPWR.n573 VGND 0.09152f
C17594 VPWR.n574 VGND 0.13913f
C17595 VPWR.n575 VGND 0.13913f
C17596 VPWR.t940 VGND 0.03331f
C17597 VPWR.t1805 VGND 0.02961f
C17598 VPWR.n576 VGND 0.09152f
C17599 VPWR.t1215 VGND 0.07849f
C17600 VPWR.t1804 VGND 0.09218f
C17601 VPWR.t757 VGND 0.03331f
C17602 VPWR.t216 VGND 0.02961f
C17603 VPWR.n577 VGND 0.09152f
C17604 VPWR.t629 VGND 0.03331f
C17605 VPWR.t324 VGND 0.02961f
C17606 VPWR.n578 VGND 0.09152f
C17607 VPWR.t1420 VGND 0.14512f
C17608 VPWR.t1446 VGND 0.07849f
C17609 VPWR.t1162 VGND 0.09218f
C17610 VPWR.t1421 VGND 0.03331f
C17611 VPWR.t1163 VGND 0.02961f
C17612 VPWR.n579 VGND 0.09152f
C17613 VPWR.n580 VGND 0.01797f
C17614 VPWR.n581 VGND 0.00728f
C17615 VPWR.n582 VGND 0.10822f
C17616 VPWR.t1152 VGND 0.11957f
C17617 VPWR.t1441 VGND 0.07849f
C17618 VPWR.t1910 VGND 0.09218f
C17619 VPWR.t1153 VGND 0.03331f
C17620 VPWR.t1911 VGND 0.02961f
C17621 VPWR.n583 VGND 0.09152f
C17622 VPWR.n584 VGND 0.01797f
C17623 VPWR.n585 VGND 0.00728f
C17624 VPWR.n586 VGND 0.10822f
C17625 VPWR.t1609 VGND 0.11957f
C17626 VPWR.t607 VGND 0.07849f
C17627 VPWR.t1350 VGND 0.09218f
C17628 VPWR.t1610 VGND 0.03331f
C17629 VPWR.t1351 VGND 0.02961f
C17630 VPWR.n587 VGND 0.09152f
C17631 VPWR.n588 VGND 0.01797f
C17632 VPWR.n589 VGND 0.00728f
C17633 VPWR.n590 VGND 0.10822f
C17634 VPWR.t1374 VGND 0.11957f
C17635 VPWR.t606 VGND 0.07849f
C17636 VPWR.t1634 VGND 0.09218f
C17637 VPWR.t1375 VGND 0.03331f
C17638 VPWR.t1635 VGND 0.02961f
C17639 VPWR.n591 VGND 0.09152f
C17640 VPWR.n592 VGND 0.01797f
C17641 VPWR.n593 VGND 0.00728f
C17642 VPWR.n594 VGND 0.10822f
C17643 VPWR.t1063 VGND 0.11957f
C17644 VPWR.t1445 VGND 0.07849f
C17645 VPWR.t1550 VGND 0.09218f
C17646 VPWR.t1064 VGND 0.03331f
C17647 VPWR.t1551 VGND 0.02961f
C17648 VPWR.n595 VGND 0.09152f
C17649 VPWR.n596 VGND 0.01797f
C17650 VPWR.n597 VGND 0.00728f
C17651 VPWR.n598 VGND 0.10822f
C17652 VPWR.t1544 VGND 0.11957f
C17653 VPWR.t1168 VGND 0.07849f
C17654 VPWR.t686 VGND 0.09218f
C17655 VPWR.t1545 VGND 0.03331f
C17656 VPWR.t687 VGND 0.02961f
C17657 VPWR.n599 VGND 0.09152f
C17658 VPWR.n600 VGND 0.01797f
C17659 VPWR.n601 VGND 0.00728f
C17660 VPWR.n602 VGND 0.10822f
C17661 VPWR.t543 VGND 0.11957f
C17662 VPWR.t1167 VGND 0.07849f
C17663 VPWR.t1790 VGND 0.09218f
C17664 VPWR.t544 VGND 0.03331f
C17665 VPWR.t1791 VGND 0.02961f
C17666 VPWR.n603 VGND 0.09152f
C17667 VPWR.n604 VGND 0.01797f
C17668 VPWR.n605 VGND 0.00728f
C17669 VPWR.n606 VGND 0.10822f
C17670 VPWR.t726 VGND 0.11957f
C17671 VPWR.t1444 VGND 0.07849f
C17672 VPWR.t911 VGND 0.09218f
C17673 VPWR.t727 VGND 0.03331f
C17674 VPWR.t912 VGND 0.02961f
C17675 VPWR.n607 VGND 0.09152f
C17676 VPWR.n608 VGND 0.01797f
C17677 VPWR.n609 VGND 0.00728f
C17678 VPWR.n610 VGND 0.10822f
C17679 VPWR.t1018 VGND 0.11957f
C17680 VPWR.t1443 VGND 0.07849f
C17681 VPWR.t1924 VGND 0.09218f
C17682 VPWR.t1019 VGND 0.03331f
C17683 VPWR.t1925 VGND 0.02961f
C17684 VPWR.n611 VGND 0.09152f
C17685 VPWR.n612 VGND 0.01797f
C17686 VPWR.n613 VGND 0.00728f
C17687 VPWR.n614 VGND 0.10822f
C17688 VPWR.t1918 VGND 0.11957f
C17689 VPWR.t1169 VGND 0.07849f
C17690 VPWR.t650 VGND 0.09218f
C17691 VPWR.t1919 VGND 0.03331f
C17692 VPWR.t651 VGND 0.02961f
C17693 VPWR.n615 VGND 0.09152f
C17694 VPWR.n616 VGND 0.01797f
C17695 VPWR.n617 VGND 0.00728f
C17696 VPWR.n618 VGND 0.10822f
C17697 VPWR.t640 VGND 0.11957f
C17698 VPWR.t1448 VGND 0.07849f
C17699 VPWR.t1102 VGND 0.09218f
C17700 VPWR.t641 VGND 0.03331f
C17701 VPWR.t1103 VGND 0.02961f
C17702 VPWR.n619 VGND 0.09152f
C17703 VPWR.n620 VGND 0.01797f
C17704 VPWR.n621 VGND 0.00728f
C17705 VPWR.n622 VGND 0.10822f
C17706 VPWR.t1055 VGND 0.11957f
C17707 VPWR.t1447 VGND 0.07849f
C17708 VPWR.t1459 VGND 0.09218f
C17709 VPWR.t1056 VGND 0.03331f
C17710 VPWR.t1460 VGND 0.02961f
C17711 VPWR.n623 VGND 0.09152f
C17712 VPWR.n624 VGND 0.01797f
C17713 VPWR.n625 VGND 0.00728f
C17714 VPWR.n626 VGND 0.10822f
C17715 VPWR.t1181 VGND 0.11957f
C17716 VPWR.t1166 VGND 0.07849f
C17717 VPWR.t1706 VGND 0.09218f
C17718 VPWR.t1182 VGND 0.03331f
C17719 VPWR.t1707 VGND 0.02961f
C17720 VPWR.n627 VGND 0.09152f
C17721 VPWR.n628 VGND 0.01797f
C17722 VPWR.n629 VGND 0.00728f
C17723 VPWR.n630 VGND 0.10822f
C17724 VPWR.t922 VGND 0.11957f
C17725 VPWR.t1165 VGND 0.07849f
C17726 VPWR.t488 VGND 0.09218f
C17727 VPWR.t923 VGND 0.03331f
C17728 VPWR.t489 VGND 0.02961f
C17729 VPWR.n631 VGND 0.09152f
C17730 VPWR.n632 VGND 0.01797f
C17731 VPWR.n633 VGND 0.00728f
C17732 VPWR.n634 VGND 0.10822f
C17733 VPWR.t680 VGND 0.11957f
C17734 VPWR.t1164 VGND 0.07849f
C17735 VPWR.t758 VGND 0.09218f
C17736 VPWR.t681 VGND 0.03331f
C17737 VPWR.t759 VGND 0.02961f
C17738 VPWR.n635 VGND 0.09152f
C17739 VPWR.n636 VGND 0.01797f
C17740 VPWR.n637 VGND 0.00728f
C17741 VPWR.n638 VGND 0.10822f
C17742 VPWR.t628 VGND 0.11957f
C17743 VPWR.t1442 VGND 0.07849f
C17744 VPWR.t323 VGND 0.13333f
C17745 VPWR.n639 VGND 0.07618f
C17746 VPWR.n640 VGND 0.01797f
C17747 VPWR.n641 VGND 0.13913f
C17748 VPWR.n642 VGND 1.01577f
C17749 VPWR.n643 VGND 0.13913f
C17750 VPWR.t1809 VGND 0.03331f
C17751 VPWR.t50 VGND 0.02961f
C17752 VPWR.n644 VGND 0.09152f
C17753 VPWR.t630 VGND 0.09218f
C17754 VPWR.t998 VGND 0.03331f
C17755 VPWR.t631 VGND 0.02961f
C17756 VPWR.n645 VGND 0.09152f
C17757 VPWR.n646 VGND 0.13913f
C17758 VPWR.n647 VGND 0.13913f
C17759 VPWR.t806 VGND 0.03331f
C17760 VPWR.t510 VGND 0.02961f
C17761 VPWR.n648 VGND 0.09152f
C17762 VPWR.t926 VGND 0.09218f
C17763 VPWR.t1206 VGND 0.03331f
C17764 VPWR.t927 VGND 0.02961f
C17765 VPWR.n649 VGND 0.09152f
C17766 VPWR.n650 VGND 0.13913f
C17767 VPWR.n651 VGND 0.13913f
C17768 VPWR.t554 VGND 0.03331f
C17769 VPWR.t1242 VGND 0.02961f
C17770 VPWR.n652 VGND 0.09152f
C17771 VPWR.t1475 VGND 0.09218f
C17772 VPWR.t1821 VGND 0.03331f
C17773 VPWR.t1476 VGND 0.02961f
C17774 VPWR.n653 VGND 0.09152f
C17775 VPWR.n654 VGND 0.13913f
C17776 VPWR.n655 VGND 0.13913f
C17777 VPWR.t1600 VGND 0.03331f
C17778 VPWR.t1827 VGND 0.02961f
C17779 VPWR.n656 VGND 0.09152f
C17780 VPWR.t1605 VGND 0.09218f
C17781 VPWR.t578 VGND 0.03331f
C17782 VPWR.t1606 VGND 0.02961f
C17783 VPWR.n657 VGND 0.09152f
C17784 VPWR.n658 VGND 0.13913f
C17785 VPWR.n659 VGND 0.13913f
C17786 VPWR.t1899 VGND 0.03331f
C17787 VPWR.t1023 VGND 0.02961f
C17788 VPWR.n660 VGND 0.09152f
C17789 VPWR.t1904 VGND 0.09218f
C17790 VPWR.t592 VGND 0.03331f
C17791 VPWR.t1905 VGND 0.02961f
C17792 VPWR.n661 VGND 0.09152f
C17793 VPWR.n662 VGND 0.13913f
C17794 VPWR.n663 VGND 0.13913f
C17795 VPWR.t1667 VGND 0.03331f
C17796 VPWR.t703 VGND 0.02961f
C17797 VPWR.n664 VGND 0.09152f
C17798 VPWR.t1559 VGND 0.09218f
C17799 VPWR.t803 VGND 0.03331f
C17800 VPWR.t1560 VGND 0.02961f
C17801 VPWR.n665 VGND 0.09152f
C17802 VPWR.n666 VGND 0.13913f
C17803 VPWR.n667 VGND 0.13913f
C17804 VPWR.t1395 VGND 0.03331f
C17805 VPWR.t1066 VGND 0.02961f
C17806 VPWR.n668 VGND 0.09152f
C17807 VPWR.t1370 VGND 0.09218f
C17808 VPWR.t1584 VGND 0.03331f
C17809 VPWR.t1371 VGND 0.02961f
C17810 VPWR.n669 VGND 0.09152f
C17811 VPWR.n670 VGND 0.13913f
C17812 VPWR.n671 VGND 0.13913f
C17813 VPWR.t1725 VGND 0.03331f
C17814 VPWR.t1590 VGND 0.02961f
C17815 VPWR.n672 VGND 0.09152f
C17816 VPWR.t1433 VGND 0.14512f
C17817 VPWR.t1506 VGND 0.07849f
C17818 VPWR.t979 VGND 0.09218f
C17819 VPWR.t1434 VGND 0.03331f
C17820 VPWR.t980 VGND 0.02961f
C17821 VPWR.n673 VGND 0.09152f
C17822 VPWR.t1440 VGND 0.03331f
C17823 VPWR.t715 VGND 0.02961f
C17824 VPWR.n674 VGND 0.09152f
C17825 VPWR.t1439 VGND 0.14512f
C17826 VPWR.t600 VGND 0.07849f
C17827 VPWR.t714 VGND 0.09218f
C17828 VPWR.t693 VGND 0.03331f
C17829 VPWR.t157 VGND 0.02961f
C17830 VPWR.n675 VGND 0.09152f
C17831 VPWR.n676 VGND 0.01797f
C17832 VPWR.n677 VGND 0.07618f
C17833 VPWR.t156 VGND 0.13333f
C17834 VPWR.t733 VGND 0.07849f
C17835 VPWR.t692 VGND 0.11957f
C17836 VPWR.t1785 VGND 0.03331f
C17837 VPWR.t1813 VGND 0.02961f
C17838 VPWR.n678 VGND 0.09152f
C17839 VPWR.n679 VGND 0.01797f
C17840 VPWR.n680 VGND 0.00728f
C17841 VPWR.n681 VGND 0.10822f
C17842 VPWR.t1812 VGND 0.09218f
C17843 VPWR.t1039 VGND 0.07849f
C17844 VPWR.t1784 VGND 0.11957f
C17845 VPWR.t452 VGND 0.03331f
C17846 VPWR.t1496 VGND 0.02961f
C17847 VPWR.n682 VGND 0.09152f
C17848 VPWR.n683 VGND 0.01797f
C17849 VPWR.n684 VGND 0.00728f
C17850 VPWR.n685 VGND 0.10822f
C17851 VPWR.t1495 VGND 0.09218f
C17852 VPWR.t1040 VGND 0.07849f
C17853 VPWR.t451 VGND 0.11957f
C17854 VPWR.t470 VGND 0.03331f
C17855 VPWR.t812 VGND 0.02961f
C17856 VPWR.n686 VGND 0.09152f
C17857 VPWR.n687 VGND 0.01797f
C17858 VPWR.n688 VGND 0.00728f
C17859 VPWR.n689 VGND 0.10822f
C17860 VPWR.t811 VGND 0.09218f
C17861 VPWR.t1041 VGND 0.07849f
C17862 VPWR.t469 VGND 0.11957f
C17863 VPWR.t1576 VGND 0.03331f
C17864 VPWR.t1755 VGND 0.02961f
C17865 VPWR.n690 VGND 0.09152f
C17866 VPWR.n691 VGND 0.01797f
C17867 VPWR.n692 VGND 0.00728f
C17868 VPWR.n693 VGND 0.10822f
C17869 VPWR.t1754 VGND 0.09218f
C17870 VPWR.t602 VGND 0.07849f
C17871 VPWR.t1575 VGND 0.11957f
C17872 VPWR.t663 VGND 0.03331f
C17873 VPWR.t1580 VGND 0.02961f
C17874 VPWR.n694 VGND 0.09152f
C17875 VPWR.n695 VGND 0.01797f
C17876 VPWR.n696 VGND 0.00728f
C17877 VPWR.n697 VGND 0.10822f
C17878 VPWR.t1579 VGND 0.09218f
C17879 VPWR.t603 VGND 0.07849f
C17880 VPWR.t662 VGND 0.11957f
C17881 VPWR.t478 VGND 0.03331f
C17882 VPWR.t669 VGND 0.02961f
C17883 VPWR.n698 VGND 0.09152f
C17884 VPWR.n699 VGND 0.01797f
C17885 VPWR.n700 VGND 0.00728f
C17886 VPWR.n701 VGND 0.10822f
C17887 VPWR.t668 VGND 0.09218f
C17888 VPWR.t1044 VGND 0.07849f
C17889 VPWR.t477 VGND 0.11957f
C17890 VPWR.t857 VGND 0.03331f
C17891 VPWR.t1115 VGND 0.02961f
C17892 VPWR.n702 VGND 0.09152f
C17893 VPWR.n703 VGND 0.01797f
C17894 VPWR.n704 VGND 0.00728f
C17895 VPWR.n705 VGND 0.10822f
C17896 VPWR.t1114 VGND 0.09218f
C17897 VPWR.t1712 VGND 0.07849f
C17898 VPWR.t856 VGND 0.11957f
C17899 VPWR.t735 VGND 0.03331f
C17900 VPWR.t869 VGND 0.02961f
C17901 VPWR.n706 VGND 0.09152f
C17902 VPWR.n707 VGND 0.01797f
C17903 VPWR.n708 VGND 0.00728f
C17904 VPWR.n709 VGND 0.10822f
C17905 VPWR.t868 VGND 0.09218f
C17906 VPWR.t598 VGND 0.07849f
C17907 VPWR.t734 VGND 0.11957f
C17908 VPWR.t962 VGND 0.03331f
C17909 VPWR.t1891 VGND 0.02961f
C17910 VPWR.n710 VGND 0.09152f
C17911 VPWR.n711 VGND 0.01797f
C17912 VPWR.n712 VGND 0.00728f
C17913 VPWR.n713 VGND 0.10822f
C17914 VPWR.t1890 VGND 0.09218f
C17915 VPWR.t1042 VGND 0.07849f
C17916 VPWR.t961 VGND 0.11957f
C17917 VPWR.t522 VGND 0.03331f
C17918 VPWR.t966 VGND 0.02961f
C17919 VPWR.n714 VGND 0.09152f
C17920 VPWR.n715 VGND 0.01797f
C17921 VPWR.n716 VGND 0.00728f
C17922 VPWR.n717 VGND 0.10822f
C17923 VPWR.t965 VGND 0.09218f
C17924 VPWR.t1043 VGND 0.07849f
C17925 VPWR.t521 VGND 0.11957f
C17926 VPWR.t1026 VGND 0.03331f
C17927 VPWR.t1570 VGND 0.02961f
C17928 VPWR.n718 VGND 0.09152f
C17929 VPWR.n719 VGND 0.01797f
C17930 VPWR.n720 VGND 0.00728f
C17931 VPWR.n721 VGND 0.10822f
C17932 VPWR.t1569 VGND 0.09218f
C17933 VPWR.t599 VGND 0.07849f
C17934 VPWR.t1025 VGND 0.11957f
C17935 VPWR.t1409 VGND 0.03331f
C17936 VPWR.t1854 VGND 0.02961f
C17937 VPWR.n722 VGND 0.09152f
C17938 VPWR.n723 VGND 0.01797f
C17939 VPWR.n724 VGND 0.00728f
C17940 VPWR.n725 VGND 0.10822f
C17941 VPWR.t1853 VGND 0.09218f
C17942 VPWR.t604 VGND 0.07849f
C17943 VPWR.t1408 VGND 0.11957f
C17944 VPWR.t840 VGND 0.03331f
C17945 VPWR.t1387 VGND 0.02961f
C17946 VPWR.n726 VGND 0.09152f
C17947 VPWR.n727 VGND 0.01797f
C17948 VPWR.n728 VGND 0.00728f
C17949 VPWR.n729 VGND 0.10822f
C17950 VPWR.t1386 VGND 0.09218f
C17951 VPWR.t605 VGND 0.07849f
C17952 VPWR.t839 VGND 0.11957f
C17953 VPWR.t902 VGND 0.03331f
C17954 VPWR.t844 VGND 0.02961f
C17955 VPWR.n730 VGND 0.09152f
C17956 VPWR.n731 VGND 0.01797f
C17957 VPWR.n732 VGND 0.00728f
C17958 VPWR.n733 VGND 0.10822f
C17959 VPWR.t843 VGND 0.09218f
C17960 VPWR.t732 VGND 0.07849f
C17961 VPWR.t901 VGND 0.11957f
C17962 VPWR.n734 VGND 0.10822f
C17963 VPWR.n735 VGND 0.00728f
C17964 VPWR.n736 VGND 0.01797f
C17965 VPWR.n737 VGND 0.13913f
C17966 VPWR.n738 VGND 1.0094f
C17967 VPWR.n739 VGND 0.13913f
C17968 VPWR.t1436 VGND 0.03331f
C17969 VPWR.t834 VGND 0.02961f
C17970 VPWR.n740 VGND 0.09152f
C17971 VPWR.t1435 VGND 0.14512f
C17972 VPWR.t789 VGND 0.07849f
C17973 VPWR.t833 VGND 0.09218f
C17974 VPWR.t1521 VGND 0.11957f
C17975 VPWR.t830 VGND 0.03331f
C17976 VPWR.t1524 VGND 0.02961f
C17977 VPWR.n741 VGND 0.09152f
C17978 VPWR.n742 VGND 0.13913f
C17979 VPWR.n743 VGND 0.13913f
C17980 VPWR.t1522 VGND 0.03331f
C17981 VPWR.t1379 VGND 0.02961f
C17982 VPWR.n744 VGND 0.09152f
C17983 VPWR.t793 VGND 0.07849f
C17984 VPWR.t1378 VGND 0.09218f
C17985 VPWR.t1029 VGND 0.11957f
C17986 VPWR.t1403 VGND 0.03331f
C17987 VPWR.t1860 VGND 0.02961f
C17988 VPWR.n745 VGND 0.09152f
C17989 VPWR.n746 VGND 0.13913f
C17990 VPWR.n747 VGND 0.13913f
C17991 VPWR.t1030 VGND 0.03331f
C17992 VPWR.t1665 VGND 0.02961f
C17993 VPWR.n748 VGND 0.09152f
C17994 VPWR.t788 VGND 0.07849f
C17995 VPWR.t1664 VGND 0.09218f
C17996 VPWR.t969 VGND 0.11957f
C17997 VPWR.t1574 VGND 0.03331f
C17998 VPWR.t590 VGND 0.02961f
C17999 VPWR.n749 VGND 0.09152f
C18000 VPWR.n750 VGND 0.13913f
C18001 VPWR.n751 VGND 0.13913f
C18002 VPWR.t970 VGND 0.03331f
C18003 VPWR.t1897 VGND 0.02961f
C18004 VPWR.n752 VGND 0.09152f
C18005 VPWR.t1075 VGND 0.07849f
C18006 VPWR.t1896 VGND 0.09218f
C18007 VPWR.t981 VGND 0.11957f
C18008 VPWR.t1895 VGND 0.03331f
C18009 VPWR.t1111 VGND 0.02961f
C18010 VPWR.n753 VGND 0.09152f
C18011 VPWR.n754 VGND 0.13913f
C18012 VPWR.n755 VGND 0.13913f
C18013 VPWR.t982 VGND 0.03331f
C18014 VPWR.t1121 VGND 0.02961f
C18015 VPWR.n756 VGND 0.09152f
C18016 VPWR.t786 VGND 0.07849f
C18017 VPWR.t1120 VGND 0.09218f
C18018 VPWR.t670 VGND 0.11957f
C18019 VPWR.t1119 VGND 0.03331f
C18020 VPWR.t675 VGND 0.02961f
C18021 VPWR.n757 VGND 0.09152f
C18022 VPWR.n758 VGND 0.13913f
C18023 VPWR.n759 VGND 0.13913f
C18024 VPWR.t671 VGND 0.03331f
C18025 VPWR.t552 VGND 0.02961f
C18026 VPWR.n760 VGND 0.09152f
C18027 VPWR.t791 VGND 0.07849f
C18028 VPWR.t551 VGND 0.09218f
C18029 VPWR.t1756 VGND 0.11957f
C18030 VPWR.t550 VGND 0.03331f
C18031 VPWR.t1204 VGND 0.02961f
C18032 VPWR.n761 VGND 0.09152f
C18033 VPWR.n762 VGND 0.13913f
C18034 VPWR.n763 VGND 0.13913f
C18035 VPWR.t1757 VGND 0.03331f
C18036 VPWR.t818 VGND 0.02961f
C18037 VPWR.n764 VGND 0.09152f
C18038 VPWR.t1074 VGND 0.07849f
C18039 VPWR.t817 VGND 0.09218f
C18040 VPWR.t1615 VGND 0.11957f
C18041 VPWR.t456 VGND 0.03331f
C18042 VPWR.t1620 VGND 0.02961f
C18043 VPWR.n765 VGND 0.09152f
C18044 VPWR.n766 VGND 0.13913f
C18045 VPWR.n767 VGND 0.13913f
C18046 VPWR.t1616 VGND 0.03331f
C18047 VPWR.t1819 VGND 0.02961f
C18048 VPWR.n768 VGND 0.09152f
C18049 VPWR.t794 VGND 0.07849f
C18050 VPWR.t1818 VGND 0.09218f
C18051 VPWR.t697 VGND 0.03331f
C18052 VPWR.t117 VGND 0.02961f
C18053 VPWR.n769 VGND 0.09152f
C18054 VPWR.t753 VGND 0.03331f
C18055 VPWR.t222 VGND 0.02961f
C18056 VPWR.n770 VGND 0.09152f
C18057 VPWR.t1414 VGND 0.14512f
C18058 VPWR.t1753 VGND 0.07849f
C18059 VPWR.t897 VGND 0.09218f
C18060 VPWR.t1415 VGND 0.03331f
C18061 VPWR.t898 VGND 0.02961f
C18062 VPWR.n771 VGND 0.09152f
C18063 VPWR.n772 VGND 0.01797f
C18064 VPWR.n773 VGND 0.00728f
C18065 VPWR.n774 VGND 0.10822f
C18066 VPWR.t531 VGND 0.11957f
C18067 VPWR.t1748 VGND 0.07849f
C18068 VPWR.t1082 VGND 0.09218f
C18069 VPWR.t532 VGND 0.03331f
C18070 VPWR.t1083 VGND 0.02961f
C18071 VPWR.n775 VGND 0.09152f
C18072 VPWR.n776 VGND 0.01797f
C18073 VPWR.n777 VGND 0.00728f
C18074 VPWR.n778 VGND 0.10822f
C18075 VPWR.t1595 VGND 0.11957f
C18076 VPWR.t1771 VGND 0.07849f
C18077 VPWR.t1398 VGND 0.09218f
C18078 VPWR.t1596 VGND 0.03331f
C18079 VPWR.t1399 VGND 0.02961f
C18080 VPWR.n779 VGND 0.09152f
C18081 VPWR.n780 VGND 0.01797f
C18082 VPWR.n781 VGND 0.00728f
C18083 VPWR.n782 VGND 0.10822f
C18084 VPWR.t1362 VGND 0.11957f
C18085 VPWR.t1770 VGND 0.07849f
C18086 VPWR.t1033 VGND 0.09218f
C18087 VPWR.t1363 VGND 0.03331f
C18088 VPWR.t1034 VGND 0.02961f
C18089 VPWR.n783 VGND 0.09152f
C18090 VPWR.n784 VGND 0.01797f
C18091 VPWR.n785 VGND 0.00728f
C18092 VPWR.n786 VGND 0.10822f
C18093 VPWR.t1628 VGND 0.11957f
C18094 VPWR.t1752 VGND 0.07849f
C18095 VPWR.t1517 VGND 0.09218f
C18096 VPWR.t1629 VGND 0.03331f
C18097 VPWR.t1518 VGND 0.02961f
C18098 VPWR.n787 VGND 0.09152f
C18099 VPWR.n788 VGND 0.01797f
C18100 VPWR.n789 VGND 0.00728f
C18101 VPWR.n790 VGND 0.10822f
C18102 VPWR.t1511 VGND 0.11957f
C18103 VPWR.t1776 VGND 0.07849f
C18104 VPWR.t563 VGND 0.09218f
C18105 VPWR.t1512 VGND 0.03331f
C18106 VPWR.t564 VGND 0.02961f
C18107 VPWR.n791 VGND 0.09152f
C18108 VPWR.n792 VGND 0.01797f
C18109 VPWR.n793 VGND 0.00728f
C18110 VPWR.n794 VGND 0.10822f
C18111 VPWR.t557 VGND 0.11957f
C18112 VPWR.t1775 VGND 0.07849f
C18113 VPWR.t738 VGND 0.09218f
C18114 VPWR.t558 VGND 0.03331f
C18115 VPWR.t739 VGND 0.02961f
C18116 VPWR.n795 VGND 0.09152f
C18117 VPWR.n796 VGND 0.01797f
C18118 VPWR.n797 VGND 0.00728f
C18119 VPWR.n798 VGND 0.10822f
C18120 VPWR.t1798 VGND 0.11957f
C18121 VPWR.t1751 VGND 0.07849f
C18122 VPWR.t571 VGND 0.09218f
C18123 VPWR.t1799 VGND 0.03331f
C18124 VPWR.t572 VGND 0.02961f
C18125 VPWR.n799 VGND 0.09152f
C18126 VPWR.n800 VGND 0.01797f
C18127 VPWR.n801 VGND 0.00728f
C18128 VPWR.n802 VGND 0.10822f
C18129 VPWR.t919 VGND 0.11957f
C18130 VPWR.t1750 VGND 0.07849f
C18131 VPWR.t955 VGND 0.09218f
C18132 VPWR.t920 VGND 0.03331f
C18133 VPWR.t956 VGND 0.02961f
C18134 VPWR.n803 VGND 0.09152f
C18135 VPWR.n804 VGND 0.01797f
C18136 VPWR.n805 VGND 0.00728f
C18137 VPWR.n806 VGND 0.10822f
C18138 VPWR.t847 VGND 0.11957f
C18139 VPWR.t1777 VGND 0.07849f
C18140 VPWR.t618 VGND 0.09218f
C18141 VPWR.t848 VGND 0.03331f
C18142 VPWR.t619 VGND 0.02961f
C18143 VPWR.n807 VGND 0.09152f
C18144 VPWR.n808 VGND 0.01797f
C18145 VPWR.n809 VGND 0.00728f
C18146 VPWR.n810 VGND 0.10822f
C18147 VPWR.t610 VGND 0.11957f
C18148 VPWR.t1769 VGND 0.07849f
C18149 VPWR.t1684 VGND 0.09218f
C18150 VPWR.t611 VGND 0.03331f
C18151 VPWR.t1685 VGND 0.02961f
C18152 VPWR.n811 VGND 0.09152f
C18153 VPWR.n812 VGND 0.01797f
C18154 VPWR.n813 VGND 0.00728f
C18155 VPWR.n814 VGND 0.10822f
C18156 VPWR.t1213 VGND 0.11957f
C18157 VPWR.t1768 VGND 0.07849f
C18158 VPWR.t465 VGND 0.09218f
C18159 VPWR.t1214 VGND 0.03331f
C18160 VPWR.t466 VGND 0.02961f
C18161 VPWR.n815 VGND 0.09152f
C18162 VPWR.n816 VGND 0.01797f
C18163 VPWR.n817 VGND 0.00728f
C18164 VPWR.n818 VGND 0.10822f
C18165 VPWR.t1760 VGND 0.11957f
C18166 VPWR.t1774 VGND 0.07849f
C18167 VPWR.t459 VGND 0.09218f
C18168 VPWR.t1761 VGND 0.03331f
C18169 VPWR.t460 VGND 0.02961f
C18170 VPWR.n819 VGND 0.09152f
C18171 VPWR.n820 VGND 0.01797f
C18172 VPWR.n821 VGND 0.00728f
C18173 VPWR.n822 VGND 0.10822f
C18174 VPWR.t1696 VGND 0.11957f
C18175 VPWR.t1773 VGND 0.07849f
C18176 VPWR.t1780 VGND 0.09218f
C18177 VPWR.t1697 VGND 0.03331f
C18178 VPWR.t1781 VGND 0.02961f
C18179 VPWR.n823 VGND 0.09152f
C18180 VPWR.n824 VGND 0.01797f
C18181 VPWR.n825 VGND 0.00728f
C18182 VPWR.n826 VGND 0.10822f
C18183 VPWR.t937 VGND 0.11957f
C18184 VPWR.t1772 VGND 0.07849f
C18185 VPWR.t700 VGND 0.09218f
C18186 VPWR.t938 VGND 0.03331f
C18187 VPWR.t701 VGND 0.02961f
C18188 VPWR.n827 VGND 0.09152f
C18189 VPWR.n828 VGND 0.01797f
C18190 VPWR.n829 VGND 0.00728f
C18191 VPWR.n830 VGND 0.10822f
C18192 VPWR.t752 VGND 0.11957f
C18193 VPWR.t1749 VGND 0.07849f
C18194 VPWR.t221 VGND 0.13333f
C18195 VPWR.n831 VGND 0.07618f
C18196 VPWR.n832 VGND 0.01797f
C18197 VPWR.n833 VGND 0.13913f
C18198 VPWR.n834 VGND 1.01577f
C18199 VPWR.n835 VGND 0.13913f
C18200 VPWR.t1811 VGND 0.03331f
C18201 VPWR.t42 VGND 0.02961f
C18202 VPWR.n836 VGND 0.09152f
C18203 VPWR.t634 VGND 0.09218f
C18204 VPWR.t1000 VGND 0.03331f
C18205 VPWR.t635 VGND 0.02961f
C18206 VPWR.n837 VGND 0.09152f
C18207 VPWR.n838 VGND 0.13913f
C18208 VPWR.n839 VGND 0.13913f
C18209 VPWR.t808 VGND 0.03331f
C18210 VPWR.t512 VGND 0.02961f
C18211 VPWR.n840 VGND 0.09152f
C18212 VPWR.t928 VGND 0.09218f
C18213 VPWR.t1208 VGND 0.03331f
C18214 VPWR.t929 VGND 0.02961f
C18215 VPWR.n841 VGND 0.09152f
C18216 VPWR.n842 VGND 0.13913f
C18217 VPWR.n843 VGND 0.13913f
C18218 VPWR.t1472 VGND 0.03331f
C18219 VPWR.t1244 VGND 0.02961f
C18220 VPWR.n844 VGND 0.09152f
C18221 VPWR.t1477 VGND 0.09218f
C18222 VPWR.t1823 VGND 0.03331f
C18223 VPWR.t1478 VGND 0.02961f
C18224 VPWR.n845 VGND 0.09152f
C18225 VPWR.n846 VGND 0.13913f
C18226 VPWR.n847 VGND 0.13913f
C18227 VPWR.t1602 VGND 0.03331f
C18228 VPWR.t1829 VGND 0.02961f
C18229 VPWR.n848 VGND 0.09152f
C18230 VPWR.t1008 VGND 0.09218f
C18231 VPWR.t865 VGND 0.03331f
C18232 VPWR.t1009 VGND 0.02961f
C18233 VPWR.n849 VGND 0.09152f
C18234 VPWR.n850 VGND 0.13913f
C18235 VPWR.n851 VGND 0.13913f
C18236 VPWR.t1901 VGND 0.03331f
C18237 VPWR.t385 VGND 0.02961f
C18238 VPWR.n852 VGND 0.09152f
C18239 VPWR.t1906 VGND 0.09218f
C18240 VPWR.t594 VGND 0.03331f
C18241 VPWR.t1907 VGND 0.02961f
C18242 VPWR.n853 VGND 0.09152f
C18243 VPWR.n854 VGND 0.13913f
C18244 VPWR.n855 VGND 0.13913f
C18245 VPWR.t1535 VGND 0.03331f
C18246 VPWR.t705 VGND 0.02961f
C18247 VPWR.n856 VGND 0.09152f
C18248 VPWR.t1561 VGND 0.09218f
C18249 VPWR.t1852 VGND 0.03331f
C18250 VPWR.t1562 VGND 0.02961f
C18251 VPWR.n857 VGND 0.09152f
C18252 VPWR.n858 VGND 0.13913f
C18253 VPWR.n859 VGND 0.13913f
C18254 VPWR.t1393 VGND 0.03331f
C18255 VPWR.t1070 VGND 0.02961f
C18256 VPWR.n860 VGND 0.09152f
C18257 VPWR.t1368 VGND 0.09218f
C18258 VPWR.t1586 VGND 0.03331f
C18259 VPWR.t1369 VGND 0.02961f
C18260 VPWR.n861 VGND 0.09152f
C18261 VPWR.n862 VGND 0.13913f
C18262 VPWR.n863 VGND 0.13913f
C18263 VPWR.t1727 VGND 0.03331f
C18264 VPWR.t1592 VGND 0.02961f
C18265 VPWR.n864 VGND 0.09152f
C18266 VPWR.t1431 VGND 0.14512f
C18267 VPWR.t1846 VGND 0.07849f
C18268 VPWR.t1122 VGND 0.09218f
C18269 VPWR.t1432 VGND 0.03331f
C18270 VPWR.t1123 VGND 0.02961f
C18271 VPWR.n865 VGND 0.09152f
C18272 VPWR.t1417 VGND 0.03331f
C18273 VPWR.t896 VGND 0.02961f
C18274 VPWR.n866 VGND 0.09152f
C18275 VPWR.t1416 VGND 0.14512f
C18276 VPWR.t1652 VGND 0.07849f
C18277 VPWR.t895 VGND 0.09218f
C18278 VPWR.t751 VGND 0.03331f
C18279 VPWR.t229 VGND 0.02961f
C18280 VPWR.n867 VGND 0.09152f
C18281 VPWR.n868 VGND 0.01797f
C18282 VPWR.n869 VGND 0.07618f
C18283 VPWR.t228 VGND 0.13333f
C18284 VPWR.t1648 VGND 0.07849f
C18285 VPWR.t750 VGND 0.11957f
C18286 VPWR.t936 VGND 0.03331f
C18287 VPWR.t699 VGND 0.02961f
C18288 VPWR.n870 VGND 0.09152f
C18289 VPWR.n871 VGND 0.01797f
C18290 VPWR.n872 VGND 0.00728f
C18291 VPWR.n873 VGND 0.10822f
C18292 VPWR.t698 VGND 0.09218f
C18293 VPWR.t1525 VGND 0.07849f
C18294 VPWR.t935 VGND 0.11957f
C18295 VPWR.t1693 VGND 0.03331f
C18296 VPWR.t1779 VGND 0.02961f
C18297 VPWR.n874 VGND 0.09152f
C18298 VPWR.n875 VGND 0.01797f
C18299 VPWR.n876 VGND 0.00728f
C18300 VPWR.n877 VGND 0.10822f
C18301 VPWR.t1778 VGND 0.09218f
C18302 VPWR.t1526 VGND 0.07849f
C18303 VPWR.t1692 VGND 0.11957f
C18304 VPWR.t1173 VGND 0.03331f
C18305 VPWR.t458 VGND 0.02961f
C18306 VPWR.n878 VGND 0.09152f
C18307 VPWR.n879 VGND 0.01797f
C18308 VPWR.n880 VGND 0.00728f
C18309 VPWR.n881 VGND 0.10822f
C18310 VPWR.t457 VGND 0.09218f
C18311 VPWR.t1527 VGND 0.07849f
C18312 VPWR.t1172 VGND 0.11957f
C18313 VPWR.t1212 VGND 0.03331f
C18314 VPWR.t1767 VGND 0.02961f
C18315 VPWR.n882 VGND 0.09152f
C18316 VPWR.n883 VGND 0.01797f
C18317 VPWR.n884 VGND 0.00728f
C18318 VPWR.n885 VGND 0.10822f
C18319 VPWR.t1766 VGND 0.09218f
C18320 VPWR.t388 VGND 0.07849f
C18321 VPWR.t1211 VGND 0.11957f
C18322 VPWR.t609 VGND 0.03331f
C18323 VPWR.t1683 VGND 0.02961f
C18324 VPWR.n886 VGND 0.09152f
C18325 VPWR.n887 VGND 0.01797f
C18326 VPWR.n888 VGND 0.00728f
C18327 VPWR.n889 VGND 0.10822f
C18328 VPWR.t1682 VGND 0.09218f
C18329 VPWR.t389 VGND 0.07849f
C18330 VPWR.t608 VGND 0.11957f
C18331 VPWR.t846 VGND 0.03331f
C18332 VPWR.t617 VGND 0.02961f
C18333 VPWR.n890 VGND 0.09152f
C18334 VPWR.n891 VGND 0.01797f
C18335 VPWR.n892 VGND 0.00728f
C18336 VPWR.n893 VGND 0.10822f
C18337 VPWR.t616 VGND 0.09218f
C18338 VPWR.t1530 VGND 0.07849f
C18339 VPWR.t845 VGND 0.11957f
C18340 VPWR.t916 VGND 0.03331f
C18341 VPWR.t954 VGND 0.02961f
C18342 VPWR.n894 VGND 0.09152f
C18343 VPWR.n895 VGND 0.01797f
C18344 VPWR.n896 VGND 0.00728f
C18345 VPWR.n897 VGND 0.10822f
C18346 VPWR.t953 VGND 0.09218f
C18347 VPWR.t1649 VGND 0.07849f
C18348 VPWR.t915 VGND 0.11957f
C18349 VPWR.t1797 VGND 0.03331f
C18350 VPWR.t984 VGND 0.02961f
C18351 VPWR.n898 VGND 0.09152f
C18352 VPWR.n899 VGND 0.01797f
C18353 VPWR.n900 VGND 0.00728f
C18354 VPWR.n901 VGND 0.10822f
C18355 VPWR.t983 VGND 0.09218f
C18356 VPWR.t1650 VGND 0.07849f
C18357 VPWR.t1796 VGND 0.11957f
C18358 VPWR.t556 VGND 0.03331f
C18359 VPWR.t1803 VGND 0.02961f
C18360 VPWR.n902 VGND 0.09152f
C18361 VPWR.n903 VGND 0.01797f
C18362 VPWR.n904 VGND 0.00728f
C18363 VPWR.n905 VGND 0.10822f
C18364 VPWR.t1802 VGND 0.09218f
C18365 VPWR.t1528 VGND 0.07849f
C18366 VPWR.t555 VGND 0.11957f
C18367 VPWR.t1510 VGND 0.03331f
C18368 VPWR.t562 VGND 0.02961f
C18369 VPWR.n906 VGND 0.09152f
C18370 VPWR.n907 VGND 0.01797f
C18371 VPWR.n908 VGND 0.00728f
C18372 VPWR.n909 VGND 0.10822f
C18373 VPWR.t561 VGND 0.09218f
C18374 VPWR.t1529 VGND 0.07849f
C18375 VPWR.t1509 VGND 0.11957f
C18376 VPWR.t1627 VGND 0.03331f
C18377 VPWR.t1516 VGND 0.02961f
C18378 VPWR.n910 VGND 0.09152f
C18379 VPWR.n911 VGND 0.01797f
C18380 VPWR.n912 VGND 0.00728f
C18381 VPWR.n913 VGND 0.10822f
C18382 VPWR.t1515 VGND 0.09218f
C18383 VPWR.t1651 VGND 0.07849f
C18384 VPWR.t1626 VGND 0.11957f
C18385 VPWR.t1365 VGND 0.03331f
C18386 VPWR.t1032 VGND 0.02961f
C18387 VPWR.n914 VGND 0.09152f
C18388 VPWR.n915 VGND 0.01797f
C18389 VPWR.n916 VGND 0.00728f
C18390 VPWR.n917 VGND 0.10822f
C18391 VPWR.t1031 VGND 0.09218f
C18392 VPWR.t390 VGND 0.07849f
C18393 VPWR.t1364 VGND 0.11957f
C18394 VPWR.t1594 VGND 0.03331f
C18395 VPWR.t1401 VGND 0.02961f
C18396 VPWR.n918 VGND 0.09152f
C18397 VPWR.n919 VGND 0.01797f
C18398 VPWR.n920 VGND 0.00728f
C18399 VPWR.n921 VGND 0.10822f
C18400 VPWR.t1400 VGND 0.09218f
C18401 VPWR.t391 VGND 0.07849f
C18402 VPWR.t1593 VGND 0.11957f
C18403 VPWR.t530 VGND 0.03331f
C18404 VPWR.t1081 VGND 0.02961f
C18405 VPWR.n922 VGND 0.09152f
C18406 VPWR.n923 VGND 0.01797f
C18407 VPWR.n924 VGND 0.00728f
C18408 VPWR.n925 VGND 0.10822f
C18409 VPWR.t1080 VGND 0.09218f
C18410 VPWR.t1647 VGND 0.07849f
C18411 VPWR.t529 VGND 0.11957f
C18412 VPWR.n926 VGND 0.10822f
C18413 VPWR.n927 VGND 0.00728f
C18414 VPWR.n928 VGND 0.01797f
C18415 VPWR.n929 VGND 0.13913f
C18416 VPWR.n930 VGND 1.0094f
C18417 VPWR.n931 VGND 0.13913f
C18418 VPWR.t1423 VGND 0.03331f
C18419 VPWR.t1161 VGND 0.02961f
C18420 VPWR.n932 VGND 0.09152f
C18421 VPWR.t1422 VGND 0.14512f
C18422 VPWR.t1487 VGND 0.07849f
C18423 VPWR.t1160 VGND 0.09218f
C18424 VPWR.t425 VGND 0.11957f
C18425 VPWR.t1740 VGND 0.03331f
C18426 VPWR.t1614 VGND 0.02961f
C18427 VPWR.n933 VGND 0.09152f
C18428 VPWR.n934 VGND 0.13913f
C18429 VPWR.n935 VGND 0.13913f
C18430 VPWR.t426 VGND 0.03331f
C18431 VPWR.t1353 VGND 0.02961f
C18432 VPWR.n936 VGND 0.09152f
C18433 VPWR.t1202 VGND 0.07849f
C18434 VPWR.t1352 VGND 0.09218f
C18435 VPWR.t1061 VGND 0.11957f
C18436 VPWR.t1377 VGND 0.03331f
C18437 VPWR.t1631 VGND 0.02961f
C18438 VPWR.n937 VGND 0.09152f
C18439 VPWR.n938 VGND 0.13913f
C18440 VPWR.n939 VGND 0.13913f
C18441 VPWR.t1062 VGND 0.03331f
C18442 VPWR.t1549 VGND 0.02961f
C18443 VPWR.n940 VGND 0.09152f
C18444 VPWR.t1486 VGND 0.07849f
C18445 VPWR.t1548 VGND 0.09218f
C18446 VPWR.t539 VGND 0.11957f
C18447 VPWR.t1718 VGND 0.03331f
C18448 VPWR.t548 VGND 0.02961f
C18449 VPWR.n941 VGND 0.09152f
C18450 VPWR.n942 VGND 0.13913f
C18451 VPWR.n943 VGND 0.13913f
C18452 VPWR.t540 VGND 0.03331f
C18453 VPWR.t731 VGND 0.02961f
C18454 VPWR.n944 VGND 0.09152f
C18455 VPWR.t431 VGND 0.07849f
C18456 VPWR.t730 VGND 0.09218f
C18457 VPWR.t1016 VGND 0.11957f
C18458 VPWR.t723 VGND 0.03331f
C18459 VPWR.t908 VGND 0.02961f
C18460 VPWR.n945 VGND 0.09152f
C18461 VPWR.n946 VGND 0.13913f
C18462 VPWR.n947 VGND 0.13913f
C18463 VPWR.t1017 VGND 0.03331f
C18464 VPWR.t1923 VGND 0.02961f
C18465 VPWR.n948 VGND 0.09152f
C18466 VPWR.t436 VGND 0.07849f
C18467 VPWR.t1922 VGND 0.09218f
C18468 VPWR.t638 VGND 0.11957f
C18469 VPWR.t1915 VGND 0.03331f
C18470 VPWR.t649 VGND 0.02961f
C18471 VPWR.n949 VGND 0.09152f
C18472 VPWR.n950 VGND 0.13913f
C18473 VPWR.n951 VGND 0.13913f
C18474 VPWR.t639 VGND 0.03331f
C18475 VPWR.t1101 VGND 0.02961f
C18476 VPWR.n952 VGND 0.09152f
C18477 VPWR.t1489 VGND 0.07849f
C18478 VPWR.t1100 VGND 0.09218f
C18479 VPWR.t1179 VGND 0.11957f
C18480 VPWR.t1052 VGND 0.03331f
C18481 VPWR.t1458 VGND 0.02961f
C18482 VPWR.n953 VGND 0.09152f
C18483 VPWR.n954 VGND 0.13913f
C18484 VPWR.n955 VGND 0.13913f
C18485 VPWR.t1180 VGND 0.03331f
C18486 VPWR.t1703 VGND 0.02961f
C18487 VPWR.n956 VGND 0.09152f
C18488 VPWR.t1456 VGND 0.07849f
C18489 VPWR.t1702 VGND 0.09218f
C18490 VPWR.t678 VGND 0.11957f
C18491 VPWR.t822 VGND 0.03331f
C18492 VPWR.t487 VGND 0.02961f
C18493 VPWR.n957 VGND 0.09152f
C18494 VPWR.n958 VGND 0.13913f
C18495 VPWR.n959 VGND 0.13913f
C18496 VPWR.t679 VGND 0.03331f
C18497 VPWR.t755 VGND 0.02961f
C18498 VPWR.n960 VGND 0.09152f
C18499 VPWR.t1454 VGND 0.07849f
C18500 VPWR.t754 VGND 0.09218f
C18501 VPWR.t627 VGND 0.03331f
C18502 VPWR.t337 VGND 0.02961f
C18503 VPWR.n961 VGND 0.09152f
C18504 VPWR.t763 VGND 0.03331f
C18505 VPWR.t189 VGND 0.02961f
C18506 VPWR.n962 VGND 0.09152f
C18507 VPWR.t1410 VGND 0.14512f
C18508 VPWR.t1260 VGND 0.07849f
C18509 VPWR.t712 VGND 0.09218f
C18510 VPWR.t1411 VGND 0.03331f
C18511 VPWR.t713 VGND 0.02961f
C18512 VPWR.n963 VGND 0.09152f
C18513 VPWR.n964 VGND 0.01797f
C18514 VPWR.n965 VGND 0.00728f
C18515 VPWR.n966 VGND 0.10822f
C18516 VPWR.t893 VGND 0.11957f
C18517 VPWR.t481 VGND 0.07849f
C18518 VPWR.t1088 VGND 0.09218f
C18519 VPWR.t894 VGND 0.03331f
C18520 VPWR.t1089 VGND 0.02961f
C18521 VPWR.n967 VGND 0.09152f
C18522 VPWR.n968 VGND 0.01797f
C18523 VPWR.n969 VGND 0.00728f
C18524 VPWR.n970 VGND 0.10822f
C18525 VPWR.t1084 VGND 0.11957f
C18526 VPWR.t525 VGND 0.07849f
C18527 VPWR.t1388 VGND 0.09218f
C18528 VPWR.t1085 VGND 0.03331f
C18529 VPWR.t1389 VGND 0.02961f
C18530 VPWR.n971 VGND 0.09152f
C18531 VPWR.n972 VGND 0.01797f
C18532 VPWR.n973 VGND 0.00728f
C18533 VPWR.n974 VGND 0.10822f
C18534 VPWR.t1354 VGND 0.11957f
C18535 VPWR.t524 VGND 0.07849f
C18536 VPWR.t1037 VGND 0.09218f
C18537 VPWR.t1355 VGND 0.03331f
C18538 VPWR.t1038 VGND 0.02961f
C18539 VPWR.n975 VGND 0.09152f
C18540 VPWR.n976 VGND 0.01797f
C18541 VPWR.n977 VGND 0.00728f
C18542 VPWR.n978 VGND 0.10822f
C18543 VPWR.t1638 VGND 0.11957f
C18544 VPWR.t796 VGND 0.07849f
C18545 VPWR.t519 VGND 0.09218f
C18546 VPWR.t1639 VGND 0.03331f
C18547 VPWR.t520 VGND 0.02961f
C18548 VPWR.n979 VGND 0.09152f
C18549 VPWR.n980 VGND 0.01797f
C18550 VPWR.n981 VGND 0.00728f
C18551 VPWR.n982 VGND 0.10822f
C18552 VPWR.t515 VGND 0.11957f
C18553 VPWR.t948 VGND 0.07849f
C18554 VPWR.t569 VGND 0.09218f
C18555 VPWR.t516 VGND 0.03331f
C18556 VPWR.t570 VGND 0.02961f
C18557 VPWR.n983 VGND 0.09152f
C18558 VPWR.n984 VGND 0.01797f
C18559 VPWR.n985 VGND 0.00728f
C18560 VPWR.n986 VGND 0.10822f
C18561 VPWR.t565 VGND 0.11957f
C18562 VPWR.t947 VGND 0.07849f
C18563 VPWR.t744 VGND 0.09218f
C18564 VPWR.t566 VGND 0.03331f
C18565 VPWR.t745 VGND 0.02961f
C18566 VPWR.n987 VGND 0.09152f
C18567 VPWR.n988 VGND 0.01797f
C18568 VPWR.n989 VGND 0.00728f
C18569 VPWR.n990 VGND 0.10822f
C18570 VPWR.t740 VGND 0.11957f
C18571 VPWR.t795 VGND 0.07849f
C18572 VPWR.t575 VGND 0.09218f
C18573 VPWR.t741 VGND 0.03331f
C18574 VPWR.t576 VGND 0.02961f
C18575 VPWR.n991 VGND 0.09152f
C18576 VPWR.n992 VGND 0.01797f
C18577 VPWR.n993 VGND 0.00728f
C18578 VPWR.n994 VGND 0.10822f
C18579 VPWR.t909 VGND 0.11957f
C18580 VPWR.t483 VGND 0.07849f
C18581 VPWR.t475 VGND 0.09218f
C18582 VPWR.t910 VGND 0.03331f
C18583 VPWR.t476 VGND 0.02961f
C18584 VPWR.n995 VGND 0.09152f
C18585 VPWR.n996 VGND 0.01797f
C18586 VPWR.n997 VGND 0.00728f
C18587 VPWR.n998 VGND 0.10822f
C18588 VPWR.t957 VGND 0.11957f
C18589 VPWR.t949 VGND 0.07849f
C18590 VPWR.t666 VGND 0.09218f
C18591 VPWR.t958 VGND 0.03331f
C18592 VPWR.t667 VGND 0.02961f
C18593 VPWR.n999 VGND 0.09152f
C18594 VPWR.n1000 VGND 0.01797f
C18595 VPWR.n1001 VGND 0.00728f
C18596 VPWR.n1002 VGND 0.10822f
C18597 VPWR.t614 VGND 0.11957f
C18598 VPWR.t523 VGND 0.07849f
C18599 VPWR.t1690 VGND 0.09218f
C18600 VPWR.t615 VGND 0.03331f
C18601 VPWR.t1691 VGND 0.02961f
C18602 VPWR.n1003 VGND 0.09152f
C18603 VPWR.n1004 VGND 0.01797f
C18604 VPWR.n1005 VGND 0.00728f
C18605 VPWR.n1006 VGND 0.10822f
C18606 VPWR.t1686 VGND 0.11957f
C18607 VPWR.t1261 VGND 0.07849f
C18608 VPWR.t473 VGND 0.09218f
C18609 VPWR.t1687 VGND 0.03331f
C18610 VPWR.t474 VGND 0.02961f
C18611 VPWR.n1007 VGND 0.09152f
C18612 VPWR.n1008 VGND 0.01797f
C18613 VPWR.n1009 VGND 0.00728f
C18614 VPWR.n1010 VGND 0.10822f
C18615 VPWR.t1764 VGND 0.11957f
C18616 VPWR.t946 VGND 0.07849f
C18617 VPWR.t463 VGND 0.09218f
C18618 VPWR.t1765 VGND 0.03331f
C18619 VPWR.t464 VGND 0.02961f
C18620 VPWR.n1011 VGND 0.09152f
C18621 VPWR.n1012 VGND 0.01797f
C18622 VPWR.n1013 VGND 0.00728f
C18623 VPWR.n1014 VGND 0.10822f
C18624 VPWR.t1704 VGND 0.11957f
C18625 VPWR.t945 VGND 0.07849f
C18626 VPWR.t1493 VGND 0.09218f
C18627 VPWR.t1705 VGND 0.03331f
C18628 VPWR.t1494 VGND 0.02961f
C18629 VPWR.n1015 VGND 0.09152f
C18630 VPWR.n1016 VGND 0.01797f
C18631 VPWR.n1017 VGND 0.00728f
C18632 VPWR.n1018 VGND 0.10822f
C18633 VPWR.t1174 VGND 0.11957f
C18634 VPWR.t526 VGND 0.07849f
C18635 VPWR.t1806 VGND 0.09218f
C18636 VPWR.t1175 VGND 0.03331f
C18637 VPWR.t1807 VGND 0.02961f
C18638 VPWR.n1019 VGND 0.09152f
C18639 VPWR.n1020 VGND 0.01797f
C18640 VPWR.n1021 VGND 0.00728f
C18641 VPWR.n1022 VGND 0.10822f
C18642 VPWR.t762 VGND 0.11957f
C18643 VPWR.t482 VGND 0.07849f
C18644 VPWR.t188 VGND 0.13333f
C18645 VPWR.n1023 VGND 0.07618f
C18646 VPWR.n1024 VGND 0.01797f
C18647 VPWR.n1025 VGND 0.13913f
C18648 VPWR.n1026 VGND 6.02311f
C18649 VPWR.n1027 VGND 0.06567f
C18650 VPWR.n1028 VGND -0.01866f
C18651 VPWR.t2061 VGND 0.01116f
C18652 VPWR.t190 VGND 0.01222f
C18653 VPWR.n1029 VGND 0.03042f
C18654 VPWR.n1030 VGND 0.00581f
C18655 VPWR.t192 VGND 0.02679f
C18656 VPWR.n1031 VGND 0.05724f
C18657 VPWR.t300 VGND 0.02961f
C18658 VPWR.n1032 VGND 0.04692f
C18659 VPWR.t764 VGND 0.09218f
C18660 VPWR.t1957 VGND 0.01116f
C18661 VPWR.t82 VGND 0.01222f
C18662 VPWR.n1033 VGND 0.03042f
C18663 VPWR.n1034 VGND 0.00581f
C18664 VPWR.t84 VGND 0.02679f
C18665 VPWR.n1035 VGND 0.05724f
C18666 VPWR.t765 VGND 0.02961f
C18667 VPWR.n1036 VGND 0.04692f
C18668 VPWR.n1037 VGND -0.01866f
C18669 VPWR.n1038 VGND 0.06567f
C18670 VPWR.t2065 VGND 0.01136f
C18671 VPWR.t38 VGND 0.0124f
C18672 VPWR.n1039 VGND 0.02769f
C18673 VPWR.n1040 VGND 0.01897f
C18674 VPWR.n1041 VGND 0.06244f
C18675 VPWR.n1042 VGND 0.09746f
C18676 VPWR.n1043 VGND 0.0544f
C18677 VPWR.n1044 VGND 0.06567f
C18678 VPWR.n1045 VGND -0.01866f
C18679 VPWR.t1967 VGND 0.01116f
C18680 VPWR.t168 VGND 0.01222f
C18681 VPWR.n1046 VGND 0.03042f
C18682 VPWR.n1047 VGND 0.00581f
C18683 VPWR.t170 VGND 0.02679f
C18684 VPWR.n1048 VGND 0.05724f
C18685 VPWR.t1171 VGND 0.02961f
C18686 VPWR.n1049 VGND 0.04692f
C18687 VPWR.t1170 VGND 0.09218f
C18688 VPWR.t46 VGND 0.11957f
C18689 VPWR.t2055 VGND 0.01116f
C18690 VPWR.t209 VGND 0.01222f
C18691 VPWR.n1050 VGND 0.03042f
C18692 VPWR.n1051 VGND 0.00581f
C18693 VPWR.t211 VGND 0.02679f
C18694 VPWR.n1052 VGND 0.05724f
C18695 VPWR.t450 VGND 0.02961f
C18696 VPWR.n1053 VGND 0.04692f
C18697 VPWR.n1054 VGND 0.00805f
C18698 VPWR.n1055 VGND 0.19371f
C18699 VPWR.n1056 VGND 0.08351f
C18700 VPWR.n1057 VGND 0.03437f
C18701 VPWR.t264 VGND 0.03331f
C18702 VPWR.t256 VGND 0.02961f
C18703 VPWR.n1058 VGND 0.09152f
C18704 VPWR.t255 VGND 0.09218f
C18705 VPWR.t11 VGND 0.11957f
C18706 VPWR.t292 VGND 0.03331f
C18707 VPWR.t284 VGND 0.02961f
C18708 VPWR.n1059 VGND 0.09152f
C18709 VPWR.n1060 VGND 0.00805f
C18710 VPWR.t12 VGND 0.03331f
C18711 VPWR.t135 VGND 0.02961f
C18712 VPWR.n1061 VGND 0.09152f
C18713 VPWR.t7 VGND 0.07849f
C18714 VPWR.t134 VGND 0.13333f
C18715 VPWR.n1062 VGND 0.07615f
C18716 VPWR.n1063 VGND 0.01698f
C18717 VPWR.t2034 VGND 0.0112f
C18718 VPWR.t133 VGND 0.01226f
C18719 VPWR.n1064 VGND 0.02993f
C18720 VPWR.n1065 VGND 0.03284f
C18721 VPWR.n1066 VGND 0.00697f
C18722 VPWR.n1067 VGND 0.01822f
C18723 VPWR.n1068 VGND 0.17585f
C18724 VPWR.t1989 VGND 0.0112f
C18725 VPWR.t254 VGND 0.01226f
C18726 VPWR.n1069 VGND 0.02993f
C18727 VPWR.n1070 VGND 0.03284f
C18728 VPWR.n1071 VGND 0.01714f
C18729 VPWR.n1072 VGND 0.00697f
C18730 VPWR.n1073 VGND 0.00805f
C18731 VPWR.n1074 VGND 0.01714f
C18732 VPWR.n1075 VGND 0.00697f
C18733 VPWR.t1988 VGND 0.01136f
C18734 VPWR.t260 VGND 0.0124f
C18735 VPWR.n1076 VGND 0.02768f
C18736 VPWR.n1077 VGND 0.02818f
C18737 VPWR.n1078 VGND 0.01822f
C18738 VPWR.n1079 VGND 0.17585f
C18739 VPWR.t1947 VGND 0.0112f
C18740 VPWR.t362 VGND 0.01226f
C18741 VPWR.n1080 VGND 0.02993f
C18742 VPWR.n1081 VGND 0.03284f
C18743 VPWR.n1082 VGND 0.01714f
C18744 VPWR.n1083 VGND 0.00697f
C18745 VPWR.n1084 VGND 0.01714f
C18746 VPWR.n1085 VGND 0.00697f
C18747 VPWR.t1945 VGND 0.01136f
C18748 VPWR.t368 VGND 0.0124f
C18749 VPWR.n1086 VGND 0.02768f
C18750 VPWR.n1087 VGND 0.02818f
C18751 VPWR.n1088 VGND 0.01822f
C18752 VPWR.n1089 VGND 0.17585f
C18753 VPWR.t1949 VGND 0.0112f
C18754 VPWR.t354 VGND 0.01226f
C18755 VPWR.n1090 VGND 0.02993f
C18756 VPWR.n1091 VGND 0.03284f
C18757 VPWR.n1092 VGND 0.01714f
C18758 VPWR.n1093 VGND 0.00697f
C18759 VPWR.n1094 VGND 0.01714f
C18760 VPWR.n1095 VGND 0.00697f
C18761 VPWR.t2049 VGND 0.01136f
C18762 VPWR.t87 VGND 0.0124f
C18763 VPWR.n1096 VGND 0.02768f
C18764 VPWR.n1097 VGND 0.02818f
C18765 VPWR.n1098 VGND 0.01822f
C18766 VPWR.n1099 VGND 0.17585f
C18767 VPWR.t2059 VGND 0.0112f
C18768 VPWR.t59 VGND 0.01226f
C18769 VPWR.n1100 VGND 0.02993f
C18770 VPWR.n1101 VGND 0.03284f
C18771 VPWR.n1102 VGND 0.01714f
C18772 VPWR.n1103 VGND 0.00697f
C18773 VPWR.n1104 VGND 0.01714f
C18774 VPWR.n1105 VGND 0.00697f
C18775 VPWR.t2014 VGND 0.01136f
C18776 VPWR.t171 VGND 0.0124f
C18777 VPWR.n1106 VGND 0.02768f
C18778 VPWR.n1107 VGND 0.02818f
C18779 VPWR.n1108 VGND 0.01822f
C18780 VPWR.n1109 VGND 0.02654f
C18781 VPWR.t2018 VGND 0.0112f
C18782 VPWR.t165 VGND 0.01226f
C18783 VPWR.n1110 VGND 0.02993f
C18784 VPWR.n1111 VGND 0.03284f
C18785 VPWR.n1112 VGND 0.01822f
C18786 VPWR.n1113 VGND 0.00697f
C18787 VPWR.t2012 VGND 0.01116f
C18788 VPWR.t311 VGND 0.01222f
C18789 VPWR.n1114 VGND 0.03115f
C18790 VPWR.n1115 VGND 0.01969f
C18791 VPWR.t1969 VGND 0.01136f
C18792 VPWR.t301 VGND 0.0124f
C18793 VPWR.n1116 VGND 0.02768f
C18794 VPWR.n1117 VGND 0.02818f
C18795 VPWR.n1118 VGND 0.01776f
C18796 VPWR.t2067 VGND 0.0112f
C18797 VPWR.t29 VGND 0.01226f
C18798 VPWR.n1119 VGND 0.02993f
C18799 VPWR.n1120 VGND 0.03284f
C18800 VPWR.n1121 VGND 0.00805f
C18801 VPWR.t313 VGND 0.03331f
C18802 VPWR.t31 VGND 0.02961f
C18803 VPWR.n1122 VGND 0.09152f
C18804 VPWR.t312 VGND 0.14512f
C18805 VPWR.t302 VGND 0.07849f
C18806 VPWR.t30 VGND 0.09218f
C18807 VPWR.t185 VGND 0.11957f
C18808 VPWR.t81 VGND 0.03331f
C18809 VPWR.t167 VGND 0.02961f
C18810 VPWR.n1123 VGND 0.09152f
C18811 VPWR.n1124 VGND 0.00833f
C18812 VPWR.t2062 VGND 0.01116f
C18813 VPWR.t184 VGND 0.01222f
C18814 VPWR.n1125 VGND 0.03115f
C18815 VPWR.n1126 VGND 0.03694f
C18816 VPWR.n1127 VGND 0.03437f
C18817 VPWR.n1128 VGND 0.13913f
C18818 VPWR.n1129 VGND 0.00805f
C18819 VPWR.n1130 VGND 0.01797f
C18820 VPWR.n1131 VGND 0.06567f
C18821 VPWR.n1132 VGND 0.0544f
C18822 VPWR.t1950 VGND 0.01136f
C18823 VPWR.t352 VGND 0.0124f
C18824 VPWR.n1133 VGND 0.02769f
C18825 VPWR.n1134 VGND 0.01897f
C18826 VPWR.n1135 VGND 0.06244f
C18827 VPWR.n1136 VGND 0.09746f
C18828 VPWR.n1137 VGND 0.06567f
C18829 VPWR.n1138 VGND 0.06567f
C18830 VPWR.n1139 VGND 0.06567f
C18831 VPWR.n1140 VGND 0.06567f
C18832 VPWR.n1141 VGND 0.06567f
C18833 VPWR.n1142 VGND 0.06567f
C18834 VPWR.n1143 VGND 0.0544f
C18835 VPWR.n1144 VGND 0.00805f
C18836 VPWR.n1145 VGND -0.01866f
C18837 VPWR.t2020 VGND 0.01116f
C18838 VPWR.t295 VGND 0.01222f
C18839 VPWR.n1146 VGND 0.03042f
C18840 VPWR.n1147 VGND 0.00581f
C18841 VPWR.t297 VGND 0.02679f
C18842 VPWR.n1148 VGND 0.05724f
C18843 VPWR.t1789 VGND 0.02961f
C18844 VPWR.n1149 VGND 0.04692f
C18845 VPWR.t1788 VGND 0.09218f
C18846 VPWR.t39 VGND 0.07849f
C18847 VPWR.t169 VGND 0.11957f
C18848 VPWR.t1975 VGND 0.01116f
C18849 VPWR.t35 VGND 0.01222f
C18850 VPWR.n1150 VGND 0.03042f
C18851 VPWR.n1151 VGND 0.00581f
C18852 VPWR.t37 VGND 0.02679f
C18853 VPWR.n1152 VGND 0.05724f
C18854 VPWR.t1107 VGND 0.02961f
C18855 VPWR.n1153 VGND 0.04692f
C18856 VPWR.n1154 VGND 0.00805f
C18857 VPWR.n1155 VGND 0.00805f
C18858 VPWR.t1927 VGND 0.01116f
C18859 VPWR.t279 VGND 0.01222f
C18860 VPWR.n1156 VGND 0.03042f
C18861 VPWR.n1157 VGND 0.00581f
C18862 VPWR.t281 VGND 0.02679f
C18863 VPWR.n1158 VGND 0.05724f
C18864 VPWR.t1484 VGND 0.02961f
C18865 VPWR.n1159 VGND 0.04692f
C18866 VPWR.t854 VGND 0.09218f
C18867 VPWR.t1938 VGND 0.01116f
C18868 VPWR.t138 VGND 0.01222f
C18869 VPWR.n1160 VGND 0.03042f
C18870 VPWR.n1161 VGND 0.00581f
C18871 VPWR.t140 VGND 0.02679f
C18872 VPWR.n1162 VGND 0.05724f
C18873 VPWR.t855 VGND 0.02961f
C18874 VPWR.n1163 VGND 0.04692f
C18875 VPWR.n1164 VGND 0.00805f
C18876 VPWR.n1165 VGND 0.00805f
C18877 VPWR.t2023 VGND 0.01116f
C18878 VPWR.t16 VGND 0.01222f
C18879 VPWR.n1166 VGND 0.03042f
C18880 VPWR.n1167 VGND 0.00581f
C18881 VPWR.t18 VGND 0.02679f
C18882 VPWR.n1168 VGND 0.05724f
C18883 VPWR.t1795 VGND 0.02961f
C18884 VPWR.n1169 VGND 0.04692f
C18885 VPWR.t690 VGND 0.09218f
C18886 VPWR.t2035 VGND 0.01116f
C18887 VPWR.t265 VGND 0.01222f
C18888 VPWR.n1170 VGND 0.03042f
C18889 VPWR.n1171 VGND 0.00581f
C18890 VPWR.t267 VGND 0.02679f
C18891 VPWR.n1172 VGND 0.05724f
C18892 VPWR.t691 VGND 0.02961f
C18893 VPWR.n1173 VGND 0.04692f
C18894 VPWR.n1174 VGND 0.00805f
C18895 VPWR.n1175 VGND 0.00833f
C18896 VPWR.t1958 VGND 0.01116f
C18897 VPWR.t76 VGND 0.01222f
C18898 VPWR.n1176 VGND 0.03115f
C18899 VPWR.n1177 VGND 0.03694f
C18900 VPWR.n1178 VGND 0.03437f
C18901 VPWR.t66 VGND 0.03331f
C18902 VPWR.t61 VGND 0.02961f
C18903 VPWR.n1179 VGND 0.09152f
C18904 VPWR.t172 VGND 0.07849f
C18905 VPWR.t179 VGND 0.09218f
C18906 VPWR.t186 VGND 0.03331f
C18907 VPWR.t180 VGND 0.02961f
C18908 VPWR.n1180 VGND 0.09152f
C18909 VPWR.n1181 VGND 0.00725f
C18910 VPWR.n1182 VGND 0.10822f
C18911 VPWR.t347 VGND 0.11957f
C18912 VPWR.t213 VGND 0.07849f
C18913 VPWR.t339 VGND 0.09218f
C18914 VPWR.t348 VGND 0.03331f
C18915 VPWR.t340 VGND 0.02961f
C18916 VPWR.n1183 VGND 0.09152f
C18917 VPWR.n1184 VGND 0.00725f
C18918 VPWR.n1185 VGND 0.10822f
C18919 VPWR.t65 VGND 0.11957f
C18920 VPWR.t321 VGND 0.07849f
C18921 VPWR.t60 VGND 0.09218f
C18922 VPWR.t137 VGND 0.07849f
C18923 VPWR.t263 VGND 0.11957f
C18924 VPWR.t26 VGND 0.03331f
C18925 VPWR.t127 VGND 0.02961f
C18926 VPWR.n1186 VGND 0.09152f
C18927 VPWR.n1187 VGND 0.00725f
C18928 VPWR.n1188 VGND 0.10822f
C18929 VPWR.t126 VGND 0.09218f
C18930 VPWR.t111 VGND 0.07849f
C18931 VPWR.t25 VGND 0.11957f
C18932 VPWR.t5 VGND 0.03331f
C18933 VPWR.t383 VGND 0.02961f
C18934 VPWR.n1189 VGND 0.09152f
C18935 VPWR.n1190 VGND 0.00725f
C18936 VPWR.n1191 VGND 0.10822f
C18937 VPWR.t382 VGND 0.09218f
C18938 VPWR.t261 VGND 0.07849f
C18939 VPWR.t4 VGND 0.11957f
C18940 VPWR.t259 VGND 0.03331f
C18941 VPWR.t364 VGND 0.02961f
C18942 VPWR.n1192 VGND 0.09152f
C18943 VPWR.n1193 VGND 0.00833f
C18944 VPWR.t2031 VGND 0.01116f
C18945 VPWR.t3 VGND 0.01222f
C18946 VPWR.n1194 VGND 0.03115f
C18947 VPWR.n1195 VGND 0.03694f
C18948 VPWR.n1196 VGND 0.03437f
C18949 VPWR.n1197 VGND 0.01714f
C18950 VPWR.n1198 VGND 0.00725f
C18951 VPWR.n1199 VGND 0.10822f
C18952 VPWR.t363 VGND 0.09218f
C18953 VPWR.t239 VGND 0.07849f
C18954 VPWR.t258 VGND 0.11957f
C18955 VPWR.t132 VGND 0.03331f
C18956 VPWR.t205 VGND 0.02961f
C18957 VPWR.n1200 VGND 0.09152f
C18958 VPWR.n1201 VGND 0.00725f
C18959 VPWR.n1202 VGND 0.10822f
C18960 VPWR.t204 VGND 0.09218f
C18961 VPWR.t86 VGND 0.07849f
C18962 VPWR.t131 VGND 0.11957f
C18963 VPWR.t106 VGND 0.03331f
C18964 VPWR.t101 VGND 0.02961f
C18965 VPWR.n1203 VGND 0.09152f
C18966 VPWR.n1204 VGND 0.00725f
C18967 VPWR.n1205 VGND 0.10822f
C18968 VPWR.t100 VGND 0.09218f
C18969 VPWR.t369 VGND 0.07849f
C18970 VPWR.t105 VGND 0.11957f
C18971 VPWR.t345 VGND 0.03331f
C18972 VPWR.t356 VGND 0.02961f
C18973 VPWR.n1206 VGND 0.09152f
C18974 VPWR.n1207 VGND 0.00833f
C18975 VPWR.t1992 VGND 0.01116f
C18976 VPWR.t104 VGND 0.01222f
C18977 VPWR.n1208 VGND 0.03115f
C18978 VPWR.n1209 VGND 0.03694f
C18979 VPWR.n1210 VGND 0.03437f
C18980 VPWR.n1211 VGND 0.01714f
C18981 VPWR.n1212 VGND 0.00725f
C18982 VPWR.n1213 VGND 0.10822f
C18983 VPWR.t355 VGND 0.09218f
C18984 VPWR.t326 VGND 0.07849f
C18985 VPWR.t344 VGND 0.11957f
C18986 VPWR.t237 VGND 0.03331f
C18987 VPWR.t316 VGND 0.02961f
C18988 VPWR.n1214 VGND 0.09152f
C18989 VPWR.n1215 VGND 0.00725f
C18990 VPWR.n1216 VGND 0.10822f
C18991 VPWR.t315 VGND 0.09218f
C18992 VPWR.t103 VGND 0.07849f
C18993 VPWR.t236 VGND 0.11957f
C18994 VPWR.t78 VGND 0.03331f
C18995 VPWR.t208 VGND 0.02961f
C18996 VPWR.n1217 VGND 0.09152f
C18997 VPWR.n1218 VGND 0.00725f
C18998 VPWR.n1219 VGND 0.10822f
C18999 VPWR.t207 VGND 0.09218f
C19000 VPWR.t88 VGND 0.07849f
C19001 VPWR.t77 VGND 0.11957f
C19002 VPWR.n1220 VGND 0.10822f
C19003 VPWR.n1221 VGND 0.00725f
C19004 VPWR.n1222 VGND 0.01714f
C19005 VPWR.n1223 VGND 0.00805f
C19006 VPWR.t2041 VGND 0.01116f
C19007 VPWR.t243 VGND 0.01222f
C19008 VPWR.n1224 VGND 0.03042f
C19009 VPWR.n1225 VGND 0.00581f
C19010 VPWR.t245 VGND 0.02679f
C19011 VPWR.n1226 VGND 0.05724f
C19012 VPWR.t1224 VGND 0.02961f
C19013 VPWR.n1227 VGND 0.04692f
C19014 VPWR.t108 VGND 0.14512f
C19015 VPWR.t93 VGND 0.07849f
C19016 VPWR.t974 VGND 0.09218f
C19017 VPWR.t1948 VGND 0.01116f
C19018 VPWR.t107 VGND 0.01222f
C19019 VPWR.n1228 VGND 0.03042f
C19020 VPWR.n1229 VGND 0.00581f
C19021 VPWR.t109 VGND 0.02679f
C19022 VPWR.n1230 VGND 0.05724f
C19023 VPWR.t975 VGND 0.02961f
C19024 VPWR.n1231 VGND 0.04692f
C19025 VPWR.n1232 VGND -0.01866f
C19026 VPWR.n1233 VGND 0.04687f
C19027 VPWR.t437 VGND 0.97566f
C19028 VPWR.n1234 VGND 0.53213f
C19029 VPWR.t443 VGND 0.97566f
C19030 VPWR.n1235 VGND 0.41384f
C19031 VPWR.n1236 VGND 0.2908f
C19032 VPWR.t506 VGND 0.05716f
C19033 VPWR.n1237 VGND 0.0092f
C19034 VPWR.t1090 VGND 0.01433f
C19035 VPWR.t874 VGND 0.01433f
C19036 VPWR.n1238 VGND 0.03146f
C19037 VPWR.t875 VGND 0.01433f
C19038 VPWR.t1710 VGND 0.01433f
C19039 VPWR.n1239 VGND 0.03141f
C19040 VPWR.t1865 VGND 0.01433f
C19041 VPWR.t1864 VGND 0.01433f
C19042 VPWR.n1240 VGND 0.03141f
C19043 VPWR.n1241 VGND 0.1042f
C19044 VPWR.n1242 VGND 0.18182f
C19045 VPWR.n1243 VGND 0.05756f
C19046 VPWR.n1244 VGND 0.04228f
C19047 VPWR.t1861 VGND 0.01433f
C19048 VPWR.t1866 VGND 0.01433f
C19049 VPWR.n1245 VGND 0.03146f
C19050 VPWR.n1246 VGND 0.12902f
C19051 VPWR.n1247 VGND 0.01119f
C19052 VPWR.n1248 VGND 0.0163f
C19053 VPWR.n1249 VGND 0.0191f
C19054 VPWR.n1250 VGND 0.02802f
C19055 VPWR.t504 VGND 0.05716f
C19056 VPWR.n1251 VGND 0.15059f
C19057 VPWR.n1252 VGND 0.01209f
C19058 VPWR.t1093 VGND 0.05714f
C19059 VPWR.t1262 VGND 0.05714f
C19060 VPWR.n1253 VGND 0.13446f
C19061 VPWR.n1254 VGND 0.33563f
C19062 VPWR.n1255 VGND 1.64092f
C19063 VPWR.n1256 VGND 0.04687f
C19064 VPWR.t442 VGND 0.97566f
C19065 VPWR.n1257 VGND 0.53213f
C19066 VPWR.t507 VGND 0.97566f
C19067 VPWR.n1258 VGND 0.41384f
C19068 VPWR.n1259 VGND 0.29342f
C19069 VPWR.n1260 VGND 0.0092f
C19070 VPWR.t782 VGND 0.01433f
C19071 VPWR.t780 VGND 0.01433f
C19072 VPWR.n1261 VGND 0.03146f
C19073 VPWR.t779 VGND 0.01433f
C19074 VPWR.t776 VGND 0.01433f
C19075 VPWR.n1262 VGND 0.03141f
C19076 VPWR.t1668 VGND 0.01433f
C19077 VPWR.t1669 VGND 0.01433f
C19078 VPWR.n1263 VGND 0.03141f
C19079 VPWR.n1264 VGND 0.1042f
C19080 VPWR.n1265 VGND 0.18182f
C19081 VPWR.n1266 VGND 0.05756f
C19082 VPWR.n1267 VGND 0.04228f
C19083 VPWR.t1177 VGND 0.01433f
C19084 VPWR.t1679 VGND 0.01433f
C19085 VPWR.n1268 VGND 0.03146f
C19086 VPWR.n1269 VGND 0.12902f
C19087 VPWR.n1270 VGND 0.01119f
C19088 VPWR.n1271 VGND 0.0163f
C19089 VPWR.n1272 VGND 0.0191f
C19090 VPWR.n1273 VGND 0.02751f
C19091 VPWR.n1274 VGND 0.00767f
C19092 VPWR.t508 VGND 0.05708f
C19093 VPWR.n1275 VGND 0.06101f
C19094 VPWR.n1276 VGND 0.00731f
C19095 VPWR.t1721 VGND 0.0572f
C19096 VPWR.n1277 VGND 0.0911f
C19097 VPWR.n1278 VGND 0.33563f
C19098 VPWR.n1279 VGND 1.64092f
C19099 VPWR.n1280 VGND 0.04687f
C19100 VPWR.t505 VGND 0.97566f
C19101 VPWR.n1281 VGND 0.53213f
C19102 VPWR.t413 VGND 0.97566f
C19103 VPWR.n1282 VGND 0.41384f
C19104 VPWR.n1283 VGND 0.29342f
C19105 VPWR.n1284 VGND 0.0092f
C19106 VPWR.t773 VGND 0.01433f
C19107 VPWR.t771 VGND 0.01433f
C19108 VPWR.n1285 VGND 0.03146f
C19109 VPWR.t770 VGND 0.01433f
C19110 VPWR.t769 VGND 0.01433f
C19111 VPWR.n1286 VGND 0.03141f
C19112 VPWR.t654 VGND 0.01433f
C19113 VPWR.t661 VGND 0.01433f
C19114 VPWR.n1287 VGND 0.03141f
C19115 VPWR.n1288 VGND 0.1042f
C19116 VPWR.n1289 VGND 0.18182f
C19117 VPWR.n1290 VGND 0.05756f
C19118 VPWR.n1291 VGND 0.04228f
C19119 VPWR.t658 VGND 0.01433f
C19120 VPWR.t655 VGND 0.01433f
C19121 VPWR.n1292 VGND 0.03146f
C19122 VPWR.n1293 VGND 0.12902f
C19123 VPWR.n1294 VGND 0.01119f
C19124 VPWR.n1295 VGND 0.0163f
C19125 VPWR.n1296 VGND 0.0191f
C19126 VPWR.n1297 VGND 0.02751f
C19127 VPWR.n1298 VGND 0.01398f
C19128 VPWR.n1299 VGND 0.01308f
C19129 VPWR.t1094 VGND 0.0572f
C19130 VPWR.t1263 VGND 0.0572f
C19131 VPWR.n1300 VGND 0.16894f
C19132 VPWR.n1301 VGND 0.33563f
C19133 VPWR.n1302 VGND 1.64092f
C19134 VPWR.t1745 VGND 0.05711f
C19135 VPWR.t987 VGND 0.0572f
C19136 VPWR.t1747 VGND 0.05672f
C19137 VPWR.n1303 VGND 0.14706f
C19138 VPWR.t588 VGND 0.05606f
C19139 VPWR.n1304 VGND 0.06775f
C19140 VPWR.n1305 VGND 0.04687f
C19141 VPWR.t873 VGND 0.05397f
C19142 VPWR.n1306 VGND 0.05133f
C19143 VPWR.t1504 VGND 0.01433f
C19144 VPWR.t934 VGND 0.01433f
C19145 VPWR.n1307 VGND 0.03131f
C19146 VPWR.t415 VGND 0.05015f
C19147 VPWR.n1308 VGND 0.07521f
C19148 VPWR.n1309 VGND 0.04687f
C19149 VPWR.t585 VGND 0.05714f
C19150 VPWR.n1310 VGND 0.07193f
C19151 VPWR.n1311 VGND 0.02751f
C19152 VPWR.n1312 VGND 0.04687f
C19153 VPWR.n1313 VGND 0.01209f
C19154 VPWR.t1539 VGND 0.01433f
C19155 VPWR.t1541 VGND 0.01433f
C19156 VPWR.n1314 VGND 0.03131f
C19157 VPWR.n1315 VGND 0.04588f
C19158 VPWR.n1316 VGND 0.01209f
C19159 VPWR.n1317 VGND 0.03515f
C19160 VPWR.n1318 VGND 0.03515f
C19161 VPWR.n1319 VGND 0.04687f
C19162 VPWR.n1320 VGND 0.0083f
C19163 VPWR.t1500 VGND 0.01433f
C19164 VPWR.t991 VGND 0.01433f
C19165 VPWR.n1321 VGND 0.03131f
C19166 VPWR.n1322 VGND 0.03605f
C19167 VPWR.t439 VGND 0.01433f
C19168 VPWR.t1743 VGND 0.01433f
C19169 VPWR.n1323 VGND 0.03131f
C19170 VPWR.n1324 VGND 0.03983f
C19171 VPWR.n1325 VGND 0.01055f
C19172 VPWR.n1326 VGND 0.04254f
C19173 VPWR.n1327 VGND 0.01605f
C19174 VPWR.n1328 VGND 0.00631f
C19175 VPWR.t950 VGND 0.04806f
C19176 VPWR.t1744 VGND 0.10812f
C19177 VPWR.t986 VGND 0.12614f
C19178 VPWR.t1746 VGND 0.23427f
C19179 VPWR.t584 VGND 0.12605f
C19180 VPWR.t1540 VGND 0.14308f
C19181 VPWR.t1538 VGND 0.1391f
C19182 VPWR.t933 VGND 0.22247f
C19183 VPWR.t1503 VGND 0.18922f
C19184 VPWR.t414 VGND 0.12614f
C19185 VPWR.t990 VGND 0.12614f
C19186 VPWR.t1742 VGND 0.12614f
C19187 VPWR.t1499 VGND 0.12614f
C19188 VPWR.t438 VGND 0.12614f
C19189 VPWR.t872 VGND 0.12614f
C19190 VPWR.t587 VGND 0.12464f
C19191 VPWR.n1329 VGND 0.4287f
C19192 VPWR.n1330 VGND 0.17419f
C19193 VPWR.n1331 VGND 0.0191f
C19194 VPWR.n1332 VGND 0.03515f
C19195 VPWR.n1333 VGND 0.04228f
C19196 VPWR.n1334 VGND 0.01083f
C19197 VPWR.n1335 VGND 0.06357f
C19198 VPWR.n1336 VGND 0.31652f
C19199 VPWR.n1337 VGND 1.64092f
C19200 VPWR.t1470 VGND 0.05619f
C19201 VPWR.t971 VGND 0.05603f
C19202 VPWR.t985 VGND 0.05714f
C19203 VPWR.n1338 VGND 0.07963f
C19204 VPWR.t876 VGND 0.05456f
C19205 VPWR.t1867 VGND 0.05456f
C19206 VPWR.n1339 VGND 0.09898f
C19207 VPWR.n1340 VGND 0.04687f
C19208 VPWR.n1341 VGND 0.00911f
C19209 VPWR.n1342 VGND 0.04687f
C19210 VPWR.t1091 VGND 0.01433f
C19211 VPWR.t1257 VGND 0.01433f
C19212 VPWR.n1343 VGND 0.03131f
C19213 VPWR.t1868 VGND 0.01433f
C19214 VPWR.t447 VGND 0.01433f
C19215 VPWR.n1344 VGND 0.03131f
C19216 VPWR.n1345 VGND 0.06379f
C19217 VPWR.t1869 VGND 0.05714f
C19218 VPWR.t1542 VGND 0.05714f
C19219 VPWR.n1346 VGND 0.13169f
C19220 VPWR.n1347 VGND 0.02751f
C19221 VPWR.n1348 VGND 0.04687f
C19222 VPWR.n1349 VGND 0.01209f
C19223 VPWR.t1259 VGND 0.01433f
C19224 VPWR.t580 VGND 0.01433f
C19225 VPWR.n1350 VGND 0.03131f
C19226 VPWR.t1872 VGND 0.01433f
C19227 VPWR.t1875 VGND 0.01433f
C19228 VPWR.n1351 VGND 0.03131f
C19229 VPWR.n1352 VGND 0.07209f
C19230 VPWR.n1353 VGND 0.01209f
C19231 VPWR.n1354 VGND 0.04687f
C19232 VPWR.n1355 VGND 0.04687f
C19233 VPWR.n1356 VGND 0.04687f
C19234 VPWR.n1357 VGND 0.01128f
C19235 VPWR.t1711 VGND 0.01433f
C19236 VPWR.t1092 VGND 0.01433f
C19237 VPWR.n1358 VGND 0.03131f
C19238 VPWR.t1863 VGND 0.01433f
C19239 VPWR.t1862 VGND 0.01433f
C19240 VPWR.n1359 VGND 0.03131f
C19241 VPWR.n1360 VGND 0.06379f
C19242 VPWR.n1361 VGND 0.01055f
C19243 VPWR.n1362 VGND 0.00983f
C19244 VPWR.n1363 VGND 0.04687f
C19245 VPWR.n1364 VGND 0.03515f
C19246 VPWR.n1365 VGND 0.00794f
C19247 VPWR.t579 VGND 0.97566f
C19248 VPWR.n1366 VGND 0.53213f
C19249 VPWR.t446 VGND 0.97566f
C19250 VPWR.n1367 VGND 0.41384f
C19251 VPWR.n1368 VGND 0.2908f
C19252 VPWR.n1369 VGND 0.0191f
C19253 VPWR.n1370 VGND 0.03515f
C19254 VPWR.n1371 VGND 0.04254f
C19255 VPWR.n1372 VGND 0.01064f
C19256 VPWR.n1373 VGND 0.05827f
C19257 VPWR.n1374 VGND 0.07893f
C19258 VPWR.n1375 VGND 0.31627f
C19259 VPWR.n1376 VGND 1.64092f
C19260 VPWR.t1024 VGND 0.05708f
C19261 VPWR.t1622 VGND 0.05708f
C19262 VPWR.n1377 VGND 0.01398f
C19263 VPWR.t778 VGND 0.05456f
C19264 VPWR.t1178 VGND 0.05456f
C19265 VPWR.n1378 VGND 0.09898f
C19266 VPWR.n1379 VGND 0.04687f
C19267 VPWR.n1380 VGND 0.00911f
C19268 VPWR.n1381 VGND 0.04687f
C19269 VPWR.t783 VGND 0.01433f
C19270 VPWR.t1870 VGND 0.01433f
C19271 VPWR.n1382 VGND 0.03131f
C19272 VPWR.t1850 VGND 0.01433f
C19273 VPWR.t1543 VGND 0.01433f
C19274 VPWR.n1383 VGND 0.03131f
C19275 VPWR.n1384 VGND 0.06379f
C19276 VPWR.t1255 VGND 0.05714f
C19277 VPWR.t445 VGND 0.05714f
C19278 VPWR.n1385 VGND 0.13169f
C19279 VPWR.n1386 VGND 0.02751f
C19280 VPWR.n1387 VGND 0.04687f
C19281 VPWR.n1388 VGND 0.01209f
C19282 VPWR.t1874 VGND 0.01433f
C19283 VPWR.t1741 VGND 0.01433f
C19284 VPWR.n1389 VGND 0.03131f
C19285 VPWR.t1256 VGND 0.01433f
C19286 VPWR.t1787 VGND 0.01433f
C19287 VPWR.n1390 VGND 0.03131f
C19288 VPWR.n1391 VGND 0.07209f
C19289 VPWR.n1392 VGND 0.01209f
C19290 VPWR.n1393 VGND 0.04687f
C19291 VPWR.n1394 VGND 0.04687f
C19292 VPWR.n1395 VGND 0.04687f
C19293 VPWR.n1396 VGND 0.01128f
C19294 VPWR.t784 VGND 0.01433f
C19295 VPWR.t781 VGND 0.01433f
C19296 VPWR.n1397 VGND 0.03131f
C19297 VPWR.t1670 VGND 0.01433f
C19298 VPWR.t1176 VGND 0.01433f
C19299 VPWR.n1398 VGND 0.03131f
C19300 VPWR.n1399 VGND 0.06379f
C19301 VPWR.n1400 VGND 0.01055f
C19302 VPWR.n1401 VGND 0.00983f
C19303 VPWR.n1402 VGND 0.04687f
C19304 VPWR.n1403 VGND 0.03515f
C19305 VPWR.n1404 VGND 0.00794f
C19306 VPWR.t777 VGND 0.97566f
C19307 VPWR.n1405 VGND 0.53213f
C19308 VPWR.t444 VGND 0.97566f
C19309 VPWR.n1406 VGND 0.41384f
C19310 VPWR.n1407 VGND 0.29342f
C19311 VPWR.n1408 VGND 0.0191f
C19312 VPWR.n1409 VGND 0.03515f
C19313 VPWR.n1410 VGND 0.04254f
C19314 VPWR.n1411 VGND 0.01083f
C19315 VPWR.n1412 VGND 0.11537f
C19316 VPWR.n1413 VGND 0.32137f
C19317 VPWR.n1414 VGND 1.64092f
C19318 VPWR.t772 VGND 0.05456f
C19319 VPWR.t656 VGND 0.05456f
C19320 VPWR.n1415 VGND 0.09898f
C19321 VPWR.n1416 VGND 0.04687f
C19322 VPWR.n1417 VGND 0.00911f
C19323 VPWR.n1418 VGND 0.04687f
C19324 VPWR.t767 VGND 0.01433f
C19325 VPWR.t1258 VGND 0.01433f
C19326 VPWR.n1419 VGND 0.03131f
C19327 VPWR.t657 VGND 0.01433f
C19328 VPWR.t583 VGND 0.01433f
C19329 VPWR.n1420 VGND 0.03131f
C19330 VPWR.n1421 VGND 0.06379f
C19331 VPWR.t1871 VGND 0.05714f
C19332 VPWR.t932 VGND 0.05714f
C19333 VPWR.n1422 VGND 0.13169f
C19334 VPWR.n1423 VGND 0.02751f
C19335 VPWR.n1424 VGND 0.04687f
C19336 VPWR.n1425 VGND 0.01209f
C19337 VPWR.t1786 VGND 0.01433f
C19338 VPWR.t582 VGND 0.01433f
C19339 VPWR.n1426 VGND 0.03131f
C19340 VPWR.t586 VGND 0.01433f
C19341 VPWR.t441 VGND 0.01433f
C19342 VPWR.n1427 VGND 0.03131f
C19343 VPWR.n1428 VGND 0.07209f
C19344 VPWR.n1429 VGND 0.01209f
C19345 VPWR.n1430 VGND 0.04687f
C19346 VPWR.n1431 VGND 0.04687f
C19347 VPWR.n1432 VGND 0.04687f
C19348 VPWR.n1433 VGND 0.01128f
C19349 VPWR.t768 VGND 0.01433f
C19350 VPWR.t766 VGND 0.01433f
C19351 VPWR.n1434 VGND 0.03131f
C19352 VPWR.t660 VGND 0.01433f
C19353 VPWR.t659 VGND 0.01433f
C19354 VPWR.n1435 VGND 0.03131f
C19355 VPWR.n1436 VGND 0.06379f
C19356 VPWR.n1437 VGND 0.01055f
C19357 VPWR.n1438 VGND 0.00983f
C19358 VPWR.n1439 VGND 0.04687f
C19359 VPWR.n1440 VGND 0.03515f
C19360 VPWR.n1441 VGND 0.00794f
C19361 VPWR.t581 VGND 0.74843f
C19362 VPWR.n1442 VGND 0.4282f
C19363 VPWR.t440 VGND 0.74843f
C19364 VPWR.n1443 VGND 0.33553f
C19365 VPWR.n1444 VGND 0.28129f
C19366 VPWR.n1445 VGND 0.43003f
C19367 VPWR.n1446 VGND 6.17638f
C19368 VPWR.n1447 VGND 9.5664f
C19369 VPWR.n1448 VGND 0.08351f
C19370 VPWR.n1449 VGND 1.09982f
C19371 VPWR.n1450 VGND 1.0094f
C19372 VPWR.n1451 VGND 0.06482f
C19373 VPWR.n1452 VGND 0.0544f
C19374 VPWR.t2045 VGND 0.01136f
C19375 VPWR.t92 VGND 0.0124f
C19376 VPWR.n1453 VGND 0.02769f
C19377 VPWR.n1454 VGND 0.01897f
C19378 VPWR.n1455 VGND 0.06244f
C19379 VPWR.n1456 VGND 0.07762f
C19380 VPWR.n1457 VGND 0.09174f
C19381 VPWR.t1996 VGND 0.01136f
C19382 VPWR.t223 VGND 0.0124f
C19383 VPWR.n1458 VGND 0.02769f
C19384 VPWR.n1459 VGND 0.01897f
C19385 VPWR.n1460 VGND 0.06244f
C19386 VPWR.n1461 VGND 0.09746f
C19387 VPWR.n1462 VGND 0.09174f
C19388 VPWR.n1463 VGND 0.06567f
C19389 VPWR.n1464 VGND 0.0544f
C19390 VPWR.n1465 VGND 0.13913f
C19391 VPWR.n1466 VGND 0.01797f
C19392 VPWR.n1467 VGND 0.00728f
C19393 VPWR.n1468 VGND 0.10822f
C19394 VPWR.t269 VGND 0.11957f
C19395 VPWR.t224 VGND 0.07849f
C19396 VPWR.t837 VGND 0.09218f
C19397 VPWR.t2044 VGND 0.01116f
C19398 VPWR.t268 VGND 0.01222f
C19399 VPWR.n1469 VGND 0.03042f
C19400 VPWR.n1470 VGND 0.00581f
C19401 VPWR.t270 VGND 0.02679f
C19402 VPWR.n1471 VGND 0.05724f
C19403 VPWR.t838 VGND 0.02961f
C19404 VPWR.n1472 VGND 0.04692f
C19405 VPWR.n1473 VGND 0.01797f
C19406 VPWR.n1474 VGND 0.00728f
C19407 VPWR.n1475 VGND 0.10822f
C19408 VPWR.t371 VGND 0.11957f
C19409 VPWR.t353 VGND 0.07849f
C19410 VPWR.t1404 VGND 0.09218f
C19411 VPWR.t1994 VGND 0.01116f
C19412 VPWR.t370 VGND 0.01222f
C19413 VPWR.n1476 VGND 0.03042f
C19414 VPWR.n1477 VGND 0.00581f
C19415 VPWR.t372 VGND 0.02679f
C19416 VPWR.n1478 VGND 0.05724f
C19417 VPWR.t1405 VGND 0.02961f
C19418 VPWR.n1479 VGND 0.04692f
C19419 VPWR.n1480 VGND 0.00728f
C19420 VPWR.n1481 VGND 0.10822f
C19421 VPWR.t142 VGND 0.11957f
C19422 VPWR.t9 VGND 0.07849f
C19423 VPWR.t1640 VGND 0.09218f
C19424 VPWR.t1982 VGND 0.01116f
C19425 VPWR.t141 VGND 0.01222f
C19426 VPWR.n1482 VGND 0.03042f
C19427 VPWR.n1483 VGND 0.00581f
C19428 VPWR.t143 VGND 0.02679f
C19429 VPWR.n1484 VGND 0.05724f
C19430 VPWR.t1641 VGND 0.02961f
C19431 VPWR.n1485 VGND 0.04692f
C19432 VPWR.n1486 VGND 0.00805f
C19433 VPWR.n1487 VGND 0.08351f
C19434 VPWR.n1488 VGND -0.01866f
C19435 VPWR.n1489 VGND 0.13913f
C19436 VPWR.n1490 VGND 0.01797f
C19437 VPWR.n1491 VGND 0.00728f
C19438 VPWR.n1492 VGND 0.10822f
C19439 VPWR.t244 VGND 0.11957f
C19440 VPWR.t119 VGND 0.07849f
C19441 VPWR.t1223 VGND 0.09218f
C19442 VPWR.t274 VGND 0.07849f
C19443 VPWR.t266 VGND 0.11957f
C19444 VPWR.n1493 VGND 0.10822f
C19445 VPWR.n1494 VGND 0.00728f
C19446 VPWR.n1495 VGND 0.01797f
C19447 VPWR.n1496 VGND 0.0544f
C19448 VPWR.n1497 VGND 0.13913f
C19449 VPWR.n1498 VGND -0.01866f
C19450 VPWR.n1499 VGND 0.08351f
C19451 VPWR.n1500 VGND 0.08351f
C19452 VPWR.n1501 VGND -0.01866f
C19453 VPWR.n1502 VGND 0.0544f
C19454 VPWR.n1503 VGND 0.13913f
C19455 VPWR.n1504 VGND 0.01797f
C19456 VPWR.n1505 VGND 0.00728f
C19457 VPWR.n1506 VGND 0.10822f
C19458 VPWR.t17 VGND 0.11957f
C19459 VPWR.t276 VGND 0.07849f
C19460 VPWR.t1794 VGND 0.09218f
C19461 VPWR.t124 VGND 0.07849f
C19462 VPWR.t139 VGND 0.11957f
C19463 VPWR.n1507 VGND 0.10822f
C19464 VPWR.n1508 VGND 0.00728f
C19465 VPWR.n1509 VGND 0.01797f
C19466 VPWR.n1510 VGND 0.0544f
C19467 VPWR.n1511 VGND 0.13913f
C19468 VPWR.n1512 VGND -0.01866f
C19469 VPWR.n1513 VGND 0.08351f
C19470 VPWR.n1514 VGND 0.08351f
C19471 VPWR.n1515 VGND -0.01866f
C19472 VPWR.n1516 VGND 0.0544f
C19473 VPWR.n1517 VGND 0.13913f
C19474 VPWR.n1518 VGND 0.01797f
C19475 VPWR.n1519 VGND 0.00728f
C19476 VPWR.n1520 VGND 0.10822f
C19477 VPWR.t280 VGND 0.11957f
C19478 VPWR.t154 VGND 0.07849f
C19479 VPWR.t1483 VGND 0.09218f
C19480 VPWR.t272 VGND 0.07849f
C19481 VPWR.t296 VGND 0.11957f
C19482 VPWR.n1521 VGND 0.10822f
C19483 VPWR.n1522 VGND 0.00728f
C19484 VPWR.n1523 VGND 0.01797f
C19485 VPWR.n1524 VGND 0.0544f
C19486 VPWR.n1525 VGND 0.13913f
C19487 VPWR.n1526 VGND -0.01866f
C19488 VPWR.n1527 VGND 0.08351f
C19489 VPWR.n1528 VGND 0.08351f
C19490 VPWR.n1529 VGND 0.08351f
C19491 VPWR.n1530 VGND 0.08351f
C19492 VPWR.n1531 VGND -0.01866f
C19493 VPWR.n1532 VGND 0.13913f
C19494 VPWR.n1533 VGND 0.01797f
C19495 VPWR.n1534 VGND 0.00728f
C19496 VPWR.n1535 VGND 0.10822f
C19497 VPWR.t1106 VGND 0.09218f
C19498 VPWR.t23 VGND 0.07849f
C19499 VPWR.t36 VGND 0.11957f
C19500 VPWR.n1536 VGND 0.10822f
C19501 VPWR.n1537 VGND 0.00728f
C19502 VPWR.n1538 VGND 0.01797f
C19503 VPWR.n1539 VGND 0.13913f
C19504 VPWR.n1540 VGND 0.0544f
C19505 VPWR.n1541 VGND 0.06567f
C19506 VPWR.n1542 VGND 0.09174f
C19507 VPWR.t1929 VGND 0.01136f
C19508 VPWR.t22 VGND 0.0124f
C19509 VPWR.n1543 VGND 0.02769f
C19510 VPWR.n1544 VGND 0.01897f
C19511 VPWR.n1545 VGND 0.06244f
C19512 VPWR.n1546 VGND 0.09746f
C19513 VPWR.n1547 VGND 0.09174f
C19514 VPWR.t1986 VGND 0.01136f
C19515 VPWR.t271 VGND 0.0124f
C19516 VPWR.n1548 VGND 0.02769f
C19517 VPWR.n1549 VGND 0.01897f
C19518 VPWR.n1550 VGND 0.06244f
C19519 VPWR.n1551 VGND 0.09746f
C19520 VPWR.n1552 VGND 0.09174f
C19521 VPWR.t2025 VGND 0.01136f
C19522 VPWR.t153 VGND 0.0124f
C19523 VPWR.n1553 VGND 0.02769f
C19524 VPWR.n1554 VGND 0.01897f
C19525 VPWR.n1555 VGND 0.06244f
C19526 VPWR.n1556 VGND 0.09746f
C19527 VPWR.n1557 VGND 0.09174f
C19528 VPWR.t2037 VGND 0.01136f
C19529 VPWR.t123 VGND 0.0124f
C19530 VPWR.n1558 VGND 0.02769f
C19531 VPWR.n1559 VGND 0.01897f
C19532 VPWR.n1560 VGND 0.06244f
C19533 VPWR.n1561 VGND 0.09746f
C19534 VPWR.n1562 VGND 0.09174f
C19535 VPWR.t1979 VGND 0.01136f
C19536 VPWR.t275 VGND 0.0124f
C19537 VPWR.n1563 VGND 0.02769f
C19538 VPWR.n1564 VGND 0.01897f
C19539 VPWR.n1565 VGND 0.06244f
C19540 VPWR.n1566 VGND 0.09746f
C19541 VPWR.n1567 VGND 0.09174f
C19542 VPWR.t1985 VGND 0.01136f
C19543 VPWR.t273 VGND 0.0124f
C19544 VPWR.n1568 VGND 0.02769f
C19545 VPWR.n1569 VGND 0.01897f
C19546 VPWR.n1570 VGND 0.06244f
C19547 VPWR.n1571 VGND 0.09746f
C19548 VPWR.n1572 VGND 0.09174f
C19549 VPWR.t2039 VGND 0.01136f
C19550 VPWR.t118 VGND 0.0124f
C19551 VPWR.n1573 VGND 0.02769f
C19552 VPWR.n1574 VGND 0.01897f
C19553 VPWR.n1575 VGND 0.06244f
C19554 VPWR.n1576 VGND 0.09746f
C19555 VPWR.n1577 VGND 0.09174f
C19556 VPWR.t1936 VGND 0.01136f
C19557 VPWR.t8 VGND 0.0124f
C19558 VPWR.n1578 VGND 0.02769f
C19559 VPWR.n1579 VGND 0.01897f
C19560 VPWR.n1580 VGND 0.06244f
C19561 VPWR.n1581 VGND 0.09746f
C19562 VPWR.n1582 VGND 0.09174f
C19563 VPWR.n1583 VGND 0.06567f
C19564 VPWR.n1584 VGND 0.0544f
C19565 VPWR.n1585 VGND 0.13913f
C19566 VPWR.n1586 VGND -0.01866f
C19567 VPWR.n1587 VGND 0.08351f
C19568 VPWR.n1588 VGND 0.08351f
C19569 VPWR.n1589 VGND -0.01866f
C19570 VPWR.n1590 VGND 0.00805f
C19571 VPWR.n1591 VGND 0.01714f
C19572 VPWR.n1592 VGND 0.00725f
C19573 VPWR.n1593 VGND 0.10822f
C19574 VPWR.t166 VGND 0.09218f
C19575 VPWR.t44 VGND 0.07849f
C19576 VPWR.t80 VGND 0.11957f
C19577 VPWR.n1594 VGND 0.10822f
C19578 VPWR.n1595 VGND 0.00725f
C19579 VPWR.n1596 VGND 0.01714f
C19580 VPWR.n1597 VGND 0.03437f
C19581 VPWR.t1966 VGND 0.01116f
C19582 VPWR.t79 VGND 0.01222f
C19583 VPWR.n1598 VGND 0.03115f
C19584 VPWR.n1599 VGND 0.03694f
C19585 VPWR.n1600 VGND 0.00833f
C19586 VPWR.t2063 VGND 0.01136f
C19587 VPWR.t43 VGND 0.0124f
C19588 VPWR.n1601 VGND 0.02768f
C19589 VPWR.n1602 VGND 0.02818f
C19590 VPWR.n1603 VGND 0.01776f
C19591 VPWR.n1604 VGND 0.00697f
C19592 VPWR.n1605 VGND 0.01822f
C19593 VPWR.n1606 VGND 0.02384f
C19594 VPWR.n1607 VGND 0.23724f
C19595 VPWR.n1608 VGND 0.17585f
C19596 VPWR.n1609 VGND 0.02384f
C19597 VPWR.n1610 VGND 0.01776f
C19598 VPWR.t2010 VGND 0.0112f
C19599 VPWR.t178 VGND 0.01226f
C19600 VPWR.n1611 VGND 0.02993f
C19601 VPWR.n1612 VGND 0.03284f
C19602 VPWR.n1613 VGND 0.03437f
C19603 VPWR.t2047 VGND 0.01116f
C19604 VPWR.t346 VGND 0.01222f
C19605 VPWR.n1614 VGND 0.03115f
C19606 VPWR.n1615 VGND 0.03694f
C19607 VPWR.n1616 VGND 0.00833f
C19608 VPWR.t2000 VGND 0.01136f
C19609 VPWR.t212 VGND 0.0124f
C19610 VPWR.n1617 VGND 0.02768f
C19611 VPWR.n1618 VGND 0.02818f
C19612 VPWR.n1619 VGND 0.01822f
C19613 VPWR.n1620 VGND 0.02384f
C19614 VPWR.n1621 VGND 0.01776f
C19615 VPWR.t1955 VGND 0.0112f
C19616 VPWR.t338 VGND 0.01226f
C19617 VPWR.n1622 VGND 0.02993f
C19618 VPWR.n1623 VGND 0.03284f
C19619 VPWR.n1624 VGND 0.03437f
C19620 VPWR.t1965 VGND 0.01116f
C19621 VPWR.t64 VGND 0.01222f
C19622 VPWR.n1625 VGND 0.03115f
C19623 VPWR.n1626 VGND 0.03694f
C19624 VPWR.n1627 VGND 0.00833f
C19625 VPWR.t1962 VGND 0.01136f
C19626 VPWR.t320 VGND 0.0124f
C19627 VPWR.n1628 VGND 0.02768f
C19628 VPWR.n1629 VGND 0.02818f
C19629 VPWR.n1630 VGND 0.01776f
C19630 VPWR.n1631 VGND 0.00697f
C19631 VPWR.n1632 VGND 0.01822f
C19632 VPWR.n1633 VGND 0.02384f
C19633 VPWR.n1634 VGND 0.17585f
C19634 VPWR.n1635 VGND 0.17585f
C19635 VPWR.n1636 VGND 0.02384f
C19636 VPWR.n1637 VGND 0.01776f
C19637 VPWR.t2002 VGND 0.0112f
C19638 VPWR.t206 VGND 0.01226f
C19639 VPWR.n1638 VGND 0.02993f
C19640 VPWR.n1639 VGND 0.03284f
C19641 VPWR.n1640 VGND 0.03437f
C19642 VPWR.t1944 VGND 0.01116f
C19643 VPWR.t235 VGND 0.01222f
C19644 VPWR.n1641 VGND 0.03115f
C19645 VPWR.n1642 VGND 0.03694f
C19646 VPWR.n1643 VGND 0.00833f
C19647 VPWR.t2042 VGND 0.01136f
C19648 VPWR.t102 VGND 0.0124f
C19649 VPWR.n1644 VGND 0.02768f
C19650 VPWR.n1645 VGND 0.02818f
C19651 VPWR.n1646 VGND 0.01822f
C19652 VPWR.n1647 VGND 0.02384f
C19653 VPWR.n1648 VGND 0.01776f
C19654 VPWR.t1964 VGND 0.0112f
C19655 VPWR.t314 VGND 0.01226f
C19656 VPWR.n1649 VGND 0.02993f
C19657 VPWR.n1650 VGND 0.03284f
C19658 VPWR.n1651 VGND 0.03437f
C19659 VPWR.t2005 VGND 0.01116f
C19660 VPWR.t343 VGND 0.01222f
C19661 VPWR.n1652 VGND 0.03115f
C19662 VPWR.n1653 VGND 0.03694f
C19663 VPWR.n1654 VGND 0.00833f
C19664 VPWR.t1959 VGND 0.01136f
C19665 VPWR.t325 VGND 0.0124f
C19666 VPWR.n1655 VGND 0.02768f
C19667 VPWR.n1656 VGND 0.02818f
C19668 VPWR.n1657 VGND 0.01776f
C19669 VPWR.n1658 VGND 0.00697f
C19670 VPWR.n1659 VGND 0.01822f
C19671 VPWR.n1660 VGND 0.02384f
C19672 VPWR.n1661 VGND 0.17585f
C19673 VPWR.n1662 VGND 0.17585f
C19674 VPWR.n1663 VGND 0.02384f
C19675 VPWR.n1664 VGND 0.01776f
C19676 VPWR.t2043 VGND 0.0112f
C19677 VPWR.t99 VGND 0.01226f
C19678 VPWR.n1665 VGND 0.02993f
C19679 VPWR.n1666 VGND 0.03284f
C19680 VPWR.n1667 VGND 0.03437f
C19681 VPWR.t1941 VGND 0.01116f
C19682 VPWR.t130 VGND 0.01222f
C19683 VPWR.n1668 VGND 0.03115f
C19684 VPWR.n1669 VGND 0.03694f
C19685 VPWR.n1670 VGND 0.00833f
C19686 VPWR.t2050 VGND 0.01136f
C19687 VPWR.t85 VGND 0.0124f
C19688 VPWR.n1671 VGND 0.02768f
C19689 VPWR.n1672 VGND 0.02818f
C19690 VPWR.n1673 VGND 0.01822f
C19691 VPWR.n1674 VGND 0.02384f
C19692 VPWR.n1675 VGND 0.01776f
C19693 VPWR.t2003 VGND 0.0112f
C19694 VPWR.t203 VGND 0.01226f
C19695 VPWR.n1676 VGND 0.02993f
C19696 VPWR.n1677 VGND 0.03284f
C19697 VPWR.n1678 VGND 0.03437f
C19698 VPWR.t2038 VGND 0.01116f
C19699 VPWR.t257 VGND 0.01222f
C19700 VPWR.n1679 VGND 0.03115f
C19701 VPWR.n1680 VGND 0.03694f
C19702 VPWR.n1681 VGND 0.00833f
C19703 VPWR.t1993 VGND 0.01136f
C19704 VPWR.t238 VGND 0.0124f
C19705 VPWR.n1682 VGND 0.02768f
C19706 VPWR.n1683 VGND 0.02818f
C19707 VPWR.n1684 VGND 0.01776f
C19708 VPWR.n1685 VGND 0.00697f
C19709 VPWR.n1686 VGND 0.01822f
C19710 VPWR.n1687 VGND 0.02384f
C19711 VPWR.n1688 VGND 0.17585f
C19712 VPWR.n1689 VGND 0.17585f
C19713 VPWR.n1690 VGND 0.02384f
C19714 VPWR.n1691 VGND 0.01776f
C19715 VPWR.t1939 VGND 0.0112f
C19716 VPWR.t381 VGND 0.01226f
C19717 VPWR.n1692 VGND 0.02993f
C19718 VPWR.n1693 VGND 0.03284f
C19719 VPWR.n1694 VGND 0.03437f
C19720 VPWR.t1978 VGND 0.01116f
C19721 VPWR.t24 VGND 0.01222f
C19722 VPWR.n1695 VGND 0.03115f
C19723 VPWR.n1696 VGND 0.03694f
C19724 VPWR.n1697 VGND 0.00833f
C19725 VPWR.t2040 VGND 0.01136f
C19726 VPWR.t110 VGND 0.0124f
C19727 VPWR.n1698 VGND 0.02768f
C19728 VPWR.n1699 VGND 0.02818f
C19729 VPWR.n1700 VGND 0.01822f
C19730 VPWR.n1701 VGND 0.02384f
C19731 VPWR.n1702 VGND 0.01776f
C19732 VPWR.t2036 VGND 0.0112f
C19733 VPWR.t125 VGND 0.01226f
C19734 VPWR.n1703 VGND 0.02993f
C19735 VPWR.n1704 VGND 0.03284f
C19736 VPWR.n1705 VGND 0.03437f
C19737 VPWR.t1935 VGND 0.01116f
C19738 VPWR.t262 VGND 0.01222f
C19739 VPWR.n1706 VGND 0.03115f
C19740 VPWR.n1707 VGND 0.03694f
C19741 VPWR.n1708 VGND 0.00833f
C19742 VPWR.t2033 VGND 0.01136f
C19743 VPWR.t136 VGND 0.0124f
C19744 VPWR.n1709 VGND 0.02768f
C19745 VPWR.n1710 VGND 0.02818f
C19746 VPWR.n1711 VGND 0.01776f
C19747 VPWR.n1712 VGND 0.00697f
C19748 VPWR.n1713 VGND 0.01822f
C19749 VPWR.n1714 VGND 0.02384f
C19750 VPWR.n1715 VGND 0.17585f
C19751 VPWR.t1977 VGND 0.0112f
C19752 VPWR.t282 VGND 0.01226f
C19753 VPWR.n1716 VGND 0.02993f
C19754 VPWR.n1717 VGND 0.03284f
C19755 VPWR.t2024 VGND 0.01116f
C19756 VPWR.t290 VGND 0.01222f
C19757 VPWR.n1718 VGND 0.03115f
C19758 VPWR.n1719 VGND 0.03694f
C19759 VPWR.n1720 VGND 0.00833f
C19760 VPWR.t2019 VGND 0.01136f
C19761 VPWR.t161 VGND 0.0124f
C19762 VPWR.n1721 VGND 0.02768f
C19763 VPWR.n1722 VGND 0.02818f
C19764 VPWR.n1723 VGND 0.01776f
C19765 VPWR.n1724 VGND 0.00697f
C19766 VPWR.n1725 VGND 0.01822f
C19767 VPWR.n1726 VGND 0.02384f
C19768 VPWR.n1727 VGND 0.21163f
C19769 VPWR.n1728 VGND 0.02541f
C19770 VPWR.n1729 VGND 0.01776f
C19771 VPWR.t1937 VGND 0.01136f
C19772 VPWR.t6 VGND 0.0124f
C19773 VPWR.n1730 VGND 0.02768f
C19774 VPWR.n1731 VGND 0.02818f
C19775 VPWR.n1732 VGND 0.00833f
C19776 VPWR.t1984 VGND 0.01116f
C19777 VPWR.t10 VGND 0.01222f
C19778 VPWR.n1733 VGND 0.03115f
C19779 VPWR.n1734 VGND 0.03694f
C19780 VPWR.n1735 VGND 0.03437f
C19781 VPWR.n1736 VGND 0.00805f
C19782 VPWR.n1737 VGND 0.01714f
C19783 VPWR.n1738 VGND 0.00725f
C19784 VPWR.n1739 VGND 0.10822f
C19785 VPWR.t283 VGND 0.09218f
C19786 VPWR.t162 VGND 0.07849f
C19787 VPWR.t291 VGND 0.11957f
C19788 VPWR.n1740 VGND 0.10822f
C19789 VPWR.n1741 VGND 0.00725f
C19790 VPWR.n1742 VGND 0.01714f
C19791 VPWR.n1743 VGND 0.00805f
C19792 VPWR.n1744 VGND 0.0544f
C19793 VPWR.t2011 VGND 0.01116f
C19794 VPWR.t45 VGND 0.01222f
C19795 VPWR.n1745 VGND 0.03042f
C19796 VPWR.n1746 VGND 0.00581f
C19797 VPWR.t47 VGND 0.02679f
C19798 VPWR.n1747 VGND 0.05724f
C19799 VPWR.t863 VGND 0.02961f
C19800 VPWR.n1748 VGND 0.04692f
C19801 VPWR.t304 VGND 0.07849f
C19802 VPWR.t862 VGND 0.09218f
C19803 VPWR.t342 VGND 0.07849f
C19804 VPWR.t83 VGND 0.11957f
C19805 VPWR.n1749 VGND 0.10822f
C19806 VPWR.n1750 VGND 0.00728f
C19807 VPWR.n1751 VGND 0.01797f
C19808 VPWR.n1752 VGND 0.13913f
C19809 VPWR.n1753 VGND -0.01866f
C19810 VPWR.n1754 VGND 0.08351f
C19811 VPWR.n1755 VGND 0.08351f
C19812 VPWR.n1756 VGND -0.01866f
C19813 VPWR.n1757 VGND 0.13913f
C19814 VPWR.n1758 VGND 0.01797f
C19815 VPWR.n1759 VGND 0.00728f
C19816 VPWR.n1760 VGND 0.10822f
C19817 VPWR.t449 VGND 0.09218f
C19818 VPWR.t286 VGND 0.07849f
C19819 VPWR.t210 VGND 0.11957f
C19820 VPWR.n1761 VGND 0.10822f
C19821 VPWR.n1762 VGND 0.00728f
C19822 VPWR.n1763 VGND 0.01797f
C19823 VPWR.n1764 VGND 0.13913f
C19824 VPWR.n1765 VGND 0.0544f
C19825 VPWR.n1766 VGND 0.06567f
C19826 VPWR.n1767 VGND 0.09174f
C19827 VPWR.t1976 VGND 0.01136f
C19828 VPWR.t285 VGND 0.0124f
C19829 VPWR.n1768 VGND 0.02769f
C19830 VPWR.n1769 VGND 0.01897f
C19831 VPWR.n1770 VGND 0.06244f
C19832 VPWR.n1771 VGND 0.09746f
C19833 VPWR.n1772 VGND 0.09174f
C19834 VPWR.t1968 VGND 0.01136f
C19835 VPWR.t303 VGND 0.0124f
C19836 VPWR.n1773 VGND 0.02769f
C19837 VPWR.n1774 VGND 0.01897f
C19838 VPWR.n1775 VGND 0.06244f
C19839 VPWR.n1776 VGND 0.09746f
C19840 VPWR.t2013 VGND 0.01136f
C19841 VPWR.t173 VGND 0.0124f
C19842 VPWR.n1777 VGND 0.02769f
C19843 VPWR.n1778 VGND 0.01897f
C19844 VPWR.n1779 VGND 0.06242f
C19845 VPWR.n1780 VGND 0.05139f
C19846 VPWR.t1953 VGND 0.01136f
C19847 VPWR.t341 VGND 0.0124f
C19848 VPWR.n1781 VGND 0.02769f
C19849 VPWR.n1782 VGND 0.01897f
C19850 VPWR.n1783 VGND 0.06244f
C19851 VPWR.n1784 VGND 0.09746f
C19852 VPWR.n1785 VGND 0.09174f
C19853 VPWR.n1786 VGND 0.06567f
C19854 VPWR.n1787 VGND 0.0544f
C19855 VPWR.n1788 VGND 0.13913f
C19856 VPWR.n1789 VGND 0.01797f
C19857 VPWR.n1790 VGND 0.00728f
C19858 VPWR.n1791 VGND 0.10822f
C19859 VPWR.t191 VGND 0.11957f
C19860 VPWR.t174 VGND 0.07849f
C19861 VPWR.t299 VGND 0.13333f
C19862 VPWR.n1792 VGND 0.07618f
C19863 VPWR.n1793 VGND 0.01797f
C19864 VPWR.n1794 VGND 0.13913f
C19865 VPWR.n1795 VGND 0.1646f
C19866 VPWR.n1796 VGND 1.01577f
C19867 VPWR.n1797 VGND 0.08351f
C19868 VPWR.n1798 VGND 0.08351f
C19869 VPWR.n1799 VGND 0.08351f
C19870 VPWR.n1800 VGND 0.08351f
C19871 VPWR.n1801 VGND 0.08351f
C19872 VPWR.n1802 VGND 0.08351f
C19873 VPWR.n1803 VGND 0.08351f
C19874 VPWR.n1804 VGND 0.08351f
C19875 VPWR.n1805 VGND 0.08351f
C19876 VPWR.n1806 VGND 0.08351f
C19877 VPWR.n1807 VGND 0.08351f
C19878 VPWR.n1808 VGND 0.08351f
C19879 VPWR.n1809 VGND 0.08351f
C19880 VPWR.n1810 VGND 0.08351f
C19881 VPWR.n1811 VGND 0.08351f
C19882 VPWR.n1812 VGND 0.19371f
C19883 VPWR.n1813 VGND 1.01577f
C19884 VPWR.n1814 VGND 1.01577f
C19885 VPWR.n1815 VGND 0.19371f
C19886 VPWR.n1816 VGND 0.13913f
C19887 VPWR.n1817 VGND 0.01797f
C19888 VPWR.n1818 VGND 0.07618f
C19889 VPWR.t336 VGND 0.13333f
C19890 VPWR.t435 VGND 0.07849f
C19891 VPWR.t626 VGND 0.11957f
C19892 VPWR.n1819 VGND 0.10822f
C19893 VPWR.n1820 VGND 0.00728f
C19894 VPWR.n1821 VGND 0.01797f
C19895 VPWR.n1822 VGND 0.13913f
C19896 VPWR.n1823 VGND 0.08351f
C19897 VPWR.n1824 VGND 0.08351f
C19898 VPWR.n1825 VGND 0.13913f
C19899 VPWR.n1826 VGND 0.01797f
C19900 VPWR.n1827 VGND 0.00728f
C19901 VPWR.n1828 VGND 0.10822f
C19902 VPWR.t486 VGND 0.09218f
C19903 VPWR.t1455 VGND 0.07849f
C19904 VPWR.t821 VGND 0.11957f
C19905 VPWR.n1829 VGND 0.10822f
C19906 VPWR.n1830 VGND 0.00728f
C19907 VPWR.n1831 VGND 0.01797f
C19908 VPWR.n1832 VGND 0.13913f
C19909 VPWR.n1833 VGND 0.08351f
C19910 VPWR.n1834 VGND 0.08351f
C19911 VPWR.n1835 VGND 0.13913f
C19912 VPWR.n1836 VGND 0.01797f
C19913 VPWR.n1837 VGND 0.00728f
C19914 VPWR.n1838 VGND 0.10822f
C19915 VPWR.t1457 VGND 0.09218f
C19916 VPWR.t1488 VGND 0.07849f
C19917 VPWR.t1051 VGND 0.11957f
C19918 VPWR.n1839 VGND 0.10822f
C19919 VPWR.n1840 VGND 0.00728f
C19920 VPWR.n1841 VGND 0.01797f
C19921 VPWR.n1842 VGND 0.13913f
C19922 VPWR.n1843 VGND 0.08351f
C19923 VPWR.n1844 VGND 0.08351f
C19924 VPWR.n1845 VGND 0.13913f
C19925 VPWR.n1846 VGND 0.01797f
C19926 VPWR.n1847 VGND 0.00728f
C19927 VPWR.n1848 VGND 0.10822f
C19928 VPWR.t648 VGND 0.09218f
C19929 VPWR.t433 VGND 0.07849f
C19930 VPWR.t1914 VGND 0.11957f
C19931 VPWR.n1849 VGND 0.10822f
C19932 VPWR.n1850 VGND 0.00728f
C19933 VPWR.n1851 VGND 0.01797f
C19934 VPWR.n1852 VGND 0.13913f
C19935 VPWR.n1853 VGND 0.08351f
C19936 VPWR.n1854 VGND 0.08351f
C19937 VPWR.n1855 VGND 0.13913f
C19938 VPWR.n1856 VGND 0.01797f
C19939 VPWR.n1857 VGND 0.00728f
C19940 VPWR.n1858 VGND 0.10822f
C19941 VPWR.t907 VGND 0.09218f
C19942 VPWR.t1485 VGND 0.07849f
C19943 VPWR.t722 VGND 0.11957f
C19944 VPWR.n1859 VGND 0.10822f
C19945 VPWR.n1860 VGND 0.00728f
C19946 VPWR.n1861 VGND 0.01797f
C19947 VPWR.n1862 VGND 0.13913f
C19948 VPWR.n1863 VGND 0.08351f
C19949 VPWR.n1864 VGND 0.08351f
C19950 VPWR.n1865 VGND 0.13913f
C19951 VPWR.n1866 VGND 0.01797f
C19952 VPWR.n1867 VGND 0.00728f
C19953 VPWR.n1868 VGND 0.10822f
C19954 VPWR.t547 VGND 0.09218f
C19955 VPWR.t432 VGND 0.07849f
C19956 VPWR.t1717 VGND 0.11957f
C19957 VPWR.n1869 VGND 0.10822f
C19958 VPWR.n1870 VGND 0.00728f
C19959 VPWR.n1871 VGND 0.01797f
C19960 VPWR.n1872 VGND 0.13913f
C19961 VPWR.n1873 VGND 0.08351f
C19962 VPWR.n1874 VGND 0.08351f
C19963 VPWR.n1875 VGND 0.13913f
C19964 VPWR.n1876 VGND 0.01797f
C19965 VPWR.n1877 VGND 0.00728f
C19966 VPWR.n1878 VGND 0.10822f
C19967 VPWR.t1630 VGND 0.09218f
C19968 VPWR.t1490 VGND 0.07849f
C19969 VPWR.t1376 VGND 0.11957f
C19970 VPWR.n1879 VGND 0.10822f
C19971 VPWR.n1880 VGND 0.00728f
C19972 VPWR.n1881 VGND 0.01797f
C19973 VPWR.n1882 VGND 0.13913f
C19974 VPWR.n1883 VGND 0.08351f
C19975 VPWR.n1884 VGND 0.08351f
C19976 VPWR.n1885 VGND 0.13913f
C19977 VPWR.n1886 VGND 0.01797f
C19978 VPWR.n1887 VGND 0.00728f
C19979 VPWR.n1888 VGND 0.10822f
C19980 VPWR.t1613 VGND 0.09218f
C19981 VPWR.t434 VGND 0.07849f
C19982 VPWR.t1739 VGND 0.11957f
C19983 VPWR.n1889 VGND 0.10822f
C19984 VPWR.n1890 VGND 0.00728f
C19985 VPWR.n1891 VGND 0.01797f
C19986 VPWR.n1892 VGND 0.13913f
C19987 VPWR.n1893 VGND 0.08351f
C19988 VPWR.n1894 VGND 1.0094f
C19989 VPWR.n1895 VGND 0.19371f
C19990 VPWR.n1896 VGND 0.08351f
C19991 VPWR.n1897 VGND 0.08351f
C19992 VPWR.n1898 VGND 0.08351f
C19993 VPWR.n1899 VGND 0.08351f
C19994 VPWR.n1900 VGND 0.08351f
C19995 VPWR.n1901 VGND 0.08351f
C19996 VPWR.n1902 VGND 0.08351f
C19997 VPWR.n1903 VGND 0.08351f
C19998 VPWR.n1904 VGND 0.08351f
C19999 VPWR.n1905 VGND 0.08351f
C20000 VPWR.n1906 VGND 0.08351f
C20001 VPWR.n1907 VGND 0.08351f
C20002 VPWR.n1908 VGND 0.08351f
C20003 VPWR.n1909 VGND 0.08351f
C20004 VPWR.n1910 VGND 0.08351f
C20005 VPWR.n1911 VGND 1.0094f
C20006 VPWR.n1912 VGND 1.0094f
C20007 VPWR.n1913 VGND 0.08351f
C20008 VPWR.n1914 VGND 0.13913f
C20009 VPWR.n1915 VGND 0.01797f
C20010 VPWR.n1916 VGND 0.00728f
C20011 VPWR.n1917 VGND 0.10822f
C20012 VPWR.t1726 VGND 0.11957f
C20013 VPWR.t852 VGND 0.07849f
C20014 VPWR.t1591 VGND 0.09218f
C20015 VPWR.t1836 VGND 0.07849f
C20016 VPWR.t1585 VGND 0.11957f
C20017 VPWR.n1918 VGND 0.10822f
C20018 VPWR.n1919 VGND 0.00728f
C20019 VPWR.n1920 VGND 0.01797f
C20020 VPWR.n1921 VGND 0.13913f
C20021 VPWR.n1922 VGND 0.08351f
C20022 VPWR.n1923 VGND 0.08351f
C20023 VPWR.n1924 VGND 0.13913f
C20024 VPWR.n1925 VGND 0.01797f
C20025 VPWR.n1926 VGND 0.00728f
C20026 VPWR.n1927 VGND 0.10822f
C20027 VPWR.t1392 VGND 0.11957f
C20028 VPWR.t1849 VGND 0.07849f
C20029 VPWR.t1069 VGND 0.09218f
C20030 VPWR.t1845 VGND 0.07849f
C20031 VPWR.t1851 VGND 0.11957f
C20032 VPWR.n1928 VGND 0.10822f
C20033 VPWR.n1929 VGND 0.00728f
C20034 VPWR.n1930 VGND 0.01797f
C20035 VPWR.n1931 VGND 0.13913f
C20036 VPWR.n1932 VGND 0.08351f
C20037 VPWR.n1933 VGND 0.08351f
C20038 VPWR.n1934 VGND 0.13913f
C20039 VPWR.n1935 VGND 0.01797f
C20040 VPWR.n1936 VGND 0.00728f
C20041 VPWR.n1937 VGND 0.10822f
C20042 VPWR.t1534 VGND 0.11957f
C20043 VPWR.t1841 VGND 0.07849f
C20044 VPWR.t704 VGND 0.09218f
C20045 VPWR.t1840 VGND 0.07849f
C20046 VPWR.t593 VGND 0.11957f
C20047 VPWR.n1938 VGND 0.10822f
C20048 VPWR.n1939 VGND 0.00728f
C20049 VPWR.n1940 VGND 0.01797f
C20050 VPWR.n1941 VGND 0.13913f
C20051 VPWR.n1942 VGND 0.08351f
C20052 VPWR.n1943 VGND 0.08351f
C20053 VPWR.n1944 VGND 0.13913f
C20054 VPWR.n1945 VGND 0.01797f
C20055 VPWR.n1946 VGND 0.00728f
C20056 VPWR.n1947 VGND 0.10822f
C20057 VPWR.t1900 VGND 0.11957f
C20058 VPWR.t1844 VGND 0.07849f
C20059 VPWR.t384 VGND 0.09218f
C20060 VPWR.t1843 VGND 0.07849f
C20061 VPWR.t864 VGND 0.11957f
C20062 VPWR.n1948 VGND 0.10822f
C20063 VPWR.n1949 VGND 0.00728f
C20064 VPWR.n1950 VGND 0.01797f
C20065 VPWR.n1951 VGND 0.13913f
C20066 VPWR.n1952 VGND 0.08351f
C20067 VPWR.n1953 VGND 0.08351f
C20068 VPWR.n1954 VGND 0.13913f
C20069 VPWR.n1955 VGND 0.01797f
C20070 VPWR.n1956 VGND 0.00728f
C20071 VPWR.n1957 VGND 0.10822f
C20072 VPWR.t1601 VGND 0.11957f
C20073 VPWR.t1842 VGND 0.07849f
C20074 VPWR.t1828 VGND 0.09218f
C20075 VPWR.t1848 VGND 0.07849f
C20076 VPWR.t1822 VGND 0.11957f
C20077 VPWR.n1958 VGND 0.10822f
C20078 VPWR.n1959 VGND 0.00728f
C20079 VPWR.n1960 VGND 0.01797f
C20080 VPWR.n1961 VGND 0.13913f
C20081 VPWR.n1962 VGND 0.08351f
C20082 VPWR.n1963 VGND 0.08351f
C20083 VPWR.n1964 VGND 0.13913f
C20084 VPWR.n1965 VGND 0.01797f
C20085 VPWR.n1966 VGND 0.00728f
C20086 VPWR.n1967 VGND 0.10822f
C20087 VPWR.t1471 VGND 0.11957f
C20088 VPWR.t1847 VGND 0.07849f
C20089 VPWR.t1243 VGND 0.09218f
C20090 VPWR.t1839 VGND 0.07849f
C20091 VPWR.t1207 VGND 0.11957f
C20092 VPWR.n1968 VGND 0.10822f
C20093 VPWR.n1969 VGND 0.00728f
C20094 VPWR.n1970 VGND 0.01797f
C20095 VPWR.n1971 VGND 0.13913f
C20096 VPWR.n1972 VGND 0.08351f
C20097 VPWR.n1973 VGND 0.08351f
C20098 VPWR.n1974 VGND 0.13913f
C20099 VPWR.n1975 VGND 0.01797f
C20100 VPWR.n1976 VGND 0.00728f
C20101 VPWR.n1977 VGND 0.10822f
C20102 VPWR.t807 VGND 0.11957f
C20103 VPWR.t1838 VGND 0.07849f
C20104 VPWR.t511 VGND 0.09218f
C20105 VPWR.t1837 VGND 0.07849f
C20106 VPWR.t999 VGND 0.11957f
C20107 VPWR.n1978 VGND 0.10822f
C20108 VPWR.n1979 VGND 0.00728f
C20109 VPWR.n1980 VGND 0.01797f
C20110 VPWR.n1981 VGND 0.13913f
C20111 VPWR.n1982 VGND 0.08351f
C20112 VPWR.n1983 VGND 0.08351f
C20113 VPWR.n1984 VGND 0.13913f
C20114 VPWR.n1985 VGND 0.01797f
C20115 VPWR.n1986 VGND 0.00728f
C20116 VPWR.n1987 VGND 0.10822f
C20117 VPWR.t1810 VGND 0.11957f
C20118 VPWR.t853 VGND 0.07849f
C20119 VPWR.t41 VGND 0.13333f
C20120 VPWR.n1988 VGND 0.07618f
C20121 VPWR.n1989 VGND 0.01797f
C20122 VPWR.n1990 VGND 0.13913f
C20123 VPWR.n1991 VGND 0.19371f
C20124 VPWR.n1992 VGND 1.01577f
C20125 VPWR.n1993 VGND 0.08351f
C20126 VPWR.n1994 VGND 0.08351f
C20127 VPWR.n1995 VGND 0.08351f
C20128 VPWR.n1996 VGND 0.08351f
C20129 VPWR.n1997 VGND 0.08351f
C20130 VPWR.n1998 VGND 0.08351f
C20131 VPWR.n1999 VGND 0.08351f
C20132 VPWR.n2000 VGND 0.08351f
C20133 VPWR.n2001 VGND 0.08351f
C20134 VPWR.n2002 VGND 0.08351f
C20135 VPWR.n2003 VGND 0.08351f
C20136 VPWR.n2004 VGND 0.08351f
C20137 VPWR.n2005 VGND 0.08351f
C20138 VPWR.n2006 VGND 0.08351f
C20139 VPWR.n2007 VGND 0.08351f
C20140 VPWR.n2008 VGND 0.19371f
C20141 VPWR.n2009 VGND 1.01577f
C20142 VPWR.n2010 VGND 1.01577f
C20143 VPWR.n2011 VGND 0.19371f
C20144 VPWR.n2012 VGND 0.13913f
C20145 VPWR.n2013 VGND 0.01797f
C20146 VPWR.n2014 VGND 0.07618f
C20147 VPWR.t116 VGND 0.13333f
C20148 VPWR.t785 VGND 0.07849f
C20149 VPWR.t696 VGND 0.11957f
C20150 VPWR.n2015 VGND 0.10822f
C20151 VPWR.n2016 VGND 0.00728f
C20152 VPWR.n2017 VGND 0.01797f
C20153 VPWR.n2018 VGND 0.13913f
C20154 VPWR.n2019 VGND 0.08351f
C20155 VPWR.n2020 VGND 0.08351f
C20156 VPWR.n2021 VGND 0.13913f
C20157 VPWR.n2022 VGND 0.01797f
C20158 VPWR.n2023 VGND 0.00728f
C20159 VPWR.n2024 VGND 0.10822f
C20160 VPWR.t1619 VGND 0.09218f
C20161 VPWR.t1073 VGND 0.07849f
C20162 VPWR.t455 VGND 0.11957f
C20163 VPWR.n2025 VGND 0.10822f
C20164 VPWR.n2026 VGND 0.00728f
C20165 VPWR.n2027 VGND 0.01797f
C20166 VPWR.n2028 VGND 0.13913f
C20167 VPWR.n2029 VGND 0.08351f
C20168 VPWR.n2030 VGND 0.08351f
C20169 VPWR.n2031 VGND 0.13913f
C20170 VPWR.n2032 VGND 0.01797f
C20171 VPWR.n2033 VGND 0.00728f
C20172 VPWR.n2034 VGND 0.10822f
C20173 VPWR.t1203 VGND 0.09218f
C20174 VPWR.t790 VGND 0.07849f
C20175 VPWR.t549 VGND 0.11957f
C20176 VPWR.n2035 VGND 0.10822f
C20177 VPWR.n2036 VGND 0.00728f
C20178 VPWR.n2037 VGND 0.01797f
C20179 VPWR.n2038 VGND 0.13913f
C20180 VPWR.n2039 VGND 0.08351f
C20181 VPWR.n2040 VGND 0.08351f
C20182 VPWR.n2041 VGND 0.13913f
C20183 VPWR.n2042 VGND 0.01797f
C20184 VPWR.n2043 VGND 0.00728f
C20185 VPWR.n2044 VGND 0.10822f
C20186 VPWR.t674 VGND 0.09218f
C20187 VPWR.t1077 VGND 0.07849f
C20188 VPWR.t1118 VGND 0.11957f
C20189 VPWR.n2045 VGND 0.10822f
C20190 VPWR.n2046 VGND 0.00728f
C20191 VPWR.n2047 VGND 0.01797f
C20192 VPWR.n2048 VGND 0.13913f
C20193 VPWR.n2049 VGND 0.08351f
C20194 VPWR.n2050 VGND 0.08351f
C20195 VPWR.n2051 VGND 0.13913f
C20196 VPWR.n2052 VGND 0.01797f
C20197 VPWR.n2053 VGND 0.00728f
C20198 VPWR.n2054 VGND 0.10822f
C20199 VPWR.t1110 VGND 0.09218f
C20200 VPWR.t787 VGND 0.07849f
C20201 VPWR.t1894 VGND 0.11957f
C20202 VPWR.n2055 VGND 0.10822f
C20203 VPWR.n2056 VGND 0.00728f
C20204 VPWR.n2057 VGND 0.01797f
C20205 VPWR.n2058 VGND 0.13913f
C20206 VPWR.n2059 VGND 0.08351f
C20207 VPWR.n2060 VGND 0.08351f
C20208 VPWR.n2061 VGND 0.13913f
C20209 VPWR.n2062 VGND 0.01797f
C20210 VPWR.n2063 VGND 0.00728f
C20211 VPWR.n2064 VGND 0.10822f
C20212 VPWR.t589 VGND 0.09218f
C20213 VPWR.t1076 VGND 0.07849f
C20214 VPWR.t1573 VGND 0.11957f
C20215 VPWR.n2065 VGND 0.10822f
C20216 VPWR.n2066 VGND 0.00728f
C20217 VPWR.n2067 VGND 0.01797f
C20218 VPWR.n2068 VGND 0.13913f
C20219 VPWR.n2069 VGND 0.08351f
C20220 VPWR.n2070 VGND 0.08351f
C20221 VPWR.n2071 VGND 0.13913f
C20222 VPWR.n2072 VGND 0.01797f
C20223 VPWR.n2073 VGND 0.00728f
C20224 VPWR.n2074 VGND 0.10822f
C20225 VPWR.t1859 VGND 0.09218f
C20226 VPWR.t792 VGND 0.07849f
C20227 VPWR.t1402 VGND 0.11957f
C20228 VPWR.n2075 VGND 0.10822f
C20229 VPWR.n2076 VGND 0.00728f
C20230 VPWR.n2077 VGND 0.01797f
C20231 VPWR.n2078 VGND 0.13913f
C20232 VPWR.n2079 VGND 0.08351f
C20233 VPWR.n2080 VGND 0.08351f
C20234 VPWR.n2081 VGND 0.13913f
C20235 VPWR.n2082 VGND 0.01797f
C20236 VPWR.n2083 VGND 0.00728f
C20237 VPWR.n2084 VGND 0.10822f
C20238 VPWR.t1523 VGND 0.09218f
C20239 VPWR.t1078 VGND 0.07849f
C20240 VPWR.t829 VGND 0.11957f
C20241 VPWR.n2085 VGND 0.10822f
C20242 VPWR.n2086 VGND 0.00728f
C20243 VPWR.n2087 VGND 0.01797f
C20244 VPWR.n2088 VGND 0.13913f
C20245 VPWR.n2089 VGND 0.08351f
C20246 VPWR.n2090 VGND 1.0094f
C20247 VPWR.n2091 VGND 0.19371f
C20248 VPWR.n2092 VGND 0.08351f
C20249 VPWR.n2093 VGND 0.08351f
C20250 VPWR.n2094 VGND 0.08351f
C20251 VPWR.n2095 VGND 0.08351f
C20252 VPWR.n2096 VGND 0.08351f
C20253 VPWR.n2097 VGND 0.08351f
C20254 VPWR.n2098 VGND 0.08351f
C20255 VPWR.n2099 VGND 0.08351f
C20256 VPWR.n2100 VGND 0.08351f
C20257 VPWR.n2101 VGND 0.08351f
C20258 VPWR.n2102 VGND 0.08351f
C20259 VPWR.n2103 VGND 0.08351f
C20260 VPWR.n2104 VGND 0.08351f
C20261 VPWR.n2105 VGND 0.08351f
C20262 VPWR.n2106 VGND 0.08351f
C20263 VPWR.n2107 VGND 1.0094f
C20264 VPWR.n2108 VGND 1.0094f
C20265 VPWR.n2109 VGND 0.08351f
C20266 VPWR.n2110 VGND 0.13913f
C20267 VPWR.n2111 VGND 0.01797f
C20268 VPWR.n2112 VGND 0.00728f
C20269 VPWR.n2113 VGND 0.10822f
C20270 VPWR.t1724 VGND 0.11957f
C20271 VPWR.t921 VGND 0.07849f
C20272 VPWR.t1589 VGND 0.09218f
C20273 VPWR.t496 VGND 0.07849f
C20274 VPWR.t1583 VGND 0.11957f
C20275 VPWR.n2114 VGND 0.10822f
C20276 VPWR.n2115 VGND 0.00728f
C20277 VPWR.n2116 VGND 0.01797f
C20278 VPWR.n2117 VGND 0.13913f
C20279 VPWR.n2118 VGND 0.08351f
C20280 VPWR.n2119 VGND 0.08351f
C20281 VPWR.n2120 VGND 0.13913f
C20282 VPWR.n2121 VGND 0.01797f
C20283 VPWR.n2122 VGND 0.00728f
C20284 VPWR.n2123 VGND 0.10822f
C20285 VPWR.t1394 VGND 0.11957f
C20286 VPWR.t495 VGND 0.07849f
C20287 VPWR.t1065 VGND 0.09218f
C20288 VPWR.t1505 VGND 0.07849f
C20289 VPWR.t802 VGND 0.11957f
C20290 VPWR.n2124 VGND 0.10822f
C20291 VPWR.n2125 VGND 0.00728f
C20292 VPWR.n2126 VGND 0.01797f
C20293 VPWR.n2127 VGND 0.13913f
C20294 VPWR.n2128 VGND 0.08351f
C20295 VPWR.n2129 VGND 0.08351f
C20296 VPWR.n2130 VGND 0.13913f
C20297 VPWR.n2131 VGND 0.01797f
C20298 VPWR.n2132 VGND 0.00728f
C20299 VPWR.n2133 VGND 0.10822f
C20300 VPWR.t1666 VGND 0.11957f
C20301 VPWR.t1565 VGND 0.07849f
C20302 VPWR.t702 VGND 0.09218f
C20303 VPWR.t1005 VGND 0.07849f
C20304 VPWR.t591 VGND 0.11957f
C20305 VPWR.n2134 VGND 0.10822f
C20306 VPWR.n2135 VGND 0.00728f
C20307 VPWR.n2136 VGND 0.01797f
C20308 VPWR.n2137 VGND 0.13913f
C20309 VPWR.n2138 VGND 0.08351f
C20310 VPWR.n2139 VGND 0.08351f
C20311 VPWR.n2140 VGND 0.13913f
C20312 VPWR.n2141 VGND 0.01797f
C20313 VPWR.n2142 VGND 0.00728f
C20314 VPWR.n2143 VGND 0.10822f
C20315 VPWR.t1898 VGND 0.11957f
C20316 VPWR.t826 VGND 0.07849f
C20317 VPWR.t1022 VGND 0.09218f
C20318 VPWR.t825 VGND 0.07849f
C20319 VPWR.t577 VGND 0.11957f
C20320 VPWR.n2144 VGND 0.10822f
C20321 VPWR.n2145 VGND 0.00728f
C20322 VPWR.n2146 VGND 0.01797f
C20323 VPWR.n2147 VGND 0.13913f
C20324 VPWR.n2148 VGND 0.08351f
C20325 VPWR.n2149 VGND 0.08351f
C20326 VPWR.n2150 VGND 0.13913f
C20327 VPWR.n2151 VGND 0.01797f
C20328 VPWR.n2152 VGND 0.00728f
C20329 VPWR.n2153 VGND 0.10822f
C20330 VPWR.t1599 VGND 0.11957f
C20331 VPWR.t1566 VGND 0.07849f
C20332 VPWR.t1826 VGND 0.09218f
C20333 VPWR.t1508 VGND 0.07849f
C20334 VPWR.t1820 VGND 0.11957f
C20335 VPWR.n2154 VGND 0.10822f
C20336 VPWR.n2155 VGND 0.00728f
C20337 VPWR.n2156 VGND 0.01797f
C20338 VPWR.n2157 VGND 0.13913f
C20339 VPWR.n2158 VGND 0.08351f
C20340 VPWR.n2159 VGND 0.08351f
C20341 VPWR.n2160 VGND 0.13913f
C20342 VPWR.n2161 VGND 0.01797f
C20343 VPWR.n2162 VGND 0.00728f
C20344 VPWR.n2163 VGND 0.10822f
C20345 VPWR.t553 VGND 0.11957f
C20346 VPWR.t1507 VGND 0.07849f
C20347 VPWR.t1241 VGND 0.09218f
C20348 VPWR.t1004 VGND 0.07849f
C20349 VPWR.t1205 VGND 0.11957f
C20350 VPWR.n2164 VGND 0.10822f
C20351 VPWR.n2165 VGND 0.00728f
C20352 VPWR.n2166 VGND 0.01797f
C20353 VPWR.n2167 VGND 0.13913f
C20354 VPWR.n2168 VGND 0.08351f
C20355 VPWR.n2169 VGND 0.08351f
C20356 VPWR.n2170 VGND 0.13913f
C20357 VPWR.n2171 VGND 0.01797f
C20358 VPWR.n2172 VGND 0.00728f
C20359 VPWR.n2173 VGND 0.10822f
C20360 VPWR.t805 VGND 0.11957f
C20361 VPWR.t1003 VGND 0.07849f
C20362 VPWR.t509 VGND 0.09218f
C20363 VPWR.t497 VGND 0.07849f
C20364 VPWR.t997 VGND 0.11957f
C20365 VPWR.n2174 VGND 0.10822f
C20366 VPWR.n2175 VGND 0.00728f
C20367 VPWR.n2176 VGND 0.01797f
C20368 VPWR.n2177 VGND 0.13913f
C20369 VPWR.n2178 VGND 0.08351f
C20370 VPWR.n2179 VGND 0.08351f
C20371 VPWR.n2180 VGND 0.13913f
C20372 VPWR.n2181 VGND 0.01797f
C20373 VPWR.n2182 VGND 0.00728f
C20374 VPWR.n2183 VGND 0.10822f
C20375 VPWR.t1808 VGND 0.11957f
C20376 VPWR.t824 VGND 0.07849f
C20377 VPWR.t49 VGND 0.13333f
C20378 VPWR.n2184 VGND 0.07618f
C20379 VPWR.n2185 VGND 0.01797f
C20380 VPWR.n2186 VGND 0.13913f
C20381 VPWR.n2187 VGND 0.19371f
C20382 VPWR.n2188 VGND 1.01577f
C20383 VPWR.n2189 VGND 0.08351f
C20384 VPWR.n2190 VGND 0.08351f
C20385 VPWR.n2191 VGND 0.08351f
C20386 VPWR.n2192 VGND 0.08351f
C20387 VPWR.n2193 VGND 0.08351f
C20388 VPWR.n2194 VGND 0.08351f
C20389 VPWR.n2195 VGND 0.08351f
C20390 VPWR.n2196 VGND 0.08351f
C20391 VPWR.n2197 VGND 0.08351f
C20392 VPWR.n2198 VGND 0.08351f
C20393 VPWR.n2199 VGND 0.08351f
C20394 VPWR.n2200 VGND 0.08351f
C20395 VPWR.n2201 VGND 0.08351f
C20396 VPWR.n2202 VGND 0.08351f
C20397 VPWR.n2203 VGND 0.08351f
C20398 VPWR.n2204 VGND 0.19371f
C20399 VPWR.n2205 VGND 1.01577f
C20400 VPWR.n2206 VGND 1.01577f
C20401 VPWR.n2207 VGND 0.19371f
C20402 VPWR.n2208 VGND 0.13913f
C20403 VPWR.n2209 VGND 0.01797f
C20404 VPWR.n2210 VGND 0.07618f
C20405 VPWR.t215 VGND 0.13333f
C20406 VPWR.t1222 VGND 0.07849f
C20407 VPWR.t756 VGND 0.11957f
C20408 VPWR.n2211 VGND 0.10822f
C20409 VPWR.n2212 VGND 0.00728f
C20410 VPWR.n2213 VGND 0.01797f
C20411 VPWR.n2214 VGND 0.13913f
C20412 VPWR.n2215 VGND 0.08351f
C20413 VPWR.n2216 VGND 0.08351f
C20414 VPWR.n2217 VGND 0.13913f
C20415 VPWR.n2218 VGND 0.01797f
C20416 VPWR.n2219 VGND 0.00728f
C20417 VPWR.n2220 VGND 0.10822f
C20418 VPWR.t1782 VGND 0.09218f
C20419 VPWR.t1216 VGND 0.07849f
C20420 VPWR.t1700 VGND 0.11957f
C20421 VPWR.n2221 VGND 0.10822f
C20422 VPWR.n2222 VGND 0.00728f
C20423 VPWR.n2223 VGND 0.01797f
C20424 VPWR.n2224 VGND 0.13913f
C20425 VPWR.n2225 VGND 0.08351f
C20426 VPWR.n2226 VGND 0.08351f
C20427 VPWR.n2227 VGND 0.13913f
C20428 VPWR.n2228 VGND 0.01797f
C20429 VPWR.n2229 VGND 0.00728f
C20430 VPWR.n2230 VGND 0.10822f
C20431 VPWR.t467 VGND 0.09218f
C20432 VPWR.t427 VGND 0.07849f
C20433 VPWR.t1680 VGND 0.11957f
C20434 VPWR.n2231 VGND 0.10822f
C20435 VPWR.n2232 VGND 0.00728f
C20436 VPWR.n2233 VGND 0.01797f
C20437 VPWR.n2234 VGND 0.13913f
C20438 VPWR.n2235 VGND 0.08351f
C20439 VPWR.n2236 VGND 0.08351f
C20440 VPWR.n2237 VGND 0.13913f
C20441 VPWR.n2238 VGND 0.01797f
C20442 VPWR.n2239 VGND 0.00728f
C20443 VPWR.n2240 VGND 0.10822f
C20444 VPWR.t620 VGND 0.09218f
C20445 VPWR.t1220 VGND 0.07849f
C20446 VPWR.t951 VGND 0.11957f
C20447 VPWR.n2241 VGND 0.10822f
C20448 VPWR.n2242 VGND 0.00728f
C20449 VPWR.n2243 VGND 0.01797f
C20450 VPWR.n2244 VGND 0.13913f
C20451 VPWR.n2245 VGND 0.08351f
C20452 VPWR.n2246 VGND 0.08351f
C20453 VPWR.n2247 VGND 0.13913f
C20454 VPWR.n2248 VGND 0.01797f
C20455 VPWR.n2249 VGND 0.00728f
C20456 VPWR.n2250 VGND 0.10822f
C20457 VPWR.t573 VGND 0.09218f
C20458 VPWR.t1272 VGND 0.07849f
C20459 VPWR.t1800 VGND 0.11957f
C20460 VPWR.n2251 VGND 0.10822f
C20461 VPWR.n2252 VGND 0.00728f
C20462 VPWR.n2253 VGND 0.01797f
C20463 VPWR.n2254 VGND 0.13913f
C20464 VPWR.n2255 VGND 0.08351f
C20465 VPWR.n2256 VGND 0.08351f
C20466 VPWR.n2257 VGND 0.13913f
C20467 VPWR.n2258 VGND 0.01797f
C20468 VPWR.n2259 VGND 0.00728f
C20469 VPWR.n2260 VGND 0.10822f
C20470 VPWR.t567 VGND 0.09218f
C20471 VPWR.t1219 VGND 0.07849f
C20472 VPWR.t1513 VGND 0.11957f
C20473 VPWR.n2261 VGND 0.10822f
C20474 VPWR.n2262 VGND 0.00728f
C20475 VPWR.n2263 VGND 0.01797f
C20476 VPWR.n2264 VGND 0.13913f
C20477 VPWR.n2265 VGND 0.08351f
C20478 VPWR.n2266 VGND 0.08351f
C20479 VPWR.n2267 VGND 0.13913f
C20480 VPWR.n2268 VGND 0.01797f
C20481 VPWR.n2269 VGND 0.00728f
C20482 VPWR.n2270 VGND 0.10822f
C20483 VPWR.t1035 VGND 0.09218f
C20484 VPWR.t429 VGND 0.07849f
C20485 VPWR.t1360 VGND 0.11957f
C20486 VPWR.n2271 VGND 0.10822f
C20487 VPWR.n2272 VGND 0.00728f
C20488 VPWR.n2273 VGND 0.01797f
C20489 VPWR.n2274 VGND 0.13913f
C20490 VPWR.n2275 VGND 0.08351f
C20491 VPWR.n2276 VGND 0.08351f
C20492 VPWR.n2277 VGND 0.13913f
C20493 VPWR.n2278 VGND 0.01797f
C20494 VPWR.n2279 VGND 0.00728f
C20495 VPWR.n2280 VGND 0.10822f
C20496 VPWR.t1086 VGND 0.09218f
C20497 VPWR.t1221 VGND 0.07849f
C20498 VPWR.t533 VGND 0.11957f
C20499 VPWR.n2281 VGND 0.10822f
C20500 VPWR.n2282 VGND 0.00728f
C20501 VPWR.n2283 VGND 0.01797f
C20502 VPWR.n2284 VGND 0.13913f
C20503 VPWR.n2285 VGND 0.08351f
C20504 VPWR.n2286 VGND 1.0094f
C20505 VPWR.n2287 VGND 0.19371f
C20506 VPWR.n2288 VGND 0.08351f
C20507 VPWR.n2289 VGND 0.08351f
C20508 VPWR.n2290 VGND 0.08351f
C20509 VPWR.n2291 VGND 0.08351f
C20510 VPWR.n2292 VGND 0.08351f
C20511 VPWR.n2293 VGND 0.08351f
C20512 VPWR.n2294 VGND 0.08351f
C20513 VPWR.n2295 VGND 0.08351f
C20514 VPWR.n2296 VGND 0.08351f
C20515 VPWR.n2297 VGND 0.08351f
C20516 VPWR.n2298 VGND 0.08351f
C20517 VPWR.n2299 VGND 0.08351f
C20518 VPWR.n2300 VGND 0.08351f
C20519 VPWR.n2301 VGND 0.08351f
C20520 VPWR.n2302 VGND 0.08351f
C20521 VPWR.n2303 VGND 1.0094f
C20522 VPWR.n2304 VGND 1.0094f
C20523 VPWR.n2305 VGND 0.08351f
C20524 VPWR.n2306 VGND 0.13913f
C20525 VPWR.n2307 VGND 0.01797f
C20526 VPWR.n2308 VGND 0.00728f
C20527 VPWR.n2309 VGND 0.10822f
C20528 VPWR.t710 VGND 0.11957f
C20529 VPWR.t1623 VGND 0.07849f
C20530 VPWR.t1519 VGND 0.09218f
C20531 VPWR.t1645 VGND 0.07849f
C20532 VPWR.t841 VGND 0.11957f
C20533 VPWR.n2310 VGND 0.10822f
C20534 VPWR.n2311 VGND 0.00728f
C20535 VPWR.n2312 VGND 0.01797f
C20536 VPWR.n2313 VGND 0.13913f
C20537 VPWR.n2314 VGND 0.08351f
C20538 VPWR.n2315 VGND 0.08351f
C20539 VPWR.n2316 VGND 0.13913f
C20540 VPWR.n2317 VGND 0.01797f
C20541 VPWR.n2318 VGND 0.00728f
C20542 VPWR.n2319 VGND 0.10822f
C20543 VPWR.t1406 VGND 0.11957f
C20544 VPWR.t1644 VGND 0.07849f
C20545 VPWR.t1857 VGND 0.09218f
C20546 VPWR.t1096 VGND 0.07849f
C20547 VPWR.t1027 VGND 0.11957f
C20548 VPWR.n2320 VGND 0.10822f
C20549 VPWR.n2321 VGND 0.00728f
C20550 VPWR.n2322 VGND 0.01797f
C20551 VPWR.n2323 VGND 0.13913f
C20552 VPWR.n2324 VGND 0.08351f
C20553 VPWR.n2325 VGND 0.08351f
C20554 VPWR.n2326 VGND 0.13913f
C20555 VPWR.n2327 VGND 0.01797f
C20556 VPWR.n2328 VGND 0.00728f
C20557 VPWR.n2329 VGND 0.10822f
C20558 VPWR.t1567 VGND 0.11957f
C20559 VPWR.t800 VGND 0.07849f
C20560 VPWR.t967 VGND 0.09218f
C20561 VPWR.t799 VGND 0.07849f
C20562 VPWR.t963 VGND 0.11957f
C20563 VPWR.n2330 VGND 0.10822f
C20564 VPWR.n2331 VGND 0.00728f
C20565 VPWR.n2332 VGND 0.01797f
C20566 VPWR.n2333 VGND 0.13913f
C20567 VPWR.n2334 VGND 0.08351f
C20568 VPWR.n2335 VGND 0.08351f
C20569 VPWR.n2336 VGND 0.13913f
C20570 VPWR.n2337 VGND 0.01797f
C20571 VPWR.n2338 VGND 0.00728f
C20572 VPWR.n2339 VGND 0.10822f
C20573 VPWR.t736 VGND 0.11957f
C20574 VPWR.t1095 VGND 0.07849f
C20575 VPWR.t870 VGND 0.09218f
C20576 VPWR.t1625 VGND 0.07849f
C20577 VPWR.t858 VGND 0.11957f
C20578 VPWR.n2340 VGND 0.10822f
C20579 VPWR.n2341 VGND 0.00728f
C20580 VPWR.n2342 VGND 0.01797f
C20581 VPWR.n2343 VGND 0.13913f
C20582 VPWR.n2344 VGND 0.08351f
C20583 VPWR.n2345 VGND 0.08351f
C20584 VPWR.n2346 VGND 0.13913f
C20585 VPWR.n2347 VGND 0.01797f
C20586 VPWR.n2348 VGND 0.00728f
C20587 VPWR.n2349 VGND 0.10822f
C20588 VPWR.t479 VGND 0.11957f
C20589 VPWR.t801 VGND 0.07849f
C20590 VPWR.t672 VGND 0.09218f
C20591 VPWR.t1643 VGND 0.07849f
C20592 VPWR.t664 VGND 0.11957f
C20593 VPWR.n2350 VGND 0.10822f
C20594 VPWR.n2351 VGND 0.00728f
C20595 VPWR.n2352 VGND 0.01797f
C20596 VPWR.n2353 VGND 0.13913f
C20597 VPWR.n2354 VGND 0.08351f
C20598 VPWR.n2355 VGND 0.08351f
C20599 VPWR.n2356 VGND 0.13913f
C20600 VPWR.n2357 VGND 0.01797f
C20601 VPWR.n2358 VGND 0.00728f
C20602 VPWR.n2359 VGND 0.10822f
C20603 VPWR.t1577 VGND 0.11957f
C20604 VPWR.t1642 VGND 0.07849f
C20605 VPWR.t1758 VGND 0.09218f
C20606 VPWR.t798 VGND 0.07849f
C20607 VPWR.t471 VGND 0.11957f
C20608 VPWR.n2360 VGND 0.10822f
C20609 VPWR.n2361 VGND 0.00728f
C20610 VPWR.n2362 VGND 0.01797f
C20611 VPWR.n2363 VGND 0.13913f
C20612 VPWR.n2364 VGND 0.08351f
C20613 VPWR.n2365 VGND 0.08351f
C20614 VPWR.n2366 VGND 0.13913f
C20615 VPWR.n2367 VGND 0.01797f
C20616 VPWR.n2368 VGND 0.00728f
C20617 VPWR.n2369 VGND 0.10822f
C20618 VPWR.t453 VGND 0.11957f
C20619 VPWR.t797 VGND 0.07849f
C20620 VPWR.t1617 VGND 0.09218f
C20621 VPWR.t1646 VGND 0.07849f
C20622 VPWR.t1491 VGND 0.11957f
C20623 VPWR.n2370 VGND 0.10822f
C20624 VPWR.n2371 VGND 0.00728f
C20625 VPWR.n2372 VGND 0.01797f
C20626 VPWR.n2373 VGND 0.13913f
C20627 VPWR.n2374 VGND 0.08351f
C20628 VPWR.n2375 VGND 0.08351f
C20629 VPWR.n2376 VGND 0.13913f
C20630 VPWR.n2377 VGND 0.01797f
C20631 VPWR.n2378 VGND 0.00728f
C20632 VPWR.n2379 VGND 0.10822f
C20633 VPWR.t694 VGND 0.11957f
C20634 VPWR.t1624 VGND 0.07849f
C20635 VPWR.t148 VGND 0.13333f
C20636 VPWR.n2380 VGND 0.07618f
C20637 VPWR.n2381 VGND 0.01797f
C20638 VPWR.n2382 VGND 0.13913f
C20639 VPWR.n2383 VGND 0.19371f
C20640 VPWR.n2384 VGND 1.01577f
C20641 VPWR.n2385 VGND 0.08351f
C20642 VPWR.n2386 VGND 0.08351f
C20643 VPWR.n2387 VGND 0.08351f
C20644 VPWR.n2388 VGND 0.08351f
C20645 VPWR.n2389 VGND 0.08351f
C20646 VPWR.n2390 VGND 0.08351f
C20647 VPWR.n2391 VGND 0.08351f
C20648 VPWR.n2392 VGND 0.08351f
C20649 VPWR.n2393 VGND 0.08351f
C20650 VPWR.n2394 VGND 0.08351f
C20651 VPWR.n2395 VGND 0.08351f
C20652 VPWR.n2396 VGND 0.08351f
C20653 VPWR.n2397 VGND 0.08351f
C20654 VPWR.n2398 VGND 0.08351f
C20655 VPWR.n2399 VGND 0.08351f
C20656 VPWR.n2400 VGND 0.19371f
C20657 VPWR.n2401 VGND 1.01577f
C20658 VPWR.n2402 VGND 1.01577f
C20659 VPWR.n2403 VGND 0.19371f
C20660 VPWR.n2404 VGND 0.13913f
C20661 VPWR.n2405 VGND 0.01797f
C20662 VPWR.n2406 VGND 0.07618f
C20663 VPWR.t318 VGND 0.13333f
C20664 VPWR.t1275 VGND 0.07849f
C20665 VPWR.t632 VGND 0.11957f
C20666 VPWR.n2407 VGND 0.10822f
C20667 VPWR.n2408 VGND 0.00728f
C20668 VPWR.n2409 VGND 0.01797f
C20669 VPWR.n2410 VGND 0.13913f
C20670 VPWR.n2411 VGND 0.08351f
C20671 VPWR.n2412 VGND 0.08351f
C20672 VPWR.n2413 VGND 0.13913f
C20673 VPWR.n2414 VGND 0.01797f
C20674 VPWR.n2415 VGND 0.00728f
C20675 VPWR.n2416 VGND 0.10822f
C20676 VPWR.t860 VGND 0.09218f
C20677 VPWR.t500 VGND 0.07849f
C20678 VPWR.t924 VGND 0.11957f
C20679 VPWR.n2417 VGND 0.10822f
C20680 VPWR.n2418 VGND 0.00728f
C20681 VPWR.n2419 VGND 0.01797f
C20682 VPWR.n2420 VGND 0.13913f
C20683 VPWR.n2421 VGND 0.08351f
C20684 VPWR.n2422 VGND 0.08351f
C20685 VPWR.n2423 VGND 0.13913f
C20686 VPWR.n2424 VGND 0.01797f
C20687 VPWR.n2425 VGND 0.00728f
C20688 VPWR.n2426 VGND 0.10822f
C20689 VPWR.t1461 VGND 0.09218f
C20690 VPWR.t1531 VGND 0.07849f
C20691 VPWR.t1098 VGND 0.11957f
C20692 VPWR.n2427 VGND 0.10822f
C20693 VPWR.n2428 VGND 0.00728f
C20694 VPWR.n2429 VGND 0.01797f
C20695 VPWR.n2430 VGND 0.13913f
C20696 VPWR.n2431 VGND 0.08351f
C20697 VPWR.n2432 VGND 0.08351f
C20698 VPWR.n2433 VGND 0.13913f
C20699 VPWR.n2434 VGND 0.01797f
C20700 VPWR.n2435 VGND 0.00728f
C20701 VPWR.n2436 VGND 0.10822f
C20702 VPWR.t652 VGND 0.09218f
C20703 VPWR.t1662 VGND 0.07849f
C20704 VPWR.t1920 VGND 0.11957f
C20705 VPWR.n2437 VGND 0.10822f
C20706 VPWR.n2438 VGND 0.00728f
C20707 VPWR.n2439 VGND 0.01797f
C20708 VPWR.n2440 VGND 0.13913f
C20709 VPWR.n2441 VGND 0.08351f
C20710 VPWR.n2442 VGND 0.08351f
C20711 VPWR.n2443 VGND 0.13913f
C20712 VPWR.n2444 VGND 0.01797f
C20713 VPWR.n2445 VGND 0.00728f
C20714 VPWR.n2446 VGND 0.10822f
C20715 VPWR.t913 VGND 0.09218f
C20716 VPWR.t1277 VGND 0.07849f
C20717 VPWR.t728 VGND 0.11957f
C20718 VPWR.n2447 VGND 0.10822f
C20719 VPWR.n2448 VGND 0.00728f
C20720 VPWR.n2449 VGND 0.01797f
C20721 VPWR.n2450 VGND 0.13913f
C20722 VPWR.n2451 VGND 0.08351f
C20723 VPWR.n2452 VGND 0.08351f
C20724 VPWR.n2453 VGND 0.13913f
C20725 VPWR.n2454 VGND 0.01797f
C20726 VPWR.n2455 VGND 0.00728f
C20727 VPWR.n2456 VGND 0.10822f
C20728 VPWR.t688 VGND 0.09218f
C20729 VPWR.t1661 VGND 0.07849f
C20730 VPWR.t1546 VGND 0.11957f
C20731 VPWR.n2457 VGND 0.10822f
C20732 VPWR.n2458 VGND 0.00728f
C20733 VPWR.n2459 VGND 0.01797f
C20734 VPWR.n2460 VGND 0.13913f
C20735 VPWR.n2461 VGND 0.08351f
C20736 VPWR.n2462 VGND 0.08351f
C20737 VPWR.n2463 VGND 0.13913f
C20738 VPWR.n2464 VGND 0.01797f
C20739 VPWR.n2465 VGND 0.00728f
C20740 VPWR.n2466 VGND 0.10822f
C20741 VPWR.t1636 VGND 0.09218f
C20742 VPWR.t1533 VGND 0.07849f
C20743 VPWR.t1372 VGND 0.11957f
C20744 VPWR.n2467 VGND 0.10822f
C20745 VPWR.n2468 VGND 0.00728f
C20746 VPWR.n2469 VGND 0.01797f
C20747 VPWR.n2470 VGND 0.13913f
C20748 VPWR.n2471 VGND 0.08351f
C20749 VPWR.n2472 VGND 0.08351f
C20750 VPWR.n2473 VGND 0.13913f
C20751 VPWR.n2474 VGND 0.01797f
C20752 VPWR.n2475 VGND 0.00728f
C20753 VPWR.n2476 VGND 0.10822f
C20754 VPWR.t835 VGND 0.09218f
C20755 VPWR.t1663 VGND 0.07849f
C20756 VPWR.t1154 VGND 0.11957f
C20757 VPWR.n2477 VGND 0.10822f
C20758 VPWR.n2478 VGND 0.00728f
C20759 VPWR.n2479 VGND 0.01797f
C20760 VPWR.n2480 VGND 0.13913f
C20761 VPWR.n2481 VGND 0.08351f
C20762 VPWR.n2482 VGND 1.0094f
C20763 VPWR.n2483 VGND 0.19371f
C20764 VPWR.n2484 VGND 0.08351f
C20765 VPWR.n2485 VGND 0.08351f
C20766 VPWR.n2486 VGND 0.08351f
C20767 VPWR.n2487 VGND 0.08351f
C20768 VPWR.n2488 VGND 0.08351f
C20769 VPWR.n2489 VGND 0.08351f
C20770 VPWR.n2490 VGND 0.08351f
C20771 VPWR.n2491 VGND 0.08351f
C20772 VPWR.n2492 VGND 0.08351f
C20773 VPWR.n2493 VGND 0.08351f
C20774 VPWR.n2494 VGND 0.08351f
C20775 VPWR.n2495 VGND 0.08351f
C20776 VPWR.n2496 VGND 0.08351f
C20777 VPWR.n2497 VGND 0.08351f
C20778 VPWR.n2498 VGND 0.08351f
C20779 VPWR.n2499 VGND 1.0094f
C20780 VPWR.n2500 VGND 0.5713f
C20781 VPWR.n2501 VGND 0.08351f
C20782 VPWR.n2502 VGND 0.08654f
C20783 VPWR.n2503 VGND 0.00805f
C20784 VPWR.n2504 VGND 0.01714f
C20785 VPWR.n2505 VGND 0.00725f
C20786 VPWR.n2506 VGND 0.10822f
C20787 VPWR.t197 VGND 0.11957f
C20788 VPWR.t164 VGND 0.07849f
C20789 VPWR.t288 VGND 0.09218f
C20790 VPWR.t294 VGND 0.07849f
C20791 VPWR.t309 VGND 0.11957f
C20792 VPWR.n2507 VGND 0.10822f
C20793 VPWR.n2508 VGND 0.00725f
C20794 VPWR.n2509 VGND 0.01714f
C20795 VPWR.n2510 VGND 0.00805f
C20796 VPWR.n2511 VGND 0.08654f
C20797 VPWR.n2512 VGND 0.08351f
C20798 VPWR.n2513 VGND 0.08351f
C20799 VPWR.n2514 VGND 0.08654f
C20800 VPWR.n2515 VGND 0.00805f
C20801 VPWR.n2516 VGND 0.01714f
C20802 VPWR.n2517 VGND 0.00725f
C20803 VPWR.n2518 VGND 0.10822f
C20804 VPWR.t74 VGND 0.11957f
C20805 VPWR.t334 VGND 0.07849f
C20806 VPWR.t68 VGND 0.09218f
C20807 VPWR.t58 VGND 0.07849f
C20808 VPWR.t182 VGND 0.11957f
C20809 VPWR.n2519 VGND 0.10822f
C20810 VPWR.n2520 VGND 0.00725f
C20811 VPWR.n2521 VGND 0.01714f
C20812 VPWR.n2522 VGND 0.00805f
C20813 VPWR.n2523 VGND 0.08654f
C20814 VPWR.n2524 VGND 0.08351f
C20815 VPWR.n2525 VGND 0.08351f
C20816 VPWR.n2526 VGND 0.08654f
C20817 VPWR.n2527 VGND 0.00805f
C20818 VPWR.n2528 VGND 0.01714f
C20819 VPWR.n2529 VGND 0.00725f
C20820 VPWR.n2530 VGND 0.10822f
C20821 VPWR.t194 VGND 0.11957f
C20822 VPWR.t202 VGND 0.07849f
C20823 VPWR.t331 VGND 0.09218f
C20824 VPWR.t226 VGND 0.07849f
C20825 VPWR.t350 VGND 0.11957f
C20826 VPWR.n2531 VGND 0.10822f
C20827 VPWR.n2532 VGND 0.00725f
C20828 VPWR.n2533 VGND 0.01714f
C20829 VPWR.n2534 VGND 0.00805f
C20830 VPWR.n2535 VGND 0.08654f
C20831 VPWR.n2536 VGND 0.08351f
C20832 VPWR.n2537 VGND 0.08351f
C20833 VPWR.n2538 VGND 0.08654f
C20834 VPWR.n2539 VGND 0.00805f
C20835 VPWR.n2540 VGND 0.01714f
C20836 VPWR.n2541 VGND 0.00725f
C20837 VPWR.n2542 VGND 0.10822f
C20838 VPWR.t71 VGND 0.11957f
C20839 VPWR.t63 VGND 0.07849f
C20840 VPWR.t90 VGND 0.09218f
C20841 VPWR.t98 VGND 0.07849f
C20842 VPWR.t231 VGND 0.11957f
C20843 VPWR.n2543 VGND 0.10822f
C20844 VPWR.n2544 VGND 0.00725f
C20845 VPWR.n2545 VGND 0.01714f
C20846 VPWR.n2546 VGND 0.00805f
C20847 VPWR.n2547 VGND 0.08654f
C20848 VPWR.n2548 VGND 0.08351f
C20849 VPWR.n2549 VGND 0.08351f
C20850 VPWR.n2550 VGND 0.08654f
C20851 VPWR.n2551 VGND 0.00805f
C20852 VPWR.n2552 VGND 0.01714f
C20853 VPWR.n2553 VGND 0.00725f
C20854 VPWR.n2554 VGND 0.10822f
C20855 VPWR.t247 VGND 0.11957f
C20856 VPWR.t200 VGND 0.07849f
C20857 VPWR.t328 VGND 0.09218f
C20858 VPWR.t361 VGND 0.07849f
C20859 VPWR.t377 VGND 0.11957f
C20860 VPWR.n2555 VGND 0.10822f
C20861 VPWR.n2556 VGND 0.00725f
C20862 VPWR.n2557 VGND 0.01714f
C20863 VPWR.n2558 VGND 0.00805f
C20864 VPWR.n2559 VGND 0.08654f
C20865 VPWR.n2560 VGND 0.08351f
C20866 VPWR.n2561 VGND 0.08351f
C20867 VPWR.n2562 VGND 0.08654f
C20868 VPWR.n2563 VGND 0.00805f
C20869 VPWR.n2564 VGND 0.01714f
C20870 VPWR.n2565 VGND 0.00725f
C20871 VPWR.n2566 VGND 0.10822f
C20872 VPWR.t121 VGND 0.11957f
C20873 VPWR.t380 VGND 0.07849f
C20874 VPWR.t113 VGND 0.09218f
C20875 VPWR.t234 VGND 0.07849f
C20876 VPWR.t151 VGND 0.11957f
C20877 VPWR.n2567 VGND 0.10822f
C20878 VPWR.n2568 VGND 0.00725f
C20879 VPWR.n2569 VGND 0.01714f
C20880 VPWR.n2570 VGND 0.00805f
C20881 VPWR.n2571 VGND 0.08654f
C20882 VPWR.n2572 VGND 0.08351f
C20883 VPWR.n2573 VGND 0.08351f
C20884 VPWR.n2574 VGND 0.08654f
C20885 VPWR.n2575 VGND 0.00805f
C20886 VPWR.n2576 VGND 0.01714f
C20887 VPWR.n2577 VGND 0.00725f
C20888 VPWR.n2578 VGND 0.10822f
C20889 VPWR.t1 VGND 0.11957f
C20890 VPWR.t253 VGND 0.07849f
C20891 VPWR.t374 VGND 0.09218f
C20892 VPWR.t278 VGND 0.07849f
C20893 VPWR.t20 VGND 0.11957f
C20894 VPWR.n2579 VGND 0.10822f
C20895 VPWR.n2580 VGND 0.00725f
C20896 VPWR.n2581 VGND 0.01714f
C20897 VPWR.n2582 VGND 0.00805f
C20898 VPWR.n2583 VGND 0.08654f
C20899 VPWR.n2584 VGND 0.08351f
C20900 VPWR.n2585 VGND 0.08351f
C20901 VPWR.n2586 VGND 0.08654f
C20902 VPWR.n2587 VGND 0.00805f
C20903 VPWR.n2588 VGND 0.01714f
C20904 VPWR.n2589 VGND 0.00725f
C20905 VPWR.n2590 VGND 0.10822f
C20906 VPWR.t145 VGND 0.11957f
C20907 VPWR.t129 VGND 0.07849f
C20908 VPWR.t250 VGND 0.13333f
C20909 VPWR.n2591 VGND 0.07615f
C20910 VPWR.n2592 VGND 0.01698f
C20911 VPWR.n2593 VGND 0.00805f
C20912 VPWR.n2594 VGND 0.10853f
C20913 VPWR.n2595 VGND 0.19371f
C20914 VPWR.n2596 VGND 2.66265f
C20915 VPWR.n2597 VGND 1.08435f
C20916 VPWR.n2598 VGND 0.45434f
C20917 VPWR.t1248 VGND 0.05456f
C20918 VPWR.t1141 VGND 0.05456f
C20919 VPWR.n2599 VGND 0.09898f
C20920 VPWR.n2600 VGND 0.04687f
C20921 VPWR.t1247 VGND 0.01433f
C20922 VPWR.t1251 VGND 0.01433f
C20923 VPWR.n2601 VGND 0.03076f
C20924 VPWR.t1151 VGND 0.01433f
C20925 VPWR.t1139 VGND 0.01433f
C20926 VPWR.n2602 VGND 0.03076f
C20927 VPWR.n2603 VGND 0.01064f
C20928 VPWR.n2604 VGND 0.04687f
C20929 VPWR.t1340 VGND 0.01433f
C20930 VPWR.t1321 VGND 0.01433f
C20931 VPWR.n2605 VGND 0.03076f
C20932 VPWR.t1304 VGND 0.01433f
C20933 VPWR.t1310 VGND 0.01433f
C20934 VPWR.n2606 VGND 0.03076f
C20935 VPWR.t1317 VGND 0.05714f
C20936 VPWR.t1296 VGND 0.05714f
C20937 VPWR.n2607 VGND 0.13176f
C20938 VPWR.n2608 VGND 0.04228f
C20939 VPWR.n2609 VGND 0.01362f
C20940 VPWR.n2610 VGND 0.06183f
C20941 VPWR.n2611 VGND 0.0092f
C20942 VPWR.t1298 VGND 0.01433f
C20943 VPWR.t1250 VGND 0.01433f
C20944 VPWR.n2612 VGND 0.03076f
C20945 VPWR.t1316 VGND 0.01433f
C20946 VPWR.t1147 VGND 0.01433f
C20947 VPWR.n2613 VGND 0.03076f
C20948 VPWR.n2614 VGND 0.06183f
C20949 VPWR.n2615 VGND 0.01425f
C20950 VPWR.n2616 VGND 0.04687f
C20951 VPWR.n2617 VGND 0.04687f
C20952 VPWR.n2618 VGND 0.04687f
C20953 VPWR.n2619 VGND 0.01281f
C20954 VPWR.n2620 VGND 0.06183f
C20955 VPWR.n2621 VGND 0.01209f
C20956 VPWR.n2622 VGND 0.00983f
C20957 VPWR.n2623 VGND 0.04687f
C20958 VPWR.n2624 VGND 0.03515f
C20959 VPWR.n2625 VGND 0.00794f
C20960 VPWR.t1295 VGND 0.1712f
C20961 VPWR.t1303 VGND 0.25229f
C20962 VPWR.t1309 VGND 0.25229f
C20963 VPWR.t1297 VGND 0.25229f
C20964 VPWR.t1146 VGND 0.25229f
C20965 VPWR.t1150 VGND 0.25229f
C20966 VPWR.t1138 VGND 0.25229f
C20967 VPWR.t1140 VGND 0.56168f
C20968 VPWR.n2626 VGND 0.61307f
C20969 VPWR.n2627 VGND 0.01783f
C20970 VPWR.n2628 VGND 1.07531f
C20971 VPWR.n2629 VGND 0.04687f
C20972 VPWR.t1293 VGND 0.1712f
C20973 VPWR.t1306 VGND 0.25229f
C20974 VPWR.t1280 VGND 0.25229f
C20975 VPWR.t1332 VGND 0.25229f
C20976 VPWR.t887 VGND 0.25229f
C20977 VPWR.t879 VGND 0.25229f
C20978 VPWR.t891 VGND 0.25229f
C20979 VPWR.t883 VGND 0.41448f
C20980 VPWR.t527 VGND 0.44001f
C20981 VPWR.n2630 VGND 0.62092f
C20982 VPWR.n2631 VGND 0.17663f
C20983 VPWR.n2632 VGND 0.04687f
C20984 VPWR.t1465 VGND 0.01433f
C20985 VPWR.t1200 VGND 0.01433f
C20986 VPWR.n2633 VGND 0.03076f
C20987 VPWR.t880 VGND 0.01433f
C20988 VPWR.t892 VGND 0.01433f
C20989 VPWR.n2634 VGND 0.03076f
C20990 VPWR.n2635 VGND 0.06183f
C20991 VPWR.n2636 VGND 0.04687f
C20992 VPWR.t1343 VGND 0.01433f
C20993 VPWR.t1201 VGND 0.01433f
C20994 VPWR.n2637 VGND 0.03076f
C20995 VPWR.t1333 VGND 0.01433f
C20996 VPWR.t888 VGND 0.01433f
C20997 VPWR.n2638 VGND 0.03076f
C20998 VPWR.n2639 VGND 0.0092f
C20999 VPWR.t1294 VGND 0.05714f
C21000 VPWR.t1342 VGND 0.05714f
C21001 VPWR.n2640 VGND 0.13176f
C21002 VPWR.t1325 VGND 0.01433f
C21003 VPWR.t1300 VGND 0.01433f
C21004 VPWR.n2641 VGND 0.03076f
C21005 VPWR.t1307 VGND 0.01433f
C21006 VPWR.t1281 VGND 0.01433f
C21007 VPWR.n2642 VGND 0.03076f
C21008 VPWR.n2643 VGND 0.06183f
C21009 VPWR.n2644 VGND 0.01362f
C21010 VPWR.n2645 VGND 0.04228f
C21011 VPWR.n2646 VGND 0.04687f
C21012 VPWR.n2647 VGND 0.04687f
C21013 VPWR.n2648 VGND 0.01425f
C21014 VPWR.n2649 VGND 0.06183f
C21015 VPWR.n2650 VGND 0.01064f
C21016 VPWR.n2651 VGND 0.01281f
C21017 VPWR.n2652 VGND 0.04687f
C21018 VPWR.n2653 VGND 0.04687f
C21019 VPWR.n2654 VGND 0.01209f
C21020 VPWR.n2655 VGND 0.00983f
C21021 VPWR.t1464 VGND 0.05456f
C21022 VPWR.t884 VGND 0.05456f
C21023 VPWR.n2656 VGND 0.09898f
C21024 VPWR.n2657 VGND 0.00794f
C21025 VPWR.n2658 VGND 0.03515f
C21026 VPWR.n2659 VGND 0.01783f
C21027 VPWR.n2660 VGND 0.03515f
C21028 VPWR.n2661 VGND 0.01398f
C21029 VPWR.n2662 VGND 0.01083f
C21030 VPWR.t528 VGND 0.05708f
C21031 VPWR.t1079 VGND 0.05708f
C21032 VPWR.n2663 VGND 0.11537f
C21033 VPWR.n2664 VGND 0.03261f
C21034 VPWR.n2665 VGND 1.63658f
C21035 VPWR.n2666 VGND 0.04687f
C21036 VPWR.t996 VGND 0.05603f
C21037 VPWR.t1327 VGND 0.1712f
C21038 VPWR.t1284 VGND 0.25229f
C21039 VPWR.t1334 VGND 0.25229f
C21040 VPWR.t1311 VGND 0.25229f
C21041 VPWR.t406 VGND 0.25229f
C21042 VPWR.t400 VGND 0.25229f
C21043 VPWR.t408 VGND 0.25229f
C21044 VPWR.t402 VGND 0.41448f
C21045 VPWR.t849 VGND 0.15918f
C21046 VPWR.t995 VGND 0.12614f
C21047 VPWR.t1269 VGND 0.28082f
C21048 VPWR.n2667 VGND 0.55034f
C21049 VPWR.n2668 VGND 0.17401f
C21050 VPWR.n2669 VGND 0.04687f
C21051 VPWR.t401 VGND 0.01433f
C21052 VPWR.t409 VGND 0.01433f
C21053 VPWR.n2670 VGND 0.03076f
C21054 VPWR.t490 VGND 0.01433f
C21055 VPWR.t597 VGND 0.01433f
C21056 VPWR.n2671 VGND 0.03076f
C21057 VPWR.n2672 VGND 0.06183f
C21058 VPWR.n2673 VGND 0.04687f
C21059 VPWR.t1329 VGND 0.01433f
C21060 VPWR.t407 VGND 0.01433f
C21061 VPWR.n2674 VGND 0.03076f
C21062 VPWR.t1312 VGND 0.01433f
C21063 VPWR.t823 VGND 0.01433f
C21064 VPWR.n2675 VGND 0.03076f
C21065 VPWR.n2676 VGND 0.0092f
C21066 VPWR.t1341 VGND 0.05714f
C21067 VPWR.t1328 VGND 0.05714f
C21068 VPWR.n2677 VGND 0.13176f
C21069 VPWR.t1301 VGND 0.01433f
C21070 VPWR.t1347 VGND 0.01433f
C21071 VPWR.n2678 VGND 0.03076f
C21072 VPWR.t1285 VGND 0.01433f
C21073 VPWR.t1335 VGND 0.01433f
C21074 VPWR.n2679 VGND 0.03076f
C21075 VPWR.n2680 VGND 0.06183f
C21076 VPWR.n2681 VGND 0.01362f
C21077 VPWR.n2682 VGND 0.04228f
C21078 VPWR.n2683 VGND 0.04687f
C21079 VPWR.n2684 VGND 0.04687f
C21080 VPWR.n2685 VGND 0.01425f
C21081 VPWR.n2686 VGND 0.06183f
C21082 VPWR.n2687 VGND 0.01064f
C21083 VPWR.n2688 VGND 0.01281f
C21084 VPWR.n2689 VGND 0.04687f
C21085 VPWR.n2690 VGND 0.04687f
C21086 VPWR.n2691 VGND 0.01209f
C21087 VPWR.n2692 VGND 0.00983f
C21088 VPWR.t403 VGND 0.05456f
C21089 VPWR.t976 VGND 0.05456f
C21090 VPWR.n2693 VGND 0.09898f
C21091 VPWR.n2694 VGND 0.00794f
C21092 VPWR.n2695 VGND 0.03515f
C21093 VPWR.n2696 VGND 0.01783f
C21094 VPWR.n2697 VGND 0.03515f
C21095 VPWR.t1270 VGND 0.05714f
C21096 VPWR.n2698 VGND 0.07963f
C21097 VPWR.n2699 VGND 0.01064f
C21098 VPWR.n2700 VGND 0.05827f
C21099 VPWR.t850 VGND 0.05618f
C21100 VPWR.n2701 VGND 0.07281f
C21101 VPWR.n2702 VGND 0.02776f
C21102 VPWR.n2703 VGND 1.63658f
C21103 VPWR.n2704 VGND 0.04687f
C21104 VPWR.t1330 VGND 0.09709f
C21105 VPWR.t1288 VGND 0.14308f
C21106 VPWR.t1336 VGND 0.1391f
C21107 VPWR.t1314 VGND 0.22247f
C21108 VPWR.t1882 VGND 0.18922f
C21109 VPWR.t1318 VGND 0.12614f
C21110 VPWR.t1888 VGND 0.12614f
C21111 VPWR.t1290 VGND 0.12614f
C21112 VPWR.t493 VGND 0.12614f
C21113 VPWR.t1322 VGND 0.12614f
C21114 VPWR.t1886 VGND 0.12614f
C21115 VPWR.t1345 VGND 0.1757f
C21116 VPWR.t1266 VGND 0.09911f
C21117 VPWR.t941 VGND 0.10812f
C21118 VPWR.t1267 VGND 0.12614f
C21119 VPWR.t943 VGND 0.23427f
C21120 VPWR.n2705 VGND 0.37764f
C21121 VPWR.n2706 VGND 0.17419f
C21122 VPWR.t944 VGND 0.05672f
C21123 VPWR.n2707 VGND 0.04687f
C21124 VPWR.t1346 VGND 0.05606f
C21125 VPWR.t1887 VGND 0.05397f
C21126 VPWR.t1291 VGND 0.01433f
C21127 VPWR.t1323 VGND 0.01433f
C21128 VPWR.n2708 VGND 0.03076f
C21129 VPWR.t1889 VGND 0.01433f
C21130 VPWR.t494 VGND 0.01433f
C21131 VPWR.n2709 VGND 0.03076f
C21132 VPWR.n2710 VGND 0.03507f
C21133 VPWR.n2711 VGND 0.04687f
C21134 VPWR.t1315 VGND 0.01433f
C21135 VPWR.t1883 VGND 0.01433f
C21136 VPWR.n2712 VGND 0.03076f
C21137 VPWR.n2713 VGND 0.0092f
C21138 VPWR.t1331 VGND 0.05714f
C21139 VPWR.n2714 VGND 0.072f
C21140 VPWR.t1289 VGND 0.01433f
C21141 VPWR.t1337 VGND 0.01433f
C21142 VPWR.n2715 VGND 0.03076f
C21143 VPWR.n2716 VGND 0.03507f
C21144 VPWR.n2717 VGND 0.01362f
C21145 VPWR.n2718 VGND 0.04228f
C21146 VPWR.n2719 VGND 0.04687f
C21147 VPWR.n2720 VGND 0.04687f
C21148 VPWR.n2721 VGND 0.01425f
C21149 VPWR.n2722 VGND 0.03425f
C21150 VPWR.t1319 VGND 0.05015f
C21151 VPWR.n2723 VGND 0.03998f
C21152 VPWR.n2724 VGND 0.00983f
C21153 VPWR.n2725 VGND 0.04687f
C21154 VPWR.n2726 VGND 0.04687f
C21155 VPWR.n2727 VGND 0.03885f
C21156 VPWR.n2728 VGND 0.01209f
C21157 VPWR.n2729 VGND 0.05142f
C21158 VPWR.n2730 VGND 0.06775f
C21159 VPWR.n2731 VGND 0.00622f
C21160 VPWR.n2732 VGND 0.02776f
C21161 VPWR.n2733 VGND 0.01783f
C21162 VPWR.n2734 VGND 0.03515f
C21163 VPWR.t1268 VGND 0.0572f
C21164 VPWR.n2735 VGND 0.14706f
C21165 VPWR.n2736 VGND 0.01083f
C21166 VPWR.t942 VGND 0.05711f
C21167 VPWR.n2737 VGND 0.06357f
C21168 VPWR.n2738 VGND 0.02751f
C21169 VPWR.n2739 VGND 1.63658f
C21170 VPWR.n2740 VGND 0.04228f
C21171 VPWR.t1324 VGND 0.66677f
C21172 VPWR.t1283 VGND 0.25229f
C21173 VPWR.t1313 VGND 0.25229f
C21174 VPWR.t1287 VGND 0.25229f
C21175 VPWR.t1144 VGND 0.25229f
C21176 VPWR.t1142 VGND 0.25229f
C21177 VPWR.t1148 VGND 0.25229f
C21178 VPWR.t1136 VGND 0.22826f
C21179 VPWR.t392 VGND 0.55264f
C21180 VPWR.t1732 VGND 0.15318f
C21181 VPWR.n2741 VGND 0.33109f
C21182 VPWR.n2742 VGND 0.17663f
C21183 VPWR.t1252 VGND 0.01433f
C21184 VPWR.t1249 VGND 0.01433f
C21185 VPWR.n2743 VGND 0.03141f
C21186 VPWR.t1145 VGND 0.01433f
C21187 VPWR.t1143 VGND 0.01433f
C21188 VPWR.n2744 VGND 0.03141f
C21189 VPWR.n2745 VGND 0.1192f
C21190 VPWR.n2746 VGND 0.09664f
C21191 VPWR.t1253 VGND 0.01433f
C21192 VPWR.t1254 VGND 0.01433f
C21193 VPWR.n2747 VGND 0.03146f
C21194 VPWR.t1149 VGND 0.01433f
C21195 VPWR.t1137 VGND 0.01433f
C21196 VPWR.n2748 VGND 0.03146f
C21197 VPWR.n2749 VGND 0.13065f
C21198 VPWR.n2750 VGND 0.01119f
C21199 VPWR.n2751 VGND 0.37741f
C21200 VPWR.n2752 VGND 0.01783f
C21201 VPWR.n2753 VGND 0.0163f
C21202 VPWR.n2754 VGND 0.01398f
C21203 VPWR.n2755 VGND 0.01308f
C21204 VPWR.t393 VGND 0.0572f
C21205 VPWR.t775 VGND 0.0572f
C21206 VPWR.n2756 VGND 0.16894f
C21207 VPWR.n2757 VGND 0.03515f
C21208 VPWR.n2758 VGND 1.63658f
C21209 VPWR.n2759 VGND 0.04228f
C21210 VPWR.t1305 VGND 0.66677f
C21211 VPWR.t1338 VGND 0.25229f
C21212 VPWR.t1292 VGND 0.25229f
C21213 VPWR.t1339 VGND 0.25229f
C21214 VPWR.t877 VGND 0.25229f
C21215 VPWR.t889 VGND 0.25229f
C21216 VPWR.t881 VGND 0.25229f
C21217 VPWR.t885 VGND 0.22826f
C21218 VPWR.t1134 VGND 0.49107f
C21219 VPWR.t1734 VGND 0.10812f
C21220 VPWR.t1738 VGND 0.10662f
C21221 VPWR.n2760 VGND 0.32959f
C21222 VPWR.n2761 VGND 0.17663f
C21223 VPWR.t1199 VGND 0.01433f
C21224 VPWR.t1463 VGND 0.01433f
C21225 VPWR.n2762 VGND 0.03141f
C21226 VPWR.t878 VGND 0.01433f
C21227 VPWR.t890 VGND 0.01433f
C21228 VPWR.n2763 VGND 0.03141f
C21229 VPWR.n2764 VGND 0.1192f
C21230 VPWR.n2765 VGND 0.09664f
C21231 VPWR.t1210 VGND 0.01433f
C21232 VPWR.t1209 VGND 0.01433f
C21233 VPWR.n2766 VGND 0.03146f
C21234 VPWR.t882 VGND 0.01433f
C21235 VPWR.t886 VGND 0.01433f
C21236 VPWR.n2767 VGND 0.03146f
C21237 VPWR.n2768 VGND 0.13065f
C21238 VPWR.n2769 VGND 0.01119f
C21239 VPWR.n2770 VGND 0.37741f
C21240 VPWR.n2771 VGND 0.01783f
C21241 VPWR.n2772 VGND 0.01605f
C21242 VPWR.n2773 VGND 0.00767f
C21243 VPWR.t1735 VGND 0.05708f
C21244 VPWR.n2774 VGND 0.06101f
C21245 VPWR.n2775 VGND 0.00731f
C21246 VPWR.t1135 VGND 0.0572f
C21247 VPWR.n2776 VGND 0.0911f
C21248 VPWR.n2777 VGND 0.03515f
C21249 VPWR.n2778 VGND 1.63658f
C21250 VPWR.n2779 VGND 0.04279f
C21251 VPWR.t1286 VGND 0.66677f
C21252 VPWR.t1299 VGND 0.25229f
C21253 VPWR.t1326 VGND 0.25229f
C21254 VPWR.t1302 VGND 0.25229f
C21255 VPWR.t410 VGND 0.25229f
C21256 VPWR.t404 VGND 0.25229f
C21257 VPWR.t396 VGND 0.25229f
C21258 VPWR.t398 VGND 0.22826f
C21259 VPWR.t394 VGND 0.5226f
C21260 VPWR.t1730 VGND 0.18021f
C21261 VPWR.n2780 VGND 0.32809f
C21262 VPWR.n2781 VGND 0.17401f
C21263 VPWR.t1733 VGND 0.05716f
C21264 VPWR.t411 VGND 0.01433f
C21265 VPWR.t405 VGND 0.01433f
C21266 VPWR.n2782 VGND 0.03141f
C21267 VPWR.t851 VGND 0.01433f
C21268 VPWR.t1621 VGND 0.01433f
C21269 VPWR.n2783 VGND 0.03141f
C21270 VPWR.n2784 VGND 0.1192f
C21271 VPWR.n2785 VGND 0.09664f
C21272 VPWR.t397 VGND 0.01433f
C21273 VPWR.t399 VGND 0.01433f
C21274 VPWR.n2786 VGND 0.03146f
C21275 VPWR.t994 VGND 0.01433f
C21276 VPWR.t601 VGND 0.01433f
C21277 VPWR.n2787 VGND 0.03146f
C21278 VPWR.n2788 VGND 0.13065f
C21279 VPWR.n2789 VGND 0.01119f
C21280 VPWR.n2790 VGND 0.37741f
C21281 VPWR.n2791 VGND 0.01783f
C21282 VPWR.n2792 VGND 0.01579f
C21283 VPWR.t1731 VGND 0.05716f
C21284 VPWR.n2793 VGND 0.15059f
C21285 VPWR.n2794 VGND 0.01209f
C21286 VPWR.t395 VGND 0.05714f
C21287 VPWR.t774 VGND 0.05714f
C21288 VPWR.n2795 VGND 0.13446f
C21289 VPWR.n2796 VGND 0.03515f
C21290 VPWR.n2797 VGND 1.63658f
C21291 VPWR.n2798 VGND 0.04279f
C21292 VPWR.t1133 VGND 0.05714f
C21293 VPWR.n2799 VGND 0.01579f
C21294 VPWR.t1737 VGND 0.05716f
C21295 VPWR.n2800 VGND 0.01783f
C21296 VPWR.t1320 VGND 0.37815f
C21297 VPWR.t1344 VGND 0.14308f
C21298 VPWR.t1308 VGND 0.14308f
C21299 VPWR.t1282 VGND 0.14308f
C21300 VPWR.t1884 VGND 0.14308f
C21301 VPWR.t676 VGND 0.14308f
C21302 VPWR.t491 VGND 0.14308f
C21303 VPWR.t417 VGND 0.12946f
C21304 VPWR.t1132 VGND 0.29639f
C21305 VPWR.t1736 VGND 0.1022f
C21306 VPWR.n2801 VGND 0.1826f
C21307 VPWR.t492 VGND 0.01433f
C21308 VPWR.t418 VGND 0.01433f
C21309 VPWR.n2802 VGND 0.03146f
C21310 VPWR.n2803 VGND 0.07742f
C21311 VPWR.t1885 VGND 0.01433f
C21312 VPWR.t677 VGND 0.01433f
C21313 VPWR.n2804 VGND 0.03274f
C21314 VPWR.n2805 VGND 0.1748f
C21315 VPWR.n2806 VGND 0.37741f
C21316 VPWR.n2807 VGND 0.01119f
C21317 VPWR.n2808 VGND 0.09661f
C21318 VPWR.n2809 VGND 0.08481f
C21319 VPWR.n2810 VGND 0.01209f
C21320 VPWR.n2811 VGND 0.0735f
C21321 VPWR.n2812 VGND 0.03515f
C21322 VPWR.n2813 VGND 2.3816f
C21323 VPWR.n2814 VGND 1.92879f
C21324 VPWR.t978 VGND 0.02906f
C21325 VPWR.n2815 VGND 0.13023f
C21326 VPWR.n2816 VGND 0.28666f
C21327 VPWR.n2817 VGND 0.0756f
C21328 VPWR.n2818 VGND 0.0359f
C21329 VPWR.n2819 VGND 0.04384f
C21330 VPWR.n2820 VGND 0.08886f
C21331 VPWR.n2821 VGND 0.11583f
C21332 VPWR.n2822 VGND 0.08886f
C21333 VPWR.t1264 VGND 2.79496f
C21334 VPWR.t977 VGND 0.88276f
C21335 VPWR.n2823 VGND 0.11674f
C21336 VPWR.n2824 VGND 0.46189f
C21337 VPWR.t1265 VGND 0.02904f
C21338 VPWR.n2825 VGND 0.17782f
C21339 VPWR.n2826 VGND 0.01795f
C21340 VPWR.n2827 VGND 0.09797f
C21341 VPWR.n2828 VGND 0.08795f
C21342 VPWR.n2829 VGND 0.11674f
C21343 VPWR.n2830 VGND 0.07352f
C21344 VPWR.t1424 VGND 0.02904f
C21345 VPWR.n2831 VGND 0.17782f
C21346 VPWR.n2832 VGND 0.01795f
C21347 VPWR.n2833 VGND 0.11674f
C21348 VPWR.n2834 VGND 0.0764f
C21349 VPWR.n2835 VGND 0.08713f
C21350 VPWR.n2836 VGND 1.67029f
C21351 VPWR.n2837 VGND 0.08713f
C21352 VPWR.n2838 VGND 0.0764f
C21353 VPWR.n2839 VGND 0.11674f
C21354 VPWR.n2840 VGND 0.09788f
C21355 VPWR.n2841 VGND 0.08096f
C21356 VPWR.n2842 VGND 1.00402f
C21357 VPWR.n2843 VGND 0.06317f
C21358 VPWR.n2844 VGND 0.08837f
C21359 VPWR.n2845 VGND 0.06143f
C21360 VPWR.n2846 VGND 0.01795f
C21361 VPWR.n2847 VGND 0.06317f
C21362 VPWR.n2848 VGND 0.04851f
C21363 VPWR.n2849 VGND 0.17356f
C21364 VPWR.n2850 VGND 0.06838f
C21365 VPWR.n2851 VGND 0.04384f
C21366 VPWR.t1130 VGND 0.34561f
C21367 VPWR.n2852 VGND 0.08096f
C21368 VPWR.n2853 VGND 0.09788f
C21369 VPWR.n2854 VGND 0.0359f
C21370 VPWR.n2855 VGND 2.02287f
C21371 VPWR.n2856 VGND 0.0359f
C21372 VPWR.n2857 VGND 0.0359f
C21373 VPWR.n2858 VGND 0.08922f
C21374 VPWR.n2859 VGND 0.04898f
C21375 VPWR.n2860 VGND 0.37936f
C21376 VPWR.n2861 VGND 0.31214f
C21377 VPWR.t1131 VGND 0.02903f
C21378 VPWR.n2862 VGND 0.21967f
C21379 VPWR.n2863 VGND 3.34958f
C21380 XThR.Tn[2].t7 VGND 0.02313f
C21381 XThR.Tn[2].t4 VGND 0.02313f
C21382 XThR.Tn[2].n0 VGND 0.04668f
C21383 XThR.Tn[2].t6 VGND 0.02313f
C21384 XThR.Tn[2].t5 VGND 0.02313f
C21385 XThR.Tn[2].n1 VGND 0.05462f
C21386 XThR.Tn[2].n2 VGND 0.16384f
C21387 XThR.Tn[2].t10 VGND 0.01503f
C21388 XThR.Tn[2].t11 VGND 0.01503f
C21389 XThR.Tn[2].n3 VGND 0.03423f
C21390 XThR.Tn[2].t9 VGND 0.01503f
C21391 XThR.Tn[2].t8 VGND 0.01503f
C21392 XThR.Tn[2].n4 VGND 0.03423f
C21393 XThR.Tn[2].t1 VGND 0.01503f
C21394 XThR.Tn[2].t2 VGND 0.01503f
C21395 XThR.Tn[2].n5 VGND 0.05704f
C21396 XThR.Tn[2].t3 VGND 0.01503f
C21397 XThR.Tn[2].t0 VGND 0.01503f
C21398 XThR.Tn[2].n6 VGND 0.03423f
C21399 XThR.Tn[2].n7 VGND 0.16303f
C21400 XThR.Tn[2].n8 VGND 0.10078f
C21401 XThR.Tn[2].n9 VGND 0.11374f
C21402 XThR.Tn[2].t21 VGND 0.01808f
C21403 XThR.Tn[2].t14 VGND 0.01979f
C21404 XThR.Tn[2].n10 VGND 0.04833f
C21405 XThR.Tn[2].n11 VGND 0.09285f
C21406 XThR.Tn[2].t40 VGND 0.01808f
C21407 XThR.Tn[2].t31 VGND 0.01979f
C21408 XThR.Tn[2].n12 VGND 0.04833f
C21409 XThR.Tn[2].t55 VGND 0.01802f
C21410 XThR.Tn[2].t66 VGND 0.01973f
C21411 XThR.Tn[2].n13 VGND 0.05029f
C21412 XThR.Tn[2].n14 VGND 0.03533f
C21413 XThR.Tn[2].n15 VGND 0.00646f
C21414 XThR.Tn[2].n16 VGND 0.11337f
C21415 XThR.Tn[2].t15 VGND 0.01808f
C21416 XThR.Tn[2].t67 VGND 0.01979f
C21417 XThR.Tn[2].n17 VGND 0.04833f
C21418 XThR.Tn[2].t30 VGND 0.01802f
C21419 XThR.Tn[2].t43 VGND 0.01973f
C21420 XThR.Tn[2].n18 VGND 0.05029f
C21421 XThR.Tn[2].n19 VGND 0.03533f
C21422 XThR.Tn[2].n20 VGND 0.00646f
C21423 XThR.Tn[2].n21 VGND 0.11337f
C21424 XThR.Tn[2].t32 VGND 0.01808f
C21425 XThR.Tn[2].t23 VGND 0.01979f
C21426 XThR.Tn[2].n22 VGND 0.04833f
C21427 XThR.Tn[2].t47 VGND 0.01802f
C21428 XThR.Tn[2].t60 VGND 0.01973f
C21429 XThR.Tn[2].n23 VGND 0.05029f
C21430 XThR.Tn[2].n24 VGND 0.03533f
C21431 XThR.Tn[2].n25 VGND 0.00646f
C21432 XThR.Tn[2].n26 VGND 0.11337f
C21433 XThR.Tn[2].t58 VGND 0.01808f
C21434 XThR.Tn[2].t50 VGND 0.01979f
C21435 XThR.Tn[2].n27 VGND 0.04833f
C21436 XThR.Tn[2].t16 VGND 0.01802f
C21437 XThR.Tn[2].t28 VGND 0.01973f
C21438 XThR.Tn[2].n28 VGND 0.05029f
C21439 XThR.Tn[2].n29 VGND 0.03533f
C21440 XThR.Tn[2].n30 VGND 0.00646f
C21441 XThR.Tn[2].n31 VGND 0.11337f
C21442 XThR.Tn[2].t34 VGND 0.01808f
C21443 XThR.Tn[2].t25 VGND 0.01979f
C21444 XThR.Tn[2].n32 VGND 0.04833f
C21445 XThR.Tn[2].t48 VGND 0.01802f
C21446 XThR.Tn[2].t62 VGND 0.01973f
C21447 XThR.Tn[2].n33 VGND 0.05029f
C21448 XThR.Tn[2].n34 VGND 0.03533f
C21449 XThR.Tn[2].n35 VGND 0.00646f
C21450 XThR.Tn[2].n36 VGND 0.11337f
C21451 XThR.Tn[2].t70 VGND 0.01808f
C21452 XThR.Tn[2].t41 VGND 0.01979f
C21453 XThR.Tn[2].n37 VGND 0.04833f
C21454 XThR.Tn[2].t22 VGND 0.01802f
C21455 XThR.Tn[2].t20 VGND 0.01973f
C21456 XThR.Tn[2].n38 VGND 0.05029f
C21457 XThR.Tn[2].n39 VGND 0.03533f
C21458 XThR.Tn[2].n40 VGND 0.00646f
C21459 XThR.Tn[2].n41 VGND 0.11337f
C21460 XThR.Tn[2].t39 VGND 0.01808f
C21461 XThR.Tn[2].t35 VGND 0.01979f
C21462 XThR.Tn[2].n42 VGND 0.04833f
C21463 XThR.Tn[2].t54 VGND 0.01802f
C21464 XThR.Tn[2].t12 VGND 0.01973f
C21465 XThR.Tn[2].n43 VGND 0.05029f
C21466 XThR.Tn[2].n44 VGND 0.03533f
C21467 XThR.Tn[2].n45 VGND 0.00646f
C21468 XThR.Tn[2].n46 VGND 0.11337f
C21469 XThR.Tn[2].t44 VGND 0.01808f
C21470 XThR.Tn[2].t49 VGND 0.01979f
C21471 XThR.Tn[2].n47 VGND 0.04833f
C21472 XThR.Tn[2].t57 VGND 0.01802f
C21473 XThR.Tn[2].t27 VGND 0.01973f
C21474 XThR.Tn[2].n48 VGND 0.05029f
C21475 XThR.Tn[2].n49 VGND 0.03533f
C21476 XThR.Tn[2].n50 VGND 0.00646f
C21477 XThR.Tn[2].n51 VGND 0.11337f
C21478 XThR.Tn[2].t61 VGND 0.01808f
C21479 XThR.Tn[2].t69 VGND 0.01979f
C21480 XThR.Tn[2].n52 VGND 0.04833f
C21481 XThR.Tn[2].t18 VGND 0.01802f
C21482 XThR.Tn[2].t45 VGND 0.01973f
C21483 XThR.Tn[2].n53 VGND 0.05029f
C21484 XThR.Tn[2].n54 VGND 0.03533f
C21485 XThR.Tn[2].n55 VGND 0.00646f
C21486 XThR.Tn[2].n56 VGND 0.11337f
C21487 XThR.Tn[2].t52 VGND 0.01808f
C21488 XThR.Tn[2].t26 VGND 0.01979f
C21489 XThR.Tn[2].n57 VGND 0.04833f
C21490 XThR.Tn[2].t68 VGND 0.01802f
C21491 XThR.Tn[2].t63 VGND 0.01973f
C21492 XThR.Tn[2].n58 VGND 0.05029f
C21493 XThR.Tn[2].n59 VGND 0.03533f
C21494 XThR.Tn[2].n60 VGND 0.00646f
C21495 XThR.Tn[2].n61 VGND 0.11337f
C21496 XThR.Tn[2].t73 VGND 0.01808f
C21497 XThR.Tn[2].t64 VGND 0.01979f
C21498 XThR.Tn[2].n62 VGND 0.04833f
C21499 XThR.Tn[2].t24 VGND 0.01802f
C21500 XThR.Tn[2].t37 VGND 0.01973f
C21501 XThR.Tn[2].n63 VGND 0.05029f
C21502 XThR.Tn[2].n64 VGND 0.03533f
C21503 XThR.Tn[2].n65 VGND 0.00646f
C21504 XThR.Tn[2].n66 VGND 0.11337f
C21505 XThR.Tn[2].t42 VGND 0.01808f
C21506 XThR.Tn[2].t36 VGND 0.01979f
C21507 XThR.Tn[2].n67 VGND 0.04833f
C21508 XThR.Tn[2].t56 VGND 0.01802f
C21509 XThR.Tn[2].t13 VGND 0.01973f
C21510 XThR.Tn[2].n68 VGND 0.05029f
C21511 XThR.Tn[2].n69 VGND 0.03533f
C21512 XThR.Tn[2].n70 VGND 0.00646f
C21513 XThR.Tn[2].n71 VGND 0.11337f
C21514 XThR.Tn[2].t59 VGND 0.01808f
C21515 XThR.Tn[2].t51 VGND 0.01979f
C21516 XThR.Tn[2].n72 VGND 0.04833f
C21517 XThR.Tn[2].t17 VGND 0.01802f
C21518 XThR.Tn[2].t29 VGND 0.01973f
C21519 XThR.Tn[2].n73 VGND 0.05029f
C21520 XThR.Tn[2].n74 VGND 0.03533f
C21521 XThR.Tn[2].n75 VGND 0.00646f
C21522 XThR.Tn[2].n76 VGND 0.11337f
C21523 XThR.Tn[2].t19 VGND 0.01808f
C21524 XThR.Tn[2].t72 VGND 0.01979f
C21525 XThR.Tn[2].n77 VGND 0.04833f
C21526 XThR.Tn[2].t33 VGND 0.01802f
C21527 XThR.Tn[2].t46 VGND 0.01973f
C21528 XThR.Tn[2].n78 VGND 0.05029f
C21529 XThR.Tn[2].n79 VGND 0.03533f
C21530 XThR.Tn[2].n80 VGND 0.00646f
C21531 XThR.Tn[2].n81 VGND 0.11337f
C21532 XThR.Tn[2].t53 VGND 0.01808f
C21533 XThR.Tn[2].t65 VGND 0.01979f
C21534 XThR.Tn[2].n82 VGND 0.04833f
C21535 XThR.Tn[2].t71 VGND 0.01802f
C21536 XThR.Tn[2].t38 VGND 0.01973f
C21537 XThR.Tn[2].n83 VGND 0.05029f
C21538 XThR.Tn[2].n84 VGND 0.03533f
C21539 XThR.Tn[2].n85 VGND 0.00646f
C21540 XThR.Tn[2].n86 VGND 0.11337f
C21541 XThR.Tn[2].n87 VGND 0.10303f
C21542 XThR.Tn[2].n88 VGND 0.22327f
.ends

