magic
tech sky130A
timestamp 1755570943
<< nwell >>
rect -440 -55 -205 35
<< pwell >>
rect -90 -60 190 185
<< nmos >>
rect -375 125 -360 175
rect -330 125 -315 175
rect -285 125 -270 175
<< pmos >>
rect -375 -35 -360 15
rect -330 -35 -315 15
rect -285 -35 -270 15
<< mvnmos >>
rect 0 75 100 125
rect 0 0 100 50
<< ndiff >>
rect -405 167 -375 175
rect -405 130 -399 167
rect -381 130 -375 167
rect -405 125 -375 130
rect -360 167 -330 175
rect -360 130 -354 167
rect -336 130 -330 167
rect -360 125 -330 130
rect -315 171 -285 175
rect -315 154 -309 171
rect -291 154 -285 171
rect -315 125 -285 154
rect -270 167 -240 175
rect -270 130 -264 167
rect -246 130 -240 167
rect -270 125 -240 130
<< pdiff >>
rect -405 -14 -375 15
rect -405 -31 -399 -14
rect -381 -31 -375 -14
rect -405 -35 -375 -31
rect -360 11 -330 15
rect -360 -6 -354 11
rect -336 -6 -330 11
rect -360 -35 -330 -6
rect -315 -35 -285 15
rect -270 5 -240 15
rect -270 -16 -263 5
rect -245 -16 -240 5
rect -270 -35 -240 -16
<< mvndiff >>
rect 0 155 100 160
rect 0 135 10 155
rect 90 135 100 155
rect 0 125 100 135
rect 0 50 100 75
rect 0 -10 100 0
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< ndiffc >>
rect -399 130 -381 167
rect -354 130 -336 167
rect -309 154 -291 171
rect -264 130 -246 167
<< pdiffc >>
rect -399 -31 -381 -14
rect -354 -6 -336 11
rect -263 -16 -245 5
<< mvndiffc >>
rect 10 135 90 155
rect 10 -30 90 -10
<< mvpsubdiff >>
rect -90 175 -40 185
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect -90 145 -40 155
rect 140 155 155 175
rect 175 155 190 175
rect 140 145 190 155
rect -90 -30 -40 -20
rect -90 -50 -75 -30
rect -55 -50 -40 -30
rect 140 -30 190 -20
rect -90 -60 -40 -50
rect 140 -50 155 -30
rect 175 -50 190 -30
rect 140 -60 190 -50
<< mvpsubdiffcont >>
rect -75 155 -55 175
rect 155 155 175 175
rect -75 -50 -55 -30
rect 155 -50 175 -30
<< poly >>
rect -375 175 -360 190
rect -330 175 -315 190
rect -285 175 -270 190
rect -375 67 -360 125
rect -330 95 -315 125
rect -285 95 -270 125
rect -45 115 0 125
rect -415 58 -360 67
rect -339 85 -306 95
rect -339 68 -331 85
rect -314 68 -306 85
rect -339 58 -306 68
rect -285 85 -252 95
rect -285 68 -277 85
rect -260 68 -252 85
rect -45 85 -40 115
rect -20 85 0 115
rect -45 75 0 85
rect 100 115 145 125
rect 100 85 120 115
rect 140 85 145 115
rect 100 75 145 85
rect -285 58 -252 68
rect -415 41 -409 58
rect -392 41 -360 58
rect -415 30 -360 41
rect -375 15 -360 30
rect -330 15 -315 58
rect -285 15 -270 58
rect -45 40 0 50
rect -45 10 -40 40
rect -20 10 0 40
rect -45 0 0 10
rect 100 40 145 50
rect 100 10 120 40
rect 140 10 145 40
rect 100 0 145 10
rect -375 -50 -360 -35
rect -330 -50 -315 -35
rect -285 -50 -270 -35
<< polycont >>
rect -331 68 -314 85
rect -277 68 -260 85
rect -40 85 -20 115
rect 120 85 140 115
rect -409 41 -392 58
rect -40 10 -20 40
rect 120 10 140 40
<< locali >>
rect -399 167 -381 177
rect -399 95 -381 130
rect -354 167 -336 177
rect -309 171 -291 188
rect -309 146 -291 154
rect -264 167 -246 177
rect -354 129 -336 130
rect -90 175 -40 185
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect 140 155 155 175
rect 175 155 190 175
rect -90 145 -40 155
rect 0 135 10 155
rect 90 135 100 155
rect 140 145 190 155
rect -264 129 -246 130
rect -354 112 -246 129
rect -45 115 -15 125
rect -399 78 -348 95
rect -424 41 -409 58
rect -392 41 -383 58
rect -365 28 -348 78
rect -331 85 -314 94
rect -331 59 -314 68
rect -277 85 -260 94
rect -45 85 -40 115
rect -20 85 -15 115
rect -45 75 -15 85
rect 115 115 145 125
rect 115 85 120 115
rect 140 85 145 115
rect 115 75 145 85
rect -277 59 -260 68
rect -45 40 -15 50
rect -365 11 -336 28
rect -399 -14 -381 -6
rect -354 -14 -336 -6
rect -263 5 -245 13
rect -399 -33 -381 -31
rect -45 10 -40 40
rect -20 10 -15 40
rect -45 0 -15 10
rect 115 40 145 50
rect 115 10 120 40
rect 140 10 145 40
rect 115 0 145 10
rect -263 -33 -245 -16
rect 0 -20 10 -10
rect -399 -50 -245 -33
rect -90 -30 10 -20
rect 90 -20 100 -10
rect 90 -30 190 -20
rect -90 -50 -75 -30
rect -55 -50 155 -30
rect 175 -50 190 -30
rect -90 -60 190 -50
<< viali >>
rect 10 135 90 155
rect -40 85 -20 115
rect 120 85 140 115
rect -40 10 -20 40
rect 120 10 140 40
rect 10 -30 90 -10
<< metal1 >>
rect 0 155 100 185
rect 0 135 10 155
rect 90 135 100 155
rect 0 130 100 135
rect -90 115 -15 125
rect 115 115 145 125
rect -90 85 -40 115
rect -20 85 120 115
rect 140 85 145 115
rect -90 75 145 85
rect -45 40 190 50
rect -45 10 -40 40
rect -20 10 120 40
rect 140 10 190 40
rect -45 0 -15 10
rect 115 0 190 10
rect 0 -10 100 -5
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< labels >>
flabel mvndiff 5 55 95 70 0 FreeSans 80 0 0 0 SM
flabel metal1 150 5 185 45 0 FreeSans 80 0 0 0 Vbias
port 1 nsew
flabel metal1 -85 80 -50 120 0 FreeSans 80 0 0 0 Ien
flabel metal1 5 165 95 180 0 FreeSans 80 0 0 0 Iout
port 2 nsew
<< end >>
