magic
tech sky130A
timestamp 1755435637
<< pwell >>
rect -90 -60 190 185
<< mvnmos >>
rect 0 75 100 125
rect 0 0 100 50
<< mvndiff >>
rect 0 155 100 160
rect 0 135 10 155
rect 90 135 100 155
rect 0 125 100 135
rect 0 50 100 75
rect 0 -10 100 0
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< mvndiffc >>
rect 10 135 90 155
rect 10 -30 90 -10
<< mvpsubdiff >>
rect -90 175 -40 185
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect -90 145 -40 155
rect 140 155 155 175
rect 175 155 190 175
rect 140 145 190 155
rect -90 -30 -40 -20
rect -90 -50 -75 -30
rect -55 -50 -40 -30
rect 140 -30 190 -20
rect -90 -60 -40 -50
rect 140 -50 155 -30
rect 175 -50 190 -30
rect 140 -60 190 -50
<< mvpsubdiffcont >>
rect -75 155 -55 175
rect 155 155 175 175
rect -75 -50 -55 -30
rect 155 -50 175 -30
<< poly >>
rect -45 115 0 125
rect -45 85 -40 115
rect -20 85 0 115
rect -45 75 0 85
rect 100 115 145 125
rect 100 85 120 115
rect 140 85 145 115
rect 100 75 145 85
rect -45 40 0 50
rect -45 10 -40 40
rect -20 10 0 40
rect -45 0 0 10
rect 100 40 145 50
rect 100 10 120 40
rect 140 10 145 40
rect 100 0 145 10
<< polycont >>
rect -40 85 -20 115
rect 120 85 140 115
rect -40 10 -20 40
rect 120 10 140 40
<< locali >>
rect -90 175 -40 185
rect -90 155 -75 175
rect -55 155 -40 175
rect 140 175 190 185
rect 140 155 155 175
rect 175 155 190 175
rect -90 145 -40 155
rect 0 135 10 155
rect 90 135 100 155
rect 140 145 190 155
rect -45 115 -15 125
rect -45 85 -40 115
rect -20 85 -15 115
rect -45 75 -15 85
rect 115 115 145 125
rect 115 85 120 115
rect 140 85 145 115
rect 115 75 145 85
rect -45 40 -15 50
rect -45 10 -40 40
rect -20 10 -15 40
rect -45 0 -15 10
rect 115 40 145 50
rect 115 10 120 40
rect 140 10 145 40
rect 115 0 145 10
rect -90 -30 -40 -20
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 140 -30 190 -20
rect -90 -50 -75 -30
rect -55 -50 -40 -30
rect -90 -60 -40 -50
rect 140 -50 155 -30
rect 175 -50 190 -30
rect 140 -60 190 -50
<< viali >>
rect 10 135 90 155
rect -40 85 -20 115
rect 120 85 140 115
rect -40 10 -20 40
rect 120 10 140 40
rect 10 -30 90 -10
<< metal1 >>
rect 0 155 100 160
rect 0 135 10 155
rect 90 135 100 155
rect 0 130 100 135
rect -45 115 -15 125
rect 115 115 145 125
rect -45 85 -40 115
rect -20 85 120 115
rect 140 85 145 115
rect -45 75 145 85
rect -45 40 145 50
rect -45 10 -40 40
rect -20 10 120 40
rect 140 10 145 40
rect -45 0 -15 10
rect 115 0 145 10
rect 0 -10 100 -5
rect 0 -30 10 -10
rect 90 -30 100 -10
rect 0 -35 100 -30
<< labels >>
flabel mvndiff 5 55 95 70 0 FreeSans 80 0 0 0 SM
<< end >>
