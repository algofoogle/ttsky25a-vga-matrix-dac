* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias bias[2] bias[1] bias[0] data[0] data[1]
+ data[2] data[3] data[4] data[5] data[6] data[7]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t203 VGND.t1965 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2 VGND.t1518 VPWR.t1926 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t1517 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X3 VGND.t151 XThC.Tn[10].t12 XA.XIR[8].XIC[10].icell.PDM VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X4 VGND.t2508 XThR.XTBN.Y a_n997_2667# VGND.t2470 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t472 XThR.Tn[14].t12 XA.XIR[15].XIC[4].icell.PUM VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X6 VPWR.t992 VPWR.t990 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t991 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X7 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1927 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t1519 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X8 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[10].icell.Ien VGND.t2640 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X9 XThC.Tn[6].t11 XThC.XTBN.Y.t4 VGND.t406 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t12 XA.XIR[15].XIC[4].icell.Ien VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X11 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t988 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t989 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X12 VGND.t407 XThC.XTBN.Y.t5 XThC.Tn[5].t7 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t54 VGND.t345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X14 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t8 VGND.t2660 VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X15 XA.XIR[15].XIC[4].icell.Ien VPWR.t985 VPWR.t987 VPWR.t986 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X16 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t227 VGND.t2248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X17 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t982 VPWR.t984 VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t177 VGND.t1806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t3 XThC.XTB5.Y VPWR.t418 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t32 VGND.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X21 VGND.t935 XThC.Tn[1].t12 XA.XIR[8].XIC[1].icell.PDM VGND.t934 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X22 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t10 VPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t178 VGND.t1807 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X24 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t1449 VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t11 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t13 XA.XIR[8].XIC[1].icell.Ien VGND.t2641 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X27 XThR.Tn[5].t3 XThR.XTBN.Y a_n1049_5611# VPWR.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t481 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VGND.t408 XThC.XTBN.Y.t8 XThC.Tn[2].t11 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 XThR.XTB2.Y XThR.XTB6.A VPWR.t558 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t589 VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X32 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t12 VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X33 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t226 VGND.t2247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X34 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t12 VGND.t1055 VGND.t1054 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X35 VGND.t1720 XThC.Tn[5].t12 XA.XIR[12].XIC[5].icell.PDM VGND.t1719 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X36 XA.XIR[14].XIC_15.icell.PDM VPWR.t1928 VGND.t1521 VGND.t1520 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X37 VGND.t1607 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t1606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X38 VGND.t1523 VPWR.t1929 XA.XIR[14].XIC_15.icell.PDM VGND.t1522 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X39 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[5].icell.Ien VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X40 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t11 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 VGND.t1609 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t1608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t13 XA.XIR[14].XIC_15.icell.Ien VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X43 VPWR.t474 XThR.Tn[14].t14 XA.XIR[15].XIC[0].icell.PUM VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X44 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t3 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t14 VGND.t2643 VGND.t2642 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X46 XThC.XTB5.Y XThC.XTB7.B VGND.t1801 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X47 XThC.Tn[7].t3 XThC.XTBN.Y.t9 VPWR.t348 VPWR.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X48 VGND.t141 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[15].XIC[0].icell.Ien VPWR.t1311 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X50 VPWR.t1783 XThR.XTBN.Y XThR.Tn[9].t11 VPWR.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X51 XThR.XTB7.Y XThR.XTB7.A VGND.t2033 VGND.t2032 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 VGND.t1722 XThC.Tn[5].t13 XA.XIR[9].XIC[5].icell.PDM VGND.t1721 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X53 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t1964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X54 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t980 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t981 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X55 XA.XIR[15].XIC[0].icell.Ien VPWR.t977 VPWR.t979 VPWR.t978 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X56 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t974 VPWR.t976 VPWR.t975 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X57 a_6243_9615# XThC.XTB7.Y VPWR.t55 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X58 VPWR.t1609 XThR.Tn[12].t13 XA.XIR[13].XIC[12].icell.PUM VPWR.t1608 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X59 XThR.Tn[7].t3 XThR.XTBN.Y VPWR.t1782 VPWR.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 VPWR.t255 XThR.Tn[11].t12 XA.XIR[12].XIC[13].icell.PUM VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X61 VPWR.t973 VPWR.t971 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t972 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X62 a_8963_9569# XThC.XTBN.Y.t10 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t12 XA.XIR[13].XIC[12].icell.Ien VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X64 VGND.t1611 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t1610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X65 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t85 VGND.t918 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1098 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X67 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t67 VGND.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X68 VGND.t2507 XThR.XTBN.Y XThR.Tn[5].t7 VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X69 VGND.t1613 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t1612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X70 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t969 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t970 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X71 VPWR.t1229 VGND.t2688 XA.XIR[0].XIC[7].icell.PUM VPWR.t1228 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X72 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t12 VPWR.t1655 VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X73 VGND.t1977 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t1976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X74 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[1].XIC[14].icell.Ien VPWR.t1533 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X75 VPWR.t968 VPWR.t966 XA.XIR[4].XIC_15.icell.PUM VPWR.t967 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X76 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t8 XA.XIR[0].XIC[7].icell.Ien VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X77 XA.XIR[4].XIC_15.icell.PUM VPWR.t964 XA.XIR[4].XIC_15.icell.Ien VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X78 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t12 VPWR.t1439 VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X79 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t13 VPWR.t480 VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X80 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t13 VPWR.t291 VPWR.t290 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X81 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t13 VPWR.t608 VPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X82 VPWR.t1876 XThR.XTB6.Y a_n1049_5611# VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X83 VGND.t1679 XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.PDM VGND.t1678 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X84 VGND.t1979 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t1978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X85 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t14 VGND.t394 VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X86 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t14 VGND.t2217 VGND.t2216 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X87 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t15 XA.XIR[12].XIC[0].icell.Ien VGND.t2218 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X88 VGND.t472 XThC.Tn[13].t12 XA.XIR[10].XIC[13].icell.PDM VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X89 a_n1049_7787# XThR.XTB2.Y VPWR.t1643 VPWR.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 VGND.t2086 XThC.Tn[14].t13 XA.XIR[13].XIC[14].icell.PDM VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X91 VPWR.t343 XThR.Tn[9].t15 XA.XIR[10].XIC[9].icell.PUM VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X92 VGND.t1981 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t1980 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X93 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t12 XA.XIR[10].XIC[13].icell.Ien VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X94 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t15 VGND.t2645 VGND.t2644 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X95 VPWR.t1611 XThR.Tn[12].t16 XA.XIR[13].XIC[10].icell.PUM VPWR.t1610 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X96 XA.XIR[0].XIC[9].icell.PDM VGND.t1465 VGND.t1467 VGND.t1466 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X97 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t13 XA.XIR[13].XIC[14].icell.Ien VGND.t2257 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X98 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[10].XIC[9].icell.Ien VPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X99 VGND.t1983 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t1982 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X100 VGND.t1525 VPWR.t1930 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t1524 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X101 VGND.t1681 XThC.Tn[0].t14 XA.XIR[9].XIC[0].icell.PDM VGND.t1680 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X102 VGND.t756 XThC.Tn[9].t13 XA.XIR[0].XIC[9].icell.PDM VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X103 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t13 XA.XIR[13].XIC[10].icell.Ien VPWR.t144 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X104 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t13 VPWR.t115 VPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X105 VPWR.t1041 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X106 VPWR.t1127 data[4].t0 a_n1335_4229# VPWR.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X107 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1931 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t1526 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X108 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t132 VGND.t1245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X109 VPWR.t1227 VGND.t2689 XA.XIR[0].XIC[11].icell.PUM VPWR.t1226 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X110 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t14 VPWR.t1657 VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X111 VGND.t2506 XThR.XTBN.Y XThR.Tn[7].t7 VGND.t2505 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X112 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t14 XA.XIR[0].XIC[9].icell.Ien VGND.t1027 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X113 a_n1319_5317# XThR.XTB7.A VPWR.t1461 VPWR.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X114 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t12 XA.XIR[0].XIC[11].icell.Ien VPWR.t1098 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X115 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t592 VPWR.t591 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X116 XThC.Tn[9].t3 XThC.XTB2.Y VPWR.t207 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X117 VGND.t1985 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t1984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X118 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t254 VGND.t2682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X119 VGND.t1987 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t1986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X120 XThC.Tn[5].t6 XThC.XTBN.Y.t11 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X121 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t1244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X122 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t16 VGND.t396 VGND.t395 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X123 VGND.t1989 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t1988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X124 VPWR.t1225 VGND.t2690 XA.XIR[0].XIC[2].icell.PUM VPWR.t1224 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X125 VGND.t1991 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t1990 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X126 VGND.t1189 XThC.Tn[11].t13 XA.XIR[10].XIC[11].icell.PDM VGND.t1188 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X127 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[10].icell.Ien VGND.t2661 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X128 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t12 XA.XIR[0].XIC[2].icell.Ien VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X129 VGND.t1464 VGND.t1462 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X130 VPWR.t257 XThR.Tn[11].t13 XA.XIR[12].XIC[6].icell.PUM VPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X131 XThR.Tn[9].t7 XThR.XTB2.Y a_n997_3755# VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X132 XThC.Tn[0].t9 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X133 XThC.Tn[5].t10 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X134 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[11].icell.Ien VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X135 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t594 VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X136 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t1528 VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X137 VGND.t480 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X138 VGND.t1993 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t1992 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X139 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t7 VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X140 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t1530 VGND.t1529 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X141 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t17 VGND.t398 VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X142 XThC.Tn[7].t7 XThC.XTBN.Y.t14 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X143 XThC.Tn[2].t10 XThC.XTBN.Y.t15 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X144 a_n997_1579# XThR.XTBN.Y VGND.t2504 VGND.t2488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 VPWR.t117 XThR.Tn[10].t15 XA.XIR[11].XIC[4].icell.PUM VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X146 VGND.t166 XThC.Tn[2].t13 XA.XIR[10].XIC[2].icell.PDM VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X147 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t81 VGND.t750 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X148 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t10 XA.XIR[7].XIC[1].icell.Ien VGND.t2662 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X149 VPWR.t963 VPWR.t961 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t962 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X150 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[11].XIC[4].icell.Ien VPWR.t325 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X151 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[2].icell.Ien VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X152 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t959 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t960 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X153 VPWR.t1613 XThR.Tn[12].t17 XA.XIR[13].XIC[5].icell.PUM VPWR.t1612 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X154 XA.XIR[0].XIC[4].icell.PDM VGND.t1459 VGND.t1461 VGND.t1460 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X155 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t14 VPWR.t259 VPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X156 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t1141 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X157 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t956 VPWR.t958 VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X158 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t126 VGND.t1207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X159 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t70 VGND.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X160 VGND.t366 XThC.Tn[4].t14 XA.XIR[0].XIC[4].icell.PDM VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X161 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[13].XIC[5].icell.Ien VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X162 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t15 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X163 VGND.t1627 XThC.Tn[12].t13 XA.XIR[4].XIC[12].icell.PDM VGND.t1626 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X164 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t95 VGND.t1053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X165 VGND.t1995 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t1994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X166 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t15 VPWR.t1659 VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X167 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[4].icell.Ien VGND.t1028 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X168 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t14 XA.XIR[4].XIC[12].icell.Ien VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X169 VGND.t11 XThC.XTBN.Y.t16 XThC.Tn[1].t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X170 VGND.t1997 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t1996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X171 VGND.t1999 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t1998 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X172 VPWR.t3 XThC.XTBN.Y.t17 XThC.Tn[10].t0 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X173 VGND.t2503 XThR.XTBN.Y XThR.Tn[3].t11 VGND.t2466 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X174 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t18 VGND.t400 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X175 XThR.Tn[0].t7 XThR.XTBN.Y a_n1049_8581# VPWR.t1780 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X176 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t18 VGND.t1850 VGND.t1849 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X177 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t125 VGND.t1194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X178 VGND.t320 XThC.Tn[6].t12 XA.XIR[10].XIC[6].icell.PDM VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X179 VPWR.t261 XThR.Tn[11].t16 XA.XIR[12].XIC[1].icell.PUM VPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X180 VPWR.t1862 XThR.Tn[7].t11 XA.XIR[8].XIC[4].icell.PUM VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X181 VPWR.t955 VPWR.t953 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t954 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X182 VPWR.t119 XThR.Tn[10].t17 XA.XIR[11].XIC[0].icell.PUM VPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X183 VGND.t215 XThC.Tn[7].t9 XA.XIR[13].XIC[7].icell.PDM VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X184 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t18 XA.XIR[10].XIC[6].icell.Ien VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X185 XThC.Tn[12].t2 XThC.XTB5.Y VPWR.t417 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 XThR.Tn[11].t11 XThR.XTBN.Y VPWR.t1779 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 VPWR.t456 XThR.Tn[14].t15 XA.XIR[15].XIC[13].icell.PUM VPWR.t455 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X188 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[8].XIC[4].icell.Ien VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X189 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t951 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t952 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X190 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t16 XA.XIR[13].XIC[7].icell.Ien VGND.t2040 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X191 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[12].XIC[12].icell.Ien VPWR.t1278 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X192 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[11].XIC[0].icell.Ien VPWR.t1312 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X193 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t1114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X194 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t16 VPWR.t1843 VPWR.t1842 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X195 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t13 XA.XIR[15].XIC[13].icell.Ien VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X196 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t19 VPWR.t1354 VPWR.t1353 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X197 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t17 VPWR.t263 VPWR.t262 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X198 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t948 VPWR.t950 VPWR.t949 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X199 XThR.Tn[2].t10 XThR.XTBN.Y VGND.t2502 VGND.t2453 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X200 VPWR.t1441 XThR.Tn[1].t13 XA.XIR[2].XIC[8].icell.PUM VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X201 XA.XIR[15].XIC[13].icell.Ien VPWR.t945 VPWR.t947 VPWR.t946 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X202 VGND.t1458 VGND.t1456 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X203 VPWR.t1778 XThR.XTBN.Y XThR.Tn[12].t11 VPWR.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X204 VPWR.t1890 XThR.Tn[8].t17 XA.XIR[9].XIC[12].icell.PUM VPWR.t1889 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X205 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[2].XIC[8].icell.Ien VPWR.t521 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X206 XThC.XTB7.A data[0].t0 VPWR.t485 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X207 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t12 VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X208 VGND.t2001 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t2000 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X209 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[9].XIC[12].icell.Ien VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X210 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t18 VGND.t301 VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X211 VGND.t2003 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t2002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X212 XThC.Tn[9].t7 XThC.XTB2.Y a_7875_9569# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X213 VGND.t1724 XThC.Tn[5].t15 XA.XIR[5].XIC[5].icell.PDM VGND.t1723 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X214 a_n1319_5611# XThR.XTB6.A VPWR.t556 VPWR.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X215 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[5].icell.Ien VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X216 VGND.t2501 XThR.XTBN.Y a_n997_3979# VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X217 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t116 VGND.t1149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X218 VGND.t2088 XThC.Tn[14].t14 XA.XIR[12].XIC[14].icell.PDM VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X219 VPWR.t5 XThC.XTBN.Y.t18 XThC.Tn[14].t11 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X220 VGND.t2560 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t2559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X221 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t20 XA.XIR[12].XIC[14].icell.Ien VGND.t1851 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X222 VGND.t2562 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t2561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X223 VPWR.t1864 XThR.Tn[7].t12 XA.XIR[8].XIC[0].icell.PUM VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X224 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t13 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X225 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[12].XIC[10].icell.Ien VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X226 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t117 VGND.t1150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X227 VGND.t2564 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t2563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X228 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[8].XIC[0].icell.Ien VPWR.t1313 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X229 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t18 VGND.t2673 VGND.t2672 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X230 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t943 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t944 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X231 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t21 VPWR.t1356 VPWR.t1355 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X232 VGND.t474 XThC.Tn[13].t14 XA.XIR[6].XIC[13].icell.PDM VGND.t473 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X233 VPWR.t1151 XThR.XTB4.Y.t2 a_n1049_6699# VPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t140 VGND.t1469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X235 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t19 VPWR.t1892 VPWR.t1891 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X236 VGND.t1748 XThC.Tn[14].t15 XA.XIR[9].XIC[14].icell.PDM VGND.t1747 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X237 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t12 XA.XIR[6].XIC[13].icell.Ien VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X238 VPWR.t47 XThR.Tn[5].t14 XA.XIR[6].XIC[9].icell.PUM VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X239 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t940 VPWR.t942 VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X240 VPWR.t1321 XThC.XTB6.Y a_5949_9615# VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 VPWR.t1153 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X242 VPWR.t1894 XThR.Tn[8].t20 XA.XIR[9].XIC[10].icell.PUM VPWR.t1893 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X243 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[6].XIC[9].icell.Ien VPWR.t1788 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X244 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[9].XIC[10].icell.Ien VPWR.t146 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X245 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t187 VGND.t1882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X246 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t13 VPWR.t165 VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X247 VGND.t2566 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t2565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X248 VGND.t1225 XThR.XTB7.B a_n1335_8107# VGND.t1219 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X249 VPWR.t1443 XThR.Tn[1].t14 XA.XIR[2].XIC[3].icell.PUM VPWR.t1442 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X250 VGND.t2568 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t2567 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X251 XThC.XTB4.Y.t0 XThC.XTB7.B VPWR.t1352 VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X252 VGND.t1455 VGND.t1453 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X253 VPWR.t458 XThR.Tn[14].t16 XA.XIR[15].XIC[6].icell.PUM VPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X254 XThR.Tn[2].t0 XThR.XTB3.Y.t3 VGND.t430 VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X255 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t12 XA.XIR[2].XIC[3].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X256 VPWR.t1481 XThR.Tn[13].t17 XA.XIR[14].XIC[7].icell.PUM VPWR.t1480 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X257 VGND.t2500 XThR.XTBN.Y a_n997_2891# VGND.t2449 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[15].XIC[6].icell.Ien VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X259 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t13 VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X260 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1934 VGND.t1532 VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X261 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t23 VGND.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X262 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t10 XA.XIR[14].XIC[7].icell.Ien VPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X263 VPWR.t1195 XThR.XTB5.Y XThR.Tn[12].t3 VPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X264 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t14 VGND.t186 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X265 VGND.t2570 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t2569 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X266 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t15 VGND.t49 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X267 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t14 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X268 VGND.t2299 XThC.Tn[0].t17 XA.XIR[5].XIC[0].icell.PDM VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X269 XA.XIR[15].XIC[6].icell.Ien VPWR.t937 VPWR.t939 VPWR.t938 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X270 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t191 VGND.t1898 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X271 VGND.t1534 VPWR.t1935 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X272 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t17 VPWR.t460 VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X273 VGND.t153 XThC.Tn[10].t16 XA.XIR[7].XIC[10].icell.PDM VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X274 VGND.t2499 XThR.XTBN.Y XThR.Tn[6].t11 VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X275 VPWR.t1777 XThR.XTBN.Y XThR.Tn[9].t10 VPWR.t1763 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X276 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t134 VGND.t1309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X277 VGND.t1191 XThC.Tn[11].t14 XA.XIR[6].XIC[11].icell.PDM VGND.t1190 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X278 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t16 XA.XIR[5].XIC[0].icell.Ien VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X279 VGND.t1452 VGND.t1450 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X280 VGND.t476 XThC.Tn[13].t15 XA.XIR[3].XIC[13].icell.PDM VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X281 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1936 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t1535 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X282 a_n997_715# XThR.XTBN.Y VGND.t2497 VGND.t2496 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X283 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t15 XA.XIR[6].XIC[11].icell.Ien VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X284 VPWR.t57 XThR.Tn[2].t15 XA.XIR[3].XIC[9].icell.PUM VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X285 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t13 XA.XIR[3].XIC[13].icell.Ien VGND.t1142 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X286 XThC.Tn[1].t10 XThC.XTBN.Y.t19 VGND.t12 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t518 VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X288 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t17 VGND.t312 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X289 XThR.Tn[14].t3 XThR.XTB7.Y VPWR.t135 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[12].XIC[5].icell.Ien VPWR.t1323 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X291 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t223 VGND.t2234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X292 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t15 XA.XIR[3].XIC[9].icell.Ien VPWR.t1789 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X293 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t236 VGND.t2408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X294 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t934 VPWR.t936 VPWR.t935 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X295 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t172 VGND.t1793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X296 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t18 VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X297 VGND.t937 XThC.Tn[1].t13 XA.XIR[7].XIC[1].icell.PDM VGND.t936 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X298 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t14 VPWR.t1057 VPWR.t1056 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X299 VGND.t168 XThC.Tn[2].t14 XA.XIR[6].XIC[2].icell.PDM VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X300 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t18 VGND.t2042 VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X301 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t22 VPWR.t1358 VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X302 VGND.t2572 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t2571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X303 VGND.t2574 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t2573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X304 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t17 XA.XIR[6].XIC[2].icell.Ien VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X305 VGND.t691 XThC.Tn[8].t13 XA.XIR[15].XIC[8].icell.PDM VGND.t690 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X306 VGND.t2518 XThC.Tn[9].t16 XA.XIR[14].XIC[9].icell.PDM VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X307 VPWR.t1194 XThR.XTB5.Y a_n1049_6405# VPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X308 VPWR.t1483 XThR.Tn[13].t19 XA.XIR[14].XIC[11].icell.PUM VPWR.t1482 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X309 XA.XIR[15].XIC[8].icell.PDM VPWR.t1937 XA.XIR[15].XIC[8].icell.Ien VGND.t1536 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X310 XThR.XTB7.B data[6].t0 VPWR.t1631 VPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X311 VPWR.t1896 XThR.Tn[8].t21 XA.XIR[9].XIC[5].icell.PUM VPWR.t1895 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X312 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t19 XA.XIR[14].XIC[9].icell.Ien VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X313 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t17 XA.XIR[9].XIC[5].icell.Ien VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X314 VPWR.t1450 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t44 VGND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X316 VGND.t2576 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t2575 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X317 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t15 XA.XIR[14].XIC[11].icell.Ien VPWR.t1099 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X318 VGND.t2252 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X319 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X320 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t20 VPWR.t462 VPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X321 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t240 VGND.t2525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X322 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X323 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t176 VGND.t1805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X324 VGND.t2578 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t2577 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X325 VGND.t553 XThC.Tn[7].t11 XA.XIR[12].XIC[7].icell.PDM VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X326 VGND.t2014 XThC.Tn[11].t16 XA.XIR[3].XIC[11].icell.PDM VGND.t2013 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X327 VPWR.t464 XThR.Tn[14].t21 XA.XIR[15].XIC[1].icell.PUM VPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X328 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t208 VGND.t2007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X329 VPWR.t1485 XThR.Tn[13].t20 XA.XIR[14].XIC[2].icell.PUM VPWR.t1484 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X330 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t15 XA.XIR[3].XIC[11].icell.Ien VGND.t1143 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X331 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[15].XIC[1].icell.Ien VPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X332 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[7].icell.Ien VGND.t1852 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X333 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t7 VPWR.t1762 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X334 VPWR.t1360 XThR.Tn[12].t24 XA.XIR[13].XIC[14].icell.PUM VPWR.t1359 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X335 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t15 XA.XIR[14].XIC[2].icell.Ien VPWR.t152 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X336 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t130 VGND.t1242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X337 VPWR.t890 VPWR.t888 XA.XIR[12].XIC_15.icell.PUM VPWR.t889 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X338 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t13 VPWR.t1866 VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X339 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t18 VGND.t314 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X340 VGND.t14 XThC.XTBN.Y.t20 XThC.Tn[4].t11 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X341 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t69 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X342 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t16 XA.XIR[13].XIC[14].icell.Ien VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X343 XA.XIR[15].XIC[1].icell.Ien VPWR.t931 VPWR.t933 VPWR.t932 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X344 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t22 VPWR.t466 VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X345 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t245 VGND.t2635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X346 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t237 VGND.t2409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X347 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t22 VGND.t2675 VGND.t2674 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X348 VGND.t322 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X349 VGND.t1449 VGND.t1447 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X350 VGND.t170 XThC.Tn[2].t16 XA.XIR[3].XIC[2].icell.PDM VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X351 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t1487 VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X352 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t14 XA.XIR[1].XIC[8].icell.Ien VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X353 VGND.t555 XThC.Tn[7].t12 XA.XIR[9].XIC[7].icell.PDM VGND.t554 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X354 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X355 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t18 XA.XIR[6].XIC[6].icell.Ien VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X356 VGND.t1643 data[1].t1 a_8739_10571# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X357 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t16 XA.XIR[3].XIC[2].icell.Ien VGND.t1144 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X358 VPWR.t1642 XThR.XTB2.Y XThR.Tn[9].t3 VPWR.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X359 VGND.t2495 XThR.XTBN.Y XThR.Tn[7].t6 VGND.t2494 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X360 VPWR.t107 XThR.Tn[10].t19 XA.XIR[11].XIC[13].icell.PUM VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X361 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t15 VPWR.t1445 VPWR.t1444 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X362 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t230 VGND.t2340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X363 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[11].XIC[13].icell.Ien VPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X364 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t23 VGND.t539 VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X365 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t22 VGND.t2044 VGND.t2043 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X366 XThR.Tn[13].t3 XThR.XTBN.Y VPWR.t1776 VPWR.t1738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X367 XA.XIR[10].XIC_15.icell.PDM VPWR.t1938 VGND.t1538 VGND.t1537 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X368 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t19 VPWR.t1505 VPWR.t1504 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X369 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t201 VGND.t1933 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X370 VGND.t2670 XThC.Tn[3].t13 XA.XIR[15].XIC[3].icell.PDM VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X371 VGND.t2580 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t2579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X372 VGND.t1446 VGND.t1444 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X373 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1939 VGND.t1540 VGND.t1539 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X374 VGND.t368 XThC.Tn[4].t16 XA.XIR[14].XIC[4].icell.PDM VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X375 VGND.t1542 VPWR.t1940 XA.XIR[10].XIC_15.icell.PDM VGND.t1541 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X376 XA.XIR[15].XIC[3].icell.PDM VPWR.t1941 XA.XIR[15].XIC[3].icell.Ien VGND.t1543 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X377 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t18 VGND.t1030 VGND.t1029 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X378 VGND.t1545 VPWR.t1942 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t1544 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X379 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[4].icell.Ien VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X380 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t20 XA.XIR[10].XIC_15.icell.Ien VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X381 VGND.t2668 XThR.XTB6.Y XThR.Tn[5].t11 VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X382 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t15 VGND.t1058 VGND.t1057 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X383 XThR.Tn[9].t6 XThR.XTB2.Y a_n997_3755# VGND.t1278 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X384 VGND.t2582 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t2581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X385 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1943 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X386 XThR.XTB6.Y XThR.XTB6.A VGND.t731 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X387 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X388 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t14 VPWR.t1868 VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X389 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t252 VGND.t2664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X390 VGND.t324 XThC.Tn[6].t15 XA.XIR[3].XIC[6].icell.PDM VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X391 a_n997_1579# XThR.XTBN.Y VGND.t2493 VGND.t2483 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t89 VGND.t1041 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X393 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t19 XA.XIR[9].XIC[13].icell.Ien VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X394 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t17 XA.XIR[3].XIC[6].icell.Ien VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X395 VPWR.t930 VPWR.t928 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t929 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X396 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X397 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t16 XA.XIR[5].XIC[12].icell.Ien VPWR.t1280 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X398 VPWR.t496 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X399 VPWR.t927 VPWR.t925 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X400 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t20 VPWR.t345 VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X401 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t19 VPWR.t277 VPWR.t276 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X402 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[8].XIC[13].icell.Ien VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X403 VGND.t2584 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t2583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X404 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[1].XIC[3].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X405 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t23 VPWR.t1898 VPWR.t1897 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X406 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t16 VPWR.t177 VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X407 VPWR.t534 XThR.XTBN.A XThR.XTBN.Y VPWR.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X408 VPWR.t109 XThR.Tn[10].t21 XA.XIR[11].XIC[6].icell.PUM VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X409 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t20 VGND.t2053 VGND.t2052 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X410 VGND.t1750 XThC.Tn[14].t17 XA.XIR[5].XIC[14].icell.PDM VGND.t1749 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X411 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t21 XA.XIR[9].XIC[11].icell.Ien VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X412 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t19 VGND.t1032 VGND.t1031 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X413 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t16 XA.XIR[11].XIC[6].icell.Ien VPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X414 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t20 XA.XIR[5].XIC[14].icell.Ien VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X415 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t175 VGND.t1804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X416 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t16 VGND.t1060 VGND.t1059 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X417 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t21 VPWR.t1507 VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X418 a_3523_10575# XThC.XTB7.B VGND.t1800 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X419 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t17 XA.XIR[5].XIC[10].icell.Ien VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X420 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t143 VGND.t1486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X421 VPWR.t7 XThC.XTBN.Y.t21 XThC.Tn[13].t11 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X422 VGND.t2586 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t2585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X423 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t21 VPWR.t279 VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X424 XThC.Tn[5].t3 XThC.XTB6.Y VGND.t1685 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X425 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t479 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X426 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t22 XA.XIR[9].XIC[2].icell.Ien VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X427 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t11 VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X428 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t22 VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X429 VGND.t1000 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t999 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X430 VGND.t1002 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t1001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X431 VGND.t693 XThC.Tn[8].t15 XA.XIR[11].XIC[8].icell.PDM VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X432 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t6 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 XThC.Tn[4].t10 XThC.XTBN.Y.t22 VGND.t15 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X434 a_n1049_5317# XThR.XTB7.Y VPWR.t133 VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X435 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t118 VGND.t1173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X436 VGND.t1004 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t1003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VGND.t1443 VGND.t1441 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t22 XA.XIR[11].XIC[8].icell.Ien VGND.t2054 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X439 XThC.XTB6.Y XThC.XTB7.B VGND.t1799 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X440 VPWR.t498 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X441 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X442 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X443 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[8].XIC[6].icell.Ien VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X444 XA.XIR[0].XIC[10].icell.PDM VGND.t1438 VGND.t1440 VGND.t1439 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X445 VPWR.t924 VPWR.t922 XA.XIR[15].XIC_15.icell.PUM VPWR.t923 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X446 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t18 XA.XIR[12].XIC[14].icell.Ien VPWR.t1339 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X447 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t199 VGND.t1911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X448 XA.XIR[15].XIC_15.icell.PUM VPWR.t920 XA.XIR[15].XIC_15.icell.Ien VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X449 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t25 VPWR.t1362 VPWR.t1361 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X450 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t24 VPWR.t1900 VPWR.t1899 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X451 XThC.Tn[13].t7 XThC.XTB6.Y VPWR.t1320 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X452 VGND.t155 XThC.Tn[10].t18 XA.XIR[0].XIC[10].icell.PDM VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X453 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t174 VGND.t1803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X454 VPWR.t111 XThR.Tn[10].t23 XA.XIR[11].XIC[1].icell.PUM VPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X455 VPWR.t426 XThR.Tn[6].t19 XA.XIR[7].XIC[4].icell.PUM VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X456 VPWR.t919 VPWR.t917 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t918 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X457 VGND.t17 XThC.XTBN.Y.t24 XThC.Tn[0].t6 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t20 XA.XIR[0].XIC[10].icell.Ien VGND.t1033 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X459 XA.XIR[15].XIC_15.icell.Ien VPWR.t914 VPWR.t916 VPWR.t915 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X460 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t23 XA.XIR[9].XIC[6].icell.Ien VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X461 XThR.Tn[3].t7 XThR.XTBN.Y a_n1049_6699# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X462 VGND.t2238 XThR.XTB4.Y.t3 XThR.Tn[3].t3 VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X463 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t15 XA.XIR[11].XIC[1].icell.Ien VPWR.t587 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X464 VPWR.t1902 XThR.Tn[8].t25 XA.XIR[9].XIC[14].icell.PUM VPWR.t1901 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X465 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[7].XIC[4].icell.Ien VPWR.t327 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X466 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t912 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t913 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X467 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t68 VGND.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X468 XA.XIR[0].XIC[1].icell.PDM VGND.t1435 VGND.t1437 VGND.t1436 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X469 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t23 VPWR.t1509 VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X470 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t909 VPWR.t911 VPWR.t910 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X471 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[5].XIC[5].icell.Ien VPWR.t1325 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X472 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[9].XIC[14].icell.Ien VPWR.t1340 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X473 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t189 VGND.t1884 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X474 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t167 VGND.t1717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X475 VGND.t939 XThC.Tn[1].t16 XA.XIR[0].XIC[1].icell.PDM VGND.t938 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X476 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t22 VPWR.t281 VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X477 VGND.t1006 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X478 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t17 VGND.t665 VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X479 VGND.t1008 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X480 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t205 VGND.t2004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X481 XThR.Tn[11].t5 XThR.XTB4.Y.t4 VPWR.t1618 VPWR.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X482 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[1].icell.Ien VGND.t1034 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X483 VGND.t695 XThC.Tn[8].t16 XA.XIR[8].XIC[8].icell.PDM VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X484 VGND.t1548 VPWR.t1944 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t1547 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X485 XThC.Tn[14].t7 XThC.XTB7.Y a_10915_9569# VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X486 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t18 VGND.t928 VGND.t927 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X487 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t26 XA.XIR[8].XIC[8].icell.Ien VGND.t2676 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X488 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1945 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X489 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t24 VGND.t122 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X490 VGND.t1726 XThC.Tn[5].t19 XA.XIR[4].XIC[5].icell.PDM VGND.t1725 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X491 XA.XIR[6].XIC_15.icell.PDM VPWR.t1946 VGND.t1551 VGND.t1550 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X492 VGND.t2012 XThC.XTB4.Y.t4 XThC.Tn[3].t3 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 VPWR.t206 XThC.XTB2.Y XThC.Tn[9].t2 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X494 VGND.t1010 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t1009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X495 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[5].icell.Ien VGND.t1502 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X496 VPWR.t1193 XThR.XTB5.Y XThR.Tn[12].t2 VPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X497 VGND.t463 XThC.Tn[3].t15 XA.XIR[11].XIC[3].icell.PDM VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X498 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1947 VGND.t1553 VGND.t1552 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X499 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t137 VGND.t1325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X500 VGND.t1555 VPWR.t1948 XA.XIR[6].XIC_15.icell.PDM VGND.t1554 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X501 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t24 XA.XIR[11].XIC[3].icell.Ien VGND.t2055 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X502 VGND.t557 XThC.Tn[7].t13 XA.XIR[5].XIC[7].icell.PDM VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X503 VGND.t1557 VPWR.t1949 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1556 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X504 VPWR.t500 XThR.Tn[7].t18 XA.XIR[8].XIC[1].icell.PUM VPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X505 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC_15.icell.Ien VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X506 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X507 VPWR.t131 XThR.XTB7.Y XThR.Tn[14].t2 VPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X508 VPWR.t428 XThR.Tn[6].t21 XA.XIR[7].XIC[0].icell.PUM VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X509 VPWR.t908 VPWR.t906 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X510 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t23 XA.XIR[5].XIC[7].icell.Ien VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X511 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t17 XA.XIR[8].XIC[1].icell.Ien VPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X512 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t18 XA.XIR[7].XIC[0].icell.Ien VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X513 XThR.Tn[8].t5 XThR.XTB1.Y.t4 a_n997_3979# VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X514 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t904 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X515 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t27 VPWR.t1904 VPWR.t1903 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X516 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t19 VPWR.t502 VPWR.t501 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X517 VPWR.t1858 data[2].t0 XThC.XTB7.B VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X518 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t901 VPWR.t903 VPWR.t902 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X519 VGND.t1434 VGND.t1432 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1433 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X520 VPWR.t596 XThR.Tn[0].t22 XA.XIR[1].XIC[12].icell.PUM VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X521 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1950 VGND.t1559 VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X522 VPWR.t1251 XThR.Tn[4].t18 XA.XIR[5].XIC[12].icell.PUM VPWR.t1250 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X523 XThC.Tn[13].t2 XThC.XTB6.Y a_10051_9569# VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X524 XThR.Tn[4].t11 XThR.XTBN.Y a_n1049_6405# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X525 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X526 VGND.t1012 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t1011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X527 XThC.Tn[8].t3 XThC.XTBN.Y.t25 VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X528 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t20 VGND.t667 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X529 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1446 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X530 VGND.t1014 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t1013 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 XA.XIR[3].XIC_15.icell.PDM VPWR.t1951 VGND.t1561 VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X532 VGND.t1016 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t1015 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X533 VGND.t1018 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t1017 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X534 XThC.Tn[8].t10 XThC.XTB1.Y.t4 a_7651_9569# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X535 XThC.Tn[13].t10 XThC.XTBN.Y.t26 VPWR.t11 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X536 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t25 VGND.t542 VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X537 VGND.t465 XThC.Tn[3].t16 XA.XIR[8].XIC[3].icell.PDM VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X538 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t75 VGND.t700 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X539 VGND.t1563 VPWR.t1952 XA.XIR[3].XIC_15.icell.PDM VGND.t1562 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X540 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t244 VGND.t2587 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X541 VGND.t1684 XThC.XTB6.Y XThC.Tn[5].t2 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X542 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t19 VGND.t930 VGND.t929 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X543 VGND.t2152 XThC.Tn[12].t17 XA.XIR[15].XIC[12].icell.PDM VGND.t2151 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X544 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[3].icell.Ien VGND.t2677 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X545 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t20 XA.XIR[3].XIC_15.icell.Ien VGND.t931 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X546 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t17 VGND.t202 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X547 VGND.t2301 XThC.Tn[0].t19 XA.XIR[4].XIC[0].icell.PDM VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X548 XA.XIR[15].XIC[12].icell.PDM VPWR.t1953 XA.XIR[15].XIC[12].icell.Ien VGND.t1564 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X549 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t23 VGND.t1036 VGND.t1035 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X550 VGND.t1020 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t1019 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X551 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t19 XA.XIR[4].XIC[0].icell.Ien VGND.t1503 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X552 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t20 VGND.t1505 VGND.t1504 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X553 VGND.t1492 XThC.Tn[13].t18 XA.XIR[2].XIC[13].icell.PDM VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X554 a_n1049_5611# XThR.XTB6.Y VPWR.t1875 VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X555 XThR.Tn[10].t4 XThR.XTB3.Y.t4 a_n997_2891# VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X556 VGND.t1022 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t1021 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X557 VPWR.t179 XThR.Tn[1].t18 XA.XIR[2].XIC[9].icell.PUM VPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X558 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[13].icell.Ien VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X559 VPWR.t155 XThC.XTBN.Y.t27 XThC.Tn[7].t2 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X560 VPWR.t1018 XThR.Tn[0].t24 XA.XIR[1].XIC[10].icell.PUM VPWR.t1017 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X561 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t17 XA.XIR[2].XIC[9].icell.Ien VPWR.t1790 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X562 VPWR.t1253 XThR.Tn[4].t21 XA.XIR[5].XIC[10].icell.PUM VPWR.t1252 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X563 VPWR.t1641 XThR.XTB2.Y XThR.Tn[9].t2 VPWR.t1640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X564 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X565 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t20 VPWR.t1268 VPWR.t1267 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X566 VGND.t1024 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t1023 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X567 VGND.t1026 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t1025 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X568 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X569 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t6 VPWR.t1722 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X570 VPWR.t350 XThR.Tn[9].t24 XA.XIR[10].XIC[7].icell.PUM VPWR.t349 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X571 XThC.Tn[0].t5 XThC.XTBN.Y.t29 VGND.t175 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X572 VGND.t972 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t971 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X573 VPWR.t1364 XThR.Tn[12].t26 XA.XIR[13].XIC[8].icell.PUM VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X574 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[10].XIC[7].icell.Ien VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X575 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t21 VPWR.t504 VPWR.t503 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X576 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t19 VGND.t204 VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X577 VGND.t974 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X578 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t7 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X579 XThR.Tn[0].t3 XThR.XTB1.Y.t5 VGND.t1277 VGND.t1276 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 VGND.t2492 XThR.XTBN.Y XThR.Tn[5].t6 VGND.t2478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X581 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t222 VGND.t2233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X582 VGND.t976 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X583 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t17 XA.XIR[13].XIC[8].icell.Ien VPWR.t523 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X585 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t25 VPWR.t113 VPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X586 VGND.t2016 XThC.Tn[11].t17 XA.XIR[2].XIC[11].icell.PDM VGND.t2015 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X587 VGND.t978 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t977 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X588 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t23 VPWR.t1081 VPWR.t1080 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X589 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t899 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t900 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X590 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t221 VGND.t2232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X591 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC[11].icell.Ien VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X592 VGND.t2491 XThR.XTBN.Y XThR.Tn[4].t7 VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X593 VPWR.t898 VPWR.t896 XA.XIR[11].XIC_15.icell.PUM VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X594 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t893 VPWR.t895 VPWR.t894 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X595 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t20 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X596 XA.XIR[11].XIC_15.icell.PUM VPWR.t891 XA.XIR[11].XIC_15.icell.Ien VPWR.t892 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X597 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t7 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X598 VGND.t980 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X599 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t66 VGND.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X600 VGND.t172 XThC.Tn[2].t17 XA.XIR[2].XIC[2].icell.PDM VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X601 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t25 VGND.t410 VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X602 VGND.t982 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X603 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t25 VPWR.t1511 VPWR.t1510 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X604 VGND.t984 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t983 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X605 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t22 XA.XIR[2].XIC[2].icell.Ien VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X606 VPWR.t1020 XThR.Tn[0].t25 XA.XIR[1].XIC[5].icell.PUM VPWR.t1019 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X607 VGND.t2520 XThC.Tn[9].t18 XA.XIR[10].XIC[9].icell.PDM VGND.t2519 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X608 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t22 XA.XIR[7].XIC[8].icell.Ien VGND.t668 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X609 VGND.t986 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t985 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X610 VGND.t177 XThC.XTBN.Y.t31 a_8739_9569# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X611 VPWR.t1255 XThR.Tn[4].t22 XA.XIR[5].XIC[5].icell.PUM VPWR.t1254 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X612 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t26 XA.XIR[10].XIC[9].icell.Ien VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X613 VPWR.t352 XThR.Tn[9].t26 XA.XIR[10].XIC[11].icell.PUM VPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X614 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[10].XIC[11].icell.Ien VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X615 VGND.t988 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t987 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X616 VGND.t990 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t989 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t27 VPWR.t103 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X618 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t13 VGND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X619 a_9827_9569# XThC.XTBN.Y.t32 VGND.t179 VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X620 VGND.t992 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t991 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t192 VGND.t1901 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X622 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t27 XA.XIR[9].XIC_15.icell.Ien VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X623 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t78 VGND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X624 VPWR.t354 XThR.Tn[9].t28 XA.XIR[10].XIC[2].icell.PUM VPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X625 VPWR.t1601 XThR.Tn[12].t27 XA.XIR[13].XIC[3].icell.PUM VPWR.t1600 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X626 VGND.t2657 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X627 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[10].XIC[2].icell.Ien VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X628 VPWR.t887 VPWR.t885 XA.XIR[8].XIC_15.icell.PUM VPWR.t886 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X629 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t23 VPWR.t506 VPWR.t505 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X630 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t21 VGND.t208 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X631 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t20 XA.XIR[5].XIC[14].icell.Ien VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X632 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t26 VGND.t1096 VGND.t1095 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X633 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t38 VGND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X634 XThR.XTB7.A data[5].t1 VPWR.t1197 VPWR.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X635 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t17 XA.XIR[13].XIC[3].icell.Ien VPWR.t396 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X636 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t28 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X637 VGND.t326 XThC.Tn[6].t18 XA.XIR[2].XIC[6].icell.PDM VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X638 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t23 VGND.t1507 VGND.t1506 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X639 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t24 VPWR.t283 VPWR.t282 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X640 XA.XIR[8].XIC_15.icell.PUM VPWR.t883 XA.XIR[8].XIC_15.icell.Ien VPWR.t884 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X641 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t24 VGND.t1169 VGND.t1168 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X642 VPWR.t1223 VGND.t2691 XA.XIR[0].XIC[4].icell.PUM VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X643 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1954 VGND.t1566 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X644 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t25 VPWR.t1083 VPWR.t1082 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X645 VPWR.t581 XThR.Tn[3].t21 XA.XIR[4].XIC[12].icell.PUM VPWR.t580 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X646 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t29 VPWR.t1906 VPWR.t1905 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X647 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t23 XA.XIR[2].XIC[6].icell.Ien VGND.t1616 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X648 VGND.t157 XThC.Tn[10].t19 XA.XIR[14].XIC[10].icell.PDM VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X649 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[0].XIC[4].icell.Ien VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X650 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[4].XIC[12].icell.Ien VPWR.t1572 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X651 VGND.t1568 VPWR.t1955 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X652 VPWR.t430 XThR.Tn[6].t22 XA.XIR[7].XIC[13].icell.PUM VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X653 VGND.t227 XThC.XTBN.A XThC.XTBN.Y.t3 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 VPWR.t1135 XThR.XTB7.B XThR.XTB1.Y.t2 VPWR.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X655 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[10].icell.Ien VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X656 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t27 VPWR.t1022 VPWR.t1021 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X657 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1956 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X658 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[7].XIC[13].icell.Ien VPWR.t1247 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X659 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t24 VPWR.t1257 VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X660 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t10 VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X661 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t26 VGND.t1171 VGND.t1170 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X662 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t29 VGND.t413 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X663 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t153 VGND.t1619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X664 VGND.t941 XThC.Tn[1].t18 XA.XIR[14].XIC[1].icell.PDM VGND.t940 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X665 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t109 VGND.t1115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X666 VGND.t370 XThC.Tn[4].t19 XA.XIR[10].XIC[4].icell.PDM VGND.t369 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X667 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[3].icell.Ien VGND.t669 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X668 VGND.t1571 VPWR.t1957 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X669 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[1].icell.Ien VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X670 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[4].icell.Ien VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X671 XThC.Tn[7].t1 XThC.XTBN.Y.t33 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X672 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X673 VGND.t1224 XThR.XTB7.B a_n1335_7243# VGND.t1223 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X674 VGND.t1494 XThC.Tn[13].t20 XA.XIR[1].XIC[13].icell.PDM VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X675 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t22 VGND.t933 VGND.t932 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X676 VGND.t1752 XThC.Tn[14].t21 XA.XIR[4].XIC[14].icell.PDM VGND.t1751 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X677 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t30 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X678 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t185 VGND.t1820 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X679 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t22 XA.XIR[1].XIC[13].icell.Ien VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X680 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t15 VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XThC.Tn[11].t3 XThC.XTB4.Y.t6 VPWR.t1009 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 VGND.t2154 XThC.Tn[12].t19 XA.XIR[11].XIC[12].icell.PDM VGND.t2153 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X683 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t19 XA.XIR[1].XIC[9].icell.Ien VPWR.t1791 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X684 VPWR.t583 XThR.Tn[3].t23 XA.XIR[4].XIC[10].icell.PUM VPWR.t582 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X685 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t25 XA.XIR[4].XIC[14].icell.Ien VGND.t1508 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X686 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t22 VGND.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X687 VPWR.t1221 VGND.t2692 XA.XIR[0].XIC[0].icell.PUM VPWR.t1220 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X688 a_n997_1803# XThR.XTBN.Y VGND.t2489 VGND.t2488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t23 VPWR.t1692 VPWR.t1691 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X690 XThR.Tn[3].t6 XThR.XTBN.Y a_n1049_6699# VPWR.t1774 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X691 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t20 XA.XIR[4].XIC[10].icell.Ien VPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X692 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[12].icell.Ien VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X693 VGND.t2487 XThR.XTBN.Y XThR.Tn[3].t10 VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X694 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t20 XA.XIR[0].XIC[0].icell.Ien VPWR.t1664 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X695 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t26 VPWR.t1701 VPWR.t1700 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X696 VGND.t994 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t993 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X697 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t28 VPWR.t1024 VPWR.t1023 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X698 XThC.Tn[2].t6 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X699 XThR.Tn[11].t6 XThR.XTB4.Y.t5 VPWR.t1619 VPWR.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 VPWR.t205 XThC.XTB2.Y a_3773_9615# VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X701 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t1155 VPWR.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t18 XA.XIR[12].XIC[8].icell.Ien VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X703 VGND.t996 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t995 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X704 VGND.t2018 XThC.Tn[11].t19 XA.XIR[1].XIC[11].icell.PDM VGND.t2017 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X705 VGND.t1431 VGND.t1429 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X706 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t28 VPWR.t1603 VPWR.t1602 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X707 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t160 VGND.t1641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X708 VPWR.t432 XThR.Tn[6].t23 XA.XIR[7].XIC[6].icell.PUM VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X709 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC[11].icell.Ien VGND.t2349 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X710 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t47 VGND.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X711 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t25 VGND.t671 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X712 VPWR.t285 XThR.Tn[5].t25 XA.XIR[6].XIC[7].icell.PUM VPWR.t284 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X713 VPWR.t454 XThC.XTB6.A a_5949_10571# VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X714 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[7].XIC[6].icell.Ien VPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X715 VPWR.t1908 XThR.Tn[8].t30 XA.XIR[9].XIC[8].icell.PUM VPWR.t1907 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X716 VGND.t2156 XThC.Tn[12].t20 XA.XIR[8].XIC[12].icell.PDM VGND.t2155 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X717 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t15 XA.XIR[6].XIC[7].icell.Ien VPWR.t476 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X718 VGND.t1905 XThR.XTB3.Y.t5 XThR.Tn[2].t2 VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X719 VGND.t1126 XThC.Tn[2].t19 XA.XIR[1].XIC[2].icell.PDM VGND.t1125 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X720 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[9].XIC[8].icell.Ien VPWR.t525 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X721 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t31 XA.XIR[8].XIC[12].icell.Ien VGND.t2678 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X722 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t63 VGND.t550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X723 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t24 VPWR.t1101 VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X724 XThC.XTBN.Y.t1 XThC.XTBN.A VPWR.t198 VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X725 VGND.t998 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X726 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t27 VGND.t484 VGND.t483 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X727 VGND.t490 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X728 XThR.Tn[8].t6 XThR.XTB1.Y.t7 a_n997_3979# VGND.t1278 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X729 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t25 XA.XIR[1].XIC[2].icell.Ien VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X730 VGND.t492 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X731 VGND.t494 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X732 VPWR.t585 XThR.Tn[3].t24 XA.XIR[4].XIC[5].icell.PUM VPWR.t584 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X733 VGND.t180 XThC.XTBN.Y.t35 a_9827_9569# VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X734 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t20 XA.XIR[4].XIC[5].icell.Ien VPWR.t1329 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X735 VPWR.t54 XThC.XTB7.Y XThC.Tn[14].t3 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X736 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t27 VPWR.t1703 VPWR.t1702 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X737 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t25 VGND.t1196 VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X738 XThR.Tn[4].t10 XThR.XTBN.Y a_n1049_6405# VPWR.t1774 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X739 VGND.t496 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X740 VGND.t498 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X741 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t26 VGND.t318 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X742 VPWR.t1620 XThR.XTB4.Y.t6 a_n1049_6699# VPWR.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X743 VGND.t500 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X744 VGND.t697 XThC.Tn[8].t20 XA.XIR[7].XIC[8].icell.PDM VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X745 VPWR.t882 VPWR.t880 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t881 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X746 VGND.t2522 XThC.Tn[9].t20 XA.XIR[6].XIC[9].icell.PDM VGND.t2521 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X747 VGND.t502 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X748 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t104 VGND.t1109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X749 VPWR.t287 XThR.Tn[5].t27 XA.XIR[6].XIC[11].icell.PUM VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X750 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t26 XA.XIR[6].XIC[9].icell.Ien VGND.t1197 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X751 VPWR.t1270 XThR.Tn[2].t24 XA.XIR[3].XIC[7].icell.PUM VPWR.t1269 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X752 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t20 XA.XIR[6].XIC[11].icell.Ien VPWR.t1452 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X753 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[3].XIC[7].icell.Ien VPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X754 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t18 XA.XIR[12].XIC[3].icell.Ien VPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X755 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t25 VGND.t728 VGND.t727 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X756 VGND.t504 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X757 VGND.t328 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t327 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X758 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t173 VGND.t1802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X759 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t27 VPWR.t1103 VPWR.t1102 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X760 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t183 VGND.t1816 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X761 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t26 VPWR.t548 VPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X762 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t29 VPWR.t1605 VPWR.t1604 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X763 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t26 XA.XIR[1].XIC[6].icell.Ien VGND.t2351 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X764 VGND.t559 XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.PDM VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X765 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t26 VPWR.t508 VPWR.t507 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X766 VPWR.t1105 XThR.Tn[6].t28 XA.XIR[7].XIC[1].icell.PUM VPWR.t1104 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X767 VPWR.t1551 XThR.Tn[5].t28 XA.XIR[6].XIC[2].icell.PUM VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X768 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t1487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X769 VGND.t506 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X770 VPWR.t1773 XThR.XTBN.Y XThR.Tn[8].t11 VPWR.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X771 VPWR.t1026 XThR.Tn[0].t29 XA.XIR[1].XIC[14].icell.PUM VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X772 XThR.Tn[10].t0 XThR.XTB3.Y.t6 a_n997_2891# VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X773 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t28 XA.XIR[4].XIC[7].icell.Ien VGND.t2407 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X774 VPWR.t1705 XThR.Tn[4].t29 XA.XIR[5].XIC[14].icell.PUM VPWR.t1704 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X775 VPWR.t1910 XThR.Tn[8].t32 XA.XIR[9].XIC[3].icell.PUM VPWR.t1909 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X776 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[7].XIC[1].icell.Ien VPWR.t589 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X777 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t20 XA.XIR[6].XIC[2].icell.Ien VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X778 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t1351 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X779 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t29 VPWR.t1107 VPWR.t1106 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X780 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t19 XA.XIR[9].XIC[3].icell.Ien VPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X781 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t51 VGND.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X782 VGND.t508 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X783 VGND.t1428 VGND.t1426 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t28 VGND.t486 VGND.t485 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X785 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t25 VGND.t1618 VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X786 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1959 VGND.t1574 VGND.t1573 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X787 VGND.t510 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X788 VPWR.t453 XThC.XTB6.A XThC.XTB2.Y VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X789 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t202 VGND.t1934 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X790 VGND.t512 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X791 VGND.t1576 VPWR.t1960 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t1575 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X792 XThR.XTB3.Y.t2 XThR.XTB7.A VPWR.t1460 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X793 VGND.t347 XThC.Tn[9].t21 XA.XIR[3].XIC[9].icell.PDM VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X794 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t119 VGND.t1174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X795 VPWR.t1272 XThR.Tn[2].t26 XA.XIR[3].XIC[11].icell.PUM VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X796 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t27 XA.XIR[3].XIC[9].icell.Ien VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X797 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1961 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1577 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X798 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t30 VGND.t1199 VGND.t1198 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X799 XA.XIR[2].XIC_15.icell.PDM VPWR.t1962 VGND.t1579 VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X800 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t29 VGND.t2127 VGND.t2126 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X801 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X802 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[3].XIC[11].icell.Ien VPWR.t1453 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X803 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1963 VGND.t1581 VGND.t1580 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X804 VGND.t514 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X805 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t8 VGND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X806 VGND.t467 XThC.Tn[3].t20 XA.XIR[7].XIC[3].icell.PDM VGND.t466 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X807 VGND.t1583 VPWR.t1964 XA.XIR[2].XIC_15.icell.PDM VGND.t1582 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X808 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t28 VPWR.t550 VPWR.t549 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X809 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t1585 VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X810 VGND.t372 XThC.Tn[4].t20 XA.XIR[6].XIC[4].icell.PDM VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X811 XThR.Tn[0].t11 XThR.XTBN.Y VGND.t2486 VGND.t2429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X812 VPWR.t1192 XThR.XTB5.Y a_n1049_6405# VPWR.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X813 VGND.t516 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X814 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t217 VGND.t2228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X815 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t31 XA.XIR[6].XIC[4].icell.Ien VGND.t1200 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X816 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t27 XA.XIR[2].XIC_15.icell.Ien VGND.t1621 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X817 XThC.Tn[10].t9 XThC.XTB3.Y.t4 VPWR.t1042 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X818 VPWR.t1274 XThR.Tn[2].t28 XA.XIR[3].XIC[2].icell.PUM VPWR.t1273 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X819 VPWR.t1771 XThR.XTBN.Y XThR.Tn[10].t8 VPWR.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X820 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t1310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X821 VPWR.t159 XThC.XTBN.Y.t36 XThC.Tn[13].t9 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X822 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[3].XIC[2].icell.Ien VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X823 a_3773_9615# XThC.XTB2.Y VPWR.t204 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 XThC.Tn[5].t1 XThC.XTB6.Y VGND.t1683 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t62 VGND.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X826 XThC.Tn[2].t0 XThC.XTB3.Y.t5 VGND.t190 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X827 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t29 VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X828 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1966 VGND.t1587 VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X829 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t144 VGND.t1488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X830 VPWR.t1085 XThR.Tn[13].t27 XA.XIR[14].XIC[4].icell.PUM VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X831 VGND.t2485 XThR.XTBN.Y a_n997_3755# VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 VGND.t1589 VPWR.t1967 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t1588 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X833 VPWR.t1219 VGND.t2693 XA.XIR[0].XIC[13].icell.PUM VPWR.t1218 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X834 VPWR.t879 VPWR.t877 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t878 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X835 VPWR.t1853 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t1852 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X836 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t21 XA.XIR[0].XIC[13].icell.Ien VPWR.t1248 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X837 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t21 XA.XIR[14].XIC[4].icell.Ien VPWR.t329 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X838 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1968 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t834 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X839 VGND.t1687 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t1686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X840 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t29 VGND.t1623 VGND.t1622 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X841 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t875 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t876 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X842 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t28 VPWR.t468 VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X843 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t121 VGND.t1185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t30 VPWR.t1028 VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X845 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t4 VGND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X846 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t2243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X847 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t216 VGND.t2057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 VGND.t374 XThC.Tn[4].t22 XA.XIR[3].XIC[4].icell.PDM VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X849 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t872 VPWR.t874 VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X850 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t1 VGND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t196 VGND.t1908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X852 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t30 XA.XIR[3].XIC[4].icell.Ien VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X853 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t157 VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X854 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t27 XA.XIR[7].XIC[12].icell.Ien VGND.t672 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X855 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t30 VPWR.t356 VPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X856 a_5155_9615# XThC.XTB5.Y VPWR.t416 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X857 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t1052 VPWR.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X858 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t29 VGND.t546 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X859 VGND.t1730 XThC.Tn[5].t21 XA.XIR[15].XIC[5].icell.PDM VGND.t1729 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X860 XA.XIR[15].XIC[5].icell.PDM VPWR.t1969 XA.XIR[15].XIC[5].icell.Ien VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X861 VPWR.t1087 XThR.Tn[13].t28 XA.XIR[14].XIC[0].icell.PUM VPWR.t1086 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X862 XThC.Tn[8].t7 XThC.XTB1.Y.t7 VPWR.t1855 VPWR.t1854 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X863 VGND.t1323 XThR.XTB5.Y XThR.Tn[4].t3 VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X864 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t7 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X865 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t21 XA.XIR[14].XIC[0].icell.Ien VPWR.t1665 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X866 XThR.XTB5.Y XThR.XTB5.A VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X867 VPWR.t871 VPWR.t869 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t870 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X868 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t30 VPWR.t470 VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X869 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t867 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t868 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X870 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[9].icell.Ien VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X871 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X872 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t838 VPWR.t840 VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X873 VPWR.t420 XThR.Tn[11].t29 XA.XIR[12].XIC[12].icell.PUM VPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X874 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[5].XIC[8].icell.Ien VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X875 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t32 VPWR.t358 VPWR.t357 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X876 VGND.t1689 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t1688 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X877 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t149 VGND.t1510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X878 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t30 VPWR.t1553 VPWR.t1552 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X879 VGND.t1691 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t1690 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X880 VPWR.t1217 VGND.t2694 XA.XIR[0].XIC[6].icell.PUM VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X881 VGND.t1693 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t1692 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X882 VPWR.t554 XThR.Tn[3].t31 XA.XIR[4].XIC[14].icell.PUM VPWR.t553 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X883 XThC.Tn[14].t6 XThC.XTB7.Y a_10915_9569# VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X884 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[0].XIC[6].icell.Ien VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X885 VPWR.t866 VPWR.t864 XA.XIR[7].XIC_15.icell.PUM VPWR.t865 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X886 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X887 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[4].XIC[14].icell.Ien VPWR.t1500 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X888 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t31 VPWR.t1030 VPWR.t1029 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X889 a_n997_1803# XThR.XTBN.Y VGND.t2484 VGND.t2483 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X890 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t33 VPWR.t360 VPWR.t359 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X891 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t30 VPWR.t1707 VPWR.t1706 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X892 XA.XIR[7].XIC_15.icell.PUM VPWR.t862 XA.XIR[7].XIC_15.icell.Ien VPWR.t863 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X893 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t31 VGND.t548 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X894 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t7 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X895 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t238 VGND.t2410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X896 VGND.t2303 XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.PDM VGND.t2302 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X897 VGND.t1695 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t1694 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X898 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t30 VGND.t2207 VGND.t2206 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X899 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t30 VGND.t488 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X900 VPWR.t182 XThC.XTB5.A XThC.XTB1.Y.t0 VPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X901 XA.XIR[15].XIC[0].icell.PDM VPWR.t1970 XA.XIR[15].XIC[0].icell.Ien VGND.t836 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X902 VGND.t1496 XThC.Tn[13].t22 XA.XIR[13].XIC[13].icell.PDM VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X903 XA.XIR[0].XIC[8].icell.PDM VGND.t1423 VGND.t1425 VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X904 VGND.t1697 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t1696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X905 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[13].icell.Ien VGND.t1172 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X906 VPWR.t1607 XThR.Tn[12].t31 XA.XIR[13].XIC[9].icell.PUM VPWR.t1606 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X907 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1971 VGND.t838 VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X908 VPWR.t422 XThR.Tn[11].t31 XA.XIR[12].XIC[10].icell.PUM VPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X909 VGND.t1699 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t1698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X910 VGND.t840 VPWR.t1972 XA.XIR[1].XIC_15.icell.PDM VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X911 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t22 XA.XIR[13].XIC[9].icell.Ien VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X912 VGND.t2626 XThC.Tn[8].t22 XA.XIR[0].XIC[8].icell.PDM VGND.t2625 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X913 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t27 XA.XIR[1].XIC_15.icell.Ien VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X914 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t115 VGND.t1138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X915 VGND.t842 VPWR.t1973 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X916 VGND.t191 XThC.XTB3.Y.t6 XThC.Tn[2].t1 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X917 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t1 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X918 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t32 XA.XIR[0].XIC[8].icell.Ien VGND.t1097 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X919 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t598 VPWR.t597 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X920 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t34 XA.XIR[9].XIC[4].icell.Ien VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X921 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1974 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X922 a_n1319_6405# XThR.XTB5.A VPWR.t35 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X923 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[5].XIC[3].icell.Ien VPWR.t381 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X924 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t35 VGND.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X925 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t1857 VPWR.t1856 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X926 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t31 VPWR.t1555 VPWR.t1554 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X927 VGND.t1701 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t1700 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X928 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t35 VGND.t360 VGND.t359 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X929 VPWR.t1215 VGND.t2695 XA.XIR[0].XIC[1].icell.PUM VPWR.t1214 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X930 VGND.t1703 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t1702 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X931 XThR.Tn[12].t10 XThR.XTBN.Y VPWR.t1769 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X932 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t1514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X933 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t74 VGND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X934 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t32 VGND.t2209 VGND.t2208 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X935 VGND.t159 XThC.Tn[10].t21 XA.XIR[10].XIC[10].icell.PDM VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X936 XThC.Tn[11].t11 XThC.XTBN.Y.t39 VPWR.t163 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X937 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[0].XIC[1].icell.Ien VPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X938 VGND.t1658 data[4].t2 XThR.XTB5.A VGND.t1657 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X939 XThR.XTBN.Y XThR.XTBN.A VGND.t711 VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X940 VGND.t2020 XThC.Tn[11].t22 XA.XIR[13].XIC[11].icell.PDM VGND.t2019 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X941 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1975 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X942 VGND.t2245 data[3].t0 XThC.XTBN.A VGND.t2244 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X943 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[10].icell.Ien VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X944 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t33 VPWR.t1032 VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X945 VGND.t1705 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t1704 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X946 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t860 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X947 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[11].icell.Ien VGND.t1042 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X948 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t36 VGND.t362 VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X949 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t7 VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X950 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t19 VGND.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X951 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t857 VPWR.t859 VPWR.t858 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X952 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t33 VGND.t2211 VGND.t2210 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X953 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t58 VGND.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 a_n997_2667# XThR.XTBN.Y VGND.t2482 VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 VGND.t610 XThC.Tn[1].t21 XA.XIR[10].XIC[1].icell.PDM VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X956 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t139 VGND.t1468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X957 VGND.t1128 XThC.Tn[2].t22 XA.XIR[13].XIC[2].icell.PDM VGND.t1127 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X958 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t32 XA.XIR[10].XIC[1].icell.Ien VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X959 VPWR.t856 VPWR.t854 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t855 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X960 XA.XIR[0].XIC[3].icell.PDM VGND.t1420 VGND.t1422 VGND.t1421 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X961 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[2].icell.Ien VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X962 VPWR.t424 XThR.Tn[11].t32 XA.XIR[12].XIC[5].icell.PUM VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X963 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t852 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X964 VGND.t446 XThC.Tn[3].t22 XA.XIR[0].XIC[3].icell.PDM VGND.t445 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X965 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t32 VGND.t2024 VGND.t2023 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X966 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t204 VGND.t1967 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X967 XThC.Tn[4].t6 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X968 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t34 XA.XIR[0].XIC[3].icell.Ien VGND.t2647 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X969 VGND.t2158 XThC.Tn[12].t21 XA.XIR[7].XIC[12].icell.PDM VGND.t2157 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X970 VPWR.t1767 XThR.XTBN.Y XThR.Tn[8].t10 VPWR.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X971 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t9 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X972 VGND.t1707 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t1706 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X973 VPWR.t415 XThC.XTB5.Y XThC.Tn[12].t1 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X974 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t33 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X975 VGND.t1709 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t1708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X976 VGND.t1732 XThC.Tn[5].t22 XA.XIR[11].XIC[5].icell.PDM VGND.t1731 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X977 VGND.t2481 XThR.XTBN.Y XThR.Tn[1].t11 VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X978 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t34 VGND.t2213 VGND.t2212 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X979 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t33 VGND.t734 VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X980 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[5].icell.Ien VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X981 VGND.t330 XThC.Tn[6].t22 XA.XIR[13].XIC[6].icell.PDM VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X982 VGND.t1711 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t1710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X983 VPWR.t434 XThR.Tn[14].t32 XA.XIR[15].XIC[12].icell.PUM VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X984 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t137 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X985 a_9827_9569# XThC.XTBN.Y.t41 VGND.t181 VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X986 VPWR.t600 XThR.Tn[13].t33 XA.XIR[14].XIC[13].icell.PUM VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X987 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t34 XA.XIR[13].XIC[6].icell.Ien VGND.t1044 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X988 XThR.Tn[9].t9 XThR.XTBN.Y VPWR.t1765 VPWR.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X989 VPWR.t851 VPWR.t849 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t850 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X990 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[15].XIC[12].icell.Ien VPWR.t1573 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X991 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[14].XIC[13].icell.Ien VPWR.t1249 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X992 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t1308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X993 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t83 VGND.t915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X994 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t847 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t848 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X995 XThC.Tn[1].t6 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X996 VPWR.t1694 XThR.Tn[1].t28 XA.XIR[2].XIC[7].icell.PUM VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X997 XA.XIR[15].XIC[12].icell.Ien VPWR.t844 VPWR.t846 VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X998 XThR.Tn[0].t10 XThR.XTBN.Y VGND.t2480 VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 VPWR.t1845 XThR.Tn[0].t35 XA.XIR[1].XIC[8].icell.PUM VPWR.t1844 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1000 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t33 VPWR.t436 VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1001 XThC.Tn[13].t1 XThC.XTB6.Y a_10051_9569# VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1002 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t841 VPWR.t843 VPWR.t842 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1003 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t18 XA.XIR[2].XIC[7].icell.Ien VPWR.t478 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1004 VPWR.t1709 XThR.Tn[4].t31 XA.XIR[5].XIC[8].icell.PUM VPWR.t1708 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1005 VPWR.t1764 XThR.XTBN.Y XThR.Tn[10].t7 VPWR.t1763 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1006 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t30 VPWR.t1276 VPWR.t1275 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1007 VGND.t1713 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t1712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1008 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t28 VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1009 VGND.t1763 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t1762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1010 VPWR.t53 XThC.XTB7.Y a_6243_9615# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1011 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t18 VGND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1012 VGND.t1734 XThC.Tn[5].t23 XA.XIR[8].XIC[5].icell.PDM VGND.t1733 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1013 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t34 VGND.t524 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1014 VGND.t1498 XThC.Tn[13].t24 XA.XIR[12].XIC[13].icell.PDM VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1015 VGND.t2047 XThC.Tn[14].t23 XA.XIR[15].XIC[14].icell.PDM VGND.t2046 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1016 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t33 XA.XIR[8].XIC[5].icell.Ien VGND.t2679 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1017 VGND.t182 XThC.XTBN.Y.t43 a_8963_9569# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1018 VGND.t1765 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t1764 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1019 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t35 XA.XIR[12].XIC[13].icell.Ien VGND.t2214 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1020 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t34 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1021 VPWR.t438 XThR.Tn[14].t35 XA.XIR[15].XIC[10].icell.PUM VPWR.t437 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1022 VPWR.t1157 XThR.XTB1.Y.t8 XThR.Tn[8].t7 VPWR.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1023 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t29 VGND.t2354 VGND.t2353 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1024 XA.XIR[15].XIC[14].icell.PDM VPWR.t1976 XA.XIR[15].XIC[14].icell.Ien VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1025 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t23 XA.XIR[12].XIC[9].icell.Ien VPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1026 VGND.t1767 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t1766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1027 VGND.t1769 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t1768 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1028 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t156 VGND.t1637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1029 VGND.t2305 XThC.Tn[0].t23 XA.XIR[11].XIC[0].icell.PDM VGND.t2304 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1030 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t34 VGND.t1294 VGND.t1293 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1031 VGND.t349 XThC.Tn[9].t24 XA.XIR[2].XIC[9].icell.PDM VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1032 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t22 XA.XIR[15].XIC[10].icell.Ien VPWR.t1302 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1033 XThR.XTBN.A data[7].t0 VPWR.t1097 VPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1034 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t36 VPWR.t1410 VPWR.t1409 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1035 VPWR.t832 VPWR.t830 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1036 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t49 VGND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1037 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[0].icell.Ien VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1038 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1039 VPWR.t1541 XThR.Tn[1].t30 XA.XIR[2].XIC[11].icell.PUM VPWR.t1540 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1040 XA.XIR[15].XIC[10].icell.Ien VPWR.t835 VPWR.t837 VPWR.t836 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1041 VGND.t1500 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t1499 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1042 VPWR.t1639 XThR.XTB2.Y a_n1049_7787# VPWR.t1638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1043 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t31 XA.XIR[2].XIC[9].icell.Ien VGND.t1624 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1044 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t833 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t834 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1045 VPWR.t1169 XThR.Tn[8].t35 XA.XIR[9].XIC[9].icell.PUM VPWR.t1168 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1046 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t23 XA.XIR[2].XIC[11].icell.Ien VPWR.t1297 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1047 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t827 VPWR.t829 VPWR.t828 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1048 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t32 VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[9].XIC[9].icell.Ien VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1050 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t106 VGND.t1111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1051 VGND.t1771 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t1770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1052 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t5 VPWR.t1762 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1053 VPWR.t1543 XThR.Tn[1].t31 XA.XIR[2].XIC[2].icell.PUM VPWR.t1542 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1054 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t194 VGND.t1903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1055 XThC.Tn[8].t6 XThC.XTB1.Y.t10 VPWR.t402 VPWR.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1056 VPWR.t1847 XThR.Tn[0].t36 XA.XIR[1].XIC[3].icell.PUM VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1057 VGND.t1645 XThC.Tn[11].t24 XA.XIR[12].XIC[11].icell.PDM VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1058 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t23 XA.XIR[2].XIC[2].icell.Ien VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1059 VPWR.t1711 XThR.Tn[4].t32 XA.XIR[5].XIC[3].icell.PUM VPWR.t1710 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1060 VPWR.t602 XThR.Tn[13].t35 XA.XIR[14].XIC[6].icell.PUM VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1061 VGND.t1419 VGND.t1417 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1062 VPWR.t826 VPWR.t824 XA.XIR[0].XIC_15.icell.PUM VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1063 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t37 XA.XIR[12].XIC[11].icell.Ien VGND.t1949 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1064 XThR.Tn[0].t0 XThR.XTB1.Y.t9 VGND.t457 VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1065 XA.XIR[0].XIC_15.icell.PUM VPWR.t822 XA.XIR[0].XIC_15.icell.Ien VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1066 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t33 VPWR.t29 VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1067 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t23 XA.XIR[14].XIC[6].icell.Ien VPWR.t297 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1068 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t32 VGND.t2129 VGND.t2128 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1069 VGND.t1773 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t1772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1070 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t29 VGND.t676 VGND.t675 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1071 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t36 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1072 VPWR.t1054 XThR.XTB3.Y.t8 XThR.Tn[10].t1 VPWR.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1977 VGND.t847 VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1074 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t37 VPWR.t1849 VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1075 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t1296 VGND.t1295 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1076 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t249 VGND.t2646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1077 VPWR.t203 XThC.XTB2.Y a_3773_9615# VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1078 VGND.t2479 XThR.XTBN.Y XThR.Tn[4].t6 VGND.t2478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1079 VGND.t2307 XThC.Tn[0].t24 XA.XIR[8].XIC[0].icell.PDM VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1080 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t56 VGND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1081 VGND.t1661 XThC.Tn[10].t23 XA.XIR[6].XIC[10].icell.PDM VGND.t1660 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1082 VGND.t1130 XThC.Tn[2].t24 XA.XIR[12].XIC[2].icell.PDM VGND.t1129 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1083 VGND.t849 VPWR.t1978 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1084 VGND.t1647 XThC.Tn[11].t25 XA.XIR[9].XIC[11].icell.PDM VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1085 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[10].icell.Ien VGND.t2025 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1086 VPWR.t1000 XThC.XTBN.Y.t44 XThC.Tn[9].t11 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1087 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t37 XA.XIR[8].XIC[0].icell.Ien VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1088 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t38 XA.XIR[12].XIC[2].icell.Ien VGND.t1950 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1089 VGND.t1074 XThC.XTBN.Y.t45 XThC.Tn[5].t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1090 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t33 VGND.t2131 VGND.t2130 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1091 VPWR.t442 XThR.Tn[14].t37 XA.XIR[15].XIC[5].icell.PUM VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1092 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t32 VGND.t2124 VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1093 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t108 VGND.t1113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1094 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t92 VGND.t1049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1095 VGND.t2477 XThR.XTBN.Y a_n997_1579# VGND.t2460 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1096 VGND.t376 XThC.Tn[4].t23 XA.XIR[2].XIC[4].icell.PDM VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1097 VGND.t612 XThC.Tn[1].t22 XA.XIR[6].XIC[1].icell.PDM VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1098 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t36 VGND.t1046 VGND.t1045 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1099 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[15].XIC[5].icell.Ien VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1100 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t38 VGND.t1299 VGND.t1298 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1101 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t250 VGND.t2658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1102 VGND.t1775 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t1774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1103 VGND.t1777 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t1776 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1104 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t8 VPWR.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1105 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[1].icell.Ien VGND.t2026 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1106 XA.XIR[15].XIC[5].icell.Ien VPWR.t819 VPWR.t821 VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1107 VGND.t1132 XThC.Tn[2].t25 XA.XIR[9].XIC[2].icell.PDM VGND.t1131 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1108 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[4].icell.Ien VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1109 VGND.t2628 XThC.Tn[8].t23 XA.XIR[14].XIC[8].icell.PDM VGND.t2627 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1110 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t38 XA.XIR[14].XIC[8].icell.Ien VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1111 XThC.Tn[12].t6 XThC.XTB5.Y a_9827_9569# VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 XThR.XTB6.A data[5].t2 VPWR.t275 VPWR.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1113 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t52 VGND.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1114 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1115 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t35 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1116 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t7 VPWR.t1760 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1117 VGND.t1779 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t1778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1118 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t61 VGND.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1119 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t206 VGND.t2005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1120 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t39 VGND.t527 VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1121 VGND.t1663 XThC.Tn[10].t24 XA.XIR[3].XIC[10].icell.PDM VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1122 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t93 VGND.t1050 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1123 VGND.t332 XThC.Tn[6].t24 XA.XIR[12].XIC[6].icell.PDM VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1124 VPWR.t1141 XThR.Tn[13].t37 XA.XIR[14].XIC[1].icell.PUM VPWR.t1140 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1125 VPWR.t315 XThR.Tn[9].t37 XA.XIR[10].XIC[4].icell.PUM VPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1126 VGND.t1161 XThC.Tn[7].t19 XA.XIR[15].XIC[7].icell.PDM VGND.t1160 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1127 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t39 XA.XIR[12].XIC[6].icell.Ien VGND.t1951 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1128 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t32 XA.XIR[3].XIC[10].icell.Ien VGND.t2034 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1129 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t23 XA.XIR[14].XIC[1].icell.Ien VPWR.t488 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1130 VPWR.t560 XThR.Tn[11].t36 XA.XIR[12].XIC[14].icell.PUM VPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1131 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t24 XA.XIR[10].XIC[4].icell.Ien VPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1132 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t817 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1133 XA.XIR[15].XIC[7].icell.PDM VPWR.t1979 XA.XIR[15].XIC[7].icell.Ien VGND.t850 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1134 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t36 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1135 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t40 VPWR.t444 VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1136 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1137 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t814 VPWR.t816 VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1138 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t39 VGND.t1301 VGND.t1300 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1139 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t57 VGND.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1140 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t103 VGND.t1108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1141 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t102 VGND.t1099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1142 VGND.t614 XThC.Tn[1].t24 XA.XIR[3].XIC[1].icell.PDM VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1143 VPWR.t1463 XThR.Tn[3].t33 XA.XIR[4].XIC[8].icell.PUM VPWR.t1462 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1144 a_6243_9615# XThC.XTB7.Y VPWR.t52 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t20 XA.XIR[1].XIC[7].icell.Ien VPWR.t1076 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1146 VGND.t1416 VGND.t1414 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1147 VGND.t334 XThC.Tn[6].t25 XA.XIR[9].XIC[6].icell.PDM VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1148 XThC.Tn[10].t8 XThC.XTBN.Y.t47 VPWR.t1002 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1149 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t34 XA.XIR[3].XIC[1].icell.Ien VGND.t2035 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1150 VPWR.t97 XThR.Tn[10].t36 XA.XIR[11].XIC[12].icell.PUM VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1151 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t33 VPWR.t1545 VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1152 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[4].XIC[8].icell.Ien VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1153 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t33 VPWR.t1713 VPWR.t1712 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1154 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t23 XA.XIR[11].XIC[12].icell.Ien VPWR.t1574 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1155 XThC.Tn[10].t2 XThC.XTB3.Y.t8 a_8739_9569# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1156 VGND.t59 XThC.XTB7.Y XThC.Tn[6].t3 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1157 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t46 VGND.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1158 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t38 VGND.t1237 VGND.t1236 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1159 XA.XIR[0].XIC[12].icell.PDM VGND.t1411 VGND.t1413 VGND.t1412 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1160 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t37 VPWR.t562 VPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 XThR.Tn[11].t10 XThR.XTBN.Y VPWR.t1761 VPWR.t1742 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1162 XA.XIR[13].XIC_15.icell.PDM VPWR.t1980 VGND.t852 VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1163 VPWR.t1003 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1164 VGND.t2160 XThC.Tn[12].t24 XA.XIR[0].XIC[12].icell.PDM VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1165 VGND.t448 XThC.Tn[3].t23 XA.XIR[14].XIC[3].icell.PDM VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1166 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1981 VGND.t854 VGND.t853 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1167 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t30 XA.XIR[7].XIC[5].icell.Ien VGND.t1968 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1168 VGND.t1781 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t1780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1169 VGND.t856 VPWR.t1982 XA.XIR[13].XIC_15.icell.PDM VGND.t855 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1170 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[3].icell.Ien VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1171 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t38 XA.XIR[0].XIC[12].icell.Ien VGND.t2648 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1172 VGND.t1783 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t1782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t39 XA.XIR[13].XIC_15.icell.Ien VGND.t1238 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1174 VPWR.t317 XThR.Tn[9].t38 XA.XIR[10].XIC[0].icell.PUM VPWR.t316 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1175 VGND.t1785 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t1784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1176 VGND.t351 XThC.Tn[9].t26 XA.XIR[1].XIC[9].icell.PDM VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1177 VGND.t1787 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t1786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1178 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[10].XIC[0].icell.Ien VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1179 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t37 VGND.t111 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1180 VGND.t2527 XThC.XTB7.A XThC.XTB7.Y VGND.t2526 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1181 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t34 XA.XIR[1].XIC[9].icell.Ien VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1182 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t6 VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1183 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t159 VGND.t1640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1184 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t38 VPWR.t99 VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1185 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t26 XA.XIR[1].XIC[11].icell.Ien VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1186 VGND.t2049 XThC.Tn[14].t24 XA.XIR[11].XIC[14].icell.PDM VGND.t2048 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1187 a_n997_2667# XThR.XTBN.Y VGND.t2476 VGND.t2431 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1188 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t811 VPWR.t813 VPWR.t812 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1189 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t38 XA.XIR[11].XIC[14].icell.Ien VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1190 VPWR.t101 XThR.Tn[10].t39 XA.XIR[11].XIC[10].icell.PUM VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1191 a_7875_9569# XThC.XTBN.Y.t49 VGND.t1075 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1192 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t35 VPWR.t1547 VPWR.t1546 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1193 VPWR.t1421 XThR.Tn[7].t31 XA.XIR[8].XIC[12].icell.PUM VPWR.t1420 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1194 VGND.t2475 XThR.XTBN.Y a_n997_3979# VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1195 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[11].XIC[10].icell.Ien VPWR.t1303 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1196 VGND.t1605 Vbias.t1 Vbias.t2 VGND.t1604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X1197 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t243 VGND.t2558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1198 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[8].XIC[12].icell.Ien VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1199 XThC.Tn[14].t10 XThC.XTBN.Y.t50 VPWR.t1004 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1200 a_n1049_6699# XThR.XTB4.Y.t7 VPWR.t1621 VPWR.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1201 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t39 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1202 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t7 VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1203 VPWR.t1465 XThR.Tn[3].t35 XA.XIR[4].XIC[3].icell.PUM VPWR.t1464 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1204 VGND.t1789 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t1788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1205 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t40 VPWR.t1171 VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1206 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t26 XA.XIR[1].XIC[2].icell.Ien VPWR.t1047 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1207 VGND.t2096 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t2095 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1208 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t36 VPWR.t1549 VPWR.t1548 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1209 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t24 XA.XIR[4].XIC[3].icell.Ien VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1210 XThC.Tn[2].t2 XThC.XTB3.Y.t9 VGND.t192 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1211 XThC.Tn[9].t10 XThC.XTBN.Y.t52 VPWR.t1006 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1212 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t34 VPWR.t1715 VPWR.t1714 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1213 XThC.Tn[5].t4 XThC.XTBN.Y.t53 VGND.t1076 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1214 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1215 VGND.t2098 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t2097 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1216 VGND.t1410 VGND.t1408 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1217 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t32 VGND.t1970 VGND.t1969 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1218 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t33 XA.XIR[7].XIC[0].icell.Ien VGND.t1971 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1219 VGND.t2136 XThC.Tn[13].t26 XA.XIR[5].XIC[13].icell.PDM VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1220 VPWR.t404 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1221 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[10].icell.Ien VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1222 XThC.Tn[0].t7 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1223 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t34 XA.XIR[5].XIC[13].icell.Ien VGND.t2132 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1224 VGND.t2051 XThC.Tn[14].t25 XA.XIR[8].XIC[14].icell.PDM VGND.t2050 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1225 XThR.Tn[12].t1 XThR.XTB5.Y VPWR.t1190 VPWR.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1226 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t41 XA.XIR[8].XIC[14].icell.Ien VGND.t1302 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1227 VPWR.t1423 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1228 VGND.t2100 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t2099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1229 VGND.t416 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1230 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t161 VGND.t1642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1231 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[5].XIC[9].icell.Ien VPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1232 XThR.Tn[6].t10 XThR.XTBN.Y VGND.t2473 VGND.t2472 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1233 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t2 VPWR.t1760 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1234 VGND.t2471 XThR.XTBN.Y a_n997_2891# VGND.t2470 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1235 VGND.t1222 XThR.XTB7.B XThR.XTB7.Y VGND.t1221 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1236 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[4].icell.Ien VGND.t1935 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1237 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t35 VPWR.t1557 VPWR.t1556 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1238 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[8].XIC[10].icell.Ien VPWR.t1304 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1239 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t129 VGND.t1213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1240 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t40 XA.XIR[9].XIC[1].icell.Ien VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1241 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t42 VPWR.t1173 VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1242 VPWR.t85 XThR.Tn[10].t40 XA.XIR[11].XIC[5].icell.PUM VPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1243 a_n997_2667# XThR.XTB4.Y.t8 XThR.Tn[11].t7 VGND.t1291 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[11].XIC[5].icell.Ien VPWR.t1331 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1245 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t220 VGND.t2231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1246 VGND.t2102 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t2101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1247 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t40 VPWR.t1489 VPWR.t1488 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1248 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t595 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1249 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t135 VGND.t1311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1250 VGND.t2104 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t2103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1251 VGND.t1077 XThC.XTBN.Y.t55 XThC.Tn[1].t9 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1252 a_n1049_6405# XThR.XTB5.Y VPWR.t1188 VPWR.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1253 VGND.t1649 XThC.Tn[11].t27 XA.XIR[5].XIC[11].icell.PDM VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1254 VGND.t2106 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t2105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1255 VGND.t1407 VGND.t1405 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1256 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t36 XA.XIR[5].XIC[11].icell.Ien VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1257 VPWR.t446 XThR.Tn[14].t42 XA.XIR[15].XIC[14].icell.PUM VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1258 VPWR.t810 VPWR.t808 XA.XIR[14].XIC_15.icell.PUM VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1259 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1983 VGND.t858 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1260 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[15].XIC[14].icell.Ien VPWR.t1501 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1261 VPWR.t389 XThR.XTB1.Y.t10 XThR.Tn[8].t0 VPWR.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1262 XA.XIR[14].XIC_15.icell.PUM VPWR.t806 XA.XIR[14].XIC_15.icell.Ien VPWR.t807 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1263 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t37 VGND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1264 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t41 VGND.t103 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1265 VPWR.t1759 XThR.XTBN.Y XThR.Tn[7].t2 VPWR.t1758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1266 VGND.t238 XThC.XTB2.Y XThC.Tn[1].t3 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 VGND.t860 VPWR.t1984 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t859 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1268 VGND.t1134 XThC.Tn[2].t27 XA.XIR[5].XIC[2].icell.PDM VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1269 VPWR.t1559 XThR.Tn[5].t37 XA.XIR[6].XIC[4].icell.PUM VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1270 XA.XIR[15].XIC[14].icell.Ien VPWR.t803 VPWR.t805 VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1271 VPWR.t802 VPWR.t800 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t801 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1272 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t43 VPWR.t448 VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1273 VGND.t1163 XThC.Tn[7].t21 XA.XIR[11].XIC[7].icell.PDM VGND.t1162 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1274 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t198 VGND.t1910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1275 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t1008 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1276 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[2].icell.Ien VGND.t2134 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1277 VPWR.t799 VPWR.t797 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1278 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[6].XIC[4].icell.Ien VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1279 VGND.t2251 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t752 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1280 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1985 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1281 XThR.Tn[1].t6 XThR.XTBN.Y a_n1049_7787# VPWR.t1737 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1282 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t41 XA.XIR[11].XIC[7].icell.Ien VGND.t2045 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1283 VPWR.t1425 XThR.Tn[7].t35 XA.XIR[8].XIC[5].icell.PUM VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1284 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t16 VGND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1285 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t35 VPWR.t1455 VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1286 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[8].XIC[5].icell.Ien VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1287 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t242 VGND.t2529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1288 VGND.t2108 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t2107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1289 VGND.t2110 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t2109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1290 VGND.t1404 VGND.t1402 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1291 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1986 VGND.t863 VGND.t862 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1292 VGND.t865 VPWR.t1987 XA.XIR[12].XIC_15.icell.PDM VGND.t864 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1293 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t43 VPWR.t1175 VPWR.t1174 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1294 XThR.Tn[9].t1 XThR.XTB2.Y VPWR.t1637 VPWR.t1636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1295 XThR.Tn[7].t5 XThR.XTBN.Y VGND.t2469 VGND.t2468 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1296 VPWR.t1055 data[1].t2 XThC.XTB6.A VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1297 VGND.t867 VPWR.t1988 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t866 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1298 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t40 XA.XIR[12].XIC_15.icell.Ien VGND.t1952 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1299 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t36 VGND.t2028 VGND.t2027 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1300 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t868 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1301 VGND.t1078 XThC.XTBN.Y.t57 a_7875_9569# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1302 VPWR.t1757 XThR.XTBN.Y XThR.Tn[13].t2 VPWR.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1303 VGND.t1736 XThC.Tn[5].t27 XA.XIR[7].XIC[5].icell.PDM VGND.t1735 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1304 XA.XIR[9].XIC_15.icell.PDM VPWR.t1990 VGND.t870 VGND.t869 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1305 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1306 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t241 VGND.t2528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1307 VGND.t2112 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t2111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1308 VPWR.t1912 XThR.XTB3.Y.t9 XThR.Tn[10].t9 VPWR.t1640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1309 VGND.t1591 XThC.Tn[6].t26 XA.XIR[5].XIC[6].icell.PDM VGND.t1590 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1310 VGND.t872 VPWR.t1991 XA.XIR[9].XIC_15.icell.PDM VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1311 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t36 VGND.t1973 VGND.t1972 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1312 XThC.Tn[3].t6 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1313 VPWR.t31 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1314 VPWR.t1561 XThR.Tn[5].t39 XA.XIR[6].XIC[0].icell.PUM VPWR.t1560 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1315 XThR.Tn[5].t10 XThR.XTB6.Y VGND.t2667 VGND.t1318 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1316 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t40 XA.XIR[5].XIC[6].icell.Ien VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1317 VGND.t1165 XThC.Tn[7].t22 XA.XIR[8].XIC[7].icell.PDM VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1318 VPWR.t1133 XThR.XTB7.B XThR.XTB4.Y.t0 VPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1319 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1320 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[3].XIC[4].icell.Ien VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1321 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[6].XIC[0].icell.Ien VPWR.t1667 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1322 VPWR.t319 XThR.Tn[9].t41 XA.XIR[10].XIC[13].icell.PUM VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1323 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t44 XA.XIR[8].XIC[7].icell.Ien VGND.t1303 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1324 VPWR.t796 VPWR.t794 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t795 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1325 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t36 VPWR.t1467 VPWR.t1466 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1326 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[10].XIC[13].icell.Ien VPWR.t1562 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1327 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t37 VPWR.t1457 VPWR.t1456 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1328 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t37 VPWR.t1427 VPWR.t1426 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1329 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t1187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1330 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t792 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t793 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1331 VGND.t2114 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t2113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1332 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t42 VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1333 VGND.t1401 VGND.t1399 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1334 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1335 VGND.t2116 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t2115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1336 VGND.t2118 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t2117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1337 VGND.t2120 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t2119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1338 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t40 VGND.t1240 VGND.t1239 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1339 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t142 VGND.t1471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1340 VGND.t2162 XThC.Tn[12].t26 XA.XIR[14].XIC[12].icell.PDM VGND.t2161 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1341 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t38 XA.XIR[7].XIC[14].icell.Ien VGND.t1974 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1342 VPWR.t13 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1343 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t38 VGND.t2030 VGND.t2029 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1344 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t39 VGND.t2650 VGND.t2649 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1345 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[12].icell.Ien VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1346 VGND.t2309 XThC.Tn[0].t27 XA.XIR[7].XIC[0].icell.PDM VGND.t2308 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1347 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t33 VGND.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1348 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t28 XA.XIR[3].XIC[0].icell.Ien VPWR.t1668 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1349 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t35 VGND.t2356 VGND.t2355 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1350 VGND.t2122 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t2121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1351 VGND.t1247 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t1246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1352 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t39 VPWR.t1429 VPWR.t1428 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1353 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t37 VPWR.t1469 VPWR.t1468 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1354 VPWR.t1851 XThR.Tn[0].t40 XA.XIR[1].XIC[9].icell.PUM VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1355 XThC.Tn[1].t8 XThC.XTBN.Y.t59 VGND.t1079 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 VPWR.t1696 XThR.Tn[4].t36 XA.XIR[5].XIC[9].icell.PUM VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1357 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t5 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1358 VGND.t1249 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t1248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1359 VGND.t1251 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t1250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1360 XThR.Tn[13].t9 XThR.XTB6.Y a_n997_1579# VGND.t1317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1361 VPWR.t321 XThR.Tn[9].t42 XA.XIR[10].XIC[6].icell.PUM VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1362 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t6 VPWR.t1756 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1363 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1364 VPWR.t1412 XThR.Tn[12].t41 XA.XIR[13].XIC[7].icell.PUM VPWR.t1411 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1365 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t27 XA.XIR[10].XIC[6].icell.Ien VPWR.t1258 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1366 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t38 VGND.t1937 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1367 VPWR.t1491 XThR.Tn[11].t42 XA.XIR[12].XIC[8].icell.PUM VPWR.t1490 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1368 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t41 VGND.t2652 VGND.t2651 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1369 VGND.t1253 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t1252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1370 VGND.t1255 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t1254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1371 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[13].XIC[7].icell.Ien VPWR.t1077 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1372 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t246 VGND.t2636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1373 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t37 VGND.t2358 VGND.t2357 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1374 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t89 VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1375 VGND.t1665 XThC.Tn[10].t27 XA.XIR[2].XIC[10].icell.PDM VGND.t1664 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1376 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t197 VGND.t1909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1377 VGND.t1257 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t1256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1378 VPWR.t791 VPWR.t789 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1379 VGND.t1259 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t1258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1380 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t41 VPWR.t1143 VPWR.t1142 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1381 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[10].icell.Ien VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1382 VGND.t726 data[2].t1 XThC.XTB7.B VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1383 VPWR.t91 XThR.Tn[10].t44 XA.XIR[11].XIC[14].icell.PUM VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1384 VGND.t2467 XThR.XTBN.Y XThR.Tn[2].t9 VGND.t2466 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1385 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t787 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t788 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1386 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t248 VGND.t2639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1387 a_n1049_5317# XThR.XTB7.Y VPWR.t129 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1388 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t39 VGND.t1939 VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1389 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t43 VPWR.t323 VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1390 VGND.t1080 XThC.XTBN.Y.t60 XThC.Tn[4].t9 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1391 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t42 VGND.t2654 VGND.t2653 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1392 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t784 VPWR.t786 VPWR.t785 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1393 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[11].XIC[14].icell.Ien VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1394 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t232 VGND.t2342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1395 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t24 VGND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1396 VGND.t616 XThC.Tn[1].t25 XA.XIR[2].XIC[1].icell.PDM VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1397 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t38 VGND.t2360 VGND.t2359 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1398 VGND.t1261 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t1260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1399 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t43 VPWR.t1493 VPWR.t1492 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1400 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t44 VGND.t217 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1401 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t40 VPWR.t1431 VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1402 VGND.t1263 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t1262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1403 VGND.t1265 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t1264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t6 VGND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1405 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[1].icell.Ien VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1406 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t42 VGND.t1954 VGND.t1953 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1407 VGND.t2630 XThC.Tn[8].t25 XA.XIR[10].XIC[8].icell.PDM VGND.t2629 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1408 XThR.Tn[3].t0 XThR.XTB4.Y.t9 VGND.t715 VGND.t714 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1409 VGND.t1267 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t1266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1410 VGND.t1922 XThC.Tn[9].t28 XA.XIR[13].XIC[9].icell.PDM VGND.t1921 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1411 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t45 XA.XIR[10].XIC[8].icell.Ien VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1412 VPWR.t51 XThC.XTB7.Y a_6243_9615# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VPWR.t1319 XThC.XTB6.Y XThC.Tn[13].t6 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1414 VPWR.t1414 XThR.Tn[12].t43 XA.XIR[13].XIC[11].icell.PUM VPWR.t1413 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1415 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[9].icell.Ien VGND.t1241 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1416 VGND.t592 data[1].t3 XThC.XTB5.A VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1417 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[13].XIC[11].icell.Ien VPWR.t1299 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1418 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t874 VGND.t873 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1419 VGND.t1269 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t1268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1420 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t151 VGND.t1512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1421 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t73 VGND.t698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1422 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t43 VPWR.t1145 VPWR.t1144 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1423 VGND.t876 VPWR.t1993 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1424 VPWR.t186 XThR.Tn[9].t45 XA.XIR[10].XIC[1].icell.PUM VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1425 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t2235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1426 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t209 VGND.t2008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1427 VGND.t253 XThC.XTBN.Y.t61 XThC.Tn[7].t6 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1428 VPWR.t1416 XThR.Tn[12].t44 XA.XIR[13].XIC[2].icell.PUM VPWR.t1415 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1429 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1994 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t877 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1430 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t169 VGND.t1790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1431 VPWR.t1495 XThR.Tn[11].t44 XA.XIR[12].XIC[3].icell.PUM VPWR.t1494 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1432 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t26 XA.XIR[10].XIC[1].icell.Ien VPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1433 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t41 XA.XIR[7].XIC[7].icell.Ien VGND.t1975 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1434 VPWR.t1433 XThR.Tn[7].t42 XA.XIR[8].XIC[14].icell.PUM VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1435 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t43 VGND.t2656 VGND.t2655 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1436 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[13].XIC[2].icell.Ien VPWR.t1048 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1437 XThR.Tn[12].t0 XThR.XTB5.Y VPWR.t1186 VPWR.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1438 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t46 VPWR.t93 VPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1439 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t39 VGND.t2362 VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1440 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t28 XA.XIR[8].XIC[14].icell.Ien VPWR.t1503 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1441 a_10915_9569# XThC.XTBN.Y.t62 VGND.t255 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t136 VGND.t1324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1443 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t46 VPWR.t188 VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1444 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t44 VPWR.t1231 VPWR.t1230 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1445 XThR.Tn[6].t9 XThR.XTBN.Y VGND.t2465 VGND.t2464 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1446 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1995 VGND.t879 VGND.t878 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1447 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t45 VPWR.t1177 VPWR.t1176 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1448 VPWR.t1459 XThR.Tn[6].t39 XA.XIR[7].XIC[12].icell.PUM VPWR.t1458 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1449 XThC.Tn[3].t2 XThC.XTB4.Y.t7 VGND.t1081 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 XThC.Tn[9].t1 XThC.XTB2.Y VPWR.t202 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1451 VGND.t881 VPWR.t1996 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t880 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1452 VPWR.t1807 XThR.Tn[5].t41 XA.XIR[6].XIC[13].icell.PUM VPWR.t1806 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1453 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[7].XIC[12].icell.Ien VPWR.t1576 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1454 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1997 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1455 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[6].XIC[13].icell.Ien VPWR.t1563 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1456 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t47 VGND.t219 VGND.t218 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1457 a_n997_2667# XThR.XTB4.Y.t10 XThR.Tn[11].t0 VGND.t716 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1458 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t40 VPWR.t265 VPWR.t264 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1459 VGND.t1271 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t1270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1460 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t45 VGND.t1754 VGND.t1753 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1461 VGND.t450 XThC.Tn[3].t25 XA.XIR[10].XIC[3].icell.PDM VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1462 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t155 VGND.t1625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1463 VGND.t884 VPWR.t1998 XA.XIR[5].XIC_15.icell.PDM VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1464 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1999 VGND.t886 VGND.t885 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1465 VGND.t418 XThC.Tn[4].t28 XA.XIR[13].XIC[4].icell.PDM VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1466 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t47 XA.XIR[10].XIC[3].icell.Ien VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1467 VGND.t888 VPWR.t2000 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t887 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1468 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC_15.icell.Ien VGND.t2599 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1469 XA.XIR[0].XIC[5].icell.PDM VGND.t1396 VGND.t1398 VGND.t1397 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1470 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t38 VGND.t2037 VGND.t2036 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1471 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t45 XA.XIR[13].XIC[4].icell.Ien VGND.t1472 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1472 VGND.t1220 XThR.XTB7.B a_n1335_8331# VGND.t1219 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1473 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2001 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t889 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1474 VGND.t1738 XThC.Tn[5].t28 XA.XIR[0].XIC[5].icell.PDM VGND.t1737 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1475 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t41 VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1476 VPWR.t225 XThC.XTBN.Y.t63 XThC.Tn[9].t9 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1477 VGND.t2138 XThC.Tn[13].t29 XA.XIR[4].XIC[13].icell.PDM VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1478 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t210 VGND.t2009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1479 a_10051_9569# XThC.XTBN.Y.t64 VGND.t257 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1480 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t44 XA.XIR[0].XIC[5].icell.Ien VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1481 VPWR.t1292 XThR.Tn[3].t39 XA.XIR[4].XIC[9].icell.PUM VPWR.t1291 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1482 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[13].icell.Ien VGND.t2363 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1483 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t152 VGND.t1513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1484 VPWR.t1755 XThR.XTBN.Y XThR.Tn[7].t1 VPWR.t1754 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1485 VGND.t2078 XThC.Tn[14].t29 XA.XIR[7].XIC[14].icell.PDM VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1486 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[4].XIC[9].icell.Ien VPWR.t1397 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1487 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t127 VGND.t1211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1488 VPWR.t267 XThR.Tn[6].t42 XA.XIR[7].XIC[10].icell.PUM VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1489 XThC.Tn[11].t2 XThC.XTB4.Y.t8 VPWR.t1010 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1490 VGND.t2463 XThR.XTBN.Y XThR.Tn[1].t10 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1491 XThR.Tn[1].t5 XThR.XTBN.Y a_n1049_7787# VPWR.t1735 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1492 VPWR.t15 XThR.Tn[2].t41 XA.XIR[3].XIC[13].icell.PUM VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1493 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[7].XIC[10].icell.Ien VPWR.t1305 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1494 a_7651_9569# XThC.XTBN.Y.t65 VGND.t259 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1495 VPWR.t783 VPWR.t781 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t782 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1496 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t41 VPWR.t1698 VPWR.t1697 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1497 VGND.t1273 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t1272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1498 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[3].XIC[13].icell.Ien VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1499 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t779 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t780 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1500 VGND.t2531 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t2530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1501 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t40 VPWR.t1294 VPWR.t1293 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1502 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t776 VPWR.t778 VPWR.t777 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1503 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t1063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1504 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1505 a_n1049_5611# XThR.XTB6.Y VPWR.t1874 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1506 XThR.Tn[9].t0 XThR.XTB2.Y VPWR.t1635 VPWR.t1634 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1507 VPWR.t450 XThR.Tn[14].t45 XA.XIR[15].XIC[8].icell.PUM VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1508 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t24 XA.XIR[12].XIC[7].icell.Ien VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1509 VGND.t1667 XThC.Tn[10].t29 XA.XIR[1].XIC[10].icell.PDM VGND.t1666 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1510 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t41 VGND.t1631 VGND.t1630 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1511 VGND.t2533 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t2532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1512 XThC.Tn[4].t8 XThC.XTBN.Y.t66 VGND.t260 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1513 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[15].XIC[8].icell.Ien VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1514 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t46 VPWR.t1343 VPWR.t1342 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VPWR.t1753 XThR.XTBN.Y XThR.Tn[13].t1 VPWR.t1731 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1516 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t40 XA.XIR[1].XIC[10].icell.Ien VGND.t1940 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1517 VGND.t1651 XThC.Tn[11].t29 XA.XIR[4].XIC[11].icell.PDM VGND.t1650 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1518 VPWR.t1809 XThR.Tn[5].t43 XA.XIR[6].XIC[6].icell.PUM VPWR.t1808 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1519 XA.XIR[15].XIC[8].icell.Ien VPWR.t773 VPWR.t775 VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1520 VGND.t1395 VGND.t1393 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1521 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t31 VGND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1522 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t42 XA.XIR[4].XIC[11].icell.Ien VGND.t2364 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1523 VPWR.t1179 XThR.Tn[8].t46 XA.XIR[9].XIC[7].icell.PUM VPWR.t1178 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1524 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t28 XA.XIR[6].XIC[6].icell.Ien VPWR.t1259 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1525 XA.XIR[0].XIC[0].icell.PDM VGND.t1390 VGND.t1392 VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1526 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t42 VGND.t1633 VGND.t1632 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1527 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t25 XA.XIR[9].XIC[7].icell.Ien VPWR.t1079 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1528 VGND.t459 XThR.XTB1.Y.t11 XThR.Tn[0].t1 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1529 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t138 VGND.t1326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1530 VGND.t618 XThC.Tn[1].t27 XA.XIR[1].XIC[1].icell.PDM VGND.t617 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1531 XThR.Tn[5].t5 XThR.XTBN.Y VGND.t2462 VGND.t2446 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1532 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t43 VPWR.t269 VPWR.t268 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1533 VGND.t1084 XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.PDM VGND.t1083 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1534 VGND.t1218 XThR.XTB7.B XThR.XTB6.Y VGND.t1216 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1535 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t41 XA.XIR[1].XIC[1].icell.Ien VGND.t1941 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1536 VGND.t1136 XThC.Tn[2].t29 XA.XIR[4].XIC[2].icell.PDM VGND.t1135 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1537 VGND.t261 XThC.XTBN.Y.t67 XThC.Tn[0].t4 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1538 VGND.t2535 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t2534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1539 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t45 XA.XIR[0].XIC[0].icell.Ien VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1540 VGND.t2537 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t2536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1541 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t43 XA.XIR[4].XIC[2].icell.Ien VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1542 VGND.t1924 XThC.Tn[9].t30 XA.XIR[12].XIC[9].icell.PDM VGND.t1923 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1543 VGND.t263 XThC.XTBN.Y.t68 XThC.Tn[3].t11 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1544 VGND.t2539 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t2538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1545 VPWR.t271 XThR.Tn[6].t44 XA.XIR[7].XIC[5].icell.PUM VPWR.t270 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1546 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t47 XA.XIR[12].XIC[9].icell.Ien VGND.t1755 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1547 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t29 XA.XIR[7].XIC[5].icell.Ien VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1548 XThC.Tn[7].t5 XThC.XTBN.Y.t69 VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1549 VPWR.t227 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1550 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[12].XIC[11].icell.Ien VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1551 VGND.t2541 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t2540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t44 VGND.t2601 VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1553 VGND.t2543 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t2542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1554 VGND.t2545 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t2544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1555 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t1305 VGND.t1304 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1556 VPWR.t1633 XThR.XTB2.Y a_n1049_7787# VPWR.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1557 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t48 VPWR.t1345 VPWR.t1344 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1558 VGND.t2632 XThC.Tn[8].t27 XA.XIR[6].XIC[8].icell.PDM VGND.t2631 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1559 VGND.t2547 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t2546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1560 VGND.t2549 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t2548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1561 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t225 VGND.t2246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1562 VGND.t267 XThC.XTBN.Y.t71 a_10915_9569# VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1563 VGND.t1926 XThC.Tn[9].t31 XA.XIR[9].XIC[9].icell.PDM VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1564 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t45 XA.XIR[6].XIC[8].icell.Ien VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1565 VPWR.t17 XThR.Tn[2].t42 XA.XIR[3].XIC[6].icell.PUM VPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1566 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t34 VGND.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1567 XThC.Tn[11].t6 XThC.XTB4.Y.t9 a_8963_9569# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1568 VPWR.t1181 XThR.Tn[8].t48 XA.XIR[9].XIC[11].icell.PUM VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1569 VPWR.t452 XThR.Tn[14].t46 XA.XIR[15].XIC[3].icell.PUM VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1570 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[12].XIC[2].icell.Ien VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1571 VGND.t1082 XThC.XTB4.Y.t10 XThC.Tn[3].t1 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1572 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[3].XIC[6].icell.Ien VPWR.t1260 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1573 VPWR.t772 VPWR.t770 XA.XIR[10].XIC_15.icell.PUM VPWR.t771 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1574 VGND.t2551 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t2550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1575 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t43 VGND.t1635 VGND.t1634 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1576 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t31 XA.XIR[9].XIC[11].icell.Ien VPWR.t482 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1577 XThR.Tn[14].t11 XThR.XTBN.Y VPWR.t1752 VPWR.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1578 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t44 VPWR.t1296 VPWR.t1295 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1579 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t26 XA.XIR[15].XIC[3].icell.Ien VPWR.t383 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1580 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t49 VPWR.t1347 VPWR.t1346 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1581 VGND.t1593 XThC.Tn[6].t30 XA.XIR[4].XIC[6].icell.PDM VGND.t1592 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1582 XA.XIR[10].XIC_15.icell.PUM VPWR.t768 XA.XIR[10].XIC_15.icell.Ien VPWR.t769 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1583 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t43 VPWR.t1435 VPWR.t1434 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1584 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t46 VGND.t307 VGND.t306 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1585 VPWR.t1401 XThR.Tn[1].t42 XA.XIR[2].XIC[4].icell.PUM VPWR.t1400 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1586 VPWR.t1811 XThR.Tn[5].t45 XA.XIR[6].XIC[1].icell.PUM VPWR.t1810 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1587 XA.XIR[15].XIC[3].icell.Ien VPWR.t765 VPWR.t767 VPWR.t766 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1588 a_7875_9569# XThC.XTBN.Y.t72 VGND.t268 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1589 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t48 VPWR.t79 VPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1590 VGND.t1167 XThC.Tn[7].t26 XA.XIR[7].XIC[7].icell.PDM VGND.t1166 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1591 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC[6].icell.Ien VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1592 VPWR.t1873 XThR.XTB6.Y XThR.Tn[13].t7 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1593 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[2].XIC[4].icell.Ien VPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1594 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t28 XA.XIR[6].XIC[1].icell.Ien VPWR.t490 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1595 VPWR.t1183 XThR.Tn[8].t49 XA.XIR[9].XIC[2].icell.PUM VPWR.t1182 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1596 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t31 XA.XIR[9].XIC[2].icell.Ien VPWR.t1158 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1597 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t5 VGND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1598 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t43 VPWR.t19 VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1599 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t47 VPWR.t273 VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1600 XThC.Tn[11].t5 XThC.XTB4.Y.t11 a_8963_9569# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1601 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t44 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1602 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t48 VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1603 VGND.t2553 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t2552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1604 VGND.t2555 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t2554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1605 VGND.t1389 VGND.t1387 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1606 XThC.Tn[0].t0 XThC.XTB1.Y.t12 VGND.t468 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1607 VGND.t2634 XThC.Tn[8].t28 XA.XIR[3].XIC[8].icell.PDM VGND.t2633 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1608 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t200 VGND.t1912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1609 VGND.t420 XThC.Tn[4].t30 XA.XIR[12].XIC[4].icell.PDM VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1610 VGND.t269 XThC.XTBN.Y.t73 a_10051_9569# VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1611 XThR.XTB1.Y.t0 XThR.XTB5.A VPWR.t33 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1612 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t45 XA.XIR[3].XIC[8].icell.Ien VGND.t1636 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1613 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t50 XA.XIR[12].XIC[4].icell.Ien VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1614 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1615 XThR.Tn[13].t8 XThR.XTB6.Y a_n997_1579# VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1616 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t46 VGND.t2603 VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1617 XA.XIR[1].XIC_15.icell.PDM VPWR.t2003 VGND.t892 VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1618 XA.XIR[5].XIC_15.icell.PDM VPWR.t2004 VGND.t894 VGND.t893 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1619 VGND.t1943 XThC.Tn[3].t27 XA.XIR[6].XIC[3].icell.PDM VGND.t1942 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1620 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t50 VGND.t1307 VGND.t1306 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1621 VGND.t270 XThC.XTBN.Y.t74 a_7651_9569# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1622 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t146 VGND.t1490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1623 XThC.XTBN.Y.t2 XThC.XTBN.A VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1624 VGND.t422 XThC.Tn[4].t31 XA.XIR[9].XIC[4].icell.PDM VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1625 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t48 XA.XIR[6].XIC[3].icell.Ien VGND.t2239 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1626 VPWR.t21 XThR.Tn[2].t45 XA.XIR[3].XIC[1].icell.PUM VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1627 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t170 VGND.t1791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1628 VPWR.t1403 XThR.Tn[1].t43 XA.XIR[2].XIC[0].icell.PUM VPWR.t1402 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1629 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1630 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1631 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[3].XIC[1].icell.Ien VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1632 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t30 XA.XIR[2].XIC[0].icell.Ien VPWR.t1011 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1633 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t6 VPWR.t1749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1634 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t46 VPWR.t137 VPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1635 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t46 VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t166 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1637 VPWR.t229 XThC.XTBN.Y.t75 XThC.Tn[7].t0 VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1638 VGND.t2461 XThR.XTBN.Y a_n997_1803# VGND.t2460 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1639 VPWR.t1213 VGND.t2696 XA.XIR[0].XIC[12].icell.PUM VPWR.t1212 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1640 XThR.Tn[3].t9 XThR.XTBN.Y VGND.t2459 VGND.t2413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1641 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t28 XA.XIR[0].XIC[12].icell.Ien VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1642 VPWR.t764 VPWR.t762 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t763 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1643 VPWR.t1820 XThC.XTB4.Y.t12 XThC.Tn[11].t1 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1644 VGND.t2557 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t2556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1645 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t47 VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1646 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t46 VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1647 VPWR.t1211 VGND.t2697 Vbias.t3 VPWR.t1210 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X1648 VGND.t1945 XThC.Tn[3].t28 XA.XIR[3].XIC[3].icell.PDM VGND.t1944 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1649 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t168 VGND.t1718 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1650 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t49 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1651 XThC.Tn[0].t3 XThC.XTBN.Y.t76 VGND.t271 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1652 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t165 VGND.t1655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t47 XA.XIR[3].XIC[3].icell.Ien VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1654 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t53 VGND.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1655 VPWR.t81 XThR.Tn[10].t49 XA.XIR[11].XIC[8].icell.PUM VPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1656 VGND.t2164 XThC.Tn[12].t29 XA.XIR[10].XIC[12].icell.PDM VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1657 XThC.Tn[3].t10 XThC.XTBN.Y.t77 VGND.t2366 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1658 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t50 VPWR.t192 VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1659 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t29 XA.XIR[11].XIC[8].icell.Ien VPWR.t1840 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1660 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t50 XA.XIR[10].XIC[12].icell.Ien VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1661 XA.XIR[0].XIC[14].icell.PDM VGND.t1384 VGND.t1386 VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1662 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t46 VGND.t1474 VGND.t1473 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1663 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t391 VPWR.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1664 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t45 VPWR.t1497 VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1665 VGND.t1854 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t1853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1666 VGND.t1740 XThC.Tn[5].t30 XA.XIR[14].XIC[5].icell.PDM VGND.t1739 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1667 VGND.t2080 XThC.Tn[14].t30 XA.XIR[0].XIC[14].icell.PDM VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1668 VPWR.t1209 VGND.t2698 XA.XIR[0].XIC[10].icell.PUM VPWR.t1208 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1669 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t47 XA.XIR[0].XIC[14].icell.Ien VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1670 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t47 XA.XIR[14].XIC[5].icell.Ien VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1671 VGND.t1856 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t1855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t30 XA.XIR[0].XIC[10].icell.Ien VPWR.t1306 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1673 XThC.XTB1.Y.t1 XThC.XTB5.A a_3299_10575# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1674 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t48 VPWR.t333 VPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VGND.t2680 XThR.XTB3.Y.t10 XThR.Tn[2].t11 VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1676 VPWR.t761 VPWR.t759 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t760 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1677 VGND.t1858 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t1857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t51 XA.XIR[9].XIC[8].icell.Ien VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1679 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t2345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1680 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t757 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t758 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1681 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t754 VPWR.t756 VPWR.t755 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1682 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t27 XA.XIR[5].XIC[7].icell.Ien VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1683 VPWR.t1437 XThR.Tn[7].t44 XA.XIR[8].XIC[8].icell.PUM VPWR.t1436 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1684 VGND.t2368 XThC.XTBN.Y.t78 XThC.Tn[6].t10 VGND.t2367 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1685 VGND.t1860 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t1859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t179 VGND.t1812 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1687 XThC.Tn[10].t3 XThC.XTB3.Y.t11 VPWR.t167 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1688 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[8].XIC[8].icell.Ien VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1689 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t47 VPWR.t1813 VPWR.t1812 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1690 VGND.t1383 VGND.t1381 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1691 VGND.t1862 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t1861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1692 VGND.t1864 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t1863 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1693 XThC.Tn[14].t2 XThC.XTB7.Y VPWR.t50 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1694 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[1].XIC[4].icell.Ien VPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1695 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t51 VPWR.t231 VPWR.t230 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1696 VPWR.t83 XThR.Tn[10].t51 XA.XIR[11].XIC[3].icell.PUM VPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1697 VPWR.t1623 XThR.Tn[6].t49 XA.XIR[7].XIC[14].icell.PUM VPWR.t1622 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1698 VGND.t469 XThC.XTB1.Y.t13 XThC.Tn[0].t1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1699 VPWR.t753 VPWR.t751 XA.XIR[6].XIC_15.icell.PUM VPWR.t752 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1700 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t44 VPWR.t1793 VPWR.t1792 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1701 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t52 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[11].XIC[3].icell.Ien VPWR.t1404 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1703 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[7].XIC[14].icell.Ien VPWR.t1530 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1704 XA.XIR[6].XIC_15.icell.PUM VPWR.t749 XA.XIR[6].XIC_15.icell.Ien VPWR.t750 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1705 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t47 VGND.t1476 VGND.t1475 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1706 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t46 VPWR.t1499 VPWR.t1498 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1707 VGND.t1866 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t1865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1708 XThR.Tn[8].t9 XThR.XTBN.Y VPWR.t1751 VPWR.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1709 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t40 VGND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1710 VGND.t1868 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t1867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1711 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t36 VGND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1712 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t50 VPWR.t1625 VPWR.t1624 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1713 VGND.t1086 XThC.Tn[0].t31 XA.XIR[14].XIC[0].icell.PDM VGND.t1085 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1714 VGND.t1928 XThC.Tn[9].t32 XA.XIR[5].XIC[9].icell.PDM VGND.t1927 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1715 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t47 VGND.t2220 VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1716 VPWR.t1207 VGND.t2699 XA.XIR[0].XIC[5].icell.PUM VPWR.t1206 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1717 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t48 XA.XIR[14].XIC[0].icell.Ien VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1718 VGND.t1870 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t1869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1719 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t48 XA.XIR[5].XIC[9].icell.Ien VGND.t2604 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1720 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t31 XA.XIR[0].XIC[5].icell.Ien VPWR.t1334 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1721 XA.XIR[4].XIC_15.icell.PDM VPWR.t2005 VGND.t896 VGND.t895 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1722 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t1 VPWR.t1749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1723 VPWR.t1615 XThR.Tn[11].t48 XA.XIR[12].XIC[9].icell.PUM VPWR.t1614 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1724 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t32 XA.XIR[5].XIC[11].icell.Ien VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1725 VGND.t1872 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t1871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t49 VPWR.t335 VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t898 VPWR.t2006 XA.XIR[4].XIC_15.icell.PDM VGND.t897 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1728 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t49 VPWR.t1815 VPWR.t1814 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1729 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2007 VGND.t900 VGND.t899 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1730 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t180 VGND.t1813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1731 XThR.XTBN.A data[7].t1 VGND.t1907 VGND.t1906 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1732 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t53 XA.XIR[9].XIC[3].icell.Ien VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1733 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t45 XA.XIR[4].XIC_15.icell.Ien VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1734 VGND.t902 VPWR.t2008 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t901 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1735 XThC.Tn[14].t1 XThC.XTB7.Y VPWR.t49 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1736 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[1].XIC[0].icell.Ien VPWR.t1012 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1737 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t32 XA.XIR[5].XIC[2].icell.Ien VPWR.t1159 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1738 VPWR.t510 XThR.Tn[7].t45 XA.XIR[8].XIC[3].icell.PUM VPWR.t509 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1739 XThC.XTB2.Y XThC.XTB7.B VPWR.t1350 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1740 VPWR.t748 VPWR.t746 XA.XIR[3].XIC_15.icell.PUM VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1741 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t45 VPWR.t1795 VPWR.t1794 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1742 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t96 VGND.t1061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1743 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t30 XA.XIR[8].XIC[3].icell.Ien VPWR.t1405 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1744 XA.XIR[3].XIC_15.icell.PUM VPWR.t744 XA.XIR[3].XIC_15.icell.Ien VPWR.t745 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1745 XThR.Tn[5].t4 XThR.XTBN.Y VGND.t2458 VGND.t2437 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1746 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t50 VPWR.t1817 VPWR.t1816 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1747 XA.XIR[0].XIC[7].icell.PDM VGND.t1378 VGND.t1380 VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1748 VGND.t1874 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t1873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1749 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t51 VGND.t1758 VGND.t1757 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1750 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2009 VGND.t904 VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1751 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t52 VPWR.t233 VPWR.t232 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1752 VGND.t1227 XThC.Tn[7].t28 XA.XIR[0].XIC[7].icell.PDM VGND.t1226 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1753 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t48 VPWR.t139 VPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1754 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t49 VGND.t2222 VGND.t2221 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1755 XThR.Tn[10].t6 XThR.XTBN.Y VPWR.t1748 VPWR.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1756 Vbias.t4 bias[1].t0 VPWR.t1860 VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X1757 VGND.t906 VPWR.t2010 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t905 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1758 a_5949_9615# XThC.XTB6.Y VPWR.t1318 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1759 VPWR.t1797 XThR.Tn[1].t46 XA.XIR[2].XIC[13].icell.PUM VPWR.t1796 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1760 VGND.t1669 XThC.Tn[10].t31 XA.XIR[13].XIC[10].icell.PDM VGND.t1668 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1761 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t50 XA.XIR[0].XIC[7].icell.Ien VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1762 VPWR.t743 VPWR.t741 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1763 VGND.t1876 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t1875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1764 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[2].XIC[13].icell.Ien VPWR.t1565 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1765 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t48 XA.XIR[13].XIC[10].icell.Ien VGND.t1477 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1766 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2011 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t907 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1767 VGND.t1878 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t1877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1768 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t163 VGND.t1653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t739 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t740 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1770 VPWR.t603 XThC.XTB3.Y.t12 XThC.Tn[10].t4 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1771 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t48 VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1772 VGND.t1377 VGND.t1375 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1773 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t98 VGND.t1064 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1774 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t52 VGND.t1760 VGND.t1759 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1775 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t9 VGND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1776 XThC.Tn[13].t8 XThC.XTBN.Y.t79 VPWR.t1699 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1777 VGND.t424 XThC.Tn[4].t33 XA.XIR[5].XIC[4].icell.PDM VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1778 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t736 VPWR.t738 VPWR.t737 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t50 VGND.t2224 VGND.t2223 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1780 a_n997_3755# XThR.XTBN.Y VGND.t2457 VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1781 VGND.t620 XThC.Tn[1].t30 XA.XIR[13].XIC[1].icell.PDM VGND.t619 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1782 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t171 VGND.t1792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1783 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t51 XA.XIR[5].XIC[4].icell.Ien VGND.t2605 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1784 VPWR.t1746 XThR.XTBN.Y XThR.Tn[14].t10 VPWR.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1785 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t88 VGND.t1038 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1786 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[1].icell.Ien VGND.t1478 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1787 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t87 VGND.t1037 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1788 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t52 VGND.t2059 VGND.t2058 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1789 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t29 VGND.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1790 XThR.Tn[7].t4 XThR.XTBN.Y VGND.t2456 VGND.t2455 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1791 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t50 VGND.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1792 VGND.t2166 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t2165 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1793 XThC.XTB4.Y.t1 XThC.XTB7.B VGND.t1798 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1794 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[12].icell.Ien VGND.t2240 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1795 VPWR.t1872 XThR.XTB6.Y XThR.Tn[13].t6 VPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t1913 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t1638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 VGND.t1880 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t1879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1798 VPWR.t1301 data[4].t3 XThR.XTB7.A VPWR.t1300 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1799 VGND.t943 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XThC.Tn[6].t9 XThC.XTBN.Y.t80 VGND.t2370 VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1801 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t51 VGND.t2226 VGND.t2225 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1802 XThR.Tn[5].t9 XThR.XTB6.Y VGND.t2666 VGND.t1314 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1803 VPWR.t414 XThC.XTB5.Y a_5155_9615# VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1804 VGND.t945 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VPWR.t1233 XThR.Tn[13].t50 XA.XIR[14].XIC[12].icell.PUM VPWR.t1232 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1806 XThR.Tn[4].t2 XThR.XTB5.Y VGND.t1319 VGND.t1318 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1807 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1821 VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1808 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t9 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1809 VGND.t947 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t946 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1810 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[14].XIC[12].icell.Ien VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1811 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t46 VPWR.t512 VPWR.t511 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t1799 XThR.Tn[1].t47 XA.XIR[2].XIC[6].icell.PUM VPWR.t1798 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1813 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t25 VGND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1814 VGND.t2371 XThC.XTBN.Y.t82 XThC.Tn[2].t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1815 VPWR.t337 XThR.Tn[0].t51 XA.XIR[1].XIC[7].icell.PUM VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1816 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t49 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1817 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t49 VPWR.t1366 VPWR.t1365 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1818 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t26 VGND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1819 VPWR.t406 XThC.XTB1.Y.t14 XThC.Tn[8].t5 VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1820 VPWR.t1593 XThR.Tn[4].t46 XA.XIR[5].XIC[7].icell.PUM VPWR.t1592 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1821 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[2].XIC[6].icell.Ien VPWR.t1261 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1822 VGND.t2325 XThC.Tn[12].t32 XA.XIR[3].XIC[12].icell.PDM VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1823 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1824 a_10915_9569# XThC.XTBN.Y.t83 VGND.t2373 VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1825 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t50 VPWR.t41 VPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1826 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t49 XA.XIR[3].XIC[12].icell.Ien VGND.t145 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1827 VGND.t949 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1828 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t54 VPWR.t299 VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1829 XThC.Tn[3].t0 XThC.XTB4.Y.t14 VGND.t2614 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t951 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1831 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t50 VGND.t1886 VGND.t1885 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1832 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t51 VGND.t2254 VGND.t2253 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1833 VGND.t2140 XThC.Tn[13].t32 XA.XIR[15].XIC[13].icell.PDM VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1834 VGND.t2082 XThC.Tn[14].t32 XA.XIR[14].XIC[14].icell.PDM VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1835 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t48 VGND.t2524 VGND.t2523 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1836 XThR.Tn[3].t8 XThR.XTBN.Y VGND.t2454 VGND.t2453 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1837 XA.XIR[15].XIC[13].icell.PDM VPWR.t2012 XA.XIR[15].XIC[13].icell.Ien VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1838 VPWR.t1368 XThR.Tn[14].t51 XA.XIR[15].XIC[9].icell.PUM VPWR.t1367 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1839 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t52 VGND.t382 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1840 VPWR.t1645 XThR.Tn[13].t52 XA.XIR[14].XIC[10].icell.PUM VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1841 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t52 XA.XIR[14].XIC[14].icell.Ien VGND.t1887 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1842 VGND.t953 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 VGND.t955 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1844 VGND.t957 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1845 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t47 VGND.t2202 VGND.t2201 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1846 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t33 XA.XIR[15].XIC[9].icell.Ien VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1847 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t5 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1848 VGND.t2287 XThC.Tn[8].t31 XA.XIR[2].XIC[8].icell.PDM VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1849 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[14].XIC[10].icell.Ien VPWR.t1307 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1850 a_4387_10575# XThC.XTB7.B VGND.t1797 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1851 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t207 VGND.t2006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1852 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t51 XA.XIR[2].XIC[8].icell.Ien VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1853 XA.XIR[15].XIC[9].icell.Ien VPWR.t733 VPWR.t735 VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1854 VPWR.t339 XThR.Tn[0].t53 XA.XIR[1].XIC[11].icell.PUM VPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1855 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t53 VPWR.t1370 VPWR.t1369 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t41 VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1857 VPWR.t1595 XThR.Tn[4].t48 XA.XIR[5].XIC[11].icell.PUM VPWR.t1594 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1858 a_10051_9569# XThC.XTBN.Y.t84 VGND.t2374 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1859 XThC.XTB1.Y.t2 XThC.XTB7.B VPWR.t1349 VPWR.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1860 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t5 VPWR.t1741 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1861 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t47 VPWR.t514 VPWR.t513 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1862 VPWR.t1801 XThR.Tn[1].t49 XA.XIR[2].XIC[1].icell.PUM VPWR.t1800 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1863 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t76 VGND.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1864 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t71 VGND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1865 VPWR.t1235 XThR.Tn[0].t54 XA.XIR[1].XIC[2].icell.PUM VPWR.t1234 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1866 VGND.t959 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1867 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t1716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1868 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t5 VPWR.t1744 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1869 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t54 VGND.t1889 VGND.t1888 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1870 VGND.t1671 XThC.Tn[10].t33 XA.XIR[12].XIC[10].icell.PDM VGND.t1670 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1871 a_7651_9569# XThC.XTBN.Y.t85 VGND.t2375 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1872 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t31 XA.XIR[2].XIC[1].icell.Ien VPWR.t492 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1873 VPWR.t1597 XThR.Tn[4].t49 XA.XIR[5].XIC[2].icell.PUM VPWR.t1596 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1874 VPWR.t1205 VGND.t2700 XA.XIR[0].XIC[14].icell.PUM VPWR.t1204 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1875 VGND.t1374 VGND.t1372 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1876 VGND.t597 XThC.Tn[11].t33 XA.XIR[15].XIC[11].icell.PDM VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1877 VPWR.t1805 XThC.XTB7.A a_6243_10571# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1878 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[1].XIC[13].icell.Ien VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1879 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[10].icell.Ien VGND.t1761 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1880 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t52 VPWR.t43 VPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1881 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[0].XIC[14].icell.Ien VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1882 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t50 VPWR.t1803 VPWR.t1802 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1883 XA.XIR[15].XIC[11].icell.PDM VPWR.t2013 XA.XIR[15].XIC[11].icell.Ien VGND.t909 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1884 XThC.Tn[10].t5 XThC.XTB3.Y.t13 a_8739_9569# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1885 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t55 VPWR.t1237 VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1886 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2014 VGND.t911 VGND.t910 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1887 VGND.t961 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t53 VGND.t273 VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1889 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t215 VGND.t2056 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1890 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t55 VGND.t1891 VGND.t1890 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1891 VGND.t622 XThC.Tn[1].t32 XA.XIR[12].XIC[1].icell.PDM VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1892 VGND.t2452 XThR.XTBN.Y XThR.Tn[2].t8 VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1893 VGND.t913 VPWR.t2015 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t912 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1894 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t235 VGND.t2406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1895 VGND.t1673 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t1672 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1896 XThR.XTB5.A data[5].t3 VGND.t309 VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1897 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t255 VGND.t2683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1898 VGND.t1280 XThC.Tn[2].t33 XA.XIR[15].XIC[2].icell.PDM VGND.t1279 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1899 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[1].icell.Ien VGND.t1208 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1900 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2016 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1901 VPWR.t732 VPWR.t730 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t731 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1902 XThR.Tn[12].t9 XThR.XTBN.Y VPWR.t1743 VPWR.t1742 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1903 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t51 VGND.t2090 VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1904 XA.XIR[15].XIC[2].icell.PDM VPWR.t2017 XA.XIR[15].XIC[2].icell.Ien VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1905 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1480 VGND.t1479 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1906 VPWR.t1647 XThR.Tn[13].t53 XA.XIR[14].XIC[5].icell.PUM VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1907 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t728 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t729 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1908 XThR.Tn[12].t5 XThR.XTB5.Y a_n997_1803# VGND.t1317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1909 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t114 VGND.t1137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1910 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t50 VGND.t2204 VGND.t2203 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1911 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t54 VGND.t275 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1912 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2018 VGND.t760 VGND.t759 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1913 VGND.t1947 XThC.Tn[3].t31 XA.XIR[2].XIC[3].icell.PDM VGND.t1946 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1914 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t32 XA.XIR[14].XIC[5].icell.Ien VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1915 XThR.Tn[3].t1 XThR.XTB4.Y.t11 VGND.t717 VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1916 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t133 VGND.t1274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1917 VGND.t2450 XThR.XTBN.Y a_n997_2667# VGND.t2449 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1918 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t725 VPWR.t727 VPWR.t726 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1919 VGND.t624 XThC.Tn[1].t33 XA.XIR[9].XIC[1].icell.PDM VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1920 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[3].icell.Ien VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1921 VGND.t762 VPWR.t2019 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1922 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t56 VPWR.t1372 VPWR.t1371 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1923 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t184 VGND.t1817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1924 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1925 VGND.t963 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1926 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2020 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1927 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t55 XA.XIR[9].XIC[12].icell.Ien VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1928 a_5155_9615# XThC.XTB5.Y VPWR.t413 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1929 VPWR.t412 XThC.XTB5.Y XThC.Tn[12].t0 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1930 XThC.Tn[5].t8 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1931 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t101 VGND.t1067 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1932 VGND.t478 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1933 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2021 VGND.t765 VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1934 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t9 VPWR.t1741 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1935 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t57 VGND.t1893 VGND.t1892 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1936 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t54 VGND.t2256 VGND.t2255 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1937 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t164 VGND.t1654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1938 XThC.Tn[2].t8 XThC.XTBN.Y.t87 VGND.t2376 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1939 VGND.t767 VPWR.t2022 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1940 VGND.t1595 XThC.Tn[6].t32 XA.XIR[15].XIC[6].icell.PDM VGND.t1594 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1941 VGND.t1229 XThC.Tn[7].t29 XA.XIR[14].XIC[7].icell.PDM VGND.t1228 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1942 VPWR.t1113 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t1112 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1943 VPWR.t724 VPWR.t722 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t723 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1944 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t5 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1945 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2023 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[6].icell.PDM VPWR.t2024 XA.XIR[15].XIC[6].icell.Ien VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1947 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t58 XA.XIR[14].XIC[7].icell.Ien VGND.t1894 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1948 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t34 XA.XIR[13].XIC[4].icell.Ien VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1949 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t720 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t721 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1950 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t42 VGND.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1951 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t2411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1952 VPWR.t1131 XThR.XTB7.B XThR.XTB2.Y VPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1953 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t1649 VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1954 Vbias.t0 bias[2].t0 VPWR.t400 VPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1955 XThC.Tn[8].t8 XThC.XTB1.Y.t15 a_7651_9569# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t33 XA.XIR[1].XIC[6].icell.Ien VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1957 VPWR.t141 XThR.Tn[3].t50 XA.XIR[4].XIC[7].icell.PUM VPWR.t140 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t30 VGND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t717 VPWR.t719 VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1960 VGND.t210 XThC.XTB5.A XThC.XTB5.Y VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t1371 VGND.t1369 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[4].XIC[7].icell.Ien VPWR.t1138 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1963 VPWR.t1627 XThR.Tn[6].t52 XA.XIR[7].XIC[8].icell.PUM VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t52 VPWR.t1535 VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1965 VGND.t131 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1966 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[7].XIC[8].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1967 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t51 VPWR.t1599 VPWR.t1598 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1968 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t56 VGND.t337 VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1969 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t113 VGND.t1120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1970 VGND.t1742 XThC.Tn[5].t33 XA.XIR[10].XIC[5].icell.PDM VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1971 XA.XIR[12].XIC_15.icell.PDM VPWR.t2025 VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1972 XThR.Tn[9].t8 XThR.XTBN.Y VPWR.t1740 VPWR.t1720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1973 VGND.t2377 XThC.XTBN.Y.t89 a_9827_9569# VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1974 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t52 XA.XIR[10].XIC[5].icell.Ien VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1975 VGND.t965 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1976 VGND.t2289 XThC.Tn[8].t33 XA.XIR[1].XIC[8].icell.PDM VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1977 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t51 VGND.t147 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1978 XThC.Tn[0].t2 XThC.XTB1.Y.t16 VGND.t470 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1979 VGND.t967 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1980 VGND.t969 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1981 VPWR.t1115 XThR.Tn[12].t56 XA.XIR[13].XIC[0].icell.PUM VPWR.t1114 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1982 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t53 VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X1983 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t0 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1984 VGND.t1930 XThC.Tn[9].t34 XA.XIR[4].XIC[9].icell.PDM VGND.t1929 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1985 VPWR.t716 VPWR.t714 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t715 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1986 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t53 XA.XIR[1].XIC[8].icell.Ien VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1987 VGND.t2168 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t2167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1988 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t33 XA.XIR[13].XIC[0].icell.Ien VPWR.t1013 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1989 VPWR.t143 XThR.Tn[3].t52 XA.XIR[4].XIC[11].icell.PUM VPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1990 VGND.t2142 XThC.Tn[13].t34 XA.XIR[11].XIC[13].icell.PDM VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1991 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t2637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1992 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t52 XA.XIR[4].XIC[9].icell.Ien VGND.t2205 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1993 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t712 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t713 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1994 XThR.Tn[14].t9 XThR.XTBN.Y VPWR.t1739 VPWR.t1738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1995 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1651 VPWR.t1650 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t52 XA.XIR[11].XIC[13].icell.Ien VGND.t2227 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X1997 VPWR.t75 XThR.Tn[10].t54 XA.XIR[11].XIC[9].icell.PUM VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1998 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t34 XA.XIR[4].XIC[11].icell.Ien VPWR.t484 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1999 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t709 VPWR.t711 VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2000 a_n997_3755# XThR.XTBN.Y VGND.t2448 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2001 XThR.Tn[8].t1 XThR.XTB1.Y.t13 VPWR.t393 VPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2002 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t53 VPWR.t1523 VPWR.t1522 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2003 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[11].XIC[9].icell.Ien VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2004 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t251 VGND.t2663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2005 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t53 VPWR.t1617 VPWR.t1616 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2006 VGND.t2170 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t2169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2007 a_n1049_7787# XThR.XTB2.Y VPWR.t1632 VPWR.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2008 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t34 XA.XIR[1].XIC[1].icell.Ien VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2009 VPWR.t577 XThR.Tn[3].t53 XA.XIR[4].XIC[2].icell.PUM VPWR.t576 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2010 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t99 VGND.t1065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2011 a_n1331_2891# data[5].t4 VGND.t1819 VGND.t1818 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2012 VGND.t2172 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t2171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2013 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t54 VPWR.t1537 VPWR.t1536 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2014 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t34 XA.XIR[4].XIC[2].icell.Ien VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2015 VPWR.t1629 XThR.Tn[6].t53 XA.XIR[7].XIC[3].icell.PUM VPWR.t1628 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2016 VPWR.t708 VPWR.t706 XA.XIR[2].XIC_15.icell.PUM VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2017 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[7].XIC[3].icell.Ien VPWR.t1406 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2018 XA.XIR[2].XIC_15.icell.PUM VPWR.t704 XA.XIR[2].XIC_15.icell.Ien VPWR.t705 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2019 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t54 VPWR.t1525 VPWR.t1524 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2020 XThR.XTB7.B data[6].t1 VGND.t1176 VGND.t1175 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2021 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t57 VGND.t339 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2022 XThR.Tn[2].t4 XThR.XTBN.Y a_n1049_7493# VPWR.t1737 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2023 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t54 VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2024 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t55 VGND.t88 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2025 VGND.t1088 XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.PDM VGND.t1087 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2026 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t79 VGND.t712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2027 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t48 VGND.t678 VGND.t677 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2028 VGND.t599 XThC.Tn[11].t35 XA.XIR[11].XIC[11].icell.PDM VGND.t598 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2029 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t56 XA.XIR[10].XIC[0].icell.Ien VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2030 VGND.t2144 XThC.Tn[13].t35 XA.XIR[8].XIC[13].icell.PDM VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2031 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2026 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2032 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t54 XA.XIR[11].XIC[11].icell.Ien VGND.t1201 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2033 VPWR.t516 XThR.Tn[7].t49 XA.XIR[8].XIC[9].icell.PUM VPWR.t515 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2034 VGND.t2174 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t2173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2035 VGND.t2607 XThC.Tn[3].t33 XA.XIR[1].XIC[3].icell.PDM VGND.t2606 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2036 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t54 VGND.t920 VGND.t919 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2037 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t55 XA.XIR[8].XIC[13].icell.Ien VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2038 VPWR.t1831 XThC.XTBN.Y.t90 XThC.Tn[8].t2 VPWR.t1830 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2039 XThR.Tn[10].t10 XThR.XTB3.Y.t12 VPWR.t1914 VPWR.t1636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2040 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t57 VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2041 XThR.Tn[4].t5 XThR.XTBN.Y VGND.t2447 VGND.t2446 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 VGND.t426 XThC.Tn[4].t35 XA.XIR[4].XIC[4].icell.PDM VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2043 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[8].XIC[9].icell.Ien VPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2044 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t55 XA.XIR[1].XIC[3].icell.Ien VGND.t2092 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t231 VGND.t2341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t1217 XThR.XTB7.B XThR.XTB5.Y VGND.t1216 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t2176 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t2175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t1282 XThC.Tn[2].t35 XA.XIR[11].XIC[2].icell.PDM VGND.t1281 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2049 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t56 VPWR.t235 VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2050 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[4].icell.Ien VGND.t2070 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2051 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t55 XA.XIR[11].XIC[2].icell.Ien VGND.t1202 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2052 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t212 VGND.t2011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2053 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t5 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2054 XThC.Tn[4].t4 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2055 VGND.t2178 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t2177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2056 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t229 VGND.t2339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2057 VGND.t2180 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t2179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2058 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t186 VGND.t1881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 VGND.t1675 XThC.Tn[10].t35 XA.XIR[5].XIC[10].icell.PDM VGND.t1674 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2060 VGND.t2182 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t2181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2061 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t680 VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2062 VGND.t2445 XThR.XTBN.Y a_n997_1579# VGND.t2427 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2063 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[10].icell.Ien VGND.t2060 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2064 VGND.t601 XThC.Tn[11].t36 XA.XIR[8].XIC[11].icell.PDM VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2065 VPWR.t1653 XThR.Tn[13].t57 XA.XIR[14].XIC[14].icell.PUM VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2066 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[12].XIC[4].icell.Ien VPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2067 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t57 XA.XIR[8].XIC[11].icell.Ien VGND.t277 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2068 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t57 VPWR.t1117 VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t34 XA.XIR[14].XIC[14].icell.Ien VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2070 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t58 VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2071 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t701 VPWR.t703 VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2072 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t39 VGND.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2073 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t107 VGND.t1112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2074 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t5 VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2075 VGND.t2616 XThC.Tn[1].t35 XA.XIR[5].XIC[1].icell.PDM VGND.t2615 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2076 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t682 VGND.t681 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2077 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t59 VPWR.t1374 VPWR.t1373 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2078 VGND.t1597 XThC.Tn[6].t34 XA.XIR[11].XIC[6].icell.PDM VGND.t1596 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2079 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t65 VGND.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2080 VPWR.t237 XThR.Tn[8].t58 XA.XIR[9].XIC[4].icell.PUM VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2081 VGND.t1284 XThC.Tn[2].t36 XA.XIR[8].XIC[2].icell.PDM VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2082 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t111 VGND.t1117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2083 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[1].icell.Ien VGND.t2061 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2084 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC[6].icell.Ien VGND.t1203 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2085 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[9].XIC[4].icell.Ien VPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2086 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[2].icell.Ien VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2087 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t56 VGND.t2094 VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2088 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t228 VGND.t2338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2089 XA.XIR[15].XIC_15.icell.PDM VPWR.t2027 VGND.t774 VGND.t773 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2090 VGND.t2327 XThC.Tn[12].t33 XA.XIR[2].XIC[12].icell.PDM VGND.t2326 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2091 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2028 VGND.t776 VGND.t775 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2092 XThR.XTBN.Y XThR.XTBN.A VPWR.t532 VPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2093 VGND.t2184 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t2183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2094 VGND.t778 VPWR.t2029 XA.XIR[15].XIC_15.icell.PDM VGND.t777 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2095 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t55 XA.XIR[2].XIC[12].icell.Ien VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2096 VGND.t780 VPWR.t2030 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t779 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2097 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t55 VGND.t2063 VGND.t2062 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2098 XA.XIR[15].XIC_15.icell.PDM VPWR.t2031 XA.XIR[15].XIC_15.icell.Ien VGND.t781 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2099 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2032 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t782 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2100 VGND.t2186 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t2185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2101 VPWR.t1736 XThR.XTBN.Y XThR.Tn[11].t9 VPWR.t1716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2102 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t35 XA.XIR[12].XIC[0].icell.Ien VPWR.t1014 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2103 VGND.t1744 XThC.Tn[5].t34 XA.XIR[6].XIC[5].icell.PDM VGND.t1743 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2104 VPWR.t1050 data[1].t4 XThC.XTB7.A VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2105 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t684 VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2106 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t58 VPWR.t1119 VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2107 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t54 XA.XIR[6].XIC[5].icell.Ien VGND.t2241 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2108 a_8739_9569# XThC.XTBN.Y.t92 VGND.t2623 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2109 VGND.t1599 XThC.Tn[6].t35 XA.XIR[8].XIC[6].icell.PDM VGND.t1598 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2110 VGND.t709 XThR.XTBN.A XThR.XTBN.Y VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2111 XThC.Tn[6].t2 XThC.XTB7.Y VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2112 VPWR.t301 XThR.Tn[9].t58 XA.XIR[10].XIC[12].icell.PUM VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2113 VPWR.t239 XThR.Tn[8].t60 XA.XIR[9].XIC[0].icell.PUM VPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2114 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t61 XA.XIR[8].XIC[6].icell.Ien VGND.t279 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2115 VPWR.t700 VPWR.t698 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2116 VPWR.t1121 XThR.Tn[12].t59 XA.XIR[13].XIC[13].icell.PUM VPWR.t1120 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2117 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t34 XA.XIR[10].XIC[12].icell.Ien VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2118 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[9].XIC[0].icell.Ien VPWR.t1015 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2119 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t696 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t697 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2120 XThR.Tn[12].t4 XThR.XTB5.Y a_n997_1803# VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t36 XA.XIR[13].XIC[13].icell.Ien VPWR.t1567 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2122 VGND.t2188 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t2187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2123 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t59 VPWR.t77 VPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2124 VPWR.t1203 VGND.t2701 XA.XIR[0].XIC[8].icell.PUM VPWR.t1202 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2125 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t693 VPWR.t695 VPWR.t694 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2126 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t58 VPWR.t1471 VPWR.t1470 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2127 VGND.t2190 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t2189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2128 XA.XIR[1].XIC_15.icell.PUM VPWR.t691 XA.XIR[1].XIC_15.icell.Ien VPWR.t692 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2129 a_n997_3979# XThR.XTBN.Y VGND.t2444 VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2130 XThC.XTB7.Y XThC.XTB7.B VGND.t1796 VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2131 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t34 XA.XIR[0].XIC[8].icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2132 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t57 VPWR.t1539 VPWR.t1538 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2133 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t56 VGND.t1069 VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2134 VGND.t2192 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t2191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2135 VGND.t2194 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t2193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2136 XThC.Tn[8].t1 XThC.XTBN.Y.t93 VPWR.t1833 VPWR.t1832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2137 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t57 VPWR.t1239 VPWR.t1238 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2138 VGND.t1822 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t1821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2139 VGND.t436 XThC.Tn[5].t35 XA.XIR[3].XIC[5].icell.PDM VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2140 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t59 VGND.t341 VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2141 a_n1049_6699# XThR.XTB4.Y.t12 VPWR.t536 VPWR.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2142 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t55 XA.XIR[3].XIC[5].icell.Ien VGND.t921 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2143 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t158 VGND.t1639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2144 VGND.t2084 XThC.Tn[14].t35 XA.XIR[10].XIC[14].icell.PDM VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2145 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC[13].icell.Ien VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2146 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t56 VGND.t2065 VGND.t2064 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2147 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t60 XA.XIR[10].XIC[14].icell.Ien VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2148 VPWR.t303 XThR.Tn[9].t60 XA.XIR[10].XIC[10].icell.PUM VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2149 VGND.t1824 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t1823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2150 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t84 VGND.t916 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2151 VGND.t1090 XThC.Tn[0].t37 XA.XIR[6].XIC[0].icell.PDM VGND.t1089 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2152 VPWR.t690 VPWR.t688 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2153 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[10].XIC[10].icell.Ien VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2154 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t54 VPWR.t518 VPWR.t517 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2155 VGND.t1826 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t1825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2156 VGND.t1828 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t1827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2157 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t55 XA.XIR[6].XIC[0].icell.Ien VGND.t2242 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2158 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t686 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2159 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t61 VPWR.t65 VPWR.t64 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2160 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t683 VPWR.t685 VPWR.t684 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2161 VGND.t294 data[1].t5 XThC.XTB6.A VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2162 a_n997_2891# XThR.XTBN.Y VGND.t2442 VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2163 VGND.t1830 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t1829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t1832 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t1831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VPWR.t1201 VGND.t2702 XA.XIR[0].XIC[3].icell.PUM VPWR.t1200 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2166 VGND.t1834 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t1833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2167 VGND.t1368 VGND.t1366 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2168 VPWR.t1123 XThR.Tn[12].t60 XA.XIR[13].XIC[6].icell.PUM VPWR.t1122 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2169 XThR.Tn[11].t1 XThR.XTB4.Y.t13 a_n997_2667# VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2170 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t55 XA.XIR[7].XIC[11].icell.Ien VGND.t686 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2171 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[0].XIC[3].icell.Ien VPWR.t1818 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2172 VPWR.t1109 XThR.Tn[11].t57 XA.XIR[12].XIC[7].icell.PUM VPWR.t1108 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2173 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t58 VGND.t1482 VGND.t1481 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2174 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t57 VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2175 VGND.t1836 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t1835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2176 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t36 XA.XIR[13].XIC[6].icell.Ien VPWR.t1263 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2177 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t59 VPWR.t1241 VPWR.t1240 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2178 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2033 VGND.t784 VGND.t783 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2179 VPWR.t411 XThC.XTB5.Y a_5155_9615# VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2180 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t56 VGND.t2072 VGND.t2071 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2181 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t17 VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2182 VGND.t1838 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t1837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2183 VGND.t1092 XThC.Tn[0].t38 XA.XIR[3].XIC[0].icell.PDM VGND.t1091 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2184 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t1473 VPWR.t1472 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2185 VGND.t786 VPWR.t2034 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t785 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2186 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t56 XA.XIR[3].XIC[0].icell.Ien VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2187 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2035 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t787 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2188 VPWR.t682 VPWR.t680 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2189 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t56 XA.XIR[7].XIC[2].icell.Ien VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2190 VGND.t2440 XThR.XTBN.Y XThR.Tn[0].t9 VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2191 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t60 VGND.t1484 VGND.t1483 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2192 VPWR.t305 XThR.Tn[9].t61 XA.XIR[10].XIC[5].icell.PUM VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2193 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t678 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t679 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2194 a_n1049_6405# XThR.XTB5.Y VPWR.t1184 VPWR.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2195 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t110 VGND.t1116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XThR.Tn[8].t2 XThR.XTB1.Y.t14 VPWR.t395 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2197 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t195 VGND.t1904 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2198 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t57 VGND.t2074 VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2199 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t36 XA.XIR[10].XIC[5].icell.Ien VPWR.t376 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2200 VGND.t1840 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t1839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2201 VGND.t2329 XThC.Tn[12].t35 XA.XIR[1].XIC[12].icell.PDM VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t59 VGND.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2203 VGND.t1842 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t1841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2204 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t61 VGND.t1210 VGND.t1209 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2205 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t58 VGND.t1205 VGND.t1204 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2206 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t62 VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2207 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[12].icell.Ien VGND.t1955 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2208 VGND.t1844 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t1843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2209 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t2250 VGND.t1276 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2210 VGND.t2291 XThC.Tn[8].t35 XA.XIR[13].XIC[8].icell.PDM VGND.t2290 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2211 VGND.t2624 XThC.XTBN.Y.t94 a_8739_9569# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2212 VGND.t1846 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2213 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[8].icell.Ien VGND.t2038 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2214 XThC.Tn[1].t2 XThC.XTB2.Y VGND.t237 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2215 VGND.t54 XThC.XTB7.Y XThC.Tn[6].t1 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2216 VPWR.t1111 XThR.Tn[11].t59 XA.XIR[12].XIC[11].icell.PUM VPWR.t1110 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2217 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2218 XA.XIR[11].XIC_15.icell.PDM VPWR.t2036 VGND.t789 VGND.t788 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2219 VGND.t1848 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t1847 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2220 VGND.t626 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2221 XThR.Tn[2].t3 XThR.XTBN.Y a_n1049_7493# VPWR.t1735 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2222 VGND.t791 VPWR.t2037 XA.XIR[11].XIC_15.icell.PDM VGND.t790 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2223 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t62 VGND.t343 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2224 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t63 XA.XIR[9].XIC[5].icell.Ien VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2225 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t55 VGND.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2226 VGND.t1231 XThC.Tn[7].t31 XA.XIR[10].XIC[7].icell.PDM VGND.t1230 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2227 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t14 VGND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2228 VPWR.t1125 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2229 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t60 XA.XIR[11].XIC_15.icell.Ien VGND.t1206 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2230 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t57 XA.XIR[7].XIC[6].icell.Ien VGND.t688 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2231 VPWR.t247 XThR.Tn[11].t61 XA.XIR[12].XIC[2].icell.PUM VPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2232 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[5].XIC[4].icell.Ien VPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2233 XThR.Tn[13].t0 XThR.XTBN.Y VPWR.t1734 VPWR.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2234 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t36 XA.XIR[13].XIC[1].icell.Ien VPWR.t1825 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2235 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t63 XA.XIR[10].XIC[7].icell.Ien VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2236 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t148 VGND.t1509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2237 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t57 VPWR.t1513 VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2238 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[12].XIC[13].icell.Ien VPWR.t1568 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2239 XThR.Tn[10].t11 XThR.XTB3.Y.t13 VPWR.t1915 VPWR.t1634 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2240 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t61 VPWR.t1475 VPWR.t1474 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[4].t4 XThR.XTBN.Y VGND.t2438 VGND.t2437 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2242 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t63 VPWR.t169 VPWR.t168 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2243 VGND.t1365 VGND.t1363 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2244 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t675 VPWR.t677 VPWR.t676 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 VGND.t2665 XThR.XTB6.Y XThR.Tn[5].t8 VGND.t1312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2246 VPWR.t1515 XThR.Tn[5].t58 XA.XIR[6].XIC[12].icell.PUM VPWR.t1514 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2247 VGND.t628 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t627 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2248 VPWR.t241 XThR.Tn[8].t62 XA.XIR[9].XIC[13].icell.PUM VPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2249 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[6].XIC[12].icell.Ien VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2250 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t5 VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2251 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[9].XIC[13].icell.Ien VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2252 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t150 VGND.t1511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2253 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t4 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2254 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t56 VPWR.t1089 VPWR.t1088 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2255 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t64 VGND.t194 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2256 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t62 VGND.t290 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2257 VGND.t630 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2258 XA.XIR[8].XIC_15.icell.PDM VPWR.t2038 VGND.t793 VGND.t792 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2259 VGND.t2609 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t2608 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2260 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t124 VGND.t1193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2261 VGND.t632 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2262 VGND.t795 VPWR.t2039 XA.XIR[8].XIC_15.icell.PDM VGND.t794 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2263 VGND.t634 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2264 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t62 XA.XIR[13].XIC[3].icell.Ien VGND.t2039 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2265 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC_15.icell.Ien VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2266 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t39 XA.XIR[5].XIC[0].icell.Ien VPWR.t1016 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2267 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t57 VGND.t1179 VGND.t1178 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2268 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t59 VGND.t2067 VGND.t2066 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2269 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t60 VPWR.t1517 VPWR.t1516 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2270 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t64 XA.XIR[9].XIC[0].icell.Ien VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2271 VGND.t2146 XThC.Tn[13].t39 XA.XIR[7].XIC[13].icell.PDM VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2272 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t166 VGND.t1715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t2317 XThC.Tn[14].t36 XA.XIR[6].XIC[14].icell.PDM VGND.t2316 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2274 VPWR.t1091 XThR.Tn[6].t58 XA.XIR[7].XIC[9].icell.PUM VPWR.t1090 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2275 VPWR.t1165 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2276 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t154 VGND.t1620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2277 VPWR.t1519 XThR.Tn[5].t61 XA.XIR[6].XIC[10].icell.PUM VPWR.t1518 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2278 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t59 XA.XIR[6].XIC[14].icell.Ien VGND.t1180 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2279 VPWR.t994 XThR.Tn[2].t58 XA.XIR[3].XIC[12].icell.PUM VPWR.t993 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2280 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[7].XIC[9].icell.Ien VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2281 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[6].XIC[10].icell.Ien VPWR.t1309 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2282 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t37 XA.XIR[3].XIC[12].icell.Ien VPWR.t1678 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2283 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t60 VPWR.t1093 VPWR.t1092 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2284 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t190 VGND.t1897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2285 VGND.t636 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2286 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t57 VPWR.t579 VPWR.t578 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2287 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2288 VGND.t638 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2289 XThR.Tn[4].t1 XThR.XTB5.Y VGND.t1315 VGND.t1314 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2290 VPWR.t1732 XThR.XTBN.Y XThR.Tn[14].t8 VPWR.t1731 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2291 XThC.Tn[13].t5 XThC.XTB6.Y VPWR.t1317 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2292 VPWR.t1376 XThR.Tn[14].t60 XA.XIR[15].XIC[7].icell.PUM VPWR.t1375 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2293 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[12].XIC[6].icell.Ien VPWR.t1264 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2294 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t58 VGND.t924 VGND.t923 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2295 VPWR.t1477 XThR.Tn[13].t63 XA.XIR[14].XIC[8].icell.PUM VPWR.t1476 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2296 VGND.t1682 XThC.XTB6.Y XThC.Tn[5].t0 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2297 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t32 XA.XIR[15].XIC[7].icell.Ien VPWR.t1139 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2298 VGND.t797 VPWR.t2040 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t796 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2299 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t36 XA.XIR[14].XIC[8].icell.Ien VPWR.t1662 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2300 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t65 VPWR.t171 VPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2301 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t61 VGND.t1182 VGND.t1181 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2302 VGND.t1677 XThC.Tn[10].t38 XA.XIR[4].XIC[10].icell.PDM VGND.t1676 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2303 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t214 VGND.t2022 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2304 VPWR.t1730 XThR.XTBN.Y XThR.Tn[11].t8 VPWR.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2305 VGND.t640 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2306 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t59 VGND.t1073 VGND.t1072 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2307 XA.XIR[15].XIC[7].icell.Ien VPWR.t672 VPWR.t674 VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2308 VGND.t1362 VGND.t1360 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2309 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t2041 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t798 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2310 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t58 XA.XIR[4].XIC[10].icell.Ien VGND.t2075 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2311 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t61 VPWR.t1378 VPWR.t1377 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2312 VGND.t745 XThC.Tn[11].t37 XA.XIR[7].XIC[11].icell.PDM VGND.t744 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2313 VPWR.t243 XThR.Tn[8].t64 XA.XIR[9].XIC[6].icell.PUM VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2314 VGND.t2319 XThC.Tn[14].t37 XA.XIR[3].XIC[14].icell.PDM VGND.t2318 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2315 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t86 VGND.t970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2316 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t59 VGND.t926 VGND.t925 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2317 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[9].XIC[6].icell.Ien VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2318 XThC.Tn[9].t4 XThC.XTB2.Y a_7875_9569# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2319 VPWR.t996 XThR.Tn[2].t60 XA.XIR[3].XIC[10].icell.PUM VPWR.t995 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2320 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[14].icell.Ien VGND.t1628 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2321 VGND.t532 XThC.XTB6.A XThC.XTB6.Y VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2322 VGND.t2618 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2617 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2323 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t62 VGND.t1184 VGND.t1183 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2324 VGND.t235 XThC.XTB2.Y XThC.Tn[1].t1 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2325 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[3].XIC[10].icell.Ien VPWR.t1310 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2326 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t12 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2327 VGND.t642 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2328 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2329 VGND.t1286 XThC.Tn[2].t37 XA.XIR[7].XIC[2].icell.PDM VGND.t1285 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2330 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t105 VGND.t1110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2331 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t59 XA.XIR[4].XIC[1].icell.Ien VGND.t2076 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2332 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t62 VGND.t1896 VGND.t1895 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2333 VGND.t2293 XThC.Tn[8].t37 XA.XIR[12].XIC[8].icell.PDM VGND.t2292 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2334 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t61 VPWR.t1282 VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2335 VGND.t644 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t646 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2337 VPWR.t127 XThR.XTB7.Y a_n1049_5317# VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2338 VPWR.t1521 XThR.Tn[5].t62 XA.XIR[6].XIC[5].icell.PUM VPWR.t1520 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2339 VGND.t353 XThC.Tn[9].t38 XA.XIR[15].XIC[9].icell.PDM VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2340 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t66 XA.XIR[12].XIC[8].icell.Ien VGND.t195 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2341 VPWR.t1316 XThC.XTB6.Y XThC.Tn[13].t4 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2342 VPWR.t1380 XThR.Tn[14].t63 XA.XIR[15].XIC[11].icell.PUM VPWR.t1379 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2343 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[6].XIC[5].icell.Ien VPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2344 XA.XIR[15].XIC[9].icell.PDM VPWR.t2042 XA.XIR[15].XIC[9].icell.Ien VGND.t799 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2345 a_n997_3979# XThR.XTBN.Y VGND.t2436 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2346 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t65 VGND.t282 VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2347 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t38 XA.XIR[15].XIC[11].icell.Ien VPWR.t569 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2348 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t63 VPWR.t1095 VPWR.t1094 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2349 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t45 VGND.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2350 VGND.t648 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t650 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t128 VGND.t1212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t720 XThR.XTB4.Y.t14 XThR.Tn[3].t2 VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t91 VGND.t1048 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t487 VPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t5 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 XA.XIR[15].XIC[11].icell.Ien VPWR.t669 VPWR.t671 VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2358 VGND.t2295 XThC.Tn[8].t38 XA.XIR[9].XIC[8].icell.PDM VGND.t2294 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t48 VGND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 VGND.t652 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2361 VGND.t1359 VGND.t1357 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VPWR.t1382 XThR.Tn[14].t64 XA.XIR[15].XIC[2].icell.PUM VPWR.t1381 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2363 VPWR.t1479 XThR.Tn[13].t64 XA.XIR[14].XIC[3].icell.PUM VPWR.t1478 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2364 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t28 VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2365 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t38 XA.XIR[12].XIC[1].icell.Ien VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2366 VPWR.t1059 XThR.Tn[9].t65 XA.XIR[10].XIC[14].icell.PUM VPWR.t1058 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2367 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t4 VPWR.t1728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2368 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t38 XA.XIR[15].XIC[2].icell.Ien VPWR.t1161 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2369 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t67 VPWR.t173 VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2370 VPWR.t668 VPWR.t666 XA.XIR[13].XIC_15.icell.PUM VPWR.t667 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2371 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t36 XA.XIR[14].XIC[3].icell.Ien VPWR.t1819 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2372 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[10].XIC[14].icell.Ien VPWR.t1672 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2373 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t64 VGND.t722 VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2374 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t11 VGND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t63 VGND.t2069 VGND.t2068 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2376 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t253 VGND.t2681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[15].XIC[2].icell.Ien VPWR.t663 VPWR.t665 VPWR.t664 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2378 XThC.Tn[3].t4 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2379 VPWR.t1243 XThR.Tn[0].t61 XA.XIR[1].XIC[4].icell.PUM VPWR.t1242 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2380 XA.XIR[13].XIC_15.icell.PUM VPWR.t661 XA.XIR[13].XIC_15.icell.Ien VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2381 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t65 VPWR.t1384 VPWR.t1383 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2382 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t64 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2383 VGND.t1601 XThC.Tn[6].t39 XA.XIR[7].XIC[6].icell.PDM VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2384 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t131 VGND.t1243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2385 VPWR.t1527 XThR.Tn[4].t60 XA.XIR[5].XIC[4].icell.PUM VPWR.t1526 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2386 VPWR.t245 XThR.Tn[8].t66 XA.XIR[9].XIC[1].icell.PUM VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2387 VGND.t1233 XThC.Tn[7].t33 XA.XIR[6].XIC[7].icell.PDM VGND.t1232 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2388 VPWR.t1911 bias[0].t0 Vbias.t5 VPWR.t1210 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X2389 XThC.XTB5.A data[0].t3 VGND.t606 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2390 VPWR.t660 VPWR.t658 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t659 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2391 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t65 VPWR.t1073 VPWR.t1072 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2392 VPWR.t1147 XThR.XTB4.Y.t15 XThR.Tn[11].t2 VPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2393 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t65 XA.XIR[6].XIC[7].icell.Ien VGND.t723 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2394 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[9].XIC[1].icell.Ien VPWR.t1827 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2395 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t656 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t657 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2396 VPWR.t998 XThR.Tn[2].t61 XA.XIR[3].XIC[5].icell.PUM VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2397 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t653 VPWR.t655 VPWR.t654 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2398 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t38 XA.XIR[3].XIC[5].icell.Ien VPWR.t378 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2399 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t66 VPWR.t1061 VPWR.t1060 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2400 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t97 VGND.t1062 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2401 VGND.t2434 XThR.XTBN.Y a_n997_715# VGND.t2433 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2402 a_n997_2891# XThR.XTBN.Y VGND.t2432 VGND.t2431 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2403 VGND.t1356 VGND.t1354 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2404 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t66 VGND.t654 VGND.t653 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2405 VGND.t2611 XThC.Tn[3].t37 XA.XIR[12].XIC[3].icell.PDM VGND.t2610 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2406 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t62 VPWR.t1284 VPWR.t1283 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2407 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2043 VGND.t801 VGND.t800 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2408 VGND.t428 XThC.Tn[4].t39 XA.XIR[15].XIC[4].icell.PDM VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2409 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[3].icell.Ien VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2410 VGND.t803 VPWR.t2044 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t802 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2411 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t58 XA.XIR[7].XIC_15.icell.Ien VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2412 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t59 VGND.t1957 VGND.t1956 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2413 XA.XIR[15].XIC[4].icell.PDM VPWR.t2045 XA.XIR[15].XIC[4].icell.Ien VGND.t804 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2414 XThR.Tn[11].t3 XThR.XTB4.Y.t16 a_n997_2667# VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2415 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2046 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t805 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2416 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t67 VGND.t284 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2417 VGND.t438 XThC.Tn[5].t39 XA.XIR[2].XIC[5].icell.PDM VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2418 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t43 VGND.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2419 VPWR.t201 XThC.XTB2.Y XThC.Tn[9].t0 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2420 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t3 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2421 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t62 XA.XIR[2].XIC[5].icell.Ien VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2422 VGND.t2613 XThC.Tn[3].t38 XA.XIR[9].XIC[3].icell.PDM VGND.t2612 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2423 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t63 VGND.t453 VGND.t452 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2424 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t181 VGND.t1814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2425 VPWR.t1835 XThC.XTBN.Y.t100 XThC.Tn[8].t0 VPWR.t1834 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2426 VPWR.t1245 XThR.Tn[0].t62 XA.XIR[1].XIC[0].icell.PUM VPWR.t1244 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2427 VGND.t1235 XThC.Tn[7].t34 XA.XIR[3].XIC[7].icell.PDM VGND.t1234 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2428 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t239 VGND.t2412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2429 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[14].icell.Ien VGND.t1147 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2430 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t1118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2431 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2432 VPWR.t1529 XThR.Tn[4].t61 XA.XIR[5].XIC[0].icell.PUM VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2433 VPWR.t652 VPWR.t650 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t651 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2434 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t63 XA.XIR[3].XIC[7].icell.Ien VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2435 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t8 VPWR.t1728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2436 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t40 XA.XIR[5].XIC[13].icell.Ien VPWR.t1570 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2437 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t648 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t649 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2438 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t68 VPWR.t1063 VPWR.t1062 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2439 XThR.Tn[7].t0 XThR.XTBN.Y VPWR.t1727 VPWR.t1726 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2440 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t64 VPWR.t209 VPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2441 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t645 VPWR.t647 VPWR.t646 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2442 VGND.t1353 VGND.t1351 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2443 XThC.Tn[9].t8 XThC.XTBN.Y.t101 VPWR.t1836 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2444 XThR.Tn[1].t9 XThR.XTBN.Y VGND.t2430 VGND.t2429 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2445 VGND.t2259 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t2258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2446 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t123 VGND.t1192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2447 VPWR.t1837 XThC.XTBN.Y.t102 XThC.Tn[11].t10 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2448 VPWR.t1871 XThR.XTB6.Y a_n1049_5611# VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2449 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t69 VGND.t198 VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2450 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t2 VGND.t1291 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2451 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t69 VGND.t603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2452 VPWR.t71 XThR.Tn[10].t65 XA.XIR[11].XIC[7].icell.PUM VPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2453 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t60 VGND.t1959 VGND.t1958 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2454 VGND.t2331 XThC.Tn[12].t38 XA.XIR[13].XIC[12].icell.PDM VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2455 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[11].XIC[7].icell.Ien VPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2456 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t90 VGND.t1047 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2457 XA.XIR[0].XIC[13].icell.PDM VGND.t1348 VGND.t1350 VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2458 VGND.t1094 XThC.Tn[0].t40 XA.XIR[2].XIC[0].icell.PDM VGND.t1093 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2459 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t66 XA.XIR[13].XIC[12].icell.Ien VGND.t1151 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2460 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t63 VPWR.t249 VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2461 VGND.t2261 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t2260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2462 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t64 XA.XIR[2].XIC[0].icell.Ien VGND.t454 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2463 VGND.t2148 XThC.Tn[13].t41 XA.XIR[0].XIC[13].icell.PDM VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2464 VGND.t2263 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t2262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2465 XThC.Tn[2].t4 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2466 VPWR.t1199 VGND.t2703 XA.XIR[0].XIC[9].icell.PUM VPWR.t1198 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2467 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t63 XA.XIR[0].XIC[13].icell.Ien VGND.t1485 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2468 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t39 XA.XIR[0].XIC[9].icell.Ien VPWR.t313 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2469 VGND.t1215 XThR.XTB7.B XThR.XTB4.Y.t1 VGND.t1214 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 VGND.t2265 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t2264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2471 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t64 VPWR.t1034 VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2472 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t66 VGND.t85 VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2473 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t69 VPWR.t1065 VPWR.t1064 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2474 VGND.t2267 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t2266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2475 VGND.t753 XThR.XTB1.Y.t16 XThR.Tn[0].t2 VGND.t752 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2476 VGND.t355 XThC.Tn[9].t40 XA.XIR[11].XIC[9].icell.PDM VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2477 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t120 VGND.t1177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2478 VPWR.t73 XThR.Tn[10].t67 XA.XIR[11].XIC[11].icell.PUM VPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2479 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t64 XA.XIR[11].XIC[9].icell.Ien VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2480 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t1516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2481 VPWR.t520 XThR.Tn[7].t59 XA.XIR[8].XIC[7].icell.PUM VPWR.t519 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2482 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t40 XA.XIR[5].XIC[6].icell.Ien VPWR.t1266 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2483 VGND.t2269 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t2268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2484 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[11].XIC[11].icell.Ien VPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2485 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t112 VGND.t1119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2486 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t65 VPWR.t211 VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2487 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[8].XIC[7].icell.Ien VPWR.t529 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2488 a_8739_9569# XThC.XTBN.Y.t104 VGND.t2509 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2489 XA.XIR[0].XIC[11].icell.PDM VGND.t1345 VGND.t1347 VGND.t1346 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2490 XA.XIR[12].XIC_15.icell.PUM VPWR.t643 XA.XIR[12].XIC_15.icell.Ien VPWR.t644 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2491 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t65 VPWR.t251 VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XThC.Tn[6].t0 XThC.XTB7.Y VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2493 VPWR.t1286 XThR.Tn[3].t64 XA.XIR[4].XIC[4].icell.PUM VPWR.t1285 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2494 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t68 VPWR.t371 VPWR.t370 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2495 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t70 VPWR.t175 VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2496 VGND.t747 XThC.Tn[11].t40 XA.XIR[0].XIC[11].icell.PDM VGND.t746 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2497 VGND.t2271 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t2270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2498 VGND.t2511 XThC.XTBN.Y.t105 XThC.Tn[7].t4 VGND.t2510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2499 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t1784 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2500 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t40 XA.XIR[4].XIC[4].icell.Ien VPWR.t341 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2501 VPWR.t59 XThR.Tn[10].t68 XA.XIR[11].XIC[2].icell.PUM VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2502 VPWR.t213 XThR.Tn[5].t66 XA.XIR[6].XIC[14].icell.PUM VPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2503 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t65 XA.XIR[0].XIC[11].icell.Ien VGND.t1100 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2504 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[7].icell.Ien VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2505 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[11].XIC[2].icell.Ien VPWR.t1162 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2506 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t62 VPWR.t1579 VPWR.t1578 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2507 VPWR.t642 VPWR.t640 XA.XIR[9].XIC_15.icell.PUM VPWR.t641 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2508 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[6].XIC[14].icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2509 XThC.Tn[12].t4 XThC.XTB5.Y a_9827_9569# VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2510 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t224 VGND.t2236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2511 XA.XIR[0].XIC[2].icell.PDM VGND.t1342 VGND.t1344 VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2512 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t66 VPWR.t253 VPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2513 XA.XIR[9].XIC_15.icell.PUM VPWR.t638 XA.XIR[9].XIC_15.icell.Ien VPWR.t639 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2514 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t4 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2515 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t211 VGND.t2010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2516 VGND.t2273 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t2272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2517 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t66 VPWR.t538 VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2518 VGND.t2275 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t2274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2519 VGND.t1288 XThC.Tn[2].t40 XA.XIR[0].XIC[2].icell.PDM VGND.t1287 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2520 XThR.Tn[13].t5 XThR.XTB6.Y VPWR.t1870 VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2521 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t60 VGND.t1914 VGND.t1913 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2522 VGND.t2297 XThC.Tn[8].t39 XA.XIR[5].XIC[8].icell.PDM VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2523 VGND.t2277 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t2276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2524 VGND.t2279 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t2278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2525 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[2].icell.Ien VGND.t1101 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2526 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t67 XA.XIR[5].XIC[8].icell.Ien VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2527 VGND.t357 XThC.Tn[9].t41 XA.XIR[8].XIC[9].icell.PDM VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2528 VGND.t440 XThC.Tn[5].t40 XA.XIR[1].XIC[5].icell.PDM VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2529 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t69 XA.XIR[8].XIC[9].icell.Ien VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2530 VPWR.t1388 XThR.Tn[7].t61 XA.XIR[8].XIC[11].icell.PUM VPWR.t1387 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2531 VGND.t2512 XThC.XTBN.Y.t107 a_7875_9569# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2532 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t69 VGND.t78 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2533 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[8].XIC[11].icell.Ien VPWR.t571 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2534 XA.XIR[7].XIC_15.icell.PDM VPWR.t2047 VGND.t807 VGND.t806 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2535 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t61 XA.XIR[1].XIC[5].icell.Ien VGND.t1960 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2536 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t2048 VGND.t809 VGND.t808 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2537 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t7 VGND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2538 VGND.t2281 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t2280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2539 VGND.t388 XThC.Tn[4].t41 XA.XIR[11].XIC[4].icell.PDM VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2540 VGND.t811 VPWR.t2049 XA.XIR[7].XIC_15.icell.PDM VGND.t810 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2541 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t373 VPWR.t372 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2542 VGND.t813 VPWR.t2050 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t812 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2543 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t141 VGND.t1470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2544 VPWR.t1288 XThR.Tn[3].t65 XA.XIR[4].XIC[0].icell.PUM VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2545 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2546 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t67 XA.XIR[11].XIC[4].icell.Ien VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2547 a_8963_9569# XThC.XTBN.Y.t108 VGND.t2513 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2548 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[5].XIC[1].icell.Ien VPWR.t1828 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2549 VPWR.t1390 XThR.Tn[7].t62 XA.XIR[8].XIC[2].icell.PUM VPWR.t1389 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2550 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t2051 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t814 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2551 VPWR.t385 XThR.Tn[2].t65 XA.XIR[3].XIC[14].icell.PUM VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2552 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[4].XIC[0].icell.Ien VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2553 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t636 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t637 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2554 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t68 VPWR.t215 VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2555 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[8].XIC[2].icell.Ien VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2556 XA.XIR[0].XIC[6].icell.PDM VGND.t1339 VGND.t1341 VGND.t1340 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2557 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t40 XA.XIR[3].XIC[14].icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2558 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t63 VPWR.t1581 VPWR.t1580 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2559 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t633 VPWR.t635 VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2560 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t375 VPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2561 VGND.t1603 XThC.Tn[6].t41 XA.XIR[0].XIC[6].icell.PDM VGND.t1602 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2562 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t66 VPWR.t1290 VPWR.t1289 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2563 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t68 VGND.t739 VGND.t738 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2564 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2052 VGND.t816 VGND.t815 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2565 VPWR.t1418 XThR.Tn[1].t62 XA.XIR[2].XIC[12].icell.PUM VPWR.t1417 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2566 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[6].icell.Ien VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2567 VPWR.t1036 XThR.Tn[0].t68 XA.XIR[1].XIC[13].icell.PUM VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2568 XThC.Tn[11].t9 XThC.XTBN.Y.t109 VPWR.t1785 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2569 VGND.t2283 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t2282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2570 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[2].XIC[12].icell.Ien VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2571 VPWR.t1583 XThR.Tn[4].t64 XA.XIR[5].XIC[13].icell.PUM VPWR.t1582 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2572 XThR.Tn[6].t5 XThR.XTBN.Y a_n1049_5317# VPWR.t1723 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2573 VGND.t818 VPWR.t2053 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t817 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2574 VPWR.t632 VPWR.t630 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t631 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2575 VPWR.t1822 XThC.XTB4.Y.t16 XThC.Tn[11].t0 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2576 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2577 VGND.t2285 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t2284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2578 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2054 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t819 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2579 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t66 VPWR.t387 VPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2580 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t628 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t629 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2581 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t741 VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2582 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t63 VGND.t1916 VGND.t1915 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2583 VGND.t2379 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t2378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2584 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2055 VGND.t821 VGND.t820 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2585 VGND.t249 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2586 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t625 VPWR.t627 VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2587 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t213 VGND.t2021 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2588 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2589 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[3].icell.Ien VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2590 VGND.t390 XThC.Tn[4].t42 XA.XIR[8].XIC[4].icell.PDM VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2591 VGND.t823 VPWR.t2056 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t822 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2592 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t147 VGND.t1501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2593 VGND.t2333 XThC.Tn[12].t40 XA.XIR[12].XIC[12].icell.PDM VGND.t2332 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2594 VPWR.t604 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2595 VGND.t1122 XThC.Tn[0].t42 XA.XIR[1].XIC[0].icell.PDM VGND.t1121 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2596 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[4].icell.Ien VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2597 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2057 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t824 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2598 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t71 XA.XIR[12].XIC[12].icell.Ien VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2599 VGND.t2428 XThR.XTBN.Y a_n997_1803# VGND.t2427 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2600 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t63 XA.XIR[1].XIC[0].icell.Ien VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2601 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t64 VGND.t1963 VGND.t1962 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2602 a_3773_9615# XThC.XTB2.Y VPWR.t199 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2603 VGND.t2381 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t2380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2604 VGND.t2321 XThC.Tn[14].t41 XA.XIR[2].XIC[14].icell.PDM VGND.t2320 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2605 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t73 VGND.t434 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2606 VGND.t2335 XThC.Tn[12].t41 XA.XIR[9].XIC[12].icell.PDM VGND.t2334 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2607 VPWR.t1682 XThR.Tn[1].t65 XA.XIR[2].XIC[10].icell.PUM VPWR.t1681 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2608 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t67 XA.XIR[2].XIC[14].icell.Ien VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2609 VPWR.t1149 XThR.XTB4.Y.t17 XThR.Tn[11].t4 VPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2610 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[2].XIC[10].icell.Ien VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2611 a_n997_715# XThR.XTBN.Y VGND.t2426 VGND.t2425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2612 VGND.t2383 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t2382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2613 VPWR.t574 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 XThR.Tn[14].t1 XThR.XTB7.Y VPWR.t125 VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2615 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t68 VPWR.t1880 VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2616 VGND.t2385 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t2384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2617 VGND.t2514 XThC.XTBN.Y.t110 XThC.Tn[3].t9 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2618 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t1714 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2619 XThC.Tn[1].t0 XThC.XTB2.Y VGND.t234 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2620 VPWR.t196 XThC.XTBN.A XThC.XTBN.Y.t0 VPWR.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2621 VGND.t2387 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t2386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2622 VPWR.t1067 XThR.Tn[9].t71 XA.XIR[10].XIC[8].icell.PUM VPWR.t1066 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2623 VGND.t2389 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t2388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2624 XThR.Tn[2].t1 XThR.XTB3.Y.t16 VGND.t1292 VGND.t714 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2625 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t40 XA.XIR[10].XIC[8].icell.Ien VPWR.t1326 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2626 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t64 VPWR.t1392 VPWR.t1391 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2627 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t182 VGND.t1815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2628 VGND.t2391 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t2390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2629 VGND.t1338 VGND.t1336 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 VGND.t2393 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t2392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2631 VPWR.t1038 XThR.Tn[0].t69 XA.XIR[1].XIC[6].icell.PUM VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2632 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t70 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2633 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t4 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2634 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t80 VGND.t732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2635 a_3299_10575# XThC.XTB7.B VGND.t1794 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2636 VPWR.t1585 XThR.Tn[4].t65 XA.XIR[5].XIC[6].icell.PUM VPWR.t1584 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2637 VGND.t2424 XThR.XTBN.Y XThR.Tn[6].t8 VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2638 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t72 VPWR.t1069 VPWR.t1068 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2639 VGND.t2395 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t2394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2640 VGND.t2397 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t2396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2641 VGND.t2399 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t2398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2642 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t67 VGND.t1153 VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2643 VGND.t2401 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t2400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VPWR.t1684 XThR.Tn[1].t66 XA.XIR[2].XIC[5].icell.PUM VPWR.t1683 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2645 VPWR.t1786 XThC.XTBN.Y.t111 XThC.Tn[10].t11 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2646 VGND.t2150 XThC.Tn[13].t42 XA.XIR[14].XIC[13].icell.PDM VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2647 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[9].icell.Ien VGND.t1917 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2648 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[2].XIC[5].icell.Ien VPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2649 VPWR.t1075 XThR.Tn[13].t68 XA.XIR[14].XIC[9].icell.PUM VPWR.t1074 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2650 VGND.t2515 XThC.XTBN.Y.t112 a_8963_9569# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2651 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t70 VGND.t1104 VGND.t1103 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2652 VGND.t2403 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t2402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2653 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t67 XA.XIR[14].XIC[13].icell.Ien VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2654 VPWR.t180 XThC.XTB5.A a_5155_10571# VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2655 VPWR.t48 XThC.XTB7.Y XThC.Tn[14].t0 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2656 XThR.Tn[1].t8 XThR.XTBN.Y VGND.t2422 VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t69 VPWR.t1882 VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2658 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t66 VGND.t2196 VGND.t2195 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2659 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t42 XA.XIR[14].XIC[9].icell.Ien VPWR.t1399 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2660 VGND.t2405 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t2404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2661 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t66 VPWR.t1394 VPWR.t1393 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2662 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t72 VGND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2663 VPWR.t1804 XThC.XTB7.A XThC.XTB3.Y.t2 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2664 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t68 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t219 VGND.t2230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2666 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t20 VGND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2667 XThR.Tn[8].t8 XThR.XTBN.Y VPWR.t1725 VPWR.t1724 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 XThR.Tn[5].t0 XThR.XTBN.Y a_n1049_5611# VPWR.t1723 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2669 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t3 VGND.t716 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2670 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2058 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t825 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2671 VPWR.t1071 XThR.Tn[9].t73 XA.XIR[10].XIC[3].icell.PUM VPWR.t1070 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2672 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2673 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t40 XA.XIR[10].XIC[3].icell.Ien VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2674 XA.XIR[5].XIC_15.icell.PUM VPWR.t623 XA.XIR[5].XIC_15.icell.Ien VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2675 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t67 VPWR.t1396 VPWR.t1395 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2676 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t2347 VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2677 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t21 VGND.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2678 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t60 VGND.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2679 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t4 VPWR.t1722 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2680 VPWR.t1040 XThR.Tn[0].t71 XA.XIR[1].XIC[1].icell.PUM VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2681 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t69 VGND.t657 VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2682 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t71 VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2683 VGND.t704 XThC.Tn[7].t37 XA.XIR[2].XIC[7].icell.PDM VGND.t703 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2684 VPWR.t1587 XThR.Tn[4].t67 XA.XIR[5].XIC[1].icell.PUM VPWR.t1586 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2685 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t70 VPWR.t217 VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2686 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t69 VGND.t1155 VGND.t1154 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2687 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t5 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2688 VPWR.t1917 XThR.Tn[3].t67 XA.XIR[4].XIC[13].icell.PUM VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2689 VGND.t827 VPWR.t2059 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t826 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2690 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t42 XA.XIR[1].XIC[12].icell.Ien VPWR.t1680 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2691 VGND.t161 XThC.Tn[10].t41 XA.XIR[15].XIC[10].icell.PDM VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2692 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[7].icell.Ien VGND.t2671 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2693 VGND.t749 XThC.Tn[11].t42 XA.XIR[14].XIC[11].icell.PDM VGND.t748 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2694 VPWR.t1129 XThR.XTB7.B XThR.XTB3.Y.t0 VPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t68 VPWR.t1686 VPWR.t1685 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2696 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t43 XA.XIR[4].XIC[13].icell.Ien VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2697 XA.XIR[15].XIC[10].icell.PDM VPWR.t2060 XA.XIR[15].XIC[10].icell.Ien VGND.t828 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2698 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2061 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t829 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2699 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t70 XA.XIR[14].XIC[11].icell.Ien VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2700 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t605 VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2701 VGND.t561 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2702 VPWR.t606 XThC.XTB3.Y.t16 XThC.Tn[10].t6 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2703 VPWR.t1787 XThC.XTBN.Y.t114 XThC.Tn[14].t9 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2704 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t68 VPWR.t1589 VPWR.t1588 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2705 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t71 VGND.t660 VGND.t659 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2706 VGND.t1335 VGND.t1333 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2707 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t70 VGND.t1157 VGND.t1156 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2708 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2062 VGND.t831 VGND.t830 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2709 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t193 VGND.t1902 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2710 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t247 VGND.t2638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2711 VGND.t2620 XThC.Tn[1].t41 XA.XIR[15].XIC[1].icell.PDM VGND.t2619 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2712 VGND.t2420 XThR.XTBN.Y XThR.Tn[0].t8 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2713 VGND.t1290 XThC.Tn[2].t42 XA.XIR[14].XIC[2].icell.PDM VGND.t1289 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2714 VGND.t833 VPWR.t2063 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t832 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2715 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t82 VGND.t914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2716 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t68 XA.XIR[7].XIC[4].icell.Ien VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2717 VGND.t1051 XThC.XTB3.Y.t17 XThC.Tn[2].t3 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2718 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t72 VGND.t1106 VGND.t1105 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2719 XA.XIR[15].XIC[1].icell.PDM VPWR.t2064 XA.XIR[15].XIC[1].icell.Ien VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2720 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t72 XA.XIR[14].XIC[2].icell.Ien VGND.t661 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2721 XThR.Tn[10].t5 XThR.XTBN.Y VPWR.t1721 VPWR.t1720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2722 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t69 VGND.t2198 VGND.t2197 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2723 XA.XIR[0].XIC_15.icell.PDM VPWR.t2065 VGND.t2590 VGND.t2589 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2724 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t162 VGND.t1652 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2725 VGND.t563 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2726 VGND.t2323 XThC.Tn[14].t42 XA.XIR[1].XIC[14].icell.PDM VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2727 VPWR.t1315 XThC.XTB6.Y a_5949_9615# VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2728 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t2249 VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2729 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t94 VGND.t1052 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2730 VGND.t2418 XThR.XTBN.Y a_n997_3755# VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2731 VGND.t2592 VPWR.t2066 XA.XIR[0].XIC_15.icell.PDM VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2732 VPWR.t1630 data[3].t1 XThC.XTBN.A VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2733 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t3 VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2734 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t408 VPWR.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2735 XThC.Tn[3].t8 XThC.XTBN.Y.t115 VGND.t2516 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2736 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t69 XA.XIR[1].XIC[14].icell.Ien VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2737 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t77 VGND.t702 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2738 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t73 XA.XIR[0].XIC_15.icell.Ien VGND.t1107 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2739 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[1].XIC[10].icell.Ien VPWR.t150 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2740 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t70 VPWR.t1688 VPWR.t1687 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2741 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t2 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2742 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2743 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t71 VGND.t1159 VGND.t1158 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2744 XThR.Tn[13].t4 XThR.XTB6.Y VPWR.t1869 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2745 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t188 VGND.t1883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2746 VGND.t386 XThC.Tn[6].t42 XA.XIR[14].XIC[6].icell.PDM VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2747 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t1167 VPWR.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2748 VPWR.t566 XThR.Tn[11].t70 XA.XIR[12].XIC[4].icell.PUM VPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2749 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t73 XA.XIR[14].XIC[6].icell.Ien VGND.t662 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2750 VGND.t1332 VGND.t1330 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2751 VGND.t565 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2752 VPWR.t1919 XThR.Tn[3].t68 XA.XIR[4].XIC[6].icell.PUM VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2753 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t218 VGND.t2229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2754 VPWR.t1448 XThC.XTB1.Y.t18 XThC.Tn[8].t4 VPWR.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2755 VPWR.t540 XThR.Tn[6].t67 XA.XIR[7].XIC[7].icell.PUM VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2756 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[4].XIC[6].icell.Ien VPWR.t340 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2757 VGND.t2337 XThC.Tn[12].t43 XA.XIR[5].XIC[12].icell.PDM VGND.t2336 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2758 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t27 VGND.t173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2759 VPWR.t219 XThR.Tn[5].t71 XA.XIR[6].XIC[8].icell.PUM VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2760 VGND.t1313 XThR.XTB5.Y XThR.Tn[4].t0 VGND.t1312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2761 XThC.Tn[10].t10 XThC.XTBN.Y.t116 VPWR.t1669 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2762 VGND.t2311 XThC.XTBN.Y.t117 XThC.Tn[6].t8 VGND.t2310 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2763 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t70 VPWR.t1591 VPWR.t1590 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2764 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[7].XIC[7].icell.Ien VPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2765 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t72 XA.XIR[5].XIC[12].icell.Ien VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2766 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[6].XIC[8].icell.Ien VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2767 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t68 VPWR.t542 VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2768 VGND.t567 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2769 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t72 VGND.t1809 VGND.t1808 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2770 VGND.t442 XThC.Tn[5].t42 XA.XIR[13].XIC[5].icell.PDM VGND.t441 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2771 VPWR.t1823 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2772 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t43 XA.XIR[1].XIC[5].icell.Ien VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2773 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC[5].icell.Ien VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2774 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t69 VGND.t2685 VGND.t2684 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2775 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t71 VPWR.t1690 VPWR.t1689 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2776 VGND.t569 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2777 XThR.Tn[6].t4 XThR.XTBN.Y a_n1049_5317# VPWR.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2778 VPWR.t568 XThR.Tn[11].t71 XA.XIR[12].XIC[0].icell.PUM VPWR.t567 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2779 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t69 VGND.t725 VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2780 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t4 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2781 VGND.t1728 XThC.Tn[8].t42 XA.XIR[4].XIC[8].icell.PDM VGND.t1727 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2782 VGND.t571 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 VGND.t2313 XThC.XTBN.Y.t118 a_10915_9569# VGND.t2312 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2784 VGND.t573 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2785 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t71 XA.XIR[4].XIC[8].icell.Ien VGND.t1745 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2786 VPWR.t622 VPWR.t620 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t621 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2787 VGND.t1932 XThC.Tn[9].t43 XA.XIR[7].XIC[9].icell.PDM VGND.t1931 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2788 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t618 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t619 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2789 VPWR.t544 XThR.Tn[6].t70 XA.XIR[7].XIC[11].icell.PUM VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2790 XThC.Tn[1].t4 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2791 VPWR.t1884 XThR.Tn[2].t71 XA.XIR[3].XIC[8].icell.PUM VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2792 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t43 XA.XIR[7].XIC[11].icell.Ien VPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2793 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t615 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2794 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t234 VGND.t2344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2795 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t43 XA.XIR[3].XIC[8].icell.Ien VPWR.t1328 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2796 VGND.t575 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2797 VGND.t706 XThC.Tn[7].t39 XA.XIR[1].XIC[7].icell.PDM VGND.t705 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2798 VPWR.t1921 XThR.Tn[3].t70 XA.XIR[4].XIC[1].icell.PUM VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2799 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t145 VGND.t1489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2800 XThC.Tn[14].t8 XThC.XTBN.Y.t120 VPWR.t1670 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2801 VGND.t577 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2802 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t71 VPWR.t1923 VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2803 VGND.t579 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2804 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t72 XA.XIR[1].XIC[7].icell.Ien VGND.t1948 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2805 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t42 XA.XIR[4].XIC[1].icell.Ien VPWR.t1829 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2806 VPWR.t546 XThR.Tn[6].t71 XA.XIR[7].XIC[2].icell.PUM VPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2807 VPWR.t1408 XThR.Tn[1].t73 XA.XIR[2].XIC[14].icell.PUM VPWR.t1407 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2808 VPWR.t221 XThR.Tn[5].t73 XA.XIR[6].XIC[3].icell.PUM VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2809 VPWR.t614 VPWR.t612 XA.XIR[1].XIC_15.icell.PUM VPWR.t613 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2810 VGND.t2416 XThR.XTBN.Y a_n997_715# VGND.t2415 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2811 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t43 XA.XIR[7].XIC[2].icell.Ien VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2812 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t72 VPWR.t1337 VPWR.t1336 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2813 VPWR.t611 VPWR.t609 XA.XIR[5].XIC_15.icell.PUM VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2814 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t43 XA.XIR[2].XIC[14].icell.Ien VPWR.t527 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2815 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t41 XA.XIR[6].XIC[3].icell.Ien VPWR.t223 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2816 VPWR.t123 XThR.XTB7.Y XThR.Tn[14].t0 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2817 VGND.t1329 VGND.t1327 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2818 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t72 VPWR.t1886 VPWR.t1885 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2819 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t72 VPWR.t1386 VPWR.t1385 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2820 VGND.t581 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2821 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t73 VGND.t1811 VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2822 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t72 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2823 XThR.XTB6.A data[5].t5 VGND.t461 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2824 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t100 VGND.t1066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2825 XThR.Tn[0].t4 XThR.XTBN.Y a_n1049_8581# VPWR.t1718 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2826 a_5949_9615# XThC.XTB6.Y VPWR.t1314 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2827 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t233 VGND.t2343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2828 VGND.t163 XThC.Tn[10].t43 XA.XIR[11].XIC[10].icell.PDM VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2829 VGND.t2314 XThC.XTBN.Y.t121 a_10051_9569# VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2830 VGND.t583 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2831 VGND.t1124 XThC.Tn[0].t43 XA.XIR[13].XIC[0].icell.PDM VGND.t1123 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2832 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t73 XA.XIR[13].XIC[0].icell.Ien VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2833 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t72 XA.XIR[11].XIC[10].icell.Ien VGND.t742 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2834 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t72 VGND.t2687 VGND.t2686 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2835 VPWR.t1671 XThC.XTBN.Y.t122 XThC.Tn[11].t8 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2836 VGND.t251 XThC.Tn[3].t42 XA.XIR[4].XIC[3].icell.PDM VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2837 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t73 VGND.t82 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2838 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t73 VGND.t1900 VGND.t1899 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2839 VGND.t2315 XThC.XTBN.Y.t123 a_7651_9569# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2840 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2067 VGND.t2594 VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
X2841 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t10 VGND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2842 XThR.Tn[2].t7 XThR.XTBN.Y VGND.t2414 VGND.t2413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2843 VGND.t2622 XThC.Tn[1].t43 XA.XIR[11].XIC[1].icell.PDM VGND.t2621 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2844 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t73 XA.XIR[4].XIC[3].icell.Ien VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2845 VPWR.t121 XThR.XTB7.Y a_n1049_5317# VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2846 VGND.t392 XThC.Tn[4].t43 XA.XIR[7].XIC[4].icell.PDM VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2847 VGND.t2596 VPWR.t2068 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2848 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2849 VGND.t585 Vbias.t260 XA.XIR[15].XIC_15.icell.SM VGND.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2850 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t7 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 VPWR.t1717 XThR.XTBN.Y XThR.Tn[12].t8 VPWR.t1716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2852 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t73 XA.XIR[11].XIC[1].icell.Ien VGND.t743 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2853 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2069 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t2597 sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.14 ps=1.56 w=0.5 l=0.15
X2854 VPWR.t1888 XThR.Tn[2].t73 XA.XIR[3].XIC[3].icell.PUM VPWR.t1887 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2855 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t64 VGND.t551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2856 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[3].XIC[3].icell.Ien VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X2857 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t122 VGND.t1186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2858 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t73 VPWR.t1925 VPWR.t1924 sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2859 VGND.t587 Vbias.t261 XA.XIR[13].XIC[2].icell.SM VGND.t586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2860 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t69 VGND.t1920 VGND.t1919 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.56 as=0.075 ps=0.8 w=0.5 l=0.15
R0 VGND.n2824 VGND.n7 32072.7
R1 VGND.n3002 VGND.n3001 21075.4
R2 VGND.n2860 VGND.n2828 13477
R3 VGND.n2828 VGND.n2827 11635.6
R4 VGND.n2995 VGND.n2994 9309.26
R5 VGND.n2893 VGND.n2860 9223.7
R6 VGND.n2894 VGND.n2893 9223.7
R7 VGND.n2947 VGND.n34 9223.7
R8 VGND.n2980 VGND.n2947 9223.7
R9 VGND.n2981 VGND.n2980 8197.04
R10 VGND.n1508 VGND.n1507 7387.65
R11 VGND.n1507 VGND.n1506 7387.65
R12 VGND.n2818 VGND.n147 7387.65
R13 VGND.n3000 VGND.n2999 7387.65
R14 VGND.n2999 VGND.n2998 7387.65
R15 VGND.n2998 VGND.n2997 7387.65
R16 VGND.n2997 VGND.n2996 7387.65
R17 VGND.n2996 VGND.n2995 7387.65
R18 VGND.n2823 VGND.n2818 7048.53
R19 VGND.n1510 VGND.t2244 6324.96
R20 VGND.n3001 VGND.n3000 5925.05
R21 VGND.n2894 VGND.n34 5231.11
R22 VGND.n1290 VGND.t759 5138.54
R23 VGND.n2994 VGND.n2993 5074.71
R24 VGND.n2827 VGND.n7 4937.78
R25 VGND.n3001 VGND.n7 4804.6
R26 VGND.n1110 VGND.n578 4542.17
R27 VGND.n2824 VGND.n2823 4343.1
R28 VGND.n2414 VGND.n273 4295.6
R29 VGND.n2994 VGND 4240.58
R30 VGND.n2415 VGND.n2414 3486.29
R31 VGND.n2416 VGND.n2415 3486.29
R32 VGND.n2417 VGND.n2416 3486.29
R33 VGND.n2418 VGND.n2417 3486.29
R34 VGND.n2419 VGND.n2418 3486.29
R35 VGND.n2420 VGND.n2419 3486.29
R36 VGND.n2421 VGND.n2420 3486.29
R37 VGND.n2422 VGND.n2421 3486.29
R38 VGND.n2423 VGND.n2422 3486.29
R39 VGND.n2424 VGND.n2423 3486.29
R40 VGND.n2425 VGND.n2424 3486.29
R41 VGND.n2426 VGND.n2425 3486.29
R42 VGND.n2427 VGND.n2426 3486.29
R43 VGND.n2427 VGND.n32 3486.29
R44 VGND.n2983 VGND.n32 3486.29
R45 VGND.n2983 VGND.n2982 3486.29
R46 VGND.n1294 VGND.n1292 3417.39
R47 VGND.n1294 VGND.n1293 3417.39
R48 VGND.n1512 VGND.n1511 3417.39
R49 VGND.n960 VGND.n580 3417.39
R50 VGND.n635 VGND.n177 3417.39
R51 VGND.n2817 VGND.n114 3417.39
R52 VGND.n2826 VGND.n2825 3417.39
R53 VGND.n1293 VGND.n578 3273.91
R54 VGND.n961 VGND.n579 3265.22
R55 VGND.n2824 VGND.n114 2756.52
R56 VGND.n2982 VGND.n2981 2723.39
R57 VGND.n2860 VGND.t2466 2655.17
R58 VGND.n2893 VGND.t2490 2655.17
R59 VGND.n2818 VGND.n2817 2517.39
R60 VGND.n2821 VGND.n5 2229.43
R61 VGND.n3003 VGND.n5 2229.43
R62 VGND.n3003 VGND.n6 2229.43
R63 VGND.n2821 VGND.n6 2229.43
R64 VGND.n1292 VGND.n1291 2130.43
R65 VGND.n2827 VGND.n2826 2082.61
R66 VGND VGND.n34 1997.7
R67 VGND.n2947 VGND 1997.7
R68 VGND.n2980 VGND 1997.7
R69 VGND.n1505 VGND.n147 1831.57
R70 VGND.t2423 VGND.n2894 1807.04
R71 VGND.n2978 VGND.t1906 1785.51
R72 VGND.n1506 VGND.n580 1691.3
R73 VGND.n2906 VGND.t1275 1618.39
R74 VGND.t718 VGND.n2946 1618.39
R75 VGND.t1317 VGND.n2979 1618.39
R76 VGND.n2828 VGND.t2439 1517.24
R77 VGND.n1509 VGND.n1508 1513.49
R78 VGND.n1510 VGND.n1509 1370.36
R79 VGND.n1291 VGND.n1290 1286.96
R80 VGND.n1509 VGND.t1466 1284.61
R81 VGND.n1083 VGND.t256 1268.93
R82 VGND.n1083 VGND.t178 1268.93
R83 VGND.n146 VGND.t262 1253.59
R84 VGND.t8 VGND.n146 1253.59
R85 VGND.n614 VGND.t4 1253.59
R86 VGND.t13 VGND.n614 1253.59
R87 VGND.n1021 VGND.t236 1253.59
R88 VGND.n1021 VGND.t258 1253.59
R89 VGND.n1052 VGND.t2 1253.59
R90 VGND.n1052 VGND.t176 1253.59
R91 VGND.n176 VGND.t10 1253.59
R92 VGND.t16 VGND.n176 1253.59
R93 VGND.n1505 VGND.t1397 1252.04
R94 VGND.n2823 VGND.n2822 1217.3
R95 VGND.n2906 VGND.t1657 1213.79
R96 VGND.n1111 VGND.n1110 1198.25
R97 VGND.n2993 VGND.n2992 1198.25
R98 VGND.n2946 VGND.t1656 1180.08
R99 VGND.n2985 VGND.n2984 1179.65
R100 VGND.n2490 VGND.n2489 1179.65
R101 VGND.n2429 VGND.n2428 1179.65
R102 VGND.n2312 VGND.n261 1179.65
R103 VGND.n2126 VGND.n262 1179.65
R104 VGND.n2121 VGND.n263 1179.65
R105 VGND.n2337 VGND.n264 1179.65
R106 VGND.n1952 VGND.n265 1179.65
R107 VGND.n1947 VGND.n266 1179.65
R108 VGND.n2362 VGND.n267 1179.65
R109 VGND.n1778 VGND.n268 1179.65
R110 VGND.n1773 VGND.n269 1179.65
R111 VGND.n2387 VGND.n270 1179.65
R112 VGND.n1604 VGND.n271 1179.65
R113 VGND.n2407 VGND.n272 1179.65
R114 VGND.n2413 VGND.n2412 1179.65
R115 VGND.n1232 VGND.n273 1179.65
R116 VGND.n2642 VGND.n33 1179.64
R117 VGND.n2645 VGND.n2644 1179.3
R118 VGND.n2647 VGND.n2646 1179.3
R119 VGND.n2652 VGND.n2651 1179.3
R120 VGND.n2654 VGND.n2653 1179.3
R121 VGND.n2659 VGND.n2658 1179.3
R122 VGND.n2661 VGND.n2660 1179.3
R123 VGND.n2666 VGND.n2665 1179.3
R124 VGND.n2668 VGND.n2667 1179.3
R125 VGND.n2673 VGND.n2672 1179.3
R126 VGND.n2675 VGND.n2674 1179.3
R127 VGND.n2680 VGND.n2679 1179.3
R128 VGND.n2682 VGND.n2681 1179.3
R129 VGND.n2687 VGND.n2686 1179.3
R130 VGND.n2688 VGND.n2570 1179.3
R131 VGND.n2690 VGND.n2689 1179.3
R132 VGND.n2766 VGND.n2765 1179.3
R133 VGND.n2764 VGND.n2763 1179.3
R134 VGND.n2759 VGND.n2758 1179.3
R135 VGND.n2754 VGND.n2753 1179.3
R136 VGND.n2749 VGND.n2748 1179.3
R137 VGND.n2744 VGND.n2743 1179.3
R138 VGND.n2739 VGND.n2738 1179.3
R139 VGND.n2734 VGND.n2733 1179.3
R140 VGND.n2729 VGND.n2728 1179.3
R141 VGND.n2724 VGND.n2723 1179.3
R142 VGND.n2719 VGND.n2718 1179.3
R143 VGND.n2714 VGND.n2713 1179.3
R144 VGND.n2709 VGND.n2708 1179.3
R145 VGND.n2704 VGND.n2703 1179.3
R146 VGND.n234 VGND.n233 1179.3
R147 VGND.n2488 VGND.n2487 1179.3
R148 VGND.n2483 VGND.n2482 1179.3
R149 VGND.n2478 VGND.n2477 1179.3
R150 VGND.n2473 VGND.n2472 1179.3
R151 VGND.n2468 VGND.n2467 1179.3
R152 VGND.n2463 VGND.n2462 1179.3
R153 VGND.n2458 VGND.n2457 1179.3
R154 VGND.n2453 VGND.n2452 1179.3
R155 VGND.n2448 VGND.n2447 1179.3
R156 VGND.n2443 VGND.n2442 1179.3
R157 VGND.n2438 VGND.n2437 1179.3
R158 VGND.n2433 VGND.n244 1179.3
R159 VGND.n2508 VGND.n2507 1179.3
R160 VGND.n2513 VGND.n2512 1179.3
R161 VGND.n2515 VGND.n2514 1179.3
R162 VGND.n2292 VGND.n2291 1179.3
R163 VGND.n2290 VGND.n2289 1179.3
R164 VGND.n2285 VGND.n2284 1179.3
R165 VGND.n2280 VGND.n2279 1179.3
R166 VGND.n2251 VGND.n2250 1179.3
R167 VGND.n2249 VGND.n2248 1179.3
R168 VGND.n2225 VGND.n2224 1179.3
R169 VGND.n2223 VGND.n2222 1179.3
R170 VGND.n2199 VGND.n2198 1179.3
R171 VGND.n2197 VGND.n2196 1179.3
R172 VGND.n2173 VGND.n2172 1179.3
R173 VGND.n2171 VGND.n2170 1179.3
R174 VGND.n373 VGND.n372 1179.3
R175 VGND.n371 VGND.n182 1179.3
R176 VGND.n2816 VGND.n2815 1179.3
R177 VGND.n2309 VGND.n2308 1179.3
R178 VGND.n2307 VGND.n2306 1179.3
R179 VGND.n2267 VGND.n2266 1179.3
R180 VGND.n2269 VGND.n2268 1179.3
R181 VGND.n2262 VGND.n2261 1179.3
R182 VGND.n2238 VGND.n2237 1179.3
R183 VGND.n2236 VGND.n2235 1179.3
R184 VGND.n2212 VGND.n2211 1179.3
R185 VGND.n2210 VGND.n2209 1179.3
R186 VGND.n2186 VGND.n2185 1179.3
R187 VGND.n2184 VGND.n2183 1179.3
R188 VGND.n2160 VGND.n2159 1179.3
R189 VGND.n2158 VGND.n2157 1179.3
R190 VGND.n1430 VGND.n1429 1179.3
R191 VGND.n1428 VGND.n1427 1179.3
R192 VGND.n2130 VGND.n2129 1179.3
R193 VGND.n2135 VGND.n2134 1179.3
R194 VGND.n2137 VGND.n2136 1179.3
R195 VGND.n1447 VGND.n1446 1179.3
R196 VGND.n1452 VGND.n1451 1179.3
R197 VGND.n1457 VGND.n1456 1179.3
R198 VGND.n1462 VGND.n1461 1179.3
R199 VGND.n1467 VGND.n1466 1179.3
R200 VGND.n1472 VGND.n1471 1179.3
R201 VGND.n1477 VGND.n1476 1179.3
R202 VGND.n1482 VGND.n1481 1179.3
R203 VGND.n1487 VGND.n1486 1179.3
R204 VGND.n1492 VGND.n1491 1179.3
R205 VGND.n1494 VGND.n1493 1179.3
R206 VGND.n1442 VGND.n1441 1179.3
R207 VGND.n2118 VGND.n2117 1179.3
R208 VGND.n2116 VGND.n2115 1179.3
R209 VGND.n2111 VGND.n2110 1179.3
R210 VGND.n2106 VGND.n2105 1179.3
R211 VGND.n2077 VGND.n2076 1179.3
R212 VGND.n2075 VGND.n2074 1179.3
R213 VGND.n2051 VGND.n2050 1179.3
R214 VGND.n2049 VGND.n2048 1179.3
R215 VGND.n2025 VGND.n2024 1179.3
R216 VGND.n2023 VGND.n2022 1179.3
R217 VGND.n1999 VGND.n1998 1179.3
R218 VGND.n1997 VGND.n1996 1179.3
R219 VGND.n628 VGND.n627 1179.3
R220 VGND.n626 VGND.n619 1179.3
R221 VGND.n1504 VGND.n1503 1179.3
R222 VGND.n2334 VGND.n2333 1179.3
R223 VGND.n2332 VGND.n2331 1179.3
R224 VGND.n2093 VGND.n2092 1179.3
R225 VGND.n2095 VGND.n2094 1179.3
R226 VGND.n2088 VGND.n2087 1179.3
R227 VGND.n2064 VGND.n2063 1179.3
R228 VGND.n2062 VGND.n2061 1179.3
R229 VGND.n2038 VGND.n2037 1179.3
R230 VGND.n2036 VGND.n2035 1179.3
R231 VGND.n2012 VGND.n2011 1179.3
R232 VGND.n2010 VGND.n2009 1179.3
R233 VGND.n1986 VGND.n1985 1179.3
R234 VGND.n1984 VGND.n1983 1179.3
R235 VGND.n654 VGND.n653 1179.3
R236 VGND.n652 VGND.n651 1179.3
R237 VGND.n1956 VGND.n1955 1179.3
R238 VGND.n1961 VGND.n1960 1179.3
R239 VGND.n1963 VGND.n1962 1179.3
R240 VGND.n904 VGND.n903 1179.3
R241 VGND.n909 VGND.n908 1179.3
R242 VGND.n914 VGND.n913 1179.3
R243 VGND.n919 VGND.n918 1179.3
R244 VGND.n924 VGND.n923 1179.3
R245 VGND.n929 VGND.n928 1179.3
R246 VGND.n934 VGND.n933 1179.3
R247 VGND.n939 VGND.n938 1179.3
R248 VGND.n944 VGND.n943 1179.3
R249 VGND.n949 VGND.n948 1179.3
R250 VGND.n954 VGND.n953 1179.3
R251 VGND.n959 VGND.n958 1179.3
R252 VGND.n1944 VGND.n1943 1179.3
R253 VGND.n1942 VGND.n1941 1179.3
R254 VGND.n1937 VGND.n1936 1179.3
R255 VGND.n1932 VGND.n1931 1179.3
R256 VGND.n1903 VGND.n1902 1179.3
R257 VGND.n1901 VGND.n1900 1179.3
R258 VGND.n1877 VGND.n1876 1179.3
R259 VGND.n1875 VGND.n1874 1179.3
R260 VGND.n1851 VGND.n1850 1179.3
R261 VGND.n1849 VGND.n1848 1179.3
R262 VGND.n1825 VGND.n1824 1179.3
R263 VGND.n1823 VGND.n1822 1179.3
R264 VGND.n1402 VGND.n1401 1179.3
R265 VGND.n1400 VGND.n1399 1179.3
R266 VGND.n1395 VGND.n1394 1179.3
R267 VGND.n2359 VGND.n2358 1179.3
R268 VGND.n2357 VGND.n2356 1179.3
R269 VGND.n1919 VGND.n1918 1179.3
R270 VGND.n1921 VGND.n1920 1179.3
R271 VGND.n1914 VGND.n1913 1179.3
R272 VGND.n1890 VGND.n1889 1179.3
R273 VGND.n1888 VGND.n1887 1179.3
R274 VGND.n1864 VGND.n1863 1179.3
R275 VGND.n1862 VGND.n1861 1179.3
R276 VGND.n1838 VGND.n1837 1179.3
R277 VGND.n1836 VGND.n1835 1179.3
R278 VGND.n1812 VGND.n1811 1179.3
R279 VGND.n1810 VGND.n1809 1179.3
R280 VGND.n1382 VGND.n1381 1179.3
R281 VGND.n1380 VGND.n1379 1179.3
R282 VGND.n1782 VGND.n1781 1179.3
R283 VGND.n1787 VGND.n1786 1179.3
R284 VGND.n1789 VGND.n1788 1179.3
R285 VGND.n1317 VGND.n1316 1179.3
R286 VGND.n1322 VGND.n1321 1179.3
R287 VGND.n1327 VGND.n1326 1179.3
R288 VGND.n1332 VGND.n1331 1179.3
R289 VGND.n1337 VGND.n1336 1179.3
R290 VGND.n1342 VGND.n1341 1179.3
R291 VGND.n1347 VGND.n1346 1179.3
R292 VGND.n1352 VGND.n1351 1179.3
R293 VGND.n1357 VGND.n1356 1179.3
R294 VGND.n1362 VGND.n1361 1179.3
R295 VGND.n1364 VGND.n1363 1179.3
R296 VGND.n1312 VGND.n1311 1179.3
R297 VGND.n1770 VGND.n1769 1179.3
R298 VGND.n1768 VGND.n1767 1179.3
R299 VGND.n1763 VGND.n1762 1179.3
R300 VGND.n1758 VGND.n1757 1179.3
R301 VGND.n1729 VGND.n1728 1179.3
R302 VGND.n1727 VGND.n1726 1179.3
R303 VGND.n1703 VGND.n1702 1179.3
R304 VGND.n1701 VGND.n1700 1179.3
R305 VGND.n1677 VGND.n1676 1179.3
R306 VGND.n1675 VGND.n1674 1179.3
R307 VGND.n1651 VGND.n1650 1179.3
R308 VGND.n1649 VGND.n1648 1179.3
R309 VGND.n1524 VGND.n1523 1179.3
R310 VGND.n1522 VGND.n1521 1179.3
R311 VGND.n1517 VGND.n1516 1179.3
R312 VGND.n2384 VGND.n2383 1179.3
R313 VGND.n2382 VGND.n2381 1179.3
R314 VGND.n1745 VGND.n1744 1179.3
R315 VGND.n1747 VGND.n1746 1179.3
R316 VGND.n1740 VGND.n1739 1179.3
R317 VGND.n1716 VGND.n1715 1179.3
R318 VGND.n1714 VGND.n1713 1179.3
R319 VGND.n1690 VGND.n1689 1179.3
R320 VGND.n1688 VGND.n1687 1179.3
R321 VGND.n1664 VGND.n1663 1179.3
R322 VGND.n1662 VGND.n1661 1179.3
R323 VGND.n1638 VGND.n1637 1179.3
R324 VGND.n1636 VGND.n1635 1179.3
R325 VGND.n1539 VGND.n1538 1179.3
R326 VGND.n1537 VGND.n1536 1179.3
R327 VGND.n1608 VGND.n1607 1179.3
R328 VGND.n1613 VGND.n1612 1179.3
R329 VGND.n1615 VGND.n1614 1179.3
R330 VGND.n1600 VGND.n1599 1179.3
R331 VGND.n1595 VGND.n1594 1179.3
R332 VGND.n1590 VGND.n1589 1179.3
R333 VGND.n1585 VGND.n1584 1179.3
R334 VGND.n1580 VGND.n1579 1179.3
R335 VGND.n1575 VGND.n1574 1179.3
R336 VGND.n1570 VGND.n1569 1179.3
R337 VGND.n1565 VGND.n1564 1179.3
R338 VGND.n1560 VGND.n1559 1179.3
R339 VGND.n1555 VGND.n1554 1179.3
R340 VGND.n1550 VGND.n1549 1179.3
R341 VGND.n1296 VGND.n1295 1179.3
R342 VGND.n2404 VGND.n2403 1179.3
R343 VGND.n2402 VGND.n2401 1179.3
R344 VGND.n845 VGND.n844 1179.3
R345 VGND.n850 VGND.n849 1179.3
R346 VGND.n855 VGND.n854 1179.3
R347 VGND.n860 VGND.n859 1179.3
R348 VGND.n865 VGND.n864 1179.3
R349 VGND.n870 VGND.n869 1179.3
R350 VGND.n875 VGND.n874 1179.3
R351 VGND.n880 VGND.n879 1179.3
R352 VGND.n885 VGND.n884 1179.3
R353 VGND.n890 VGND.n889 1179.3
R354 VGND.n892 VGND.n891 1179.3
R355 VGND.n840 VGND.n839 1179.3
R356 VGND.n835 VGND.n834 1179.3
R357 VGND.n1229 VGND.n1228 1179.3
R358 VGND.n1227 VGND.n1226 1179.3
R359 VGND.n1210 VGND.n1209 1179.3
R360 VGND.n1208 VGND.n1207 1179.3
R361 VGND.n1197 VGND.n1196 1179.3
R362 VGND.n1195 VGND.n1194 1179.3
R363 VGND.n1178 VGND.n1177 1179.3
R364 VGND.n1176 VGND.n1175 1179.3
R365 VGND.n1165 VGND.n1164 1179.3
R366 VGND.n1163 VGND.n1162 1179.3
R367 VGND.n1146 VGND.n1145 1179.3
R368 VGND.n1144 VGND.n1143 1179.3
R369 VGND.n1133 VGND.n1132 1179.3
R370 VGND.n1131 VGND.n1130 1179.3
R371 VGND.n1123 VGND.n1122 1179.3
R372 VGND.n782 VGND.n781 1179.3
R373 VGND.n780 VGND.n779 1179.3
R374 VGND.n775 VGND.n774 1179.3
R375 VGND.n770 VGND.n769 1179.3
R376 VGND.n765 VGND.n764 1179.3
R377 VGND.n760 VGND.n759 1179.3
R378 VGND.n755 VGND.n754 1179.3
R379 VGND.n750 VGND.n749 1179.3
R380 VGND.n745 VGND.n744 1179.3
R381 VGND.n740 VGND.n739 1179.3
R382 VGND.n735 VGND.n734 1179.3
R383 VGND.n730 VGND.n729 1179.3
R384 VGND.n725 VGND.n724 1179.3
R385 VGND.n720 VGND.n679 1179.3
R386 VGND.n1289 VGND.n1288 1179.3
R387 VGND.n1511 VGND.n1510 1169.57
R388 VGND.n2998 VGND.t33 1146.36
R389 VGND.n3000 VGND.t32 1112.64
R390 VGND.n2999 VGND.t2031 1112.64
R391 VGND.n2981 VGND 1081.89
R392 VGND.n1506 VGND.n1505 1052.29
R393 VGND.t405 VGND.n961 1032.59
R394 VGND.n2689 VGND.t1527 1017.59
R395 VGND.n2688 VGND.t783 1017.59
R396 VGND.n2687 VGND.t764 1017.59
R397 VGND.n2681 VGND.t1531 1017.59
R398 VGND.n2680 VGND.t1529 1017.59
R399 VGND.n2674 VGND.t910 1017.59
R400 VGND.n2673 VGND.t846 1017.59
R401 VGND.n2667 VGND.t1586 1017.59
R402 VGND.n2666 VGND.t830 1017.59
R403 VGND.n2660 VGND.t903 1017.59
R404 VGND.n2659 VGND.t1573 1017.59
R405 VGND.n2653 VGND.t1558 1017.59
R406 VGND.n2652 VGND.t815 1017.59
R407 VGND.n2646 VGND.t878 1017.59
R408 VGND.n2645 VGND.t1565 1017.59
R409 VGND.n233 VGND.t1031 1017.59
R410 VGND.t1958 VGND.n2704 1017.59
R411 VGND.t1070 VGND.n2709 1017.59
R412 VGND.t929 VGND.n2714 1017.59
R413 VGND.t1059 VGND.n2719 1017.59
R414 VGND.t2064 VGND.n2724 1017.59
R415 VGND.t2029 VGND.n2729 1017.59
R416 VGND.t675 VGND.n2734 1017.59
R417 VGND.t2644 VGND.n2739 1017.59
R418 VGND.t338 VGND.n2744 1017.59
R419 VGND.t108 VGND.n2749 1017.59
R420 VGND.t485 VGND.n2754 1017.59
R421 VGND.t1810 VGND.n2759 1017.59
R422 VGND.t1475 VGND.n2764 1017.59
R423 VGND.n2765 VGND.t547 1017.59
R424 VGND.n2514 VGND.t1483 1017.59
R425 VGND.n2513 VGND.t1938 1017.59
R426 VGND.n2508 VGND.t30 1017.59
R427 VGND.t925 VGND.n2433 1017.59
R428 VGND.t2073 VGND.n2438 1017.59
R429 VGND.t2130 VGND.n2443 1017.59
R430 VGND.t517 VGND.n2448 1017.59
R431 VGND.t2659 VGND.n2453 1017.59
R432 VGND.t274 VGND.n2458 1017.59
R433 VGND.t361 VGND.n2463 1017.59
R434 VGND.t81 VGND.n2468 1017.59
R435 VGND.t740 VGND.n2473 1017.59
R436 VGND.t1759 VGND.n2478 1017.59
R437 VGND.t1170 VGND.n2483 1017.59
R438 VGND.t659 VGND.n2488 1017.59
R439 VGND.n2816 VGND.t2653 1017.59
R440 VGND.t205 VGND.n371 1017.59
R441 VGND.n372 VGND.t68 1017.59
R442 VGND.t1632 VGND.n2171 1017.59
R443 VGND.n2172 VGND.t2359 1017.59
R444 VGND.t311 VGND.n2197 1017.59
R445 VGND.n2198 VGND.t1183 1017.59
R446 VGND.t681 VGND.n2223 1017.59
R447 VGND.n2224 VGND.t1298 1017.59
R448 VGND.t397 VGND.n2249 1017.59
R449 VGND.n2250 VGND.t90 1017.59
R450 VGND.t2223 VGND.n2280 1017.59
R451 VGND.t2210 VGND.n2285 1017.59
R452 VGND.t1156 VGND.n2290 1017.59
R453 VGND.n2291 VGND.t1890 1017.59
R454 VGND.t1105 VGND.n1428 1017.59
R455 VGND.n1429 VGND.t2089 1017.59
R456 VGND.t23 VGND.n2158 1017.59
R457 VGND.n2159 VGND.t2686 1017.59
R458 VGND.t2197 VGND.n2184 1017.59
R459 VGND.n2185 VGND.t2602 1017.59
R460 VGND.t1198 VGND.n2210 1017.59
R461 VGND.n2211 VGND.t666 1017.59
R462 VGND.t283 VGND.n2236 1017.59
R463 VGND.n2237 VGND.t218 1017.59
R464 VGND.t121 VGND.n2262 1017.59
R465 VGND.n2268 VGND.t300 1017.59
R466 VGND.n2267 VGND.t193 1017.59
R467 VGND.t1236 VGND.n2307 1017.59
R468 VGND.n2308 VGND.t538 1017.59
R469 VGND.t1479 VGND.n1442 1017.59
R470 VGND.n1493 VGND.t2123 1017.59
R471 VGND.n1492 VGND.t1622 1017.59
R472 VGND.n1487 VGND.t919 1017.59
R473 VGND.n1482 VGND.t2203 1017.59
R474 VGND.n1477 VGND.t2126 1017.59
R475 VGND.n1472 VGND.t1899 1017.59
R476 VGND.n1467 VGND.t1915 1017.59
R477 VGND.n1462 VGND.t1306 1017.59
R478 VGND.n1457 VGND.t412 1017.59
R479 VGND.n1452 VGND.t77 1017.59
R480 VGND.n1447 VGND.t289 1017.59
R481 VGND.n2136 VGND.t1753 1017.59
R482 VGND.n2135 VGND.t2043 1017.59
R483 VGND.n2130 VGND.t653 1017.59
R484 VGND.n1504 VGND.t1029 1017.59
R485 VGND.t1956 VGND.n626 1017.59
R486 VGND.n627 VGND.t1068 1017.59
R487 VGND.t927 VGND.n1997 1017.59
R488 VGND.n1998 VGND.t1057 1017.59
R489 VGND.t2062 VGND.n2023 1017.59
R490 VGND.n2024 VGND.t2027 1017.59
R491 VGND.t673 VGND.n2049 1017.59
R492 VGND.n2050 VGND.t2642 1017.59
R493 VGND.t336 VGND.n2075 1017.59
R494 VGND.n2076 VGND.t106 1017.59
R495 VGND.t483 VGND.n2106 1017.59
R496 VGND.t1808 VGND.n2111 1017.59
R497 VGND.t1473 VGND.n2116 1017.59
R498 VGND.n2117 VGND.t545 1017.59
R499 VGND.t2655 VGND.n652 1017.59
R500 VGND.n653 VGND.t207 1017.59
R501 VGND.t70 VGND.n1984 1017.59
R502 VGND.n1985 VGND.t1634 1017.59
R503 VGND.t2361 VGND.n2010 1017.59
R504 VGND.n2011 VGND.t313 1017.59
R505 VGND.t721 VGND.n2036 1017.59
R506 VGND.n2037 VGND.t683 1017.59
R507 VGND.t1300 VGND.n2062 1017.59
R508 VGND.n2063 VGND.t399 1017.59
R509 VGND.t92 VGND.n2088 1017.59
R510 VGND.n2094 VGND.t2225 1017.59
R511 VGND.n2093 VGND.t2212 1017.59
R512 VGND.t1158 VGND.n2332 1017.59
R513 VGND.n2333 VGND.t1892 1017.59
R514 VGND.n959 VGND.t1095 1017.59
R515 VGND.n954 VGND.t2346 1017.59
R516 VGND.n949 VGND.t452 1017.59
R517 VGND.n944 VGND.t727 1017.59
R518 VGND.n939 VGND.t1506 1017.59
R519 VGND.n934 VGND.t2068 1017.59
R520 VGND.n929 VGND.t306 1017.59
R521 VGND.n924 VGND.t1972 1017.59
R522 VGND.n919 VGND.t2674 1017.59
R523 VGND.n914 VGND.t342 1017.59
R524 VGND.n909 VGND.t102 1017.59
R525 VGND.n904 VGND.t733 1017.59
R526 VGND.n1962 VGND.t1849 1017.59
R527 VGND.n1961 VGND.t2255 1017.59
R528 VGND.n1956 VGND.t526 1017.59
R529 VGND.t1103 VGND.n1395 1017.59
R530 VGND.t2523 VGND.n1400 1017.59
R531 VGND.n1401 VGND.t21 1017.59
R532 VGND.t2684 VGND.n1823 1017.59
R533 VGND.n1824 VGND.t2195 1017.59
R534 VGND.t2600 VGND.n1849 1017.59
R535 VGND.n1850 VGND.t1195 1017.59
R536 VGND.t664 VGND.n1875 1017.59
R537 VGND.n1876 VGND.t281 1017.59
R538 VGND.t216 VGND.n1901 1017.59
R539 VGND.n1902 VGND.t119 1017.59
R540 VGND.t298 VGND.n1932 1017.59
R541 VGND.t1209 VGND.n1937 1017.59
R542 VGND.t1045 VGND.n1942 1017.59
R543 VGND.n1943 VGND.t535 1017.59
R544 VGND.t381 VGND.n1380 1017.59
R545 VGND.n1381 VGND.t2353 1017.59
R546 VGND.t1617 VGND.n1810 1017.59
R547 VGND.n1811 VGND.t146 1017.59
R548 VGND.t2201 VGND.n1836 1017.59
R549 VGND.n1837 VGND.t317 1017.59
R550 VGND.t724 VGND.n1862 1017.59
R551 VGND.n1863 VGND.t1913 1017.59
R552 VGND.t1304 VGND.n1888 1017.59
R553 VGND.n1889 VGND.t409 1017.59
R554 VGND.t84 VGND.n1914 1017.59
R555 VGND.n1920 VGND.t1204 1017.59
R556 VGND.n1919 VGND.t1953 1017.59
R557 VGND.t2041 VGND.n2357 1017.59
R558 VGND.n2358 VGND.t1895 1017.59
R559 VGND.t1481 VGND.n1312 1017.59
R560 VGND.n1363 VGND.t1936 1017.59
R561 VGND.n1362 VGND.t28 1017.59
R562 VGND.n1357 VGND.t923 1017.59
R563 VGND.n1352 VGND.t2071 1017.59
R564 VGND.n1347 VGND.t2128 1017.59
R565 VGND.n1342 VGND.t185 1017.59
R566 VGND.n1337 VGND.t1919 1017.59
R567 VGND.n1332 VGND.t272 1017.59
R568 VGND.n1327 VGND.t359 1017.59
R569 VGND.n1322 VGND.t79 1017.59
R570 VGND.n1317 VGND.t738 1017.59
R571 VGND.n1788 VGND.t1757 1017.59
R572 VGND.n1787 VGND.t1168 1017.59
R573 VGND.n1782 VGND.t656 1017.59
R574 VGND.t2651 VGND.n1517 1017.59
R575 VGND.t203 VGND.n1522 1017.59
R576 VGND.n1523 VGND.t66 1017.59
R577 VGND.t1630 VGND.n1649 1017.59
R578 VGND.n1650 VGND.t2357 1017.59
R579 VGND.t48 VGND.n1675 1017.59
R580 VGND.n1676 VGND.t1181 1017.59
R581 VGND.t679 VGND.n1701 1017.59
R582 VGND.n1702 VGND.t1295 1017.59
R583 VGND.t395 VGND.n1727 1017.59
R584 VGND.n1728 VGND.t87 1017.59
R585 VGND.t2221 VGND.n1758 1017.59
R586 VGND.t2208 VGND.n1763 1017.59
R587 VGND.t1154 VGND.n1768 1017.59
R588 VGND.n1769 VGND.t1888 1017.59
R589 VGND.t588 VGND.n1537 1017.59
R590 VGND.n1538 VGND.t2093 1017.59
R591 VGND.t25 VGND.n1636 1017.59
R592 VGND.n1637 VGND.t1140 1017.59
R593 VGND.t1054 VGND.n1662 1017.59
R594 VGND.n1663 VGND.t2058 1017.59
R595 VGND.t2023 VGND.n1688 1017.59
R596 VGND.n1689 VGND.t670 1017.59
R597 VGND.t433 VGND.n1714 1017.59
R598 VGND.n1715 VGND.t220 1017.59
R599 VGND.t114 VGND.n1740 1017.59
R600 VGND.n1746 VGND.t2052 1017.59
R601 VGND.n1745 VGND.t197 1017.59
R602 VGND.t1239 VGND.n2382 1017.59
R603 VGND.n2383 VGND.t541 1017.59
R604 VGND.n1295 VGND.t2649 1017.59
R605 VGND.t201 VGND.n1550 1017.59
R606 VGND.t64 VGND.n1555 1017.59
R607 VGND.t2036 VGND.n1560 1017.59
R608 VGND.t2355 VGND.n1565 1017.59
R609 VGND.t46 VGND.n1570 1017.59
R610 VGND.t1178 VGND.n1575 1017.59
R611 VGND.t677 VGND.n1580 1017.59
R612 VGND.t1293 VGND.n1585 1017.59
R613 VGND.t393 VGND.n1590 1017.59
R614 VGND.t100 VGND.n1595 1017.59
R615 VGND.t2219 VGND.n1600 1017.59
R616 VGND.n1614 VGND.t2206 1017.59
R617 VGND.n1613 VGND.t1152 1017.59
R618 VGND.n1608 VGND.t1885 1017.59
R619 VGND.t1035 VGND.n835 1017.59
R620 VGND.t1962 VGND.n840 1017.59
R621 VGND.n891 VGND.t1072 1017.59
R622 VGND.n890 VGND.t932 1017.59
R623 VGND.n885 VGND.t1504 1017.59
R624 VGND.n880 VGND.t2066 1017.59
R625 VGND.n875 VGND.t303 1017.59
R626 VGND.n870 VGND.t1969 1017.59
R627 VGND.n865 VGND.t2672 1017.59
R628 VGND.n860 VGND.t340 1017.59
R629 VGND.n855 VGND.t110 1017.59
R630 VGND.n850 VGND.t487 1017.59
R631 VGND.n845 VGND.t2216 1017.59
R632 VGND.t2253 VGND.n2402 1017.59
R633 VGND.n2403 VGND.t523 1017.59
R634 VGND.n1289 VGND.t891 1017.59
R635 VGND.t1578 VGND.n720 1017.59
R636 VGND.t1560 VGND.n725 1017.59
R637 VGND.t895 VGND.n730 1017.59
R638 VGND.t893 VGND.n735 1017.59
R639 VGND.t1550 VGND.n740 1017.59
R640 VGND.t806 VGND.n745 1017.59
R641 VGND.t792 VGND.n750 1017.59
R642 VGND.t869 VGND.n755 1017.59
R643 VGND.t1537 VGND.n760 1017.59
R644 VGND.t788 VGND.n765 1017.59
R645 VGND.t770 VGND.n770 1017.59
R646 VGND.t851 VGND.n775 1017.59
R647 VGND.t1520 VGND.n780 1017.59
R648 VGND.n781 VGND.t773 1017.59
R649 VGND.n1508 VGND.n579 934.784
R650 VGND.n2892 VGND 927.203
R651 VGND.n2895 VGND 927.203
R652 VGND.n962 VGND 918.774
R653 VGND.n113 VGND 910.346
R654 VGND.n2859 VGND 910.346
R655 VGND.n2993 VGND.t139 909.365
R656 VGND.n2818 VGND.n177 900
R657 VGND.n1507 VGND 851.341
R658 VGND.n2689 VGND.t1187 838.438
R659 VGND.t1114 VGND.n2688 838.438
R660 VGND.t1098 VGND.n2687 838.438
R661 VGND.n2681 VGND.t2637 838.438
R662 VGND.t1308 VGND.n2680 838.438
R663 VGND.n2674 VGND.t1964 838.438
R664 VGND.t2411 VGND.n2673 838.438
R665 VGND.n2667 VGND.t2345 838.438
R666 VGND.t590 VGND.n2666 838.438
R667 VGND.n2660 VGND.t1714 838.438
R668 VGND.t1516 VGND.n2659 838.438
R669 VGND.n2653 VGND.t2243 838.438
R670 VGND.t1659 VGND.n2652 838.438
R671 VGND.n2646 VGND.t296 838.438
R672 VGND.t1063 VGND.n2645 838.438
R673 VGND.t917 VGND.n33 838.438
R674 VGND.n233 VGND.t38 838.438
R675 VGND.n2704 VGND.t602 838.438
R676 VGND.n2709 VGND.t2340 838.438
R677 VGND.n2714 VGND.t1509 838.438
R678 VGND.n2719 VGND.t95 838.438
R679 VGND.n2724 VGND.t1242 838.438
R680 VGND.n2729 VGND.t1116 838.438
R681 VGND.n2734 VGND.t244 838.438
R682 VGND.n2739 VGND.t443 838.438
R683 VGND.n2744 VGND.t345 838.438
R684 VGND.n2749 VGND.t2229 838.438
R685 VGND.n2754 VGND.t1113 838.438
R686 VGND.n2759 VGND.t1185 838.438
R687 VGND.n2764 VGND.t286 838.438
R688 VGND.n2765 VGND.t1653 838.438
R689 VGND.n2984 VGND.t1718 838.438
R690 VGND.n2514 VGND.t295 838.438
R691 VGND.t2236 VGND.n2513 838.438
R692 VGND.t1062 VGND.n2508 838.438
R693 VGND.n2433 VGND.t1324 838.438
R694 VGND.n2438 VGND.t1717 838.438
R695 VGND.n2443 VGND.t73 838.438
R696 VGND.n2448 VGND.t2342 838.438
R697 VGND.n2453 VGND.t1099 838.438
R698 VGND.n2458 VGND.t2635 838.438
R699 VGND.n2463 VGND.t1112 838.438
R700 VGND.n2468 VGND.t188 838.438
R701 VGND.n2473 VGND.t2408 838.438
R702 VGND.n2478 VGND.t2248 838.438
R703 VGND.n2483 VGND.t173 838.438
R704 VGND.n2488 VGND.t123 838.438
R705 VGND.n2489 VGND.t18 838.438
R706 VGND.t297 VGND.n2816 838.438
R707 VGND.n371 VGND.t551 838.438
R708 VGND.n372 VGND.t35 838.438
R709 VGND.n2171 VGND.t1037 838.438
R710 VGND.n2172 VGND.t534 838.438
R711 VGND.n2197 VGND.t1652 838.438
R712 VGND.n2198 VGND.t1061 838.438
R713 VGND.n2223 VGND.t2009 838.438
R714 VGND.n2224 VGND.t1820 838.438
R715 VGND.n2249 VGND.t245 838.438
R716 VGND.n2250 VGND.t1715 838.438
R717 VGND.n2280 VGND.t232 838.438
R718 VGND.n2285 VGND.t2664 838.438
R719 VGND.n2290 VGND.t1469 838.438
R720 VGND.n2291 VGND.t2528 838.438
R721 VGND.n2428 VGND.t1640 838.438
R722 VGND.n1428 VGND.t246 838.438
R723 VGND.n1429 VGND.t2011 838.438
R724 VGND.n2158 VGND.t1067 838.438
R725 VGND.n2159 VGND.t1967 838.438
R726 VGND.n2184 VGND.t1186 838.438
R727 VGND.n2185 VGND.t1274 838.438
R728 VGND.n2210 VGND.t228 838.438
R729 VGND.n2211 VGND.t86 838.438
R730 VGND.n2236 VGND.t36 838.438
R731 VGND.n2237 VGND.t1490 838.438
R732 VGND.n2262 VGND.t1513 838.438
R733 VGND.n2268 VGND.t522 838.438
R734 VGND.t1814 VGND.n2267 838.438
R735 VGND.n2307 VGND.t1620 838.438
R736 VGND.n2308 VGND.t1325 838.438
R737 VGND.t1041 VGND.n261 838.438
R738 VGND.n1442 VGND.t247 838.438
R739 VGND.n1493 VGND.t2231 838.438
R740 VGND.t533 VGND.n1492 838.438
R741 VGND.t1053 VGND.n1487 838.438
R742 VGND.t2339 VGND.n1482 838.438
R743 VGND.t2658 VGND.n1477 838.438
R744 VGND.t2682 VGND.n1472 838.438
R745 VGND.t702 VGND.n1467 838.438
R746 VGND.t1817 VGND.n1462 838.438
R747 VGND.t2228 VGND.n1457 838.438
R748 VGND.t142 VGND.n1452 838.438
R749 VGND.t607 VGND.n1447 838.438
R750 VGND.n2136 VGND.t1791 838.438
R751 VGND.t1211 VGND.n2135 838.438
R752 VGND.t1470 VGND.n2130 838.438
R753 VGND.t2412 VGND.n262 838.438
R754 VGND.t1326 VGND.n1504 838.438
R755 VGND.n626 VGND.t1804 838.438
R756 VGND.n627 VGND.t2234 838.438
R757 VGND.n1997 VGND.t96 838.438
R758 VGND.n1998 VGND.t1642 838.438
R759 VGND.n2023 VGND.t143 838.438
R760 VGND.n2024 VGND.t916 838.438
R761 VGND.n2049 VGND.t2056 838.438
R762 VGND.n2050 VGND.t2646 838.438
R763 VGND.n2075 VGND.t1066 838.438
R764 VGND.n2076 VGND.t1902 838.438
R765 VGND.n2106 VGND.t1637 838.438
R766 VGND.n2111 VGND.t1934 838.438
R767 VGND.n2116 VGND.t1115 838.438
R768 VGND.n2117 VGND.t229 838.438
R769 VGND.t1912 VGND.n263 838.438
R770 VGND.n652 VGND.t550 838.438
R771 VGND.n653 VGND.t1047 838.438
R772 VGND.n1984 VGND.t74 838.438
R773 VGND.n1985 VGND.t1909 838.438
R774 VGND.n2010 VGND.t1486 838.438
R775 VGND.n2011 VGND.t2022 838.438
R776 VGND.n2036 VGND.t211 838.438
R777 VGND.n2037 VGND.t384 838.438
R778 VGND.n2062 VGND.t1309 838.438
R779 VGND.n2063 VGND.t712 838.438
R780 VGND.n2088 VGND.t2406 838.438
R781 VGND.n2094 VGND.t1150 838.438
R782 VGND.t2343 VGND.n2093 838.438
R783 VGND.n2332 VGND.t914 838.438
R784 VGND.n2333 VGND.t2410 838.438
R785 VGND.t1174 VGND.n264 838.438
R786 VGND.t1111 VGND.n959 838.438
R787 VGND.t2344 VGND.n954 838.438
R788 VGND.t129 VGND.n949 838.438
R789 VGND.t1813 VGND.n944 838.438
R790 VGND.t1802 VGND.n939 838.438
R791 VGND.t608 VGND.n934 838.438
R792 VGND.t1812 VGND.n929 838.438
R793 VGND.t1512 VGND.n924 838.438
R794 VGND.t75 VGND.n919 838.438
R795 VGND.t1212 VGND.n914 838.438
R796 VGND.t383 VGND.n909 838.438
R797 VGND.t2233 VGND.n904 838.438
R798 VGND.n1962 VGND.t2525 838.438
R799 VGND.t1194 VGND.n1961 838.438
R800 VGND.t1311 VGND.n1956 838.438
R801 VGND.t1050 VGND.n265 838.438
R802 VGND.n1395 VGND.t1882 838.438
R803 VGND.n1400 VGND.t2663 838.438
R804 VGND.n1401 VGND.t701 838.438
R805 VGND.n1823 VGND.t1138 838.438
R806 VGND.n1824 VGND.t1489 838.438
R807 VGND.n1849 VGND.t2006 838.438
R808 VGND.n1850 VGND.t1510 838.438
R809 VGND.n1875 VGND.t1901 838.438
R810 VGND.n1876 VGND.t2230 838.438
R811 VGND.n1901 VGND.t2246 838.438
R812 VGND.n1902 VGND.t2008 838.438
R813 VGND.n1932 VGND.t1815 838.438
R814 VGND.n1937 VGND.t287 838.438
R815 VGND.n1942 VGND.t76 838.438
R816 VGND.n1943 VGND.t1173 838.438
R817 VGND.t2007 VGND.n266 838.438
R818 VGND.n1380 VGND.t1897 838.438
R819 VGND.n1381 VGND.t2558 838.438
R820 VGND.n1810 VGND.t1903 838.438
R821 VGND.n1811 VGND.t1245 838.438
R822 VGND.n1836 VGND.t1065 838.438
R823 VGND.n1837 VGND.t288 838.438
R824 VGND.n1862 VGND.t918 838.438
R825 VGND.n1863 VGND.t128 838.438
R826 VGND.n1888 VGND.t240 838.438
R827 VGND.n1889 VGND.t1109 838.438
R828 VGND.n1914 VGND.t707 838.438
R829 VGND.n1920 VGND.t149 838.438
R830 VGND.t212 VGND.n1919 838.438
R831 VGND.n2357 VGND.t1790 838.438
R832 VGND.n2358 VGND.t1177 838.438
R833 VGND.t174 VGND.n267 838.438
R834 VGND.n1312 VGND.t1816 838.438
R835 VGND.n1363 VGND.t1119 838.438
R836 VGND.t2681 VGND.n1362 838.438
R837 VGND.t698 VGND.n1357 838.438
R838 VGND.t1911 VGND.n1352 838.438
R839 VGND.t1048 VGND.n1347 838.438
R840 VGND.t2636 VGND.n1342 838.438
R841 VGND.t2005 VGND.n1337 838.438
R842 VGND.t1805 VGND.n1332 838.438
R843 VGND.t1881 VGND.n1327 838.438
R844 VGND.t1654 VGND.n1322 838.438
R845 VGND.t1898 VGND.n1317 838.438
R846 VGND.n1788 VGND.t1965 838.438
R847 VGND.t1883 VGND.n1787 838.438
R848 VGND.t699 VGND.n1782 838.438
R849 VGND.t1488 VGND.n268 838.438
R850 VGND.n1517 VGND.t1511 838.438
R851 VGND.n1522 VGND.t285 838.438
R852 VGND.n1523 VGND.t105 838.438
R853 VGND.n1649 VGND.t594 838.438
R854 VGND.n1650 VGND.t1120 838.438
R855 VGND.n1675 VGND.t915 838.438
R856 VGND.n1676 VGND.t2247 838.438
R857 VGND.n1701 VGND.t732 838.438
R858 VGND.n1702 VGND.t164 838.438
R859 VGND.n1727 VGND.t1641 838.438
R860 VGND.n1728 VGND.t2232 838.438
R861 VGND.n1758 VGND.t183 838.438
R862 VGND.n1763 VGND.t189 838.438
R863 VGND.n1768 VGND.t2639 838.438
R864 VGND.n1769 VGND.t1192 838.438
R865 VGND.t970 VGND.n269 838.438
R866 VGND.n1537 VGND.t1884 838.438
R867 VGND.n1538 VGND.t1904 838.438
R868 VGND.n1636 VGND.t2338 838.438
R869 VGND.n1637 VGND.t1108 838.438
R870 VGND.n1662 VGND.t605 838.438
R871 VGND.n1663 VGND.t233 838.438
R872 VGND.n1688 VGND.t1049 838.438
R873 VGND.n1689 VGND.t2057 838.438
R874 VGND.n1714 VGND.t1806 838.438
R875 VGND.n1715 VGND.t62 838.438
R876 VGND.n1740 VGND.t1655 838.438
R877 VGND.n1746 VGND.t63 838.438
R878 VGND.t2021 VGND.n1745 838.438
R879 VGND.n2382 VGND.t603 838.438
R880 VGND.n2383 VGND.t1619 838.438
R881 VGND.t2587 VGND.n270 838.438
R882 VGND.n1295 VGND.t2010 838.438
R883 VGND.n1550 VGND.t148 838.438
R884 VGND.n1555 VGND.t2529 838.438
R885 VGND.n1560 VGND.t2409 838.438
R886 VGND.n1565 VGND.t477 838.438
R887 VGND.n1570 VGND.t230 838.438
R888 VGND.n1575 VGND.t1793 838.438
R889 VGND.n1580 VGND.t200 838.438
R890 VGND.n1585 VGND.t591 838.438
R891 VGND.n1590 VGND.t444 838.438
R892 VGND.n1595 VGND.t1908 838.438
R893 VGND.n1600 VGND.t2341 838.438
R894 VGND.n1614 VGND.t1792 838.438
R895 VGND.t302 VGND.n1613 838.438
R896 VGND.t2638 VGND.n1608 838.438
R897 VGND.t1501 VGND.n271 838.438
R898 VGND.n835 VGND.t239 838.438
R899 VGND.n840 VGND.t593 838.438
R900 VGND.n891 VGND.t2004 838.438
R901 VGND.t1243 VGND.n890 838.438
R902 VGND.t39 VGND.n885 838.438
R903 VGND.t1803 VGND.n880 838.438
R904 VGND.t1110 VGND.n875 838.438
R905 VGND.t1117 VGND.n870 838.438
R906 VGND.t1910 VGND.n865 838.438
R907 VGND.t750 VGND.n860 838.438
R908 VGND.t1807 VGND.n855 838.438
R909 VGND.t1213 VGND.n850 838.438
R910 VGND.t1468 VGND.n845 838.438
R911 VGND.n2402 VGND.t1638 838.438
R912 VGND.n2403 VGND.t2683 838.438
R913 VGND.t1038 VGND.n272 838.438
R914 VGND.t1207 VGND.n1289 838.438
R915 VGND.n720 VGND.t1137 838.438
R916 VGND.n725 VGND.t293 838.438
R917 VGND.n730 VGND.t37 838.438
R918 VGND.n735 VGND.t1052 838.438
R919 VGND.n740 VGND.t1064 838.438
R920 VGND.n745 VGND.t41 838.438
R921 VGND.n750 VGND.t700 838.438
R922 VGND.n755 VGND.t0 838.438
R923 VGND.n760 VGND.t1625 838.438
R924 VGND.n765 VGND.t1471 838.438
R925 VGND.n770 VGND.t40 838.438
R926 VGND.n775 VGND.t1193 838.438
R927 VGND.n780 VGND.t1639 838.438
R928 VGND.n781 VGND.t1933 838.438
R929 VGND.n2413 VGND.t1149 838.438
R930 VGND.n2826 VGND.t857 824.105
R931 VGND.n2825 VGND.t1391 824.105
R932 VGND.t1436 VGND.n114 824.105
R933 VGND.n2817 VGND.t1343 824.105
R934 VGND.t1421 VGND.n177 824.105
R935 VGND.t1460 VGND.n635 824.105
R936 VGND.t1340 VGND.n580 824.105
R937 VGND.n960 VGND.t1379 824.105
R938 VGND.t1424 VGND.n579 824.105
R939 VGND.n1511 VGND.t1439 824.105
R940 VGND.t1346 VGND.n1512 824.105
R941 VGND.n1293 VGND.t1412 824.105
R942 VGND.t1349 VGND.n1294 824.105
R943 VGND.n1292 VGND.t1385 824.105
R944 VGND.n1290 VGND.t2589 824.105
R945 VGND.n2982 VGND.n33 738.111
R946 VGND.n2984 VGND.n2983 738.111
R947 VGND.n2489 VGND.n32 738.111
R948 VGND.n2428 VGND.n2427 738.111
R949 VGND.n2426 VGND.n261 738.111
R950 VGND.n2425 VGND.n262 738.111
R951 VGND.n2424 VGND.n263 738.111
R952 VGND.n2423 VGND.n264 738.111
R953 VGND.n2422 VGND.n265 738.111
R954 VGND.n2421 VGND.n266 738.111
R955 VGND.n2420 VGND.n267 738.111
R956 VGND.n2419 VGND.n268 738.111
R957 VGND.n2418 VGND.n269 738.111
R958 VGND.n2417 VGND.n270 738.111
R959 VGND.n2416 VGND.n271 738.111
R960 VGND.n2415 VGND.n272 738.111
R961 VGND.n2414 VGND.n2413 738.111
R962 VGND.t2439 VGND.t2421 708.047
R963 VGND.t2421 VGND.t2419 708.047
R964 VGND.t2419 VGND.t2429 708.047
R965 VGND.t2429 VGND.t752 708.047
R966 VGND.t752 VGND.t1276 708.047
R967 VGND.t1276 VGND.t458 708.047
R968 VGND.t458 VGND.t456 708.047
R969 VGND.t1219 VGND.t32 708.047
R970 VGND.t2466 VGND.t2453 708.047
R971 VGND.t2453 VGND.t2451 708.047
R972 VGND.t2451 VGND.t2413 708.047
R973 VGND.t2413 VGND.t2237 708.047
R974 VGND.t2237 VGND.t714 708.047
R975 VGND.t714 VGND.t719 708.047
R976 VGND.t719 VGND.t429 708.047
R977 VGND.t2490 VGND.t2437 708.047
R978 VGND.t2437 VGND.t2478 708.047
R979 VGND.t2478 VGND.t2446 708.047
R980 VGND.t2446 VGND.t1322 708.047
R981 VGND.t1322 VGND.t1318 708.047
R982 VGND.t1318 VGND.t1312 708.047
R983 VGND.t1312 VGND.t1314 708.047
R984 VGND.t1216 VGND.t33 708.047
R985 VGND.t2474 VGND.t2435 708.047
R986 VGND.t2443 VGND.t2474 708.047
R987 VGND.t2417 VGND.t2443 708.047
R988 VGND.t754 VGND.t2417 708.047
R989 VGND.t1278 VGND.t754 708.047
R990 VGND.t751 VGND.t1278 708.047
R991 VGND.t1275 VGND.t751 708.047
R992 VGND.t2431 VGND.t2470 708.047
R993 VGND.t2470 VGND.t2441 708.047
R994 VGND.t2441 VGND.t2449 708.047
R995 VGND.t2449 VGND.t716 708.047
R996 VGND.t716 VGND.t1139 708.047
R997 VGND.t1139 VGND.t1291 708.047
R998 VGND.t1291 VGND.t718 708.047
R999 VGND.t2483 VGND.t2427 708.047
R1000 VGND.t2427 VGND.t2488 708.047
R1001 VGND.t2488 VGND.t2460 708.047
R1002 VGND.t2460 VGND.t1320 708.047
R1003 VGND.t1320 VGND.t1316 708.047
R1004 VGND.t1316 VGND.t1321 708.047
R1005 VGND.t1321 VGND.t1317 708.047
R1006 VGND.n2979 VGND.n2978 708.047
R1007 VGND.t224 VGND.t2526 691.188
R1008 VGND.t708 VGND.t2032 691.188
R1009 VGND.n2822 VGND.t1604 685.545
R1010 VGND.n3002 VGND.t1604 685.545
R1011 VGND.n2825 VGND.n2824 660.87
R1012 VGND.t252 VGND.t55 657.471
R1013 VGND.t264 VGND.t53 657.471
R1014 VGND.t2510 VGND.t51 657.471
R1015 VGND.t6 VGND.t2367 657.471
R1016 VGND.t2494 VGND.t2472 657.471
R1017 VGND.t2468 VGND.t140 657.471
R1018 VGND.t2505 VGND.t136 657.471
R1019 VGND.t2455 VGND.t130 657.471
R1020 VGND.t2367 VGND.t2369 654.197
R1021 VGND.t2472 VGND.t2498 654.197
R1022 VGND.t861 VGND.t859 644.952
R1023 VGND.t796 VGND.t798 644.952
R1024 VGND.t785 VGND.t787 644.952
R1025 VGND.t768 VGND.t766 644.952
R1026 VGND.t1533 VGND.t1535 644.952
R1027 VGND.t1519 VGND.t1517 644.952
R1028 VGND.t912 VGND.t757 644.952
R1029 VGND.t844 VGND.t848 644.952
R1030 VGND.t1588 VGND.t834 644.952
R1031 VGND.t772 VGND.t832 644.952
R1032 VGND.t905 VGND.t907 644.952
R1033 VGND.t1577 VGND.t1575 644.952
R1034 VGND.t826 VGND.t829 644.952
R1035 VGND.t819 VGND.t817 644.952
R1036 VGND.t880 VGND.t882 644.952
R1037 VGND.t1567 VGND.t1569 644.952
R1038 VGND.t378 VGND.t1083 644.952
R1039 VGND.t1121 VGND.t1961 644.952
R1040 VGND.t454 VGND.t1093 644.952
R1041 VGND.t922 VGND.t1091 644.952
R1042 VGND.t1503 VGND.t2300 644.952
R1043 VGND.t310 VGND.t2298 644.952
R1044 VGND.t2242 VGND.t1089 644.952
R1045 VGND.t1971 VGND.t2308 644.952
R1046 VGND.t1297 VGND.t2306 644.952
R1047 VGND.t1146 VGND.t1680 644.952
R1048 VGND.t89 VGND.t1087 644.952
R1049 VGND.t736 VGND.t2304 644.952
R1050 VGND.t2218 VGND.t1678 644.952
R1051 VGND.t1040 VGND.t1123 644.952
R1052 VGND.t531 VGND.t1085 644.952
R1053 VGND.t2302 VGND.t836 644.952
R1054 VGND.t1034 VGND.t938 644.952
R1055 VGND.t617 VGND.t1941 644.952
R1056 VGND.t615 VGND.t20 644.952
R1057 VGND.t2035 VGND.t613 644.952
R1058 VGND.t2076 VGND.t2617 644.952
R1059 VGND.t2061 VGND.t2615 644.952
R1060 VGND.t2026 VGND.t611 644.952
R1061 VGND.t2662 VGND.t936 644.952
R1062 VGND.t2641 VGND.t934 644.952
R1063 VGND.t364 VGND.t623 644.952
R1064 VGND.t117 VGND.t609 644.952
R1065 VGND.t743 VGND.t2621 644.952
R1066 VGND.t1208 VGND.t621 644.952
R1067 VGND.t1478 VGND.t619 644.952
R1068 VGND.t544 VGND.t940 644.952
R1069 VGND.t2588 VGND.t2619 644.952
R1070 VGND.t1287 VGND.t1101 644.952
R1071 VGND.t2350 VGND.t1125 644.952
R1072 VGND.t1615 VGND.t171 644.952
R1073 VGND.t169 VGND.t1144 644.952
R1074 VGND.t2365 VGND.t1135 644.952
R1075 VGND.t1133 VGND.t2134 644.952
R1076 VGND.t519 VGND.t167 644.952
R1077 VGND.t1285 VGND.t687 644.952
R1078 VGND.t278 VGND.t1283 644.952
R1079 VGND.t1131 VGND.t403 644.952
R1080 VGND.t126 VGND.t165 644.952
R1081 VGND.t1281 VGND.t1202 644.952
R1082 VGND.t1950 VGND.t1129 644.952
R1083 VGND.t1043 VGND.t1127 644.952
R1084 VGND.t661 VGND.t1289 644.952
R1085 VGND.t1279 VGND.t758 644.952
R1086 VGND.t2647 VGND.t445 644.952
R1087 VGND.t2092 VGND.t2606 644.952
R1088 VGND.t1946 VGND.t43 644.952
R1089 VGND.t144 VGND.t1944 644.952
R1090 VGND.t250 VGND.t1746 644.952
R1091 VGND.t242 VGND.t248 644.952
R1092 VGND.t1942 VGND.t2239 644.952
R1093 VGND.t669 VGND.t466 644.952
R1094 VGND.t464 VGND.t2677 644.952
R1095 VGND.t223 VGND.t2612 644.952
R1096 VGND.t449 VGND.t97 644.952
R1097 VGND.t2055 VGND.t462 644.952
R1098 VGND.t2610 VGND.t196 644.952
R1099 VGND.t2608 VGND.t2039 644.952
R1100 VGND.t528 VGND.t447 644.952
R1101 VGND.t2669 VGND.t1543 644.952
R1102 VGND.t1028 VGND.t365 644.952
R1103 VGND.t1935 VGND.t415 644.952
R1104 VGND.t375 VGND.t27 644.952
R1105 VGND.t373 VGND.t730 644.952
R1106 VGND.t425 VGND.t2070 644.952
R1107 VGND.t423 VGND.t2605 644.952
R1108 VGND.t371 VGND.t1200 644.952
R1109 VGND.t391 VGND.t1918 644.952
R1110 VGND.t389 VGND.t432 644.952
R1111 VGND.t421 VGND.t358 644.952
R1112 VGND.t369 VGND.t113 644.952
R1113 VGND.t387 VGND.t292 644.952
R1114 VGND.t419 VGND.t1756 644.952
R1115 VGND.t417 VGND.t1472 644.952
R1116 VGND.t367 VGND.t540 644.952
R1117 VGND.t427 VGND.t804 644.952
R1118 VGND.t1737 VGND.t377 644.952
R1119 VGND.t1960 VGND.t439 644.952
R1120 VGND.t451 VGND.t437 644.952
R1121 VGND.t435 VGND.t921 644.952
R1122 VGND.t1502 VGND.t1725 644.952
R1123 VGND.t1723 VGND.t45 644.952
R1124 VGND.t2241 VGND.t1743 644.952
R1125 VGND.t1735 VGND.t1968 644.952
R1126 VGND.t2679 VGND.t1733 644.952
R1127 VGND.t1721 VGND.t344 644.952
R1128 VGND.t99 VGND.t1741 644.952
R1129 VGND.t1731 VGND.t735 644.952
R1130 VGND.t2215 VGND.t1719 644.952
R1131 VGND.t1039 VGND.t441 644.952
R1132 VGND.t530 VGND.t1739 644.952
R1133 VGND.t1729 VGND.t835 644.952
R1134 VGND.t1102 VGND.t1602 644.952
R1135 VGND.t2351 VGND.t327 644.952
R1136 VGND.t325 VGND.t1616 644.952
R1137 VGND.t1145 VGND.t323 644.952
R1138 VGND.t1592 VGND.t2199 644.952
R1139 VGND.t2598 VGND.t1590 644.952
R1140 VGND.t321 VGND.t520 644.952
R1141 VGND.t688 VGND.t1600 644.952
R1142 VGND.t1598 VGND.t279 644.952
R1143 VGND.t404 VGND.t333 644.952
R1144 VGND.t319 VGND.t127 644.952
R1145 VGND.t1203 VGND.t1596 644.952
R1146 VGND.t331 VGND.t1951 644.952
R1147 VGND.t329 VGND.t1044 644.952
R1148 VGND.t662 VGND.t385 644.952
R1149 VGND.t1594 VGND.t769 644.952
R1150 VGND.t1226 VGND.t380 644.952
R1151 VGND.t705 VGND.t1948 644.952
R1152 VGND.t703 VGND.t2671 644.952
R1153 VGND.t1234 VGND.t1629 644.952
R1154 VGND.t558 VGND.t2407 644.952
R1155 VGND.t556 VGND.t316 644.952
R1156 VGND.t1232 VGND.t723 644.952
R1157 VGND.t1166 VGND.t1975 644.952
R1158 VGND.t1164 VGND.t1303 644.952
R1159 VGND.t554 VGND.t1148 644.952
R1160 VGND.t1230 VGND.t83 644.952
R1161 VGND.t1162 VGND.t2045 644.952
R1162 VGND.t552 VGND.t1852 644.952
R1163 VGND.t214 VGND.t2040 644.952
R1164 VGND.t1228 VGND.t1894 644.952
R1165 VGND.t1160 VGND.t850 644.952
R1166 VGND.t1097 VGND.t2625 644.952
R1167 VGND.t2091 VGND.t2288 644.952
R1168 VGND.t42 VGND.t2286 644.952
R1169 VGND.t2633 VGND.t1636 644.952
R1170 VGND.t1745 VGND.t1727 644.952
R1171 VGND.t2296 VGND.t241 644.952
R1172 VGND.t305 VGND.t2631 644.952
R1173 VGND.t696 VGND.t668 644.952
R1174 VGND.t2676 VGND.t694 644.952
R1175 VGND.t2294 VGND.t222 644.952
R1176 VGND.t104 VGND.t2629 644.952
R1177 VGND.t692 VGND.t2054 644.952
R1178 VGND.t195 VGND.t2292 644.952
R1179 VGND.t2038 VGND.t2290 644.952
R1180 VGND.t525 VGND.t2627 644.952
R1181 VGND.t690 VGND.t1536 644.952
R1182 VGND.t1027 VGND.t755 644.952
R1183 VGND.t2125 VGND.t350 644.952
R1184 VGND.t348 VGND.t1624 644.952
R1185 VGND.t729 VGND.t346 644.952
R1186 VGND.t1929 VGND.t2205 644.952
R1187 VGND.t2604 VGND.t1927 644.952
R1188 VGND.t2521 VGND.t1197 644.952
R1189 VGND.t1917 VGND.t1931 644.952
R1190 VGND.t356 VGND.t431 644.952
R1191 VGND.t414 VGND.t1925 644.952
R1192 VGND.t2519 VGND.t112 644.952
R1193 VGND.t291 VGND.t354 644.952
R1194 VGND.t1923 VGND.t1755 644.952
R1195 VGND.t1921 VGND.t1241 644.952
R1196 VGND.t537 VGND.t2517 644.952
R1197 VGND.t352 VGND.t799 644.952
R1198 VGND.t1033 VGND.t154 644.952
R1199 VGND.t1940 VGND.t1666 644.952
R1200 VGND.t1664 VGND.t19 644.952
R1201 VGND.t1662 VGND.t2034 644.952
R1202 VGND.t1676 VGND.t2075 644.952
R1203 VGND.t1674 VGND.t2060 644.952
R1204 VGND.t1660 VGND.t2025 644.952
R1205 VGND.t152 VGND.t2661 644.952
R1206 VGND.t150 VGND.t2640 644.952
R1207 VGND.t1672 VGND.t363 644.952
R1208 VGND.t158 VGND.t116 644.952
R1209 VGND.t162 VGND.t742 644.952
R1210 VGND.t1670 VGND.t1761 644.952
R1211 VGND.t1668 VGND.t1477 644.952
R1212 VGND.t156 VGND.t543 644.952
R1213 VGND.t160 VGND.t828 644.952
R1214 VGND.t1100 VGND.t746 644.952
R1215 VGND.t2349 VGND.t2017 644.952
R1216 VGND.t1614 VGND.t2015 644.952
R1217 VGND.t2013 VGND.t1143 644.952
R1218 VGND.t2364 VGND.t1650 644.952
R1219 VGND.t1648 VGND.t2133 644.952
R1220 VGND.t187 VGND.t1190 644.952
R1221 VGND.t744 VGND.t686 644.952
R1222 VGND.t277 VGND.t600 644.952
R1223 VGND.t1646 VGND.t402 644.952
R1224 VGND.t125 VGND.t1188 644.952
R1225 VGND.t598 VGND.t1201 644.952
R1226 VGND.t1949 VGND.t1644 644.952
R1227 VGND.t1042 VGND.t2019 644.952
R1228 VGND.t658 VGND.t748 644.952
R1229 VGND.t596 VGND.t909 644.952
R1230 VGND.t2159 VGND.t2648 644.952
R1231 VGND.t1955 VGND.t2328 644.952
R1232 VGND.t2326 VGND.t44 644.952
R1233 VGND.t145 VGND.t2324 644.952
R1234 VGND.t1626 VGND.t1056 644.952
R1235 VGND.t243 VGND.t2336 644.952
R1236 VGND.t2165 VGND.t2240 644.952
R1237 VGND.t672 VGND.t2157 644.952
R1238 VGND.t2155 VGND.t2678 644.952
R1239 VGND.t335 VGND.t2334 644.952
R1240 VGND.t2163 VGND.t98 644.952
R1241 VGND.t482 VGND.t2153 644.952
R1242 VGND.t2332 VGND.t199 644.952
R1243 VGND.t2330 VGND.t1151 644.952
R1244 VGND.t529 VGND.t2161 644.952
R1245 VGND.t2151 VGND.t1564 644.952
R1246 VGND.t1485 VGND.t2147 644.952
R1247 VGND.t1493 VGND.t209 644.952
R1248 VGND.t72 VGND.t1491 644.952
R1249 VGND.t1142 VGND.t475 644.952
R1250 VGND.t2363 VGND.t2137 644.952
R1251 VGND.t2132 VGND.t2135 644.952
R1252 VGND.t184 VGND.t473 644.952
R1253 VGND.t685 VGND.t2145 644.952
R1254 VGND.t276 VGND.t2143 644.952
R1255 VGND.t401 VGND.t1499 644.952
R1256 VGND.t124 VGND.t471 644.952
R1257 VGND.t2227 VGND.t2141 644.952
R1258 VGND.t2214 VGND.t1497 644.952
R1259 VGND.t1495 VGND.t1172 644.952
R1260 VGND.t2149 VGND.t655 644.952
R1261 VGND.t2139 VGND.t908 644.952
R1262 VGND.t379 VGND.t2079 644.952
R1263 VGND.t2348 VGND.t2322 644.952
R1264 VGND.t455 VGND.t2320 644.952
R1265 VGND.t2318 VGND.t1628 644.952
R1266 VGND.t1751 VGND.t1508 644.952
R1267 VGND.t1749 VGND.t315 644.952
R1268 VGND.t2316 VGND.t1180 644.952
R1269 VGND.t2077 VGND.t1974 644.952
R1270 VGND.t2050 VGND.t1302 644.952
R1271 VGND.t1747 VGND.t1147 644.952
R1272 VGND.t2083 VGND.t94 644.952
R1273 VGND.t2048 VGND.t737 644.952
R1274 VGND.t2087 VGND.t1851 644.952
R1275 VGND.t2085 VGND.t2257 644.952
R1276 VGND.t1887 VGND.t2081 644.952
R1277 VGND.t2046 VGND.t845 644.952
R1278 VGND.t2591 VGND.t1107 644.952
R1279 VGND.t2352 VGND.t839 644.952
R1280 VGND.t1621 VGND.t1582 644.952
R1281 VGND.t931 VGND.t1562 644.952
R1282 VGND.t2200 VGND.t897 644.952
R1283 VGND.t2599 VGND.t883 644.952
R1284 VGND.t521 VGND.t1554 644.952
R1285 VGND.t689 VGND.t810 644.952
R1286 VGND.t280 VGND.t794 644.952
R1287 VGND.t411 VGND.t871 644.952
R1288 VGND.t118 VGND.t1541 644.952
R1289 VGND.t1206 VGND.t790 644.952
R1290 VGND.t1952 VGND.t864 644.952
R1291 VGND.t1238 VGND.t855 644.952
R1292 VGND.t549 VGND.t1522 644.952
R1293 VGND.t777 VGND.t781 644.952
R1294 VGND.n962 VGND 640.614
R1295 VGND VGND.n113 640.614
R1296 VGND VGND.n2859 640.614
R1297 VGND VGND.n2892 640.614
R1298 VGND.n2895 VGND 632.184
R1299 VGND.n990 VGND.n962 599.125
R1300 VGND.n113 VGND.n112 599.125
R1301 VGND.n2859 VGND.n2858 599.125
R1302 VGND.n2892 VGND.n2891 599.125
R1303 VGND.n2896 VGND.n2895 599.125
R1304 VGND.n2907 VGND.n2906 599.125
R1305 VGND.n2979 VGND.n2977 599.125
R1306 VGND.n2946 VGND.n2945 599.125
R1307 VGND.t1818 VGND 581.61
R1308 VGND.t456 VGND 573.181
R1309 VGND.t429 VGND 573.181
R1310 VGND.t1314 VGND 573.181
R1311 VGND VGND.t132 573.181
R1312 VGND.t710 VGND 564.751
R1313 VGND.n2997 VGND 564.751
R1314 VGND.n2996 VGND 564.751
R1315 VGND.n2995 VGND 556.322
R1316 VGND VGND.t1795 539.465
R1317 VGND.t308 VGND 539.465
R1318 VGND.n1122 VGND.t1580 514.663
R1319 VGND.t2593 VGND.n1131 514.663
R1320 VGND.n1132 VGND.t820 514.663
R1321 VGND.t837 VGND.n1144 514.663
R1322 VGND.n1145 VGND.t1584 514.663
R1323 VGND.t808 VGND.n1163 514.663
R1324 VGND.n1164 VGND.t899 514.663
R1325 VGND.t885 VGND.n1176 514.663
R1326 VGND.n1177 VGND.t1552 514.663
R1327 VGND.t800 VGND.n1195 514.663
R1328 VGND.n1196 VGND.t873 514.663
R1329 VGND.t853 VGND.n1208 514.663
R1330 VGND.n1209 VGND.t1539 514.663
R1331 VGND.t775 VGND.n1227 514.663
R1332 VGND.n1228 VGND.t862 514.663
R1333 VGND.t256 VGND.n578 494.779
R1334 VGND.t2369 VGND.t2310 481.877
R1335 VGND.t2310 VGND.t405 481.877
R1336 VGND.t2464 VGND.t2423 481.877
R1337 VGND.t2498 VGND.t2464 481.877
R1338 VGND.t2244 VGND 452.382
R1339 VGND.n1122 VGND.t595 424.053
R1340 VGND.n1131 VGND.t1244 424.053
R1341 VGND.n1132 VGND.t1966 424.053
R1342 VGND.n1144 VGND.t713 424.053
R1343 VGND.n1145 VGND.t1514 424.053
R1344 VGND.n1163 VGND.t1 424.053
R1345 VGND.n1164 VGND.t1716 424.053
R1346 VGND.n1176 VGND.t1515 424.053
R1347 VGND.n1177 VGND.t1310 424.053
R1348 VGND.n1195 VGND.t663 424.053
R1349 VGND.n1196 VGND.t1118 424.053
R1350 VGND.n1208 VGND.t1487 424.053
R1351 VGND.n1209 VGND.t231 424.053
R1352 VGND.n1227 VGND.t213 424.053
R1353 VGND.n1228 VGND.t2235 424.053
R1354 VGND.t604 VGND.n273 424.053
R1355 VGND.t178 VGND 419.68
R1356 VGND.n635 VGND.n147 413.043
R1357 VGND.t2496 VGND.t2415 397.848
R1358 VGND.t2415 VGND.t2425 397.848
R1359 VGND.t2425 VGND.t2433 397.848
R1360 VGND.t2433 VGND.t134 397.848
R1361 VGND.t134 VGND.t135 397.848
R1362 VGND.t135 VGND.t138 397.848
R1363 VGND.t138 VGND.t139 397.848
R1364 VGND.t1214 VGND.t2031 396.17
R1365 VGND.t1656 VGND.t1175 396.17
R1366 VGND.t1376 VGND.t857 394.137
R1367 VGND.t1527 VGND.t1328 394.137
R1368 VGND.t783 VGND.t1334 394.137
R1369 VGND.t1352 VGND.t764 394.137
R1370 VGND.t1531 VGND.t1427 394.137
R1371 VGND.t1433 VGND.t1529 394.137
R1372 VGND.t910 VGND.t1355 394.137
R1373 VGND.t1388 VGND.t846 394.137
R1374 VGND.t1586 VGND.t1400 394.137
R1375 VGND.t1445 VGND.t830 394.137
R1376 VGND.t903 VGND.t1364 394.137
R1377 VGND.t1403 VGND.t1573 394.137
R1378 VGND.t1558 VGND.t1448 394.137
R1379 VGND.t1457 VGND.t815 394.137
R1380 VGND.t878 VGND.t1370 394.137
R1381 VGND.t1565 VGND.t1415 394.137
R1382 VGND.t2173 VGND.t1391 394.137
R1383 VGND.t1031 VGND.t2559 394.137
R1384 VGND.t1980 VGND.t1958 394.137
R1385 VGND.t560 VGND.t1070 394.137
R1386 VGND.t1764 VGND.t929 394.137
R1387 VGND.t507 VGND.t1059 394.137
R1388 VGND.t2402 VGND.t2064 394.137
R1389 VGND.t952 VGND.t2029 394.137
R1390 VGND.t2552 VGND.t675 394.137
R1391 VGND.t987 VGND.t2644 394.137
R1392 VGND.t2272 VGND.t338 394.137
R1393 VGND.t2540 VGND.t108 394.137
R1394 VGND.t979 VGND.t485 394.137
R1395 VGND.t1005 VGND.t1810 394.137
R1396 VGND.t1839 VGND.t1475 394.137
R1397 VGND.t547 VGND.t1260 394.137
R1398 VGND.t2099 VGND.t1436 394.137
R1399 VGND.t1483 VGND.t633 394.137
R1400 VGND.t1938 VGND.t1823 394.137
R1401 VGND.t960 VGND.t30 394.137
R1402 VGND.t2561 VGND.t925 394.137
R1403 VGND.t580 VGND.t2073 394.137
R1404 VGND.t956 VGND.t2130 394.137
R1405 VGND.t1766 VGND.t517 394.137
R1406 VGND.t509 VGND.t2659 394.137
R1407 VGND.t2404 VGND.t274 394.137
R1408 VGND.t1865 VGND.t361 394.137
R1409 VGND.t495 VGND.t81 394.137
R1410 VGND.t2394 VGND.t740 394.137
R1411 VGND.t2276 VGND.t1759 394.137
R1412 VGND.t1262 VGND.t1170 394.137
R1413 VGND.t981 VGND.t659 394.137
R1414 VGND.t1343 VGND.t2550 394.137
R1415 VGND.t2386 VGND.t2653 394.137
R1416 VGND.t2268 VGND.t205 394.137
R1417 VGND.t68 VGND.t1847 394.137
R1418 VGND.t971 VGND.t1632 394.137
R1419 VGND.t2359 VGND.t2575 394.137
R1420 VGND.t1835 VGND.t311 394.137
R1421 VGND.t1183 VGND.t1252 394.137
R1422 VGND.t1778 VGND.t681 394.137
R1423 VGND.t1298 VGND.t1992 394.137
R1424 VGND.t2177 VGND.t397 394.137
R1425 VGND.t90 VGND.t1772 394.137
R1426 VGND.t1984 VGND.t2223 394.137
R1427 VGND.t586 VGND.t2210 394.137
R1428 VGND.t1873 VGND.t1156 394.137
R1429 VGND.t1890 VGND.t1700 394.137
R1430 VGND.t503 VGND.t1421 394.137
R1431 VGND.t944 VGND.t1105 394.137
R1432 VGND.t2089 VGND.t1859 394.137
R1433 VGND.t1268 VGND.t23 394.137
R1434 VGND.t2686 VGND.t2388 394.137
R1435 VGND.t647 VGND.t2197 394.137
R1436 VGND.t2602 VGND.t1254 394.137
R1437 VGND.t973 VGND.t1198 394.137
R1438 VGND.t666 VGND.t2577 394.137
R1439 VGND.t1837 VGND.t283 394.137
R1440 VGND.t218 VGND.t2103 394.137
R1441 VGND.t2569 VGND.t121 394.137
R1442 VGND.t300 VGND.t1829 394.137
R1443 VGND.t193 VGND.t2181 394.137
R1444 VGND.t1702 VGND.t1236 394.137
R1445 VGND.t538 VGND.t1988 394.137
R1446 VGND.t574 VGND.t1460 394.137
R1447 VGND.t1710 VGND.t1479 394.137
R1448 VGND.t2123 VGND.t1688 394.137
R1449 VGND.t1622 VGND.t991 394.137
R1450 VGND.t919 VGND.t946 394.137
R1451 VGND.t2203 VGND.t2546 394.137
R1452 VGND.t2126 VGND.t975 394.137
R1453 VGND.t1899 VGND.t2390 394.137
R1454 VGND.t1915 VGND.t651 394.137
R1455 VGND.t1306 VGND.t1256 394.137
R1456 VGND.t412 VGND.t1003 394.137
R1457 VGND.t77 VGND.t639 394.137
R1458 VGND.t289 VGND.t1250 394.137
R1459 VGND.t1753 VGND.t2105 394.137
R1460 VGND.t2043 VGND.t1990 394.137
R1461 VGND.t653 VGND.t1833 394.137
R1462 VGND.t1397 VGND.t966 394.137
R1463 VGND.t1996 VGND.t1029 394.137
R1464 VGND.t1608 VGND.t1956 394.137
R1465 VGND.t1068 VGND.t2396 394.137
R1466 VGND.t1706 VGND.t927 394.137
R1467 VGND.t1057 VGND.t997 394.137
R1468 VGND.t2382 VGND.t2062 394.137
R1469 VGND.t2027 VGND.t1879 394.137
R1470 VGND.t2534 VGND.t673 394.137
R1471 VGND.t2642 VGND.t1023 394.137
R1472 VGND.t2260 VGND.t336 394.137
R1473 VGND.t106 VGND.t1272 394.137
R1474 VGND.t1019 VGND.t483 394.137
R1475 VGND.t2585 VGND.t1808 394.137
R1476 VGND.t1827 VGND.t1473 394.137
R1477 VGND.t545 VGND.t2121 394.137
R1478 VGND.t1784 VGND.t1340 394.137
R1479 VGND.t1845 VGND.t2655 394.137
R1480 VGND.t207 VGND.t2185 394.137
R1481 VGND.t950 VGND.t70 394.137
R1482 VGND.t1634 VGND.t1998 394.137
R1483 VGND.t566 VGND.t2361 394.137
R1484 VGND.t313 VGND.t942 394.137
R1485 VGND.t1708 VGND.t721 394.137
R1486 VGND.t683 VGND.t493 394.137
R1487 VGND.t2384 VGND.t1300 394.137
R1488 VGND.t399 VGND.t1853 394.137
R1489 VGND.t993 VGND.t92 394.137
R1490 VGND.t2225 VGND.t2380 394.137
R1491 VGND.t2212 VGND.t2262 394.137
R1492 VGND.t1246 VGND.t1158 394.137
R1493 VGND.t1892 VGND.t1021 394.137
R1494 VGND.t1379 VGND.t2532 394.137
R1495 VGND.t1095 VGND.t2282 394.137
R1496 VGND.t2346 VGND.t2258 394.137
R1497 VGND.t452 VGND.t1831 394.137
R1498 VGND.t727 VGND.t1011 394.137
R1499 VGND.t1506 VGND.t2565 394.137
R1500 VGND.t2068 VGND.t2191 394.137
R1501 VGND.t306 VGND.t2115 394.137
R1502 VGND.t1972 VGND.t1770 394.137
R1503 VGND.t2674 VGND.t1978 394.137
R1504 VGND.t342 VGND.t2169 394.137
R1505 VGND.t102 VGND.t1712 394.137
R1506 VGND.t733 VGND.t1610 394.137
R1507 VGND.t1849 VGND.t578 394.137
R1508 VGND.t2255 VGND.t1861 394.137
R1509 VGND.t526 VGND.t1690 394.137
R1510 VGND.t995 VGND.t1424 394.137
R1511 VGND.t1875 VGND.t1103 394.137
R1512 VGND.t2556 VGND.t2523 394.137
R1513 VGND.t21 VGND.t1248 394.137
R1514 VGND.t2284 VGND.t2684 394.137
R1515 VGND.t2195 VGND.t635 394.137
R1516 VGND.t2117 VGND.t2600 394.137
R1517 VGND.t1195 VGND.t1013 394.137
R1518 VGND.t2567 VGND.t664 394.137
R1519 VGND.t281 VGND.t1821 394.137
R1520 VGND.t1788 VGND.t216 394.137
R1521 VGND.t119 VGND.t2002 394.137
R1522 VGND.t2187 VGND.t298 394.137
R1523 VGND.t2171 VGND.t1209 394.137
R1524 VGND.t1692 VGND.t1045 394.137
R1525 VGND.t535 VGND.t1612 394.137
R1526 VGND.t564 VGND.t1466 394.137
R1527 VGND.t1704 VGND.t381 394.137
R1528 VGND.t2353 VGND.t1686 394.137
R1529 VGND.t1025 VGND.t1617 394.137
R1530 VGND.t146 VGND.t1877 394.137
R1531 VGND.t2530 VGND.t2201 394.137
R1532 VGND.t317 VGND.t1015 394.137
R1533 VGND.t2378 VGND.t724 394.137
R1534 VGND.t1913 VGND.t637 394.137
R1535 VGND.t2119 VGND.t1304 394.137
R1536 VGND.t409 VGND.t2583 394.137
R1537 VGND.t629 VGND.t84 394.137
R1538 VGND.t1204 VGND.t2113 394.137
R1539 VGND.t1953 VGND.t2095 394.137
R1540 VGND.t1976 VGND.t2041 394.137
R1541 VGND.t1895 VGND.t2189 394.137
R1542 VGND.t2097 VGND.t1439 394.137
R1543 VGND.t627 VGND.t1481 394.137
R1544 VGND.t1936 VGND.t2193 394.137
R1545 VGND.t28 VGND.t958 394.137
R1546 VGND.t923 VGND.t2000 394.137
R1547 VGND.t2071 VGND.t576 394.137
R1548 VGND.t2128 VGND.t948 394.137
R1549 VGND.t185 VGND.t1762 394.137
R1550 VGND.t1919 VGND.t505 394.137
R1551 VGND.t272 VGND.t2398 394.137
R1552 VGND.t359 VGND.t1863 394.137
R1553 VGND.t79 VGND.t489 394.137
R1554 VGND.t738 VGND.t2392 394.137
R1555 VGND.t1757 VGND.t2270 394.137
R1556 VGND.t1168 VGND.t1258 394.137
R1557 VGND.t656 VGND.t977 394.137
R1558 VGND.t562 VGND.t1346 394.137
R1559 VGND.t1696 VGND.t2651 394.137
R1560 VGND.t513 VGND.t203 394.137
R1561 VGND.t66 VGND.t1017 394.137
R1562 VGND.t1871 VGND.t1630 394.137
R1563 VGND.t2357 VGND.t1270 394.137
R1564 VGND.t1009 VGND.t48 394.137
R1565 VGND.t1181 VGND.t2280 394.137
R1566 VGND.t631 VGND.t679 394.137
R1567 VGND.t1295 VGND.t2111 394.137
R1568 VGND.t2579 VGND.t395 394.137
R1569 VGND.t87 VGND.t625 394.137
R1570 VGND.t2109 VGND.t2221 394.137
R1571 VGND.t1780 VGND.t2208 394.137
R1572 VGND.t1606 VGND.t1154 394.137
R1573 VGND.t1888 VGND.t2183 394.137
R1574 VGND.t1412 VGND.t1698 394.137
R1575 VGND.t964 VGND.t588 394.137
R1576 VGND.t2093 VGND.t954 394.137
R1577 VGND.t2554 VGND.t25 394.137
R1578 VGND.t1140 VGND.t568 394.137
R1579 VGND.t2274 VGND.t1054 394.137
R1580 VGND.t2058 VGND.t2544 394.137
R1581 VGND.t497 VGND.t2023 394.137
R1582 VGND.t670 VGND.t1007 394.137
R1583 VGND.t649 VGND.t433 394.137
R1584 VGND.t220 VGND.t1264 394.137
R1585 VGND.t999 VGND.t114 394.137
R1586 VGND.t2052 VGND.t641 394.137
R1587 VGND.t197 VGND.t1843 394.137
R1588 VGND.t1774 VGND.t1239 394.137
R1589 VGND.t541 VGND.t2571 394.137
R1590 VGND.t1982 VGND.t1349 394.137
R1591 VGND.t2649 VGND.t1782 394.137
R1592 VGND.t1768 VGND.t201 394.137
R1593 VGND.t511 VGND.t64 394.137
R1594 VGND.t968 VGND.t2036 394.137
R1595 VGND.t1867 VGND.t2355 394.137
R1596 VGND.t499 VGND.t46 394.137
R1597 VGND.t570 VGND.t1178 394.137
R1598 VGND.t2278 VGND.t677 394.137
R1599 VGND.t2548 VGND.t1293 394.137
R1600 VGND.t983 VGND.t393 394.137
R1601 VGND.t2266 VGND.t100 394.137
R1602 VGND.t2536 VGND.t2219 394.137
R1603 VGND.t2206 VGND.t1266 394.137
R1604 VGND.t1152 VGND.t2573 394.137
R1605 VGND.t1885 VGND.t643 394.137
R1606 VGND.t1825 VGND.t1385 394.137
R1607 VGND.t2581 VGND.t1035 394.137
R1608 VGND.t2563 VGND.t1962 394.137
R1609 VGND.t1072 VGND.t582 394.137
R1610 VGND.t932 VGND.t1786 394.137
R1611 VGND.t1504 VGND.t1694 394.137
R1612 VGND.t2066 VGND.t572 394.137
R1613 VGND.t303 VGND.t2167 394.137
R1614 VGND.t1969 VGND.t1869 394.137
R1615 VGND.t2672 VGND.t501 394.137
R1616 VGND.t340 VGND.t2400 394.137
R1617 VGND.t110 VGND.t1857 394.137
R1618 VGND.t487 VGND.t491 394.137
R1619 VGND.t2216 VGND.t985 394.137
R1620 VGND.t645 VGND.t2253 394.137
R1621 VGND.t523 VGND.t2538 394.137
R1622 VGND.t2589 VGND.t989 394.137
R1623 VGND.t1855 VGND.t891 394.137
R1624 VGND.t2542 VGND.t1578 394.137
R1625 VGND.t2107 VGND.t1560 394.137
R1626 VGND.t2264 VGND.t895 394.137
R1627 VGND.t1841 VGND.t893 394.137
R1628 VGND.t2101 VGND.t1550 394.137
R1629 VGND.t1001 VGND.t806 394.137
R1630 VGND.t1994 VGND.t792 394.137
R1631 VGND.t2179 VGND.t869 394.137
R1632 VGND.t1776 VGND.t1537 394.137
R1633 VGND.t1986 VGND.t788 394.137
R1634 VGND.t2175 VGND.t770 394.137
R1635 VGND.t962 VGND.t851 394.137
R1636 VGND.t515 VGND.t1520 394.137
R1637 VGND.t773 VGND.t584 394.137
R1638 VGND.n147 VGND.t262 387.421
R1639 VGND.n1506 VGND.t4 387.421
R1640 VGND.n1508 VGND.t236 387.421
R1641 VGND.n1510 VGND.t2 387.421
R1642 VGND.n2818 VGND.t10 387.421
R1643 VGND.t1657 VGND.t460 362.452
R1644 VGND.t460 VGND.t308 345.594
R1645 VGND VGND.t8 328.616
R1646 VGND VGND.t13 328.616
R1647 VGND.t258 VGND 328.616
R1648 VGND.t176 VGND 328.616
R1649 VGND VGND.t16 328.616
R1650 VGND.t763 VGND.t761 326.195
R1651 VGND.t1524 VGND.t1526 326.195
R1652 VGND.t2597 VGND.t2595 326.195
R1653 VGND.t822 VGND.t824 326.195
R1654 VGND.t843 VGND.t841 326.195
R1655 VGND.t1570 VGND.t1572 326.195
R1656 VGND.t814 VGND.t812 326.195
R1657 VGND.t901 VGND.t890 326.195
R1658 VGND.t889 VGND.t887 326.195
R1659 VGND.t1556 VGND.t825 326.195
R1660 VGND.t805 VGND.t802 326.195
R1661 VGND.t875 VGND.t877 326.195
R1662 VGND.t1549 VGND.t1547 326.195
R1663 VGND.t1544 VGND.t1546 326.195
R1664 VGND.t782 VGND.t779 326.195
R1665 VGND.t866 VGND.t868 326.195
R1666 VGND.t1223 VGND.t1214 311.877
R1667 VGND.t1175 VGND.t1818 311.877
R1668 VGND VGND.t1219 303.449
R1669 VGND VGND.t1223 295.019
R1670 VGND.n70 VGND.t2424 287.832
R1671 VGND VGND.t58 286.591
R1672 VGND.n964 VGND.t253 282.327
R1673 VGND.n62 VGND.t2456 282.327
R1674 VGND.n969 VGND.t7 281.13
R1675 VGND.n73 VGND.t2495 281.13
R1676 VGND.n126 VGND.t9 280.978
R1677 VGND.n126 VGND.t2516 280.978
R1678 VGND.n594 VGND.t260 280.978
R1679 VGND.n594 VGND.t1076 280.978
R1680 VGND.n974 VGND.t406 280.978
R1681 VGND.n156 VGND.t271 280.978
R1682 VGND.n156 VGND.t1079 280.978
R1683 VGND.n96 VGND.t2440 280.978
R1684 VGND.n96 VGND.t2481 280.978
R1685 VGND.n2840 VGND.t2467 280.978
R1686 VGND.n2840 VGND.t2503 280.978
R1687 VGND.n2872 VGND.t2491 280.978
R1688 VGND.n2872 VGND.t2507 280.978
R1689 VGND.t226 VGND 278.161
R1690 VGND.n2978 VGND 271.014
R1691 VGND.n3004 VGND.n4 259.389
R1692 VGND.n2820 VGND.n4 259.389
R1693 VGND.n3005 VGND.n3 252.988
R1694 VGND VGND.t1216 252.875
R1695 VGND VGND.t1221 252.875
R1696 VGND.t2435 VGND 252.875
R1697 VGND VGND.t2431 252.875
R1698 VGND VGND.t2483 252.875
R1699 VGND.t859 VGND.t1376 250.815
R1700 VGND.t1328 VGND.t796 250.815
R1701 VGND.t1334 VGND.t785 250.815
R1702 VGND.t766 VGND.t1352 250.815
R1703 VGND.t1427 VGND.t1533 250.815
R1704 VGND.t1517 VGND.t1433 250.815
R1705 VGND.t1355 VGND.t912 250.815
R1706 VGND.t848 VGND.t1388 250.815
R1707 VGND.t1400 VGND.t1588 250.815
R1708 VGND.t832 VGND.t1445 250.815
R1709 VGND.t1364 VGND.t905 250.815
R1710 VGND.t1575 VGND.t1403 250.815
R1711 VGND.t1448 VGND.t826 250.815
R1712 VGND.t817 VGND.t1457 250.815
R1713 VGND.t1370 VGND.t880 250.815
R1714 VGND.t1415 VGND.t1567 250.815
R1715 VGND.t1083 VGND.t2173 250.815
R1716 VGND.t2559 VGND.t1121 250.815
R1717 VGND.t1093 VGND.t1980 250.815
R1718 VGND.t1091 VGND.t560 250.815
R1719 VGND.t2300 VGND.t1764 250.815
R1720 VGND.t2298 VGND.t507 250.815
R1721 VGND.t1089 VGND.t2402 250.815
R1722 VGND.t2308 VGND.t952 250.815
R1723 VGND.t2306 VGND.t2552 250.815
R1724 VGND.t1680 VGND.t987 250.815
R1725 VGND.t1087 VGND.t2272 250.815
R1726 VGND.t2304 VGND.t2540 250.815
R1727 VGND.t1678 VGND.t979 250.815
R1728 VGND.t1123 VGND.t1005 250.815
R1729 VGND.t1085 VGND.t1839 250.815
R1730 VGND.t1260 VGND.t2302 250.815
R1731 VGND.t938 VGND.t2099 250.815
R1732 VGND.t633 VGND.t617 250.815
R1733 VGND.t1823 VGND.t615 250.815
R1734 VGND.t613 VGND.t960 250.815
R1735 VGND.t2617 VGND.t2561 250.815
R1736 VGND.t2615 VGND.t580 250.815
R1737 VGND.t611 VGND.t956 250.815
R1738 VGND.t936 VGND.t1766 250.815
R1739 VGND.t934 VGND.t509 250.815
R1740 VGND.t623 VGND.t2404 250.815
R1741 VGND.t609 VGND.t1865 250.815
R1742 VGND.t2621 VGND.t495 250.815
R1743 VGND.t621 VGND.t2394 250.815
R1744 VGND.t619 VGND.t2276 250.815
R1745 VGND.t940 VGND.t1262 250.815
R1746 VGND.t2619 VGND.t981 250.815
R1747 VGND.t2550 VGND.t1287 250.815
R1748 VGND.t1125 VGND.t2386 250.815
R1749 VGND.t171 VGND.t2268 250.815
R1750 VGND.t1847 VGND.t169 250.815
R1751 VGND.t1135 VGND.t971 250.815
R1752 VGND.t2575 VGND.t1133 250.815
R1753 VGND.t167 VGND.t1835 250.815
R1754 VGND.t1252 VGND.t1285 250.815
R1755 VGND.t1283 VGND.t1778 250.815
R1756 VGND.t1992 VGND.t1131 250.815
R1757 VGND.t165 VGND.t2177 250.815
R1758 VGND.t1772 VGND.t1281 250.815
R1759 VGND.t1129 VGND.t1984 250.815
R1760 VGND.t1127 VGND.t586 250.815
R1761 VGND.t1289 VGND.t1873 250.815
R1762 VGND.t1700 VGND.t1279 250.815
R1763 VGND.t445 VGND.t503 250.815
R1764 VGND.t2606 VGND.t944 250.815
R1765 VGND.t1859 VGND.t1946 250.815
R1766 VGND.t1944 VGND.t1268 250.815
R1767 VGND.t2388 VGND.t250 250.815
R1768 VGND.t248 VGND.t647 250.815
R1769 VGND.t1254 VGND.t1942 250.815
R1770 VGND.t466 VGND.t973 250.815
R1771 VGND.t2577 VGND.t464 250.815
R1772 VGND.t2612 VGND.t1837 250.815
R1773 VGND.t2103 VGND.t449 250.815
R1774 VGND.t462 VGND.t2569 250.815
R1775 VGND.t1829 VGND.t2610 250.815
R1776 VGND.t2181 VGND.t2608 250.815
R1777 VGND.t447 VGND.t1702 250.815
R1778 VGND.t1988 VGND.t2669 250.815
R1779 VGND.t365 VGND.t574 250.815
R1780 VGND.t415 VGND.t1710 250.815
R1781 VGND.t1688 VGND.t375 250.815
R1782 VGND.t991 VGND.t373 250.815
R1783 VGND.t946 VGND.t425 250.815
R1784 VGND.t2546 VGND.t423 250.815
R1785 VGND.t975 VGND.t371 250.815
R1786 VGND.t2390 VGND.t391 250.815
R1787 VGND.t651 VGND.t389 250.815
R1788 VGND.t1256 VGND.t421 250.815
R1789 VGND.t1003 VGND.t369 250.815
R1790 VGND.t639 VGND.t387 250.815
R1791 VGND.t1250 VGND.t419 250.815
R1792 VGND.t2105 VGND.t417 250.815
R1793 VGND.t1990 VGND.t367 250.815
R1794 VGND.t1833 VGND.t427 250.815
R1795 VGND.t966 VGND.t1737 250.815
R1796 VGND.t439 VGND.t1996 250.815
R1797 VGND.t437 VGND.t1608 250.815
R1798 VGND.t2396 VGND.t435 250.815
R1799 VGND.t1725 VGND.t1706 250.815
R1800 VGND.t997 VGND.t1723 250.815
R1801 VGND.t1743 VGND.t2382 250.815
R1802 VGND.t1879 VGND.t1735 250.815
R1803 VGND.t1733 VGND.t2534 250.815
R1804 VGND.t1023 VGND.t1721 250.815
R1805 VGND.t1741 VGND.t2260 250.815
R1806 VGND.t1272 VGND.t1731 250.815
R1807 VGND.t1719 VGND.t1019 250.815
R1808 VGND.t441 VGND.t2585 250.815
R1809 VGND.t1739 VGND.t1827 250.815
R1810 VGND.t2121 VGND.t1729 250.815
R1811 VGND.t1602 VGND.t1784 250.815
R1812 VGND.t327 VGND.t1845 250.815
R1813 VGND.t2185 VGND.t325 250.815
R1814 VGND.t323 VGND.t950 250.815
R1815 VGND.t1998 VGND.t1592 250.815
R1816 VGND.t1590 VGND.t566 250.815
R1817 VGND.t942 VGND.t321 250.815
R1818 VGND.t1600 VGND.t1708 250.815
R1819 VGND.t493 VGND.t1598 250.815
R1820 VGND.t333 VGND.t2384 250.815
R1821 VGND.t1853 VGND.t319 250.815
R1822 VGND.t1596 VGND.t993 250.815
R1823 VGND.t2380 VGND.t331 250.815
R1824 VGND.t2262 VGND.t329 250.815
R1825 VGND.t385 VGND.t1246 250.815
R1826 VGND.t1021 VGND.t1594 250.815
R1827 VGND.t2532 VGND.t1226 250.815
R1828 VGND.t2282 VGND.t705 250.815
R1829 VGND.t2258 VGND.t703 250.815
R1830 VGND.t1831 VGND.t1234 250.815
R1831 VGND.t1011 VGND.t558 250.815
R1832 VGND.t2565 VGND.t556 250.815
R1833 VGND.t2191 VGND.t1232 250.815
R1834 VGND.t2115 VGND.t1166 250.815
R1835 VGND.t1770 VGND.t1164 250.815
R1836 VGND.t1978 VGND.t554 250.815
R1837 VGND.t2169 VGND.t1230 250.815
R1838 VGND.t1712 VGND.t1162 250.815
R1839 VGND.t1610 VGND.t552 250.815
R1840 VGND.t578 VGND.t214 250.815
R1841 VGND.t1861 VGND.t1228 250.815
R1842 VGND.t1690 VGND.t1160 250.815
R1843 VGND.t2625 VGND.t995 250.815
R1844 VGND.t2288 VGND.t1875 250.815
R1845 VGND.t2286 VGND.t2556 250.815
R1846 VGND.t1248 VGND.t2633 250.815
R1847 VGND.t1727 VGND.t2284 250.815
R1848 VGND.t635 VGND.t2296 250.815
R1849 VGND.t2631 VGND.t2117 250.815
R1850 VGND.t1013 VGND.t696 250.815
R1851 VGND.t694 VGND.t2567 250.815
R1852 VGND.t1821 VGND.t2294 250.815
R1853 VGND.t2629 VGND.t1788 250.815
R1854 VGND.t2002 VGND.t692 250.815
R1855 VGND.t2292 VGND.t2187 250.815
R1856 VGND.t2290 VGND.t2171 250.815
R1857 VGND.t2627 VGND.t1692 250.815
R1858 VGND.t1612 VGND.t690 250.815
R1859 VGND.t755 VGND.t564 250.815
R1860 VGND.t350 VGND.t1704 250.815
R1861 VGND.t1686 VGND.t348 250.815
R1862 VGND.t346 VGND.t1025 250.815
R1863 VGND.t1877 VGND.t1929 250.815
R1864 VGND.t1927 VGND.t2530 250.815
R1865 VGND.t1015 VGND.t2521 250.815
R1866 VGND.t1931 VGND.t2378 250.815
R1867 VGND.t637 VGND.t356 250.815
R1868 VGND.t1925 VGND.t2119 250.815
R1869 VGND.t2583 VGND.t2519 250.815
R1870 VGND.t354 VGND.t629 250.815
R1871 VGND.t2113 VGND.t1923 250.815
R1872 VGND.t2095 VGND.t1921 250.815
R1873 VGND.t2517 VGND.t1976 250.815
R1874 VGND.t2189 VGND.t352 250.815
R1875 VGND.t154 VGND.t2097 250.815
R1876 VGND.t1666 VGND.t627 250.815
R1877 VGND.t2193 VGND.t1664 250.815
R1878 VGND.t958 VGND.t1662 250.815
R1879 VGND.t2000 VGND.t1676 250.815
R1880 VGND.t576 VGND.t1674 250.815
R1881 VGND.t948 VGND.t1660 250.815
R1882 VGND.t1762 VGND.t152 250.815
R1883 VGND.t505 VGND.t150 250.815
R1884 VGND.t2398 VGND.t1672 250.815
R1885 VGND.t1863 VGND.t158 250.815
R1886 VGND.t489 VGND.t162 250.815
R1887 VGND.t2392 VGND.t1670 250.815
R1888 VGND.t2270 VGND.t1668 250.815
R1889 VGND.t1258 VGND.t156 250.815
R1890 VGND.t977 VGND.t160 250.815
R1891 VGND.t746 VGND.t562 250.815
R1892 VGND.t2017 VGND.t1696 250.815
R1893 VGND.t2015 VGND.t513 250.815
R1894 VGND.t1017 VGND.t2013 250.815
R1895 VGND.t1650 VGND.t1871 250.815
R1896 VGND.t1270 VGND.t1648 250.815
R1897 VGND.t1190 VGND.t1009 250.815
R1898 VGND.t2280 VGND.t744 250.815
R1899 VGND.t600 VGND.t631 250.815
R1900 VGND.t2111 VGND.t1646 250.815
R1901 VGND.t1188 VGND.t2579 250.815
R1902 VGND.t625 VGND.t598 250.815
R1903 VGND.t1644 VGND.t2109 250.815
R1904 VGND.t2019 VGND.t1780 250.815
R1905 VGND.t748 VGND.t1606 250.815
R1906 VGND.t2183 VGND.t596 250.815
R1907 VGND.t1698 VGND.t2159 250.815
R1908 VGND.t2328 VGND.t964 250.815
R1909 VGND.t954 VGND.t2326 250.815
R1910 VGND.t2324 VGND.t2554 250.815
R1911 VGND.t568 VGND.t1626 250.815
R1912 VGND.t2336 VGND.t2274 250.815
R1913 VGND.t2544 VGND.t2165 250.815
R1914 VGND.t2157 VGND.t497 250.815
R1915 VGND.t1007 VGND.t2155 250.815
R1916 VGND.t2334 VGND.t649 250.815
R1917 VGND.t1264 VGND.t2163 250.815
R1918 VGND.t2153 VGND.t999 250.815
R1919 VGND.t641 VGND.t2332 250.815
R1920 VGND.t1843 VGND.t2330 250.815
R1921 VGND.t2161 VGND.t1774 250.815
R1922 VGND.t2571 VGND.t2151 250.815
R1923 VGND.t2147 VGND.t1982 250.815
R1924 VGND.t1782 VGND.t1493 250.815
R1925 VGND.t1491 VGND.t1768 250.815
R1926 VGND.t475 VGND.t511 250.815
R1927 VGND.t2137 VGND.t968 250.815
R1928 VGND.t2135 VGND.t1867 250.815
R1929 VGND.t473 VGND.t499 250.815
R1930 VGND.t2145 VGND.t570 250.815
R1931 VGND.t2143 VGND.t2278 250.815
R1932 VGND.t1499 VGND.t2548 250.815
R1933 VGND.t471 VGND.t983 250.815
R1934 VGND.t2141 VGND.t2266 250.815
R1935 VGND.t1497 VGND.t2536 250.815
R1936 VGND.t1266 VGND.t1495 250.815
R1937 VGND.t2573 VGND.t2149 250.815
R1938 VGND.t643 VGND.t2139 250.815
R1939 VGND.t2079 VGND.t1825 250.815
R1940 VGND.t2322 VGND.t2581 250.815
R1941 VGND.t2320 VGND.t2563 250.815
R1942 VGND.t582 VGND.t2318 250.815
R1943 VGND.t1786 VGND.t1751 250.815
R1944 VGND.t1694 VGND.t1749 250.815
R1945 VGND.t572 VGND.t2316 250.815
R1946 VGND.t2167 VGND.t2077 250.815
R1947 VGND.t1869 VGND.t2050 250.815
R1948 VGND.t501 VGND.t1747 250.815
R1949 VGND.t2400 VGND.t2083 250.815
R1950 VGND.t1857 VGND.t2048 250.815
R1951 VGND.t491 VGND.t2087 250.815
R1952 VGND.t985 VGND.t2085 250.815
R1953 VGND.t2081 VGND.t645 250.815
R1954 VGND.t2538 VGND.t2046 250.815
R1955 VGND.t989 VGND.t2591 250.815
R1956 VGND.t839 VGND.t1855 250.815
R1957 VGND.t1582 VGND.t2542 250.815
R1958 VGND.t1562 VGND.t2107 250.815
R1959 VGND.t897 VGND.t2264 250.815
R1960 VGND.t883 VGND.t1841 250.815
R1961 VGND.t1554 VGND.t2101 250.815
R1962 VGND.t810 VGND.t1001 250.815
R1963 VGND.t794 VGND.t1994 250.815
R1964 VGND.t871 VGND.t2179 250.815
R1965 VGND.t1541 VGND.t1776 250.815
R1966 VGND.t790 VGND.t1986 250.815
R1967 VGND.t864 VGND.t2175 250.815
R1968 VGND.t855 VGND.t962 250.815
R1969 VGND.t1522 VGND.t515 250.815
R1970 VGND.t584 VGND.t777 250.815
R1971 VGND.n2573 VGND.t1377 241.405
R1972 VGND.n229 VGND.t2174 241.405
R1973 VGND.n239 VGND.t2100 241.405
R1974 VGND.n179 VGND.t2551 241.405
R1975 VGND.n1419 VGND.t504 241.405
R1976 VGND.n637 VGND.t575 241.405
R1977 VGND.n616 VGND.t967 241.405
R1978 VGND.n643 VGND.t1785 241.405
R1979 VGND.n659 VGND.t2533 241.405
R1980 VGND.n668 VGND.t996 241.405
R1981 VGND.n1371 VGND.t565 241.405
R1982 VGND.n1303 VGND.t2098 241.405
R1983 VGND.n572 VGND.t563 241.405
R1984 VGND.n568 VGND.t1699 241.405
R1985 VGND.n671 VGND.t1983 241.405
R1986 VGND.n825 VGND.t1826 241.405
R1987 VGND.n815 VGND.t1383 241.405
R1988 VGND.n676 VGND.t990 241.405
R1989 VGND.n2691 VGND.t1329 241.284
R1990 VGND.n2621 VGND.t1335 241.284
R1991 VGND.n2685 VGND.t1353 241.284
R1992 VGND.n2623 VGND.t1428 241.284
R1993 VGND.n2678 VGND.t1434 241.284
R1994 VGND.n2626 VGND.t1356 241.284
R1995 VGND.n2671 VGND.t1389 241.284
R1996 VGND.n2629 VGND.t1401 241.284
R1997 VGND.n2664 VGND.t1446 241.284
R1998 VGND.n2632 VGND.t1365 241.284
R1999 VGND.n2657 VGND.t1404 241.284
R2000 VGND.n2635 VGND.t1449 241.284
R2001 VGND.n2650 VGND.t1458 241.284
R2002 VGND.n2638 VGND.t1371 241.284
R2003 VGND.n2643 VGND.t1416 241.284
R2004 VGND.n232 VGND.t2560 241.284
R2005 VGND.n2702 VGND.t1981 241.284
R2006 VGND.n2707 VGND.t561 241.284
R2007 VGND.n2712 VGND.t1765 241.284
R2008 VGND.n2717 VGND.t508 241.284
R2009 VGND.n2722 VGND.t2403 241.284
R2010 VGND.n2727 VGND.t953 241.284
R2011 VGND.n2732 VGND.t2553 241.284
R2012 VGND.n2737 VGND.t988 241.284
R2013 VGND.n2742 VGND.t2273 241.284
R2014 VGND.n2747 VGND.t2541 241.284
R2015 VGND.n2752 VGND.t980 241.284
R2016 VGND.n2757 VGND.t1006 241.284
R2017 VGND.n2762 VGND.t1840 241.284
R2018 VGND.n227 VGND.t1261 241.284
R2019 VGND.n242 VGND.t634 241.284
R2020 VGND.n2511 VGND.t1824 241.284
R2021 VGND.n2506 VGND.t961 241.284
R2022 VGND.n246 VGND.t2562 241.284
R2023 VGND.n2436 VGND.t581 241.284
R2024 VGND.n2441 VGND.t957 241.284
R2025 VGND.n2446 VGND.t1767 241.284
R2026 VGND.n2451 VGND.t510 241.284
R2027 VGND.n2456 VGND.t2405 241.284
R2028 VGND.n2461 VGND.t1866 241.284
R2029 VGND.n2466 VGND.t496 241.284
R2030 VGND.n2471 VGND.t2395 241.284
R2031 VGND.n2476 VGND.t2277 241.284
R2032 VGND.n2481 VGND.t1263 241.284
R2033 VGND.n2486 VGND.t982 241.284
R2034 VGND.n2814 VGND.t2387 241.284
R2035 VGND.n366 VGND.t2269 241.284
R2036 VGND.n370 VGND.t1848 241.284
R2037 VGND.n2169 VGND.t972 241.284
R2038 VGND.n364 VGND.t2576 241.284
R2039 VGND.n2195 VGND.t1836 241.284
R2040 VGND.n356 VGND.t1253 241.284
R2041 VGND.n2221 VGND.t1779 241.284
R2042 VGND.n348 VGND.t1993 241.284
R2043 VGND.n2247 VGND.t2178 241.284
R2044 VGND.n340 VGND.t1773 241.284
R2045 VGND.n2278 VGND.t1985 241.284
R2046 VGND.n2283 VGND.t587 241.284
R2047 VGND.n2288 VGND.t1874 241.284
R2048 VGND.n332 VGND.t1701 241.284
R2049 VGND.n1426 VGND.t945 241.284
R2050 VGND.n1423 VGND.t1860 241.284
R2051 VGND.n2156 VGND.t1269 241.284
R2052 VGND.n379 VGND.t2389 241.284
R2053 VGND.n2182 VGND.t648 241.284
R2054 VGND.n360 VGND.t1255 241.284
R2055 VGND.n2208 VGND.t974 241.284
R2056 VGND.n352 VGND.t2578 241.284
R2057 VGND.n2234 VGND.t1838 241.284
R2058 VGND.n344 VGND.t2104 241.284
R2059 VGND.n2260 VGND.t2570 241.284
R2060 VGND.n336 VGND.t1830 241.284
R2061 VGND.n2265 VGND.t2182 241.284
R2062 VGND.n2305 VGND.t1703 241.284
R2063 VGND.n2310 VGND.t1989 241.284
R2064 VGND.n1440 VGND.t1711 241.284
R2065 VGND.n634 VGND.t1689 241.284
R2066 VGND.n1490 VGND.t992 241.284
R2067 VGND.n1485 VGND.t947 241.284
R2068 VGND.n1480 VGND.t2547 241.284
R2069 VGND.n1475 VGND.t976 241.284
R2070 VGND.n1470 VGND.t2391 241.284
R2071 VGND.n1465 VGND.t652 241.284
R2072 VGND.n1460 VGND.t1257 241.284
R2073 VGND.n1455 VGND.t1004 241.284
R2074 VGND.n1450 VGND.t640 241.284
R2075 VGND.n1445 VGND.t1251 241.284
R2076 VGND.n393 VGND.t2106 241.284
R2077 VGND.n2133 VGND.t1991 241.284
R2078 VGND.n2128 VGND.t1834 241.284
R2079 VGND.n1502 VGND.t1997 241.284
R2080 VGND.n621 VGND.t1609 241.284
R2081 VGND.n625 VGND.t2397 241.284
R2082 VGND.n1995 VGND.t1707 241.284
R2083 VGND.n431 VGND.t998 241.284
R2084 VGND.n2021 VGND.t2383 241.284
R2085 VGND.n423 VGND.t1880 241.284
R2086 VGND.n2047 VGND.t2535 241.284
R2087 VGND.n415 VGND.t1024 241.284
R2088 VGND.n2073 VGND.t2261 241.284
R2089 VGND.n407 VGND.t1273 241.284
R2090 VGND.n2104 VGND.t1020 241.284
R2091 VGND.n2109 VGND.t2586 241.284
R2092 VGND.n2114 VGND.t1828 241.284
R2093 VGND.n2119 VGND.t2122 241.284
R2094 VGND.n650 VGND.t1846 241.284
R2095 VGND.n647 VGND.t2186 241.284
R2096 VGND.n1982 VGND.t951 241.284
R2097 VGND.n435 VGND.t1999 241.284
R2098 VGND.n2008 VGND.t567 241.284
R2099 VGND.n427 VGND.t943 241.284
R2100 VGND.n2034 VGND.t1709 241.284
R2101 VGND.n419 VGND.t494 241.284
R2102 VGND.n2060 VGND.t2385 241.284
R2103 VGND.n411 VGND.t1854 241.284
R2104 VGND.n2086 VGND.t994 241.284
R2105 VGND.n403 VGND.t2381 241.284
R2106 VGND.n2091 VGND.t2263 241.284
R2107 VGND.n2330 VGND.t1247 241.284
R2108 VGND.n2335 VGND.t1022 241.284
R2109 VGND.n957 VGND.t2283 241.284
R2110 VGND.n952 VGND.t2259 241.284
R2111 VGND.n947 VGND.t1832 241.284
R2112 VGND.n942 VGND.t1012 241.284
R2113 VGND.n937 VGND.t2566 241.284
R2114 VGND.n932 VGND.t2192 241.284
R2115 VGND.n927 VGND.t2116 241.284
R2116 VGND.n922 VGND.t1771 241.284
R2117 VGND.n917 VGND.t1979 241.284
R2118 VGND.n912 VGND.t2170 241.284
R2119 VGND.n907 VGND.t1713 241.284
R2120 VGND.n902 VGND.t1611 241.284
R2121 VGND.n449 VGND.t579 241.284
R2122 VGND.n1959 VGND.t1862 241.284
R2123 VGND.n1954 VGND.t1691 241.284
R2124 VGND.n1393 VGND.t1876 241.284
R2125 VGND.n1398 VGND.t2557 241.284
R2126 VGND.n666 VGND.t1249 241.284
R2127 VGND.n1821 VGND.t2285 241.284
R2128 VGND.n487 VGND.t636 241.284
R2129 VGND.n1847 VGND.t2118 241.284
R2130 VGND.n479 VGND.t1014 241.284
R2131 VGND.n1873 VGND.t2568 241.284
R2132 VGND.n471 VGND.t1822 241.284
R2133 VGND.n1899 VGND.t1789 241.284
R2134 VGND.n463 VGND.t2003 241.284
R2135 VGND.n1930 VGND.t2188 241.284
R2136 VGND.n1935 VGND.t2172 241.284
R2137 VGND.n1940 VGND.t1693 241.284
R2138 VGND.n1945 VGND.t1613 241.284
R2139 VGND.n1378 VGND.t1705 241.284
R2140 VGND.n1375 VGND.t1687 241.284
R2141 VGND.n1808 VGND.t1026 241.284
R2142 VGND.n491 VGND.t1878 241.284
R2143 VGND.n1834 VGND.t2531 241.284
R2144 VGND.n483 VGND.t1016 241.284
R2145 VGND.n1860 VGND.t2379 241.284
R2146 VGND.n475 VGND.t638 241.284
R2147 VGND.n1886 VGND.t2120 241.284
R2148 VGND.n467 VGND.t2584 241.284
R2149 VGND.n1912 VGND.t630 241.284
R2150 VGND.n459 VGND.t2114 241.284
R2151 VGND.n1917 VGND.t2096 241.284
R2152 VGND.n2355 VGND.t1977 241.284
R2153 VGND.n2360 VGND.t2190 241.284
R2154 VGND.n1310 VGND.t628 241.284
R2155 VGND.n1307 VGND.t2194 241.284
R2156 VGND.n1360 VGND.t959 241.284
R2157 VGND.n1355 VGND.t2001 241.284
R2158 VGND.n1350 VGND.t577 241.284
R2159 VGND.n1345 VGND.t949 241.284
R2160 VGND.n1340 VGND.t1763 241.284
R2161 VGND.n1335 VGND.t506 241.284
R2162 VGND.n1330 VGND.t2399 241.284
R2163 VGND.n1325 VGND.t1864 241.284
R2164 VGND.n1320 VGND.t490 241.284
R2165 VGND.n1315 VGND.t2393 241.284
R2166 VGND.n505 VGND.t2271 241.284
R2167 VGND.n1785 VGND.t1259 241.284
R2168 VGND.n1780 VGND.t978 241.284
R2169 VGND.n1515 VGND.t1697 241.284
R2170 VGND.n1520 VGND.t514 241.284
R2171 VGND.n577 VGND.t1018 241.284
R2172 VGND.n1647 VGND.t1872 241.284
R2173 VGND.n543 VGND.t1271 241.284
R2174 VGND.n1673 VGND.t1010 241.284
R2175 VGND.n535 VGND.t2281 241.284
R2176 VGND.n1699 VGND.t632 241.284
R2177 VGND.n527 VGND.t2112 241.284
R2178 VGND.n1725 VGND.t2580 241.284
R2179 VGND.n519 VGND.t626 241.284
R2180 VGND.n1756 VGND.t2110 241.284
R2181 VGND.n1761 VGND.t1781 241.284
R2182 VGND.n1766 VGND.t1607 241.284
R2183 VGND.n1771 VGND.t2184 241.284
R2184 VGND.n1535 VGND.t965 241.284
R2185 VGND.n566 VGND.t955 241.284
R2186 VGND.n1634 VGND.t2555 241.284
R2187 VGND.n547 VGND.t569 241.284
R2188 VGND.n1660 VGND.t2275 241.284
R2189 VGND.n539 VGND.t2545 241.284
R2190 VGND.n1686 VGND.t498 241.284
R2191 VGND.n531 VGND.t1008 241.284
R2192 VGND.n1712 VGND.t650 241.284
R2193 VGND.n523 VGND.t1265 241.284
R2194 VGND.n1738 VGND.t1000 241.284
R2195 VGND.n515 VGND.t642 241.284
R2196 VGND.n1743 VGND.t1844 241.284
R2197 VGND.n2380 VGND.t1775 241.284
R2198 VGND.n2385 VGND.t2572 241.284
R2199 VGND.n674 VGND.t1783 241.284
R2200 VGND.n1548 VGND.t1769 241.284
R2201 VGND.n1553 VGND.t512 241.284
R2202 VGND.n1558 VGND.t969 241.284
R2203 VGND.n1563 VGND.t1868 241.284
R2204 VGND.n1568 VGND.t500 241.284
R2205 VGND.n1573 VGND.t571 241.284
R2206 VGND.n1578 VGND.t2279 241.284
R2207 VGND.n1583 VGND.t2549 241.284
R2208 VGND.n1588 VGND.t984 241.284
R2209 VGND.n1593 VGND.t2267 241.284
R2210 VGND.n1598 VGND.t2537 241.284
R2211 VGND.n561 VGND.t1267 241.284
R2212 VGND.n1611 VGND.t2574 241.284
R2213 VGND.n1606 VGND.t644 241.284
R2214 VGND.n833 VGND.t2582 241.284
R2215 VGND.n838 VGND.t2564 241.284
R2216 VGND.n830 VGND.t583 241.284
R2217 VGND.n888 VGND.t1787 241.284
R2218 VGND.n883 VGND.t1695 241.284
R2219 VGND.n878 VGND.t573 241.284
R2220 VGND.n873 VGND.t2168 241.284
R2221 VGND.n868 VGND.t1870 241.284
R2222 VGND.n863 VGND.t502 241.284
R2223 VGND.n858 VGND.t2401 241.284
R2224 VGND.n853 VGND.t1858 241.284
R2225 VGND.n848 VGND.t492 241.284
R2226 VGND.n843 VGND.t986 241.284
R2227 VGND.n2400 VGND.t646 241.284
R2228 VGND.n2405 VGND.t2539 241.284
R2229 VGND.n1124 VGND.t1332 241.284
R2230 VGND.n1129 VGND.t1338 241.284
R2231 VGND.n1134 VGND.t1359 241.284
R2232 VGND.n1142 VGND.t1431 241.284
R2233 VGND.n810 VGND.t1443 241.284
R2234 VGND.n1161 VGND.t1362 241.284
R2235 VGND.n1166 VGND.t1395 241.284
R2236 VGND.n1174 VGND.t1407 241.284
R2237 VGND.n802 VGND.t1452 241.284
R2238 VGND.n1193 VGND.t1368 241.284
R2239 VGND.n1198 VGND.t1410 241.284
R2240 VGND.n1206 VGND.t1455 241.284
R2241 VGND.n794 VGND.t1464 241.284
R2242 VGND.n1225 VGND.t1374 241.284
R2243 VGND.n1230 VGND.t1419 241.284
R2244 VGND.n1287 VGND.t1856 241.284
R2245 VGND.n683 VGND.t2543 241.284
R2246 VGND.n723 VGND.t2108 241.284
R2247 VGND.n728 VGND.t2265 241.284
R2248 VGND.n733 VGND.t1842 241.284
R2249 VGND.n738 VGND.t2102 241.284
R2250 VGND.n743 VGND.t1002 241.284
R2251 VGND.n748 VGND.t1995 241.284
R2252 VGND.n753 VGND.t2180 241.284
R2253 VGND.n758 VGND.t1777 241.284
R2254 VGND.n763 VGND.t1987 241.284
R2255 VGND.n768 VGND.t2176 241.284
R2256 VGND.n773 VGND.t963 241.284
R2257 VGND.n778 VGND.t516 241.284
R2258 VGND.n719 VGND.t585 241.284
R2259 VGND.n2819 VGND.n3 218.73
R2260 VGND.n133 VGND.n131 214.365
R2261 VGND.n133 VGND.n132 214.365
R2262 VGND.n123 VGND.n121 214.365
R2263 VGND.n123 VGND.n122 214.365
R2264 VGND.n141 VGND.n139 214.365
R2265 VGND.n141 VGND.n140 214.365
R2266 VGND.n601 VGND.n599 214.365
R2267 VGND.n601 VGND.n600 214.365
R2268 VGND.n591 VGND.n589 214.365
R2269 VGND.n591 VGND.n590 214.365
R2270 VGND.n609 VGND.n607 214.365
R2271 VGND.n609 VGND.n608 214.365
R2272 VGND.n971 VGND.n970 214.365
R2273 VGND.n163 VGND.n161 214.365
R2274 VGND.n163 VGND.n162 214.365
R2275 VGND.n153 VGND.n151 214.365
R2276 VGND.n153 VGND.n152 214.365
R2277 VGND.n171 VGND.n169 214.365
R2278 VGND.n171 VGND.n170 214.365
R2279 VGND.n1096 VGND.n1095 213.613
R2280 VGND.n1098 VGND.n1097 213.613
R2281 VGND.n1068 VGND.n1066 213.613
R2282 VGND.n1068 VGND.n1067 213.613
R2283 VGND.n1071 VGND.n1069 213.613
R2284 VGND.n1071 VGND.n1070 213.613
R2285 VGND.n1006 VGND.n1004 213.613
R2286 VGND.n1006 VGND.n1005 213.613
R2287 VGND.n1009 VGND.n1007 213.613
R2288 VGND.n1009 VGND.n1008 213.613
R2289 VGND.n1037 VGND.n1035 213.613
R2290 VGND.n1037 VGND.n1036 213.613
R2291 VGND.n1040 VGND.n1038 213.613
R2292 VGND.n1040 VGND.n1039 213.613
R2293 VGND.n1110 VGND.t50 212.422
R2294 VGND.n968 VGND.n967 207.965
R2295 VGND.n985 VGND.n965 207.965
R2296 VGND.n98 VGND.n94 207.965
R2297 VGND.n98 VGND.n95 207.965
R2298 VGND.n92 VGND.n90 207.965
R2299 VGND.n92 VGND.n91 207.965
R2300 VGND.n105 VGND.n88 207.965
R2301 VGND.n105 VGND.n89 207.965
R2302 VGND.n2842 VGND.n2838 207.965
R2303 VGND.n2842 VGND.n2839 207.965
R2304 VGND.n2836 VGND.n2834 207.965
R2305 VGND.n2836 VGND.n2835 207.965
R2306 VGND.n2849 VGND.n2832 207.965
R2307 VGND.n2849 VGND.n2833 207.965
R2308 VGND.n2874 VGND.n2870 207.965
R2309 VGND.n2874 VGND.n2871 207.965
R2310 VGND.n2868 VGND.n2866 207.965
R2311 VGND.n2868 VGND.n2867 207.965
R2312 VGND.n2881 VGND.n2864 207.965
R2313 VGND.n2881 VGND.n2865 207.965
R2314 VGND.n67 VGND.n66 207.965
R2315 VGND.n79 VGND.n64 207.965
R2316 VGND.n71 VGND.n69 207.965
R2317 VGND.n984 VGND.n966 207.213
R2318 VGND.n14 VGND.n13 207.213
R2319 VGND.n18 VGND.n12 207.213
R2320 VGND.n43 VGND.n41 207.213
R2321 VGND.n43 VGND.n42 207.213
R2322 VGND.n47 VGND.n39 207.213
R2323 VGND.n47 VGND.n40 207.213
R2324 VGND.n78 VGND.n65 207.213
R2325 VGND.n2916 VGND.n2914 207.213
R2326 VGND.n2916 VGND.n2915 207.213
R2327 VGND.n2920 VGND.n2911 207.213
R2328 VGND.n2920 VGND.n2912 207.213
R2329 VGND.n2956 VGND.n2954 207.213
R2330 VGND.n2956 VGND.n2955 207.213
R2331 VGND.n2960 VGND.n2952 207.213
R2332 VGND.n2960 VGND.n2953 207.213
R2333 VGND.t1382 VGND.t759 199.341
R2334 VGND.t1580 VGND.t1331 199.341
R2335 VGND.t1337 VGND.t2593 199.341
R2336 VGND.t820 VGND.t1358 199.341
R2337 VGND.t1430 VGND.t837 199.341
R2338 VGND.t1584 VGND.t1442 199.341
R2339 VGND.t1361 VGND.t808 199.341
R2340 VGND.t899 VGND.t1394 199.341
R2341 VGND.t1406 VGND.t885 199.341
R2342 VGND.t1552 VGND.t1451 199.341
R2343 VGND.t1367 VGND.t800 199.341
R2344 VGND.t873 VGND.t1409 199.341
R2345 VGND.t1454 VGND.t853 199.341
R2346 VGND.t1539 VGND.t1463 199.341
R2347 VGND.t1373 VGND.t775 199.341
R2348 VGND.t862 VGND.t1418 199.341
R2349 VGND VGND.n2641 194.423
R2350 VGND VGND.n2639 194.423
R2351 VGND VGND.n2648 194.423
R2352 VGND VGND.n2636 194.423
R2353 VGND VGND.n2655 194.423
R2354 VGND VGND.n2633 194.423
R2355 VGND VGND.n2662 194.423
R2356 VGND VGND.n2630 194.423
R2357 VGND VGND.n2669 194.423
R2358 VGND VGND.n2627 194.423
R2359 VGND VGND.n2676 194.423
R2360 VGND VGND.n2624 194.423
R2361 VGND VGND.n2683 194.423
R2362 VGND VGND.n2620 194.423
R2363 VGND VGND.n2571 194.423
R2364 VGND.n2573 VGND.n2572 194.405
R2365 VGND.n226 VGND.n225 194.405
R2366 VGND.n2761 VGND.n2760 194.405
R2367 VGND.n2756 VGND.n2755 194.405
R2368 VGND.n2751 VGND.n2750 194.405
R2369 VGND.n2746 VGND.n2745 194.405
R2370 VGND.n2741 VGND.n2740 194.405
R2371 VGND.n2736 VGND.n2735 194.405
R2372 VGND.n2731 VGND.n2730 194.405
R2373 VGND.n2726 VGND.n2725 194.405
R2374 VGND.n2721 VGND.n2720 194.405
R2375 VGND.n2716 VGND.n2715 194.405
R2376 VGND.n2711 VGND.n2710 194.405
R2377 VGND.n2706 VGND.n2705 194.405
R2378 VGND.n2701 VGND.n2700 194.405
R2379 VGND.n231 VGND.n230 194.405
R2380 VGND.n229 VGND.n228 194.405
R2381 VGND.n2485 VGND.n2484 194.405
R2382 VGND.n2480 VGND.n2479 194.405
R2383 VGND.n2475 VGND.n2474 194.405
R2384 VGND.n2470 VGND.n2469 194.405
R2385 VGND.n2465 VGND.n2464 194.405
R2386 VGND.n2460 VGND.n2459 194.405
R2387 VGND.n2455 VGND.n2454 194.405
R2388 VGND.n2450 VGND.n2449 194.405
R2389 VGND.n2445 VGND.n2444 194.405
R2390 VGND.n2440 VGND.n2439 194.405
R2391 VGND.n2435 VGND.n2434 194.405
R2392 VGND.n247 VGND.n245 194.405
R2393 VGND.n2505 VGND.n243 194.405
R2394 VGND.n2510 VGND.n2509 194.405
R2395 VGND.n241 VGND.n240 194.405
R2396 VGND.n239 VGND.n238 194.405
R2397 VGND.n331 VGND.n330 194.405
R2398 VGND.n2287 VGND.n2286 194.405
R2399 VGND.n2282 VGND.n2281 194.405
R2400 VGND.n2277 VGND.n2276 194.405
R2401 VGND.n339 VGND.n338 194.405
R2402 VGND.n2246 VGND.n2245 194.405
R2403 VGND.n347 VGND.n346 194.405
R2404 VGND.n2220 VGND.n2219 194.405
R2405 VGND.n355 VGND.n354 194.405
R2406 VGND.n2194 VGND.n2193 194.405
R2407 VGND.n363 VGND.n362 194.405
R2408 VGND.n2168 VGND.n2167 194.405
R2409 VGND.n369 VGND.n368 194.405
R2410 VGND.n367 VGND.n365 194.405
R2411 VGND.n2813 VGND.n181 194.405
R2412 VGND.n179 VGND.n178 194.405
R2413 VGND.n2311 VGND.n326 194.405
R2414 VGND.n2304 VGND.n2303 194.405
R2415 VGND.n2264 VGND.n2263 194.405
R2416 VGND.n335 VGND.n334 194.405
R2417 VGND.n2259 VGND.n2258 194.405
R2418 VGND.n343 VGND.n342 194.405
R2419 VGND.n2233 VGND.n2232 194.405
R2420 VGND.n351 VGND.n350 194.405
R2421 VGND.n2207 VGND.n2206 194.405
R2422 VGND.n359 VGND.n358 194.405
R2423 VGND.n2181 VGND.n2180 194.405
R2424 VGND.n378 VGND.n377 194.405
R2425 VGND.n2155 VGND.n2154 194.405
R2426 VGND.n1422 VGND.n1421 194.405
R2427 VGND.n1425 VGND.n1424 194.405
R2428 VGND.n1419 VGND.n1418 194.405
R2429 VGND.n2127 VGND.n394 194.405
R2430 VGND.n2132 VGND.n2131 194.405
R2431 VGND.n392 VGND.n391 194.405
R2432 VGND.n1444 VGND.n1443 194.405
R2433 VGND.n1449 VGND.n1448 194.405
R2434 VGND.n1454 VGND.n1453 194.405
R2435 VGND.n1459 VGND.n1458 194.405
R2436 VGND.n1464 VGND.n1463 194.405
R2437 VGND.n1469 VGND.n1468 194.405
R2438 VGND.n1474 VGND.n1473 194.405
R2439 VGND.n1479 VGND.n1478 194.405
R2440 VGND.n1484 VGND.n1483 194.405
R2441 VGND.n1489 VGND.n1488 194.405
R2442 VGND.n633 VGND.n632 194.405
R2443 VGND.n1439 VGND.n1438 194.405
R2444 VGND.n637 VGND.n636 194.405
R2445 VGND.n2120 VGND.n397 194.405
R2446 VGND.n2113 VGND.n2112 194.405
R2447 VGND.n2108 VGND.n2107 194.405
R2448 VGND.n2103 VGND.n2102 194.405
R2449 VGND.n406 VGND.n405 194.405
R2450 VGND.n2072 VGND.n2071 194.405
R2451 VGND.n414 VGND.n413 194.405
R2452 VGND.n2046 VGND.n2045 194.405
R2453 VGND.n422 VGND.n421 194.405
R2454 VGND.n2020 VGND.n2019 194.405
R2455 VGND.n430 VGND.n429 194.405
R2456 VGND.n1994 VGND.n1993 194.405
R2457 VGND.n624 VGND.n623 194.405
R2458 VGND.n622 VGND.n620 194.405
R2459 VGND.n1501 VGND.n618 194.405
R2460 VGND.n616 VGND.n615 194.405
R2461 VGND.n2336 VGND.n315 194.405
R2462 VGND.n2329 VGND.n2328 194.405
R2463 VGND.n2090 VGND.n2089 194.405
R2464 VGND.n402 VGND.n401 194.405
R2465 VGND.n2085 VGND.n2084 194.405
R2466 VGND.n410 VGND.n409 194.405
R2467 VGND.n2059 VGND.n2058 194.405
R2468 VGND.n418 VGND.n417 194.405
R2469 VGND.n2033 VGND.n2032 194.405
R2470 VGND.n426 VGND.n425 194.405
R2471 VGND.n2007 VGND.n2006 194.405
R2472 VGND.n434 VGND.n433 194.405
R2473 VGND.n1981 VGND.n1980 194.405
R2474 VGND.n646 VGND.n645 194.405
R2475 VGND.n649 VGND.n648 194.405
R2476 VGND.n643 VGND.n642 194.405
R2477 VGND.n1953 VGND.n450 194.405
R2478 VGND.n1958 VGND.n1957 194.405
R2479 VGND.n448 VGND.n447 194.405
R2480 VGND.n901 VGND.n900 194.405
R2481 VGND.n906 VGND.n905 194.405
R2482 VGND.n911 VGND.n910 194.405
R2483 VGND.n916 VGND.n915 194.405
R2484 VGND.n921 VGND.n920 194.405
R2485 VGND.n926 VGND.n925 194.405
R2486 VGND.n931 VGND.n930 194.405
R2487 VGND.n936 VGND.n935 194.405
R2488 VGND.n941 VGND.n940 194.405
R2489 VGND.n946 VGND.n945 194.405
R2490 VGND.n951 VGND.n950 194.405
R2491 VGND.n956 VGND.n955 194.405
R2492 VGND.n659 VGND.n658 194.405
R2493 VGND.n1946 VGND.n453 194.405
R2494 VGND.n1939 VGND.n1938 194.405
R2495 VGND.n1934 VGND.n1933 194.405
R2496 VGND.n1929 VGND.n1928 194.405
R2497 VGND.n462 VGND.n461 194.405
R2498 VGND.n1898 VGND.n1897 194.405
R2499 VGND.n470 VGND.n469 194.405
R2500 VGND.n1872 VGND.n1871 194.405
R2501 VGND.n478 VGND.n477 194.405
R2502 VGND.n1846 VGND.n1845 194.405
R2503 VGND.n486 VGND.n485 194.405
R2504 VGND.n1820 VGND.n1819 194.405
R2505 VGND.n665 VGND.n664 194.405
R2506 VGND.n1397 VGND.n1396 194.405
R2507 VGND.n1392 VGND.n1391 194.405
R2508 VGND.n668 VGND.n667 194.405
R2509 VGND.n2361 VGND.n303 194.405
R2510 VGND.n2354 VGND.n2353 194.405
R2511 VGND.n1916 VGND.n1915 194.405
R2512 VGND.n458 VGND.n457 194.405
R2513 VGND.n1911 VGND.n1910 194.405
R2514 VGND.n466 VGND.n465 194.405
R2515 VGND.n1885 VGND.n1884 194.405
R2516 VGND.n474 VGND.n473 194.405
R2517 VGND.n1859 VGND.n1858 194.405
R2518 VGND.n482 VGND.n481 194.405
R2519 VGND.n1833 VGND.n1832 194.405
R2520 VGND.n490 VGND.n489 194.405
R2521 VGND.n1807 VGND.n1806 194.405
R2522 VGND.n1374 VGND.n1373 194.405
R2523 VGND.n1377 VGND.n1376 194.405
R2524 VGND.n1371 VGND.n1370 194.405
R2525 VGND.n1779 VGND.n506 194.405
R2526 VGND.n1784 VGND.n1783 194.405
R2527 VGND.n504 VGND.n503 194.405
R2528 VGND.n1314 VGND.n1313 194.405
R2529 VGND.n1319 VGND.n1318 194.405
R2530 VGND.n1324 VGND.n1323 194.405
R2531 VGND.n1329 VGND.n1328 194.405
R2532 VGND.n1334 VGND.n1333 194.405
R2533 VGND.n1339 VGND.n1338 194.405
R2534 VGND.n1344 VGND.n1343 194.405
R2535 VGND.n1349 VGND.n1348 194.405
R2536 VGND.n1354 VGND.n1353 194.405
R2537 VGND.n1359 VGND.n1358 194.405
R2538 VGND.n1306 VGND.n1305 194.405
R2539 VGND.n1309 VGND.n1308 194.405
R2540 VGND.n1303 VGND.n1302 194.405
R2541 VGND.n1772 VGND.n509 194.405
R2542 VGND.n1765 VGND.n1764 194.405
R2543 VGND.n1760 VGND.n1759 194.405
R2544 VGND.n1755 VGND.n1754 194.405
R2545 VGND.n518 VGND.n517 194.405
R2546 VGND.n1724 VGND.n1723 194.405
R2547 VGND.n526 VGND.n525 194.405
R2548 VGND.n1698 VGND.n1697 194.405
R2549 VGND.n534 VGND.n533 194.405
R2550 VGND.n1672 VGND.n1671 194.405
R2551 VGND.n542 VGND.n541 194.405
R2552 VGND.n1646 VGND.n1645 194.405
R2553 VGND.n576 VGND.n575 194.405
R2554 VGND.n1519 VGND.n1518 194.405
R2555 VGND.n1514 VGND.n1513 194.405
R2556 VGND.n572 VGND.n571 194.405
R2557 VGND.n2386 VGND.n290 194.405
R2558 VGND.n2379 VGND.n2378 194.405
R2559 VGND.n1742 VGND.n1741 194.405
R2560 VGND.n514 VGND.n513 194.405
R2561 VGND.n1737 VGND.n1736 194.405
R2562 VGND.n522 VGND.n521 194.405
R2563 VGND.n1711 VGND.n1710 194.405
R2564 VGND.n530 VGND.n529 194.405
R2565 VGND.n1685 VGND.n1684 194.405
R2566 VGND.n538 VGND.n537 194.405
R2567 VGND.n1659 VGND.n1658 194.405
R2568 VGND.n546 VGND.n545 194.405
R2569 VGND.n1633 VGND.n1632 194.405
R2570 VGND.n565 VGND.n564 194.405
R2571 VGND.n1534 VGND.n1533 194.405
R2572 VGND.n568 VGND.n567 194.405
R2573 VGND.n1605 VGND.n1601 194.405
R2574 VGND.n1610 VGND.n1609 194.405
R2575 VGND.n560 VGND.n559 194.405
R2576 VGND.n1597 VGND.n1596 194.405
R2577 VGND.n1592 VGND.n1591 194.405
R2578 VGND.n1587 VGND.n1586 194.405
R2579 VGND.n1582 VGND.n1581 194.405
R2580 VGND.n1577 VGND.n1576 194.405
R2581 VGND.n1572 VGND.n1571 194.405
R2582 VGND.n1567 VGND.n1566 194.405
R2583 VGND.n1562 VGND.n1561 194.405
R2584 VGND.n1557 VGND.n1556 194.405
R2585 VGND.n1552 VGND.n1551 194.405
R2586 VGND.n1547 VGND.n1546 194.405
R2587 VGND.n673 VGND.n672 194.405
R2588 VGND.n671 VGND.n670 194.405
R2589 VGND.n2406 VGND.n278 194.405
R2590 VGND.n2399 VGND.n2398 194.405
R2591 VGND.n842 VGND.n841 194.405
R2592 VGND.n847 VGND.n846 194.405
R2593 VGND.n852 VGND.n851 194.405
R2594 VGND.n857 VGND.n856 194.405
R2595 VGND.n862 VGND.n861 194.405
R2596 VGND.n867 VGND.n866 194.405
R2597 VGND.n872 VGND.n871 194.405
R2598 VGND.n877 VGND.n876 194.405
R2599 VGND.n882 VGND.n881 194.405
R2600 VGND.n887 VGND.n886 194.405
R2601 VGND.n829 VGND.n828 194.405
R2602 VGND.n837 VGND.n836 194.405
R2603 VGND.n832 VGND.n831 194.405
R2604 VGND.n825 VGND.n824 194.405
R2605 VGND.n1231 VGND.n787 194.405
R2606 VGND.n1224 VGND.n1223 194.405
R2607 VGND.n793 VGND.n792 194.405
R2608 VGND.n1205 VGND.n1204 194.405
R2609 VGND.n1199 VGND.n795 194.405
R2610 VGND.n1192 VGND.n1191 194.405
R2611 VGND.n801 VGND.n800 194.405
R2612 VGND.n1173 VGND.n1172 194.405
R2613 VGND.n1167 VGND.n803 194.405
R2614 VGND.n1160 VGND.n1159 194.405
R2615 VGND.n809 VGND.n808 194.405
R2616 VGND.n1141 VGND.n1140 194.405
R2617 VGND.n1135 VGND.n811 194.405
R2618 VGND.n1128 VGND.n1127 194.405
R2619 VGND.n1125 VGND.n813 194.405
R2620 VGND.n815 VGND.n814 194.405
R2621 VGND.n718 VGND.n717 194.405
R2622 VGND.n777 VGND.n776 194.405
R2623 VGND.n772 VGND.n771 194.405
R2624 VGND.n767 VGND.n766 194.405
R2625 VGND.n762 VGND.n761 194.405
R2626 VGND.n757 VGND.n756 194.405
R2627 VGND.n752 VGND.n751 194.405
R2628 VGND.n747 VGND.n746 194.405
R2629 VGND.n742 VGND.n741 194.405
R2630 VGND.n737 VGND.n736 194.405
R2631 VGND.n732 VGND.n731 194.405
R2632 VGND.n727 VGND.n726 194.405
R2633 VGND.n722 VGND.n721 194.405
R2634 VGND.n684 VGND.n682 194.405
R2635 VGND.n1286 VGND.n678 194.405
R2636 VGND.n676 VGND.n675 194.405
R2637 VGND.t1187 VGND.t861 179.154
R2638 VGND.t798 VGND.t1114 179.154
R2639 VGND.t787 VGND.t1098 179.154
R2640 VGND.t2637 VGND.t768 179.154
R2641 VGND.t1535 VGND.t1308 179.154
R2642 VGND.t1964 VGND.t1519 179.154
R2643 VGND.t757 VGND.t2411 179.154
R2644 VGND.t2345 VGND.t844 179.154
R2645 VGND.t834 VGND.t590 179.154
R2646 VGND.t1714 VGND.t772 179.154
R2647 VGND.t907 VGND.t1516 179.154
R2648 VGND.t2243 VGND.t1577 179.154
R2649 VGND.t829 VGND.t1659 179.154
R2650 VGND.t296 VGND.t819 179.154
R2651 VGND.t882 VGND.t1063 179.154
R2652 VGND.t1569 VGND.t917 179.154
R2653 VGND.t38 VGND.t378 179.154
R2654 VGND.t1961 VGND.t602 179.154
R2655 VGND.t2340 VGND.t454 179.154
R2656 VGND.t1509 VGND.t922 179.154
R2657 VGND.t95 VGND.t1503 179.154
R2658 VGND.t1242 VGND.t310 179.154
R2659 VGND.t1116 VGND.t2242 179.154
R2660 VGND.t244 VGND.t1971 179.154
R2661 VGND.t443 VGND.t1297 179.154
R2662 VGND.t345 VGND.t1146 179.154
R2663 VGND.t2229 VGND.t89 179.154
R2664 VGND.t1113 VGND.t736 179.154
R2665 VGND.t1185 VGND.t2218 179.154
R2666 VGND.t286 VGND.t1040 179.154
R2667 VGND.t1653 VGND.t531 179.154
R2668 VGND.t836 VGND.t1718 179.154
R2669 VGND.t295 VGND.t1034 179.154
R2670 VGND.t1941 VGND.t2236 179.154
R2671 VGND.t20 VGND.t1062 179.154
R2672 VGND.t1324 VGND.t2035 179.154
R2673 VGND.t1717 VGND.t2076 179.154
R2674 VGND.t73 VGND.t2061 179.154
R2675 VGND.t2342 VGND.t2026 179.154
R2676 VGND.t1099 VGND.t2662 179.154
R2677 VGND.t2635 VGND.t2641 179.154
R2678 VGND.t1112 VGND.t364 179.154
R2679 VGND.t188 VGND.t117 179.154
R2680 VGND.t2408 VGND.t743 179.154
R2681 VGND.t2248 VGND.t1208 179.154
R2682 VGND.t173 VGND.t1478 179.154
R2683 VGND.t123 VGND.t544 179.154
R2684 VGND.t18 VGND.t2588 179.154
R2685 VGND.t1101 VGND.t297 179.154
R2686 VGND.t551 VGND.t2350 179.154
R2687 VGND.t35 VGND.t1615 179.154
R2688 VGND.t1144 VGND.t1037 179.154
R2689 VGND.t534 VGND.t2365 179.154
R2690 VGND.t2134 VGND.t1652 179.154
R2691 VGND.t1061 VGND.t519 179.154
R2692 VGND.t687 VGND.t2009 179.154
R2693 VGND.t1820 VGND.t278 179.154
R2694 VGND.t403 VGND.t245 179.154
R2695 VGND.t1715 VGND.t126 179.154
R2696 VGND.t1202 VGND.t232 179.154
R2697 VGND.t2664 VGND.t1950 179.154
R2698 VGND.t1469 VGND.t1043 179.154
R2699 VGND.t2528 VGND.t661 179.154
R2700 VGND.t758 VGND.t1640 179.154
R2701 VGND.t246 VGND.t2647 179.154
R2702 VGND.t2011 VGND.t2092 179.154
R2703 VGND.t43 VGND.t1067 179.154
R2704 VGND.t1967 VGND.t144 179.154
R2705 VGND.t1746 VGND.t1186 179.154
R2706 VGND.t1274 VGND.t242 179.154
R2707 VGND.t2239 VGND.t228 179.154
R2708 VGND.t86 VGND.t669 179.154
R2709 VGND.t2677 VGND.t36 179.154
R2710 VGND.t1490 VGND.t223 179.154
R2711 VGND.t97 VGND.t1513 179.154
R2712 VGND.t522 VGND.t2055 179.154
R2713 VGND.t196 VGND.t1814 179.154
R2714 VGND.t2039 VGND.t1620 179.154
R2715 VGND.t1325 VGND.t528 179.154
R2716 VGND.t1543 VGND.t1041 179.154
R2717 VGND.t247 VGND.t1028 179.154
R2718 VGND.t2231 VGND.t1935 179.154
R2719 VGND.t27 VGND.t533 179.154
R2720 VGND.t730 VGND.t1053 179.154
R2721 VGND.t2070 VGND.t2339 179.154
R2722 VGND.t2605 VGND.t2658 179.154
R2723 VGND.t1200 VGND.t2682 179.154
R2724 VGND.t1918 VGND.t702 179.154
R2725 VGND.t432 VGND.t1817 179.154
R2726 VGND.t358 VGND.t2228 179.154
R2727 VGND.t113 VGND.t142 179.154
R2728 VGND.t292 VGND.t607 179.154
R2729 VGND.t1756 VGND.t1791 179.154
R2730 VGND.t1472 VGND.t1211 179.154
R2731 VGND.t540 VGND.t1470 179.154
R2732 VGND.t804 VGND.t2412 179.154
R2733 VGND.t377 VGND.t1326 179.154
R2734 VGND.t1804 VGND.t1960 179.154
R2735 VGND.t2234 VGND.t451 179.154
R2736 VGND.t921 VGND.t96 179.154
R2737 VGND.t1642 VGND.t1502 179.154
R2738 VGND.t45 VGND.t143 179.154
R2739 VGND.t916 VGND.t2241 179.154
R2740 VGND.t1968 VGND.t2056 179.154
R2741 VGND.t2646 VGND.t2679 179.154
R2742 VGND.t344 VGND.t1066 179.154
R2743 VGND.t1902 VGND.t99 179.154
R2744 VGND.t735 VGND.t1637 179.154
R2745 VGND.t1934 VGND.t2215 179.154
R2746 VGND.t1115 VGND.t1039 179.154
R2747 VGND.t229 VGND.t530 179.154
R2748 VGND.t835 VGND.t1912 179.154
R2749 VGND.t550 VGND.t1102 179.154
R2750 VGND.t1047 VGND.t2351 179.154
R2751 VGND.t1616 VGND.t74 179.154
R2752 VGND.t1909 VGND.t1145 179.154
R2753 VGND.t2199 VGND.t1486 179.154
R2754 VGND.t2022 VGND.t2598 179.154
R2755 VGND.t520 VGND.t211 179.154
R2756 VGND.t384 VGND.t688 179.154
R2757 VGND.t279 VGND.t1309 179.154
R2758 VGND.t712 VGND.t404 179.154
R2759 VGND.t127 VGND.t2406 179.154
R2760 VGND.t1150 VGND.t1203 179.154
R2761 VGND.t1951 VGND.t2343 179.154
R2762 VGND.t1044 VGND.t914 179.154
R2763 VGND.t2410 VGND.t662 179.154
R2764 VGND.t769 VGND.t1174 179.154
R2765 VGND.t380 VGND.t1111 179.154
R2766 VGND.t1948 VGND.t2344 179.154
R2767 VGND.t2671 VGND.t129 179.154
R2768 VGND.t1629 VGND.t1813 179.154
R2769 VGND.t2407 VGND.t1802 179.154
R2770 VGND.t316 VGND.t608 179.154
R2771 VGND.t723 VGND.t1812 179.154
R2772 VGND.t1975 VGND.t1512 179.154
R2773 VGND.t1303 VGND.t75 179.154
R2774 VGND.t1148 VGND.t1212 179.154
R2775 VGND.t83 VGND.t383 179.154
R2776 VGND.t2045 VGND.t2233 179.154
R2777 VGND.t1852 VGND.t2525 179.154
R2778 VGND.t2040 VGND.t1194 179.154
R2779 VGND.t1894 VGND.t1311 179.154
R2780 VGND.t850 VGND.t1050 179.154
R2781 VGND.t1882 VGND.t1097 179.154
R2782 VGND.t2663 VGND.t2091 179.154
R2783 VGND.t701 VGND.t42 179.154
R2784 VGND.t1636 VGND.t1138 179.154
R2785 VGND.t1489 VGND.t1745 179.154
R2786 VGND.t241 VGND.t2006 179.154
R2787 VGND.t1510 VGND.t305 179.154
R2788 VGND.t668 VGND.t1901 179.154
R2789 VGND.t2230 VGND.t2676 179.154
R2790 VGND.t222 VGND.t2246 179.154
R2791 VGND.t2008 VGND.t104 179.154
R2792 VGND.t2054 VGND.t1815 179.154
R2793 VGND.t287 VGND.t195 179.154
R2794 VGND.t76 VGND.t2038 179.154
R2795 VGND.t1173 VGND.t525 179.154
R2796 VGND.t1536 VGND.t2007 179.154
R2797 VGND.t1897 VGND.t1027 179.154
R2798 VGND.t2558 VGND.t2125 179.154
R2799 VGND.t1624 VGND.t1903 179.154
R2800 VGND.t1245 VGND.t729 179.154
R2801 VGND.t2205 VGND.t1065 179.154
R2802 VGND.t288 VGND.t2604 179.154
R2803 VGND.t1197 VGND.t918 179.154
R2804 VGND.t128 VGND.t1917 179.154
R2805 VGND.t431 VGND.t240 179.154
R2806 VGND.t1109 VGND.t414 179.154
R2807 VGND.t112 VGND.t707 179.154
R2808 VGND.t149 VGND.t291 179.154
R2809 VGND.t1755 VGND.t212 179.154
R2810 VGND.t1241 VGND.t1790 179.154
R2811 VGND.t1177 VGND.t537 179.154
R2812 VGND.t799 VGND.t174 179.154
R2813 VGND.t1816 VGND.t1033 179.154
R2814 VGND.t1119 VGND.t1940 179.154
R2815 VGND.t19 VGND.t2681 179.154
R2816 VGND.t2034 VGND.t698 179.154
R2817 VGND.t2075 VGND.t1911 179.154
R2818 VGND.t2060 VGND.t1048 179.154
R2819 VGND.t2025 VGND.t2636 179.154
R2820 VGND.t2661 VGND.t2005 179.154
R2821 VGND.t2640 VGND.t1805 179.154
R2822 VGND.t363 VGND.t1881 179.154
R2823 VGND.t116 VGND.t1654 179.154
R2824 VGND.t742 VGND.t1898 179.154
R2825 VGND.t1761 VGND.t1965 179.154
R2826 VGND.t1477 VGND.t1883 179.154
R2827 VGND.t543 VGND.t699 179.154
R2828 VGND.t828 VGND.t1488 179.154
R2829 VGND.t1511 VGND.t1100 179.154
R2830 VGND.t285 VGND.t2349 179.154
R2831 VGND.t105 VGND.t1614 179.154
R2832 VGND.t1143 VGND.t594 179.154
R2833 VGND.t1120 VGND.t2364 179.154
R2834 VGND.t2133 VGND.t915 179.154
R2835 VGND.t2247 VGND.t187 179.154
R2836 VGND.t686 VGND.t732 179.154
R2837 VGND.t164 VGND.t277 179.154
R2838 VGND.t402 VGND.t1641 179.154
R2839 VGND.t2232 VGND.t125 179.154
R2840 VGND.t1201 VGND.t183 179.154
R2841 VGND.t189 VGND.t1949 179.154
R2842 VGND.t2639 VGND.t1042 179.154
R2843 VGND.t1192 VGND.t658 179.154
R2844 VGND.t909 VGND.t970 179.154
R2845 VGND.t2648 VGND.t1884 179.154
R2846 VGND.t1904 VGND.t1955 179.154
R2847 VGND.t44 VGND.t2338 179.154
R2848 VGND.t1108 VGND.t145 179.154
R2849 VGND.t1056 VGND.t605 179.154
R2850 VGND.t233 VGND.t243 179.154
R2851 VGND.t2240 VGND.t1049 179.154
R2852 VGND.t2057 VGND.t672 179.154
R2853 VGND.t2678 VGND.t1806 179.154
R2854 VGND.t62 VGND.t335 179.154
R2855 VGND.t98 VGND.t1655 179.154
R2856 VGND.t63 VGND.t482 179.154
R2857 VGND.t199 VGND.t2021 179.154
R2858 VGND.t1151 VGND.t603 179.154
R2859 VGND.t1619 VGND.t529 179.154
R2860 VGND.t1564 VGND.t2587 179.154
R2861 VGND.t2010 VGND.t1485 179.154
R2862 VGND.t209 VGND.t148 179.154
R2863 VGND.t2529 VGND.t72 179.154
R2864 VGND.t2409 VGND.t1142 179.154
R2865 VGND.t477 VGND.t2363 179.154
R2866 VGND.t230 VGND.t2132 179.154
R2867 VGND.t1793 VGND.t184 179.154
R2868 VGND.t200 VGND.t685 179.154
R2869 VGND.t591 VGND.t276 179.154
R2870 VGND.t444 VGND.t401 179.154
R2871 VGND.t1908 VGND.t124 179.154
R2872 VGND.t2341 VGND.t2227 179.154
R2873 VGND.t1792 VGND.t2214 179.154
R2874 VGND.t1172 VGND.t302 179.154
R2875 VGND.t655 VGND.t2638 179.154
R2876 VGND.t908 VGND.t1501 179.154
R2877 VGND.t239 VGND.t379 179.154
R2878 VGND.t593 VGND.t2348 179.154
R2879 VGND.t2004 VGND.t455 179.154
R2880 VGND.t1628 VGND.t1243 179.154
R2881 VGND.t1508 VGND.t39 179.154
R2882 VGND.t315 VGND.t1803 179.154
R2883 VGND.t1180 VGND.t1110 179.154
R2884 VGND.t1974 VGND.t1117 179.154
R2885 VGND.t1302 VGND.t1910 179.154
R2886 VGND.t1147 VGND.t750 179.154
R2887 VGND.t94 VGND.t1807 179.154
R2888 VGND.t737 VGND.t1213 179.154
R2889 VGND.t1851 VGND.t1468 179.154
R2890 VGND.t2257 VGND.t1638 179.154
R2891 VGND.t2683 VGND.t1887 179.154
R2892 VGND.t845 VGND.t1038 179.154
R2893 VGND.t1107 VGND.t1207 179.154
R2894 VGND.t1137 VGND.t2352 179.154
R2895 VGND.t293 VGND.t1621 179.154
R2896 VGND.t37 VGND.t931 179.154
R2897 VGND.t1052 VGND.t2200 179.154
R2898 VGND.t1064 VGND.t2599 179.154
R2899 VGND.t41 VGND.t521 179.154
R2900 VGND.t700 VGND.t689 179.154
R2901 VGND.t0 VGND.t280 179.154
R2902 VGND.t1625 VGND.t411 179.154
R2903 VGND.t1471 VGND.t118 179.154
R2904 VGND.t40 VGND.t1206 179.154
R2905 VGND.t1193 VGND.t1952 179.154
R2906 VGND.t1639 VGND.t1238 179.154
R2907 VGND.t1933 VGND.t549 179.154
R2908 VGND.t781 VGND.t1149 179.154
R2909 VGND.n2564 VGND.n2563 161.303
R2910 VGND.n2561 VGND.n2560 161.303
R2911 VGND.n2558 VGND.n2557 161.303
R2912 VGND.n2555 VGND.n2554 161.303
R2913 VGND.n2552 VGND.n2551 161.303
R2914 VGND.n2549 VGND.n2548 161.303
R2915 VGND.n2546 VGND.n2545 161.303
R2916 VGND.n2543 VGND.n2542 161.303
R2917 VGND.n2540 VGND.n2539 161.303
R2918 VGND.n2537 VGND.n2536 161.303
R2919 VGND.n2534 VGND.n2533 161.303
R2920 VGND.n2531 VGND.n2530 161.303
R2921 VGND.n2528 VGND.n2527 161.303
R2922 VGND.n2525 VGND.n2524 161.303
R2923 VGND.n2522 VGND.n2521 161.303
R2924 VGND.n2563 VGND.t2692 161.106
R2925 VGND.n2560 VGND.t2695 161.106
R2926 VGND.n2557 VGND.t2690 161.106
R2927 VGND.n2554 VGND.t2702 161.106
R2928 VGND.n2551 VGND.t2691 161.106
R2929 VGND.n2548 VGND.t2699 161.106
R2930 VGND.n2545 VGND.t2694 161.106
R2931 VGND.n2542 VGND.t2688 161.106
R2932 VGND.n2539 VGND.t2701 161.106
R2933 VGND.n2536 VGND.t2703 161.106
R2934 VGND.n2533 VGND.t2698 161.106
R2935 VGND.n2530 VGND.t2689 161.106
R2936 VGND.n2527 VGND.t2696 161.106
R2937 VGND.n2524 VGND.t2693 161.106
R2938 VGND.n2521 VGND.t2700 161.106
R2939 VGND.n996 VGND.t227 159.315
R2940 VGND.n2902 VGND.t711 159.315
R2941 VGND.n1088 VGND.t2245 158.361
R2942 VGND.n2972 VGND.t1907 158.361
R2943 VGND.n898 VGND.t225 157.291
R2944 VGND.n2900 VGND.t709 157.291
R2945 VGND.n582 VGND.t1801 156.915
R2946 VGND.n2862 VGND.t1217 156.915
R2947 VGND.n582 VGND.t1799 156.915
R2948 VGND.n2862 VGND.t1218 156.915
R2949 VGND.n2563 VGND.t1390 154.679
R2950 VGND.n2560 VGND.t1435 154.679
R2951 VGND.n2557 VGND.t1342 154.679
R2952 VGND.n2554 VGND.t1420 154.679
R2953 VGND.n2551 VGND.t1459 154.679
R2954 VGND.n2548 VGND.t1396 154.679
R2955 VGND.n2545 VGND.t1339 154.679
R2956 VGND.n2542 VGND.t1378 154.679
R2957 VGND.n2539 VGND.t1423 154.679
R2958 VGND.n2536 VGND.t1465 154.679
R2959 VGND.n2533 VGND.t1438 154.679
R2960 VGND.n2530 VGND.t1345 154.679
R2961 VGND.n2527 VGND.t1411 154.679
R2962 VGND.n2524 VGND.t1348 154.679
R2963 VGND.n2521 VGND.t1384 154.679
R2964 VGND.n584 VGND.t210 154.131
R2965 VGND.n584 VGND.t532 154.131
R2966 VGND.n996 VGND.t2527 154.131
R2967 VGND.n999 VGND.t606 154.131
R2968 VGND.n2886 VGND.t731 154.131
R2969 VGND.n2886 VGND.t34 154.131
R2970 VGND.n2902 VGND.t2033 154.131
R2971 VGND.n2932 VGND.t1658 154.131
R2972 VGND.n118 VGND.t1798 153.631
R2973 VGND.n1026 VGND.t294 153.631
R2974 VGND.n1057 VGND.t726 153.631
R2975 VGND.n2854 VGND.t1215 153.631
R2976 VGND.n2934 VGND.t461 153.631
R2977 VGND.n2939 VGND.t1176 153.631
R2978 VGND.n1027 VGND.t592 152.757
R2979 VGND.n2935 VGND.t309 152.757
R2980 VGND.n991 VGND.t1796 152.381
R2981 VGND.n61 VGND.t1222 152.381
R2982 VGND.n961 VGND.n960 152.174
R2983 VGND.n149 VGND.t1800 150.922
R2984 VGND.n149 VGND.t1794 150.922
R2985 VGND.n86 VGND.t1225 150.922
R2986 VGND.n86 VGND.t1220 150.922
R2987 VGND.n116 VGND.t2012 150.922
R2988 VGND.n581 VGND.t1682 150.922
R2989 VGND.n148 VGND.t238 150.922
R2990 VGND.n85 VGND.t2249 150.922
R2991 VGND.n2829 VGND.t717 150.922
R2992 VGND.n2861 VGND.t2666 150.922
R2993 VGND.n116 VGND.t1051 150.922
R2994 VGND.n581 VGND.t478 150.922
R2995 VGND.n148 VGND.t2657 150.922
R2996 VGND.n85 VGND.t457 150.922
R2997 VGND.n2829 VGND.t430 150.922
R2998 VGND.n2861 VGND.t1315 150.922
R2999 VGND.n117 VGND.t1797 147.411
R3000 VGND.n1058 VGND.t1643 147.411
R3001 VGND.n2853 VGND.t1224 147.411
R3002 VGND.n2940 VGND.t1819 147.411
R3003 VGND.n899 VGND.t59 146.964
R3004 VGND.n84 VGND.t133 146.964
R3005 VGND.n1512 VGND.n578 143.478
R3006 VGND VGND.t2496 142.089
R3007 VGND.t761 VGND.t1382 126.853
R3008 VGND.t1331 VGND.t1524 126.853
R3009 VGND.t2595 VGND.t1337 126.853
R3010 VGND.t1358 VGND.t822 126.853
R3011 VGND.t841 VGND.t1430 126.853
R3012 VGND.t1442 VGND.t1570 126.853
R3013 VGND.t812 VGND.t1361 126.853
R3014 VGND.t1394 VGND.t901 126.853
R3015 VGND.t887 VGND.t1406 126.853
R3016 VGND.t1451 VGND.t1556 126.853
R3017 VGND.t802 VGND.t1367 126.853
R3018 VGND.t1409 VGND.t875 126.853
R3019 VGND.t1547 VGND.t1454 126.853
R3020 VGND.t1463 VGND.t1544 126.853
R3021 VGND.t779 VGND.t1373 126.853
R3022 VGND.t1418 VGND.t866 126.853
R3023 VGND.n822 VGND.t1381 119.309
R3024 VGND.n785 VGND.t1417 119.309
R3025 VGND.n2579 VGND.t1414 119.309
R3026 VGND.n2576 VGND.t1375 119.309
R3027 VGND.n2581 VGND.t1369 119.309
R3028 VGND.n2584 VGND.t1456 119.309
R3029 VGND.n2587 VGND.t1447 119.309
R3030 VGND.n2590 VGND.t1402 119.309
R3031 VGND.n2593 VGND.t1363 119.309
R3032 VGND.n2596 VGND.t1444 119.309
R3033 VGND.n2599 VGND.t1399 119.309
R3034 VGND.n2602 VGND.t1387 119.309
R3035 VGND.n2605 VGND.t1354 119.309
R3036 VGND.n2608 VGND.t1432 119.309
R3037 VGND.n2611 VGND.t1426 119.309
R3038 VGND.n2614 VGND.t1351 119.309
R3039 VGND.n2575 VGND.t1333 119.309
R3040 VGND.n2568 VGND.t1327 119.309
R3041 VGND.n819 VGND.t1330 119.309
R3042 VGND.n816 VGND.t1336 119.309
R3043 VGND.n1136 VGND.t1357 119.309
R3044 VGND.n807 VGND.t1429 119.309
R3045 VGND.n805 VGND.t1441 119.309
R3046 VGND.n1151 VGND.t1360 119.309
R3047 VGND.n1168 VGND.t1393 119.309
R3048 VGND.n799 VGND.t1405 119.309
R3049 VGND.n797 VGND.t1450 119.309
R3050 VGND.n1183 VGND.t1366 119.309
R3051 VGND.n1200 VGND.t1408 119.309
R3052 VGND.n791 VGND.t1453 119.309
R3053 VGND.n789 VGND.t1462 119.309
R3054 VGND.n1215 VGND.t1372 119.309
R3055 VGND.n6 VGND.n4 117.001
R3056 VGND.t1604 VGND.n6 117.001
R3057 VGND.n5 VGND.n3 117.001
R3058 VGND.t1604 VGND.n5 117.001
R3059 VGND.t50 VGND.t60 92.9349
R3060 VGND.t60 VGND.t57 92.9349
R3061 VGND.t57 VGND.t61 92.9349
R3062 VGND.t61 VGND.t254 92.9349
R3063 VGND.t254 VGND.t266 92.9349
R3064 VGND.t266 VGND.t2372 92.9349
R3065 VGND.t2372 VGND.t2312 92.9349
R3066 VGND.t595 VGND.t763 90.6101
R3067 VGND.t1526 VGND.t1244 90.6101
R3068 VGND.t1966 VGND.t2597 90.6101
R3069 VGND.t824 VGND.t713 90.6101
R3070 VGND.t1514 VGND.t843 90.6101
R3071 VGND.t1572 VGND.t1 90.6101
R3072 VGND.t1716 VGND.t814 90.6101
R3073 VGND.t890 VGND.t1515 90.6101
R3074 VGND.t1310 VGND.t889 90.6101
R3075 VGND.t825 VGND.t663 90.6101
R3076 VGND.t1118 VGND.t805 90.6101
R3077 VGND.t877 VGND.t1487 90.6101
R3078 VGND.t231 VGND.t1549 90.6101
R3079 VGND.t1546 VGND.t213 90.6101
R3080 VGND.t2235 VGND.t782 90.6101
R3081 VGND.t868 VGND.t604 90.6101
R3082 VGND VGND.n578 80.9529
R3083 VGND.n1291 VGND 75.2331
R3084 VGND VGND.n578 75.1009
R3085 VGND.t2312 VGND 70.8076
R3086 VGND.n147 VGND 58.8055
R3087 VGND.n1506 VGND 58.8055
R3088 VGND.n1508 VGND 58.8055
R3089 VGND.n1510 VGND 58.8055
R3090 VGND.n2818 VGND 58.8055
R3091 VGND.n2821 VGND.n2820 53.1823
R3092 VGND.n2822 VGND.n2821 53.1823
R3093 VGND.n3004 VGND.n3003 53.1823
R3094 VGND.n3003 VGND.n3002 53.1823
R3095 VGND.t58 VGND.t252 50.5752
R3096 VGND.t55 VGND.t264 50.5752
R3097 VGND.t53 VGND.t2510 50.5752
R3098 VGND.t51 VGND.t6 50.5752
R3099 VGND.t140 VGND.t2494 50.5752
R3100 VGND.t136 VGND.t2468 50.5752
R3101 VGND.t130 VGND.t2505 50.5752
R3102 VGND.t132 VGND.t2455 50.5752
R3103 VGND VGND.n14 43.2063
R3104 VGND VGND.n43 43.2063
R3105 VGND VGND.n2916 43.2063
R3106 VGND VGND.n2956 43.2063
R3107 VGND.n2820 VGND.n2819 40.6593
R3108 VGND.n2572 VGND.t858 36.0005
R3109 VGND.n2572 VGND.t860 36.0005
R3110 VGND.n2641 VGND.t1566 36.0005
R3111 VGND.n2641 VGND.t1568 36.0005
R3112 VGND.n2639 VGND.t879 36.0005
R3113 VGND.n2639 VGND.t881 36.0005
R3114 VGND.n2648 VGND.t816 36.0005
R3115 VGND.n2648 VGND.t818 36.0005
R3116 VGND.n2636 VGND.t1559 36.0005
R3117 VGND.n2636 VGND.t827 36.0005
R3118 VGND.n2655 VGND.t1574 36.0005
R3119 VGND.n2655 VGND.t1576 36.0005
R3120 VGND.n2633 VGND.t904 36.0005
R3121 VGND.n2633 VGND.t906 36.0005
R3122 VGND.n2662 VGND.t831 36.0005
R3123 VGND.n2662 VGND.t833 36.0005
R3124 VGND.n2630 VGND.t1587 36.0005
R3125 VGND.n2630 VGND.t1589 36.0005
R3126 VGND.n2669 VGND.t847 36.0005
R3127 VGND.n2669 VGND.t849 36.0005
R3128 VGND.n2627 VGND.t911 36.0005
R3129 VGND.n2627 VGND.t913 36.0005
R3130 VGND.n2676 VGND.t1530 36.0005
R3131 VGND.n2676 VGND.t1518 36.0005
R3132 VGND.n2624 VGND.t1532 36.0005
R3133 VGND.n2624 VGND.t1534 36.0005
R3134 VGND.n2683 VGND.t765 36.0005
R3135 VGND.n2683 VGND.t767 36.0005
R3136 VGND.n2620 VGND.t784 36.0005
R3137 VGND.n2620 VGND.t786 36.0005
R3138 VGND.n2571 VGND.t1528 36.0005
R3139 VGND.n2571 VGND.t797 36.0005
R3140 VGND.n225 VGND.t548 36.0005
R3141 VGND.n225 VGND.t2303 36.0005
R3142 VGND.n2760 VGND.t1476 36.0005
R3143 VGND.n2760 VGND.t1086 36.0005
R3144 VGND.n2755 VGND.t1811 36.0005
R3145 VGND.n2755 VGND.t1124 36.0005
R3146 VGND.n2750 VGND.t486 36.0005
R3147 VGND.n2750 VGND.t1679 36.0005
R3148 VGND.n2745 VGND.t109 36.0005
R3149 VGND.n2745 VGND.t2305 36.0005
R3150 VGND.n2740 VGND.t339 36.0005
R3151 VGND.n2740 VGND.t1088 36.0005
R3152 VGND.n2735 VGND.t2645 36.0005
R3153 VGND.n2735 VGND.t1681 36.0005
R3154 VGND.n2730 VGND.t676 36.0005
R3155 VGND.n2730 VGND.t2307 36.0005
R3156 VGND.n2725 VGND.t2030 36.0005
R3157 VGND.n2725 VGND.t2309 36.0005
R3158 VGND.n2720 VGND.t2065 36.0005
R3159 VGND.n2720 VGND.t1090 36.0005
R3160 VGND.n2715 VGND.t1060 36.0005
R3161 VGND.n2715 VGND.t2299 36.0005
R3162 VGND.n2710 VGND.t930 36.0005
R3163 VGND.n2710 VGND.t2301 36.0005
R3164 VGND.n2705 VGND.t1071 36.0005
R3165 VGND.n2705 VGND.t1092 36.0005
R3166 VGND.n2700 VGND.t1959 36.0005
R3167 VGND.n2700 VGND.t1094 36.0005
R3168 VGND.n230 VGND.t1032 36.0005
R3169 VGND.n230 VGND.t1122 36.0005
R3170 VGND.n228 VGND.t1392 36.0005
R3171 VGND.n228 VGND.t1084 36.0005
R3172 VGND.n2484 VGND.t660 36.0005
R3173 VGND.n2484 VGND.t2620 36.0005
R3174 VGND.n2479 VGND.t1171 36.0005
R3175 VGND.n2479 VGND.t941 36.0005
R3176 VGND.n2474 VGND.t1760 36.0005
R3177 VGND.n2474 VGND.t620 36.0005
R3178 VGND.n2469 VGND.t741 36.0005
R3179 VGND.n2469 VGND.t622 36.0005
R3180 VGND.n2464 VGND.t82 36.0005
R3181 VGND.n2464 VGND.t2622 36.0005
R3182 VGND.n2459 VGND.t362 36.0005
R3183 VGND.n2459 VGND.t610 36.0005
R3184 VGND.n2454 VGND.t275 36.0005
R3185 VGND.n2454 VGND.t624 36.0005
R3186 VGND.n2449 VGND.t2660 36.0005
R3187 VGND.n2449 VGND.t935 36.0005
R3188 VGND.n2444 VGND.t518 36.0005
R3189 VGND.n2444 VGND.t937 36.0005
R3190 VGND.n2439 VGND.t2131 36.0005
R3191 VGND.n2439 VGND.t612 36.0005
R3192 VGND.n2434 VGND.t2074 36.0005
R3193 VGND.n2434 VGND.t2616 36.0005
R3194 VGND.n245 VGND.t926 36.0005
R3195 VGND.n245 VGND.t2618 36.0005
R3196 VGND.n243 VGND.t31 36.0005
R3197 VGND.n243 VGND.t614 36.0005
R3198 VGND.n2509 VGND.t1939 36.0005
R3199 VGND.n2509 VGND.t616 36.0005
R3200 VGND.n240 VGND.t1484 36.0005
R3201 VGND.n240 VGND.t618 36.0005
R3202 VGND.n238 VGND.t1437 36.0005
R3203 VGND.n238 VGND.t939 36.0005
R3204 VGND.n330 VGND.t1891 36.0005
R3205 VGND.n330 VGND.t1280 36.0005
R3206 VGND.n2286 VGND.t1157 36.0005
R3207 VGND.n2286 VGND.t1290 36.0005
R3208 VGND.n2281 VGND.t2211 36.0005
R3209 VGND.n2281 VGND.t1128 36.0005
R3210 VGND.n2276 VGND.t2224 36.0005
R3211 VGND.n2276 VGND.t1130 36.0005
R3212 VGND.n338 VGND.t91 36.0005
R3213 VGND.n338 VGND.t1282 36.0005
R3214 VGND.n2245 VGND.t398 36.0005
R3215 VGND.n2245 VGND.t166 36.0005
R3216 VGND.n346 VGND.t1299 36.0005
R3217 VGND.n346 VGND.t1132 36.0005
R3218 VGND.n2219 VGND.t682 36.0005
R3219 VGND.n2219 VGND.t1284 36.0005
R3220 VGND.n354 VGND.t1184 36.0005
R3221 VGND.n354 VGND.t1286 36.0005
R3222 VGND.n2193 VGND.t312 36.0005
R3223 VGND.n2193 VGND.t168 36.0005
R3224 VGND.n362 VGND.t2360 36.0005
R3225 VGND.n362 VGND.t1134 36.0005
R3226 VGND.n2167 VGND.t1633 36.0005
R3227 VGND.n2167 VGND.t1136 36.0005
R3228 VGND.n368 VGND.t69 36.0005
R3229 VGND.n368 VGND.t170 36.0005
R3230 VGND.n365 VGND.t206 36.0005
R3231 VGND.n365 VGND.t172 36.0005
R3232 VGND.n181 VGND.t2654 36.0005
R3233 VGND.n181 VGND.t1126 36.0005
R3234 VGND.n178 VGND.t1344 36.0005
R3235 VGND.n178 VGND.t1288 36.0005
R3236 VGND.n326 VGND.t539 36.0005
R3237 VGND.n326 VGND.t2670 36.0005
R3238 VGND.n2303 VGND.t1237 36.0005
R3239 VGND.n2303 VGND.t448 36.0005
R3240 VGND.n2263 VGND.t194 36.0005
R3241 VGND.n2263 VGND.t2609 36.0005
R3242 VGND.n334 VGND.t301 36.0005
R3243 VGND.n334 VGND.t2611 36.0005
R3244 VGND.n2258 VGND.t122 36.0005
R3245 VGND.n2258 VGND.t463 36.0005
R3246 VGND.n342 VGND.t219 36.0005
R3247 VGND.n342 VGND.t450 36.0005
R3248 VGND.n2232 VGND.t284 36.0005
R3249 VGND.n2232 VGND.t2613 36.0005
R3250 VGND.n350 VGND.t667 36.0005
R3251 VGND.n350 VGND.t465 36.0005
R3252 VGND.n2206 VGND.t1199 36.0005
R3253 VGND.n2206 VGND.t467 36.0005
R3254 VGND.n358 VGND.t2603 36.0005
R3255 VGND.n358 VGND.t1943 36.0005
R3256 VGND.n2180 VGND.t2198 36.0005
R3257 VGND.n2180 VGND.t249 36.0005
R3258 VGND.n377 VGND.t2687 36.0005
R3259 VGND.n377 VGND.t251 36.0005
R3260 VGND.n2154 VGND.t24 36.0005
R3261 VGND.n2154 VGND.t1945 36.0005
R3262 VGND.n1421 VGND.t2090 36.0005
R3263 VGND.n1421 VGND.t1947 36.0005
R3264 VGND.n1424 VGND.t1106 36.0005
R3265 VGND.n1424 VGND.t2607 36.0005
R3266 VGND.n1418 VGND.t1422 36.0005
R3267 VGND.n1418 VGND.t446 36.0005
R3268 VGND.n394 VGND.t654 36.0005
R3269 VGND.n394 VGND.t428 36.0005
R3270 VGND.n2131 VGND.t2044 36.0005
R3271 VGND.n2131 VGND.t368 36.0005
R3272 VGND.n391 VGND.t1754 36.0005
R3273 VGND.n391 VGND.t418 36.0005
R3274 VGND.n1443 VGND.t290 36.0005
R3275 VGND.n1443 VGND.t420 36.0005
R3276 VGND.n1448 VGND.t78 36.0005
R3277 VGND.n1448 VGND.t388 36.0005
R3278 VGND.n1453 VGND.t413 36.0005
R3279 VGND.n1453 VGND.t370 36.0005
R3280 VGND.n1458 VGND.t1307 36.0005
R3281 VGND.n1458 VGND.t422 36.0005
R3282 VGND.n1463 VGND.t1916 36.0005
R3283 VGND.n1463 VGND.t390 36.0005
R3284 VGND.n1468 VGND.t1900 36.0005
R3285 VGND.n1468 VGND.t392 36.0005
R3286 VGND.n1473 VGND.t2127 36.0005
R3287 VGND.n1473 VGND.t372 36.0005
R3288 VGND.n1478 VGND.t2204 36.0005
R3289 VGND.n1478 VGND.t424 36.0005
R3290 VGND.n1483 VGND.t920 36.0005
R3291 VGND.n1483 VGND.t426 36.0005
R3292 VGND.n1488 VGND.t1623 36.0005
R3293 VGND.n1488 VGND.t374 36.0005
R3294 VGND.n632 VGND.t2124 36.0005
R3295 VGND.n632 VGND.t376 36.0005
R3296 VGND.n1438 VGND.t1480 36.0005
R3297 VGND.n1438 VGND.t416 36.0005
R3298 VGND.n636 VGND.t1461 36.0005
R3299 VGND.n636 VGND.t366 36.0005
R3300 VGND.n397 VGND.t546 36.0005
R3301 VGND.n397 VGND.t1730 36.0005
R3302 VGND.n2112 VGND.t1474 36.0005
R3303 VGND.n2112 VGND.t1740 36.0005
R3304 VGND.n2107 VGND.t1809 36.0005
R3305 VGND.n2107 VGND.t442 36.0005
R3306 VGND.n2102 VGND.t484 36.0005
R3307 VGND.n2102 VGND.t1720 36.0005
R3308 VGND.n405 VGND.t107 36.0005
R3309 VGND.n405 VGND.t1732 36.0005
R3310 VGND.n2071 VGND.t337 36.0005
R3311 VGND.n2071 VGND.t1742 36.0005
R3312 VGND.n413 VGND.t2643 36.0005
R3313 VGND.n413 VGND.t1722 36.0005
R3314 VGND.n2045 VGND.t674 36.0005
R3315 VGND.n2045 VGND.t1734 36.0005
R3316 VGND.n421 VGND.t2028 36.0005
R3317 VGND.n421 VGND.t1736 36.0005
R3318 VGND.n2019 VGND.t2063 36.0005
R3319 VGND.n2019 VGND.t1744 36.0005
R3320 VGND.n429 VGND.t1058 36.0005
R3321 VGND.n429 VGND.t1724 36.0005
R3322 VGND.n1993 VGND.t928 36.0005
R3323 VGND.n1993 VGND.t1726 36.0005
R3324 VGND.n623 VGND.t1069 36.0005
R3325 VGND.n623 VGND.t436 36.0005
R3326 VGND.n620 VGND.t1957 36.0005
R3327 VGND.n620 VGND.t438 36.0005
R3328 VGND.n618 VGND.t1030 36.0005
R3329 VGND.n618 VGND.t440 36.0005
R3330 VGND.n615 VGND.t1398 36.0005
R3331 VGND.n615 VGND.t1738 36.0005
R3332 VGND.n315 VGND.t1893 36.0005
R3333 VGND.n315 VGND.t1595 36.0005
R3334 VGND.n2328 VGND.t1159 36.0005
R3335 VGND.n2328 VGND.t386 36.0005
R3336 VGND.n2089 VGND.t2213 36.0005
R3337 VGND.n2089 VGND.t330 36.0005
R3338 VGND.n401 VGND.t2226 36.0005
R3339 VGND.n401 VGND.t332 36.0005
R3340 VGND.n2084 VGND.t93 36.0005
R3341 VGND.n2084 VGND.t1597 36.0005
R3342 VGND.n409 VGND.t400 36.0005
R3343 VGND.n409 VGND.t320 36.0005
R3344 VGND.n2058 VGND.t1301 36.0005
R3345 VGND.n2058 VGND.t334 36.0005
R3346 VGND.n417 VGND.t684 36.0005
R3347 VGND.n417 VGND.t1599 36.0005
R3348 VGND.n2032 VGND.t722 36.0005
R3349 VGND.n2032 VGND.t1601 36.0005
R3350 VGND.n425 VGND.t314 36.0005
R3351 VGND.n425 VGND.t322 36.0005
R3352 VGND.n2006 VGND.t2362 36.0005
R3353 VGND.n2006 VGND.t1591 36.0005
R3354 VGND.n433 VGND.t1635 36.0005
R3355 VGND.n433 VGND.t1593 36.0005
R3356 VGND.n1980 VGND.t71 36.0005
R3357 VGND.n1980 VGND.t324 36.0005
R3358 VGND.n645 VGND.t208 36.0005
R3359 VGND.n645 VGND.t326 36.0005
R3360 VGND.n648 VGND.t2656 36.0005
R3361 VGND.n648 VGND.t328 36.0005
R3362 VGND.n642 VGND.t1341 36.0005
R3363 VGND.n642 VGND.t1603 36.0005
R3364 VGND.n450 VGND.t527 36.0005
R3365 VGND.n450 VGND.t1161 36.0005
R3366 VGND.n1957 VGND.t2256 36.0005
R3367 VGND.n1957 VGND.t1229 36.0005
R3368 VGND.n447 VGND.t1850 36.0005
R3369 VGND.n447 VGND.t215 36.0005
R3370 VGND.n900 VGND.t734 36.0005
R3371 VGND.n900 VGND.t553 36.0005
R3372 VGND.n905 VGND.t103 36.0005
R3373 VGND.n905 VGND.t1163 36.0005
R3374 VGND.n910 VGND.t343 36.0005
R3375 VGND.n910 VGND.t1231 36.0005
R3376 VGND.n915 VGND.t2675 36.0005
R3377 VGND.n915 VGND.t555 36.0005
R3378 VGND.n920 VGND.t1973 36.0005
R3379 VGND.n920 VGND.t1165 36.0005
R3380 VGND.n925 VGND.t307 36.0005
R3381 VGND.n925 VGND.t1167 36.0005
R3382 VGND.n930 VGND.t2069 36.0005
R3383 VGND.n930 VGND.t1233 36.0005
R3384 VGND.n935 VGND.t1507 36.0005
R3385 VGND.n935 VGND.t557 36.0005
R3386 VGND.n940 VGND.t728 36.0005
R3387 VGND.n940 VGND.t559 36.0005
R3388 VGND.n945 VGND.t453 36.0005
R3389 VGND.n945 VGND.t1235 36.0005
R3390 VGND.n950 VGND.t2347 36.0005
R3391 VGND.n950 VGND.t704 36.0005
R3392 VGND.n955 VGND.t1096 36.0005
R3393 VGND.n955 VGND.t706 36.0005
R3394 VGND.n658 VGND.t1380 36.0005
R3395 VGND.n658 VGND.t1227 36.0005
R3396 VGND.n453 VGND.t536 36.0005
R3397 VGND.n453 VGND.t691 36.0005
R3398 VGND.n1938 VGND.t1046 36.0005
R3399 VGND.n1938 VGND.t2628 36.0005
R3400 VGND.n1933 VGND.t1210 36.0005
R3401 VGND.n1933 VGND.t2291 36.0005
R3402 VGND.n1928 VGND.t299 36.0005
R3403 VGND.n1928 VGND.t2293 36.0005
R3404 VGND.n461 VGND.t120 36.0005
R3405 VGND.n461 VGND.t693 36.0005
R3406 VGND.n1897 VGND.t217 36.0005
R3407 VGND.n1897 VGND.t2630 36.0005
R3408 VGND.n469 VGND.t282 36.0005
R3409 VGND.n469 VGND.t2295 36.0005
R3410 VGND.n1871 VGND.t665 36.0005
R3411 VGND.n1871 VGND.t695 36.0005
R3412 VGND.n477 VGND.t1196 36.0005
R3413 VGND.n477 VGND.t697 36.0005
R3414 VGND.n1845 VGND.t2601 36.0005
R3415 VGND.n1845 VGND.t2632 36.0005
R3416 VGND.n485 VGND.t2196 36.0005
R3417 VGND.n485 VGND.t2297 36.0005
R3418 VGND.n1819 VGND.t2685 36.0005
R3419 VGND.n1819 VGND.t1728 36.0005
R3420 VGND.n664 VGND.t22 36.0005
R3421 VGND.n664 VGND.t2634 36.0005
R3422 VGND.n1396 VGND.t2524 36.0005
R3423 VGND.n1396 VGND.t2287 36.0005
R3424 VGND.n1391 VGND.t1104 36.0005
R3425 VGND.n1391 VGND.t2289 36.0005
R3426 VGND.n667 VGND.t1425 36.0005
R3427 VGND.n667 VGND.t2626 36.0005
R3428 VGND.n303 VGND.t1896 36.0005
R3429 VGND.n303 VGND.t353 36.0005
R3430 VGND.n2353 VGND.t2042 36.0005
R3431 VGND.n2353 VGND.t2518 36.0005
R3432 VGND.n1915 VGND.t1954 36.0005
R3433 VGND.n1915 VGND.t1922 36.0005
R3434 VGND.n457 VGND.t1205 36.0005
R3435 VGND.n457 VGND.t1924 36.0005
R3436 VGND.n1910 VGND.t85 36.0005
R3437 VGND.n1910 VGND.t355 36.0005
R3438 VGND.n465 VGND.t410 36.0005
R3439 VGND.n465 VGND.t2520 36.0005
R3440 VGND.n1884 VGND.t1305 36.0005
R3441 VGND.n1884 VGND.t1926 36.0005
R3442 VGND.n473 VGND.t1914 36.0005
R3443 VGND.n473 VGND.t357 36.0005
R3444 VGND.n1858 VGND.t725 36.0005
R3445 VGND.n1858 VGND.t1932 36.0005
R3446 VGND.n481 VGND.t318 36.0005
R3447 VGND.n481 VGND.t2522 36.0005
R3448 VGND.n1832 VGND.t2202 36.0005
R3449 VGND.n1832 VGND.t1928 36.0005
R3450 VGND.n489 VGND.t147 36.0005
R3451 VGND.n489 VGND.t1930 36.0005
R3452 VGND.n1806 VGND.t1618 36.0005
R3453 VGND.n1806 VGND.t347 36.0005
R3454 VGND.n1373 VGND.t2354 36.0005
R3455 VGND.n1373 VGND.t349 36.0005
R3456 VGND.n1376 VGND.t382 36.0005
R3457 VGND.n1376 VGND.t351 36.0005
R3458 VGND.n1370 VGND.t1467 36.0005
R3459 VGND.n1370 VGND.t756 36.0005
R3460 VGND.n506 VGND.t657 36.0005
R3461 VGND.n506 VGND.t161 36.0005
R3462 VGND.n1783 VGND.t1169 36.0005
R3463 VGND.n1783 VGND.t157 36.0005
R3464 VGND.n503 VGND.t1758 36.0005
R3465 VGND.n503 VGND.t1669 36.0005
R3466 VGND.n1313 VGND.t739 36.0005
R3467 VGND.n1313 VGND.t1671 36.0005
R3468 VGND.n1318 VGND.t80 36.0005
R3469 VGND.n1318 VGND.t163 36.0005
R3470 VGND.n1323 VGND.t360 36.0005
R3471 VGND.n1323 VGND.t159 36.0005
R3472 VGND.n1328 VGND.t273 36.0005
R3473 VGND.n1328 VGND.t1673 36.0005
R3474 VGND.n1333 VGND.t1920 36.0005
R3475 VGND.n1333 VGND.t151 36.0005
R3476 VGND.n1338 VGND.t186 36.0005
R3477 VGND.n1338 VGND.t153 36.0005
R3478 VGND.n1343 VGND.t2129 36.0005
R3479 VGND.n1343 VGND.t1661 36.0005
R3480 VGND.n1348 VGND.t2072 36.0005
R3481 VGND.n1348 VGND.t1675 36.0005
R3482 VGND.n1353 VGND.t924 36.0005
R3483 VGND.n1353 VGND.t1677 36.0005
R3484 VGND.n1358 VGND.t29 36.0005
R3485 VGND.n1358 VGND.t1663 36.0005
R3486 VGND.n1305 VGND.t1937 36.0005
R3487 VGND.n1305 VGND.t1665 36.0005
R3488 VGND.n1308 VGND.t1482 36.0005
R3489 VGND.n1308 VGND.t1667 36.0005
R3490 VGND.n1302 VGND.t1440 36.0005
R3491 VGND.n1302 VGND.t155 36.0005
R3492 VGND.n509 VGND.t1889 36.0005
R3493 VGND.n509 VGND.t597 36.0005
R3494 VGND.n1764 VGND.t1155 36.0005
R3495 VGND.n1764 VGND.t749 36.0005
R3496 VGND.n1759 VGND.t2209 36.0005
R3497 VGND.n1759 VGND.t2020 36.0005
R3498 VGND.n1754 VGND.t2222 36.0005
R3499 VGND.n1754 VGND.t1645 36.0005
R3500 VGND.n517 VGND.t88 36.0005
R3501 VGND.n517 VGND.t599 36.0005
R3502 VGND.n1723 VGND.t396 36.0005
R3503 VGND.n1723 VGND.t1189 36.0005
R3504 VGND.n525 VGND.t1296 36.0005
R3505 VGND.n525 VGND.t1647 36.0005
R3506 VGND.n1697 VGND.t680 36.0005
R3507 VGND.n1697 VGND.t601 36.0005
R3508 VGND.n533 VGND.t1182 36.0005
R3509 VGND.n533 VGND.t745 36.0005
R3510 VGND.n1671 VGND.t49 36.0005
R3511 VGND.n1671 VGND.t1191 36.0005
R3512 VGND.n541 VGND.t2358 36.0005
R3513 VGND.n541 VGND.t1649 36.0005
R3514 VGND.n1645 VGND.t1631 36.0005
R3515 VGND.n1645 VGND.t1651 36.0005
R3516 VGND.n575 VGND.t67 36.0005
R3517 VGND.n575 VGND.t2014 36.0005
R3518 VGND.n1518 VGND.t204 36.0005
R3519 VGND.n1518 VGND.t2016 36.0005
R3520 VGND.n1513 VGND.t2652 36.0005
R3521 VGND.n1513 VGND.t2018 36.0005
R3522 VGND.n571 VGND.t1347 36.0005
R3523 VGND.n571 VGND.t747 36.0005
R3524 VGND.n290 VGND.t542 36.0005
R3525 VGND.n290 VGND.t2152 36.0005
R3526 VGND.n2378 VGND.t1240 36.0005
R3527 VGND.n2378 VGND.t2162 36.0005
R3528 VGND.n1741 VGND.t198 36.0005
R3529 VGND.n1741 VGND.t2331 36.0005
R3530 VGND.n513 VGND.t2053 36.0005
R3531 VGND.n513 VGND.t2333 36.0005
R3532 VGND.n1736 VGND.t115 36.0005
R3533 VGND.n1736 VGND.t2154 36.0005
R3534 VGND.n521 VGND.t221 36.0005
R3535 VGND.n521 VGND.t2164 36.0005
R3536 VGND.n1710 VGND.t434 36.0005
R3537 VGND.n1710 VGND.t2335 36.0005
R3538 VGND.n529 VGND.t671 36.0005
R3539 VGND.n529 VGND.t2156 36.0005
R3540 VGND.n1684 VGND.t2024 36.0005
R3541 VGND.n1684 VGND.t2158 36.0005
R3542 VGND.n537 VGND.t2059 36.0005
R3543 VGND.n537 VGND.t2166 36.0005
R3544 VGND.n1658 VGND.t1055 36.0005
R3545 VGND.n1658 VGND.t2337 36.0005
R3546 VGND.n545 VGND.t1141 36.0005
R3547 VGND.n545 VGND.t1627 36.0005
R3548 VGND.n1632 VGND.t26 36.0005
R3549 VGND.n1632 VGND.t2325 36.0005
R3550 VGND.n564 VGND.t2094 36.0005
R3551 VGND.n564 VGND.t2327 36.0005
R3552 VGND.n1533 VGND.t589 36.0005
R3553 VGND.n1533 VGND.t2329 36.0005
R3554 VGND.n567 VGND.t1413 36.0005
R3555 VGND.n567 VGND.t2160 36.0005
R3556 VGND.n1601 VGND.t1886 36.0005
R3557 VGND.n1601 VGND.t2140 36.0005
R3558 VGND.n1609 VGND.t1153 36.0005
R3559 VGND.n1609 VGND.t2150 36.0005
R3560 VGND.n559 VGND.t2207 36.0005
R3561 VGND.n559 VGND.t1496 36.0005
R3562 VGND.n1596 VGND.t2220 36.0005
R3563 VGND.n1596 VGND.t1498 36.0005
R3564 VGND.n1591 VGND.t101 36.0005
R3565 VGND.n1591 VGND.t2142 36.0005
R3566 VGND.n1586 VGND.t394 36.0005
R3567 VGND.n1586 VGND.t472 36.0005
R3568 VGND.n1581 VGND.t1294 36.0005
R3569 VGND.n1581 VGND.t1500 36.0005
R3570 VGND.n1576 VGND.t678 36.0005
R3571 VGND.n1576 VGND.t2144 36.0005
R3572 VGND.n1571 VGND.t1179 36.0005
R3573 VGND.n1571 VGND.t2146 36.0005
R3574 VGND.n1566 VGND.t47 36.0005
R3575 VGND.n1566 VGND.t474 36.0005
R3576 VGND.n1561 VGND.t2356 36.0005
R3577 VGND.n1561 VGND.t2136 36.0005
R3578 VGND.n1556 VGND.t2037 36.0005
R3579 VGND.n1556 VGND.t2138 36.0005
R3580 VGND.n1551 VGND.t65 36.0005
R3581 VGND.n1551 VGND.t476 36.0005
R3582 VGND.n1546 VGND.t202 36.0005
R3583 VGND.n1546 VGND.t1492 36.0005
R3584 VGND.n672 VGND.t2650 36.0005
R3585 VGND.n672 VGND.t1494 36.0005
R3586 VGND.n670 VGND.t1350 36.0005
R3587 VGND.n670 VGND.t2148 36.0005
R3588 VGND.n278 VGND.t524 36.0005
R3589 VGND.n278 VGND.t2047 36.0005
R3590 VGND.n2398 VGND.t2254 36.0005
R3591 VGND.n2398 VGND.t2082 36.0005
R3592 VGND.n841 VGND.t2217 36.0005
R3593 VGND.n841 VGND.t2086 36.0005
R3594 VGND.n846 VGND.t488 36.0005
R3595 VGND.n846 VGND.t2088 36.0005
R3596 VGND.n851 VGND.t111 36.0005
R3597 VGND.n851 VGND.t2049 36.0005
R3598 VGND.n856 VGND.t341 36.0005
R3599 VGND.n856 VGND.t2084 36.0005
R3600 VGND.n861 VGND.t2673 36.0005
R3601 VGND.n861 VGND.t1748 36.0005
R3602 VGND.n866 VGND.t1970 36.0005
R3603 VGND.n866 VGND.t2051 36.0005
R3604 VGND.n871 VGND.t304 36.0005
R3605 VGND.n871 VGND.t2078 36.0005
R3606 VGND.n876 VGND.t2067 36.0005
R3607 VGND.n876 VGND.t2317 36.0005
R3608 VGND.n881 VGND.t1505 36.0005
R3609 VGND.n881 VGND.t1750 36.0005
R3610 VGND.n886 VGND.t933 36.0005
R3611 VGND.n886 VGND.t1752 36.0005
R3612 VGND.n828 VGND.t1073 36.0005
R3613 VGND.n828 VGND.t2319 36.0005
R3614 VGND.n836 VGND.t1963 36.0005
R3615 VGND.n836 VGND.t2321 36.0005
R3616 VGND.n831 VGND.t1036 36.0005
R3617 VGND.n831 VGND.t2323 36.0005
R3618 VGND.n824 VGND.t1386 36.0005
R3619 VGND.n824 VGND.t2080 36.0005
R3620 VGND.n787 VGND.t863 36.0005
R3621 VGND.n787 VGND.t867 36.0005
R3622 VGND.n1223 VGND.t776 36.0005
R3623 VGND.n1223 VGND.t780 36.0005
R3624 VGND.n792 VGND.t1540 36.0005
R3625 VGND.n792 VGND.t1545 36.0005
R3626 VGND.n1204 VGND.t854 36.0005
R3627 VGND.n1204 VGND.t1548 36.0005
R3628 VGND.n795 VGND.t874 36.0005
R3629 VGND.n795 VGND.t876 36.0005
R3630 VGND.n1191 VGND.t801 36.0005
R3631 VGND.n1191 VGND.t803 36.0005
R3632 VGND.n800 VGND.t1553 36.0005
R3633 VGND.n800 VGND.t1557 36.0005
R3634 VGND.n1172 VGND.t886 36.0005
R3635 VGND.n1172 VGND.t888 36.0005
R3636 VGND.n803 VGND.t900 36.0005
R3637 VGND.n803 VGND.t902 36.0005
R3638 VGND.n1159 VGND.t809 36.0005
R3639 VGND.n1159 VGND.t813 36.0005
R3640 VGND.n808 VGND.t1585 36.0005
R3641 VGND.n808 VGND.t1571 36.0005
R3642 VGND.n1140 VGND.t838 36.0005
R3643 VGND.n1140 VGND.t842 36.0005
R3644 VGND.n811 VGND.t821 36.0005
R3645 VGND.n811 VGND.t823 36.0005
R3646 VGND.n1127 VGND.t2594 36.0005
R3647 VGND.n1127 VGND.t2596 36.0005
R3648 VGND.n813 VGND.t1581 36.0005
R3649 VGND.n813 VGND.t1525 36.0005
R3650 VGND.n814 VGND.t760 36.0005
R3651 VGND.n814 VGND.t762 36.0005
R3652 VGND.n717 VGND.t774 36.0005
R3653 VGND.n717 VGND.t778 36.0005
R3654 VGND.n776 VGND.t1521 36.0005
R3655 VGND.n776 VGND.t1523 36.0005
R3656 VGND.n771 VGND.t852 36.0005
R3657 VGND.n771 VGND.t856 36.0005
R3658 VGND.n766 VGND.t771 36.0005
R3659 VGND.n766 VGND.t865 36.0005
R3660 VGND.n761 VGND.t789 36.0005
R3661 VGND.n761 VGND.t791 36.0005
R3662 VGND.n756 VGND.t1538 36.0005
R3663 VGND.n756 VGND.t1542 36.0005
R3664 VGND.n751 VGND.t870 36.0005
R3665 VGND.n751 VGND.t872 36.0005
R3666 VGND.n746 VGND.t793 36.0005
R3667 VGND.n746 VGND.t795 36.0005
R3668 VGND.n741 VGND.t807 36.0005
R3669 VGND.n741 VGND.t811 36.0005
R3670 VGND.n736 VGND.t1551 36.0005
R3671 VGND.n736 VGND.t1555 36.0005
R3672 VGND.n731 VGND.t894 36.0005
R3673 VGND.n731 VGND.t884 36.0005
R3674 VGND.n726 VGND.t896 36.0005
R3675 VGND.n726 VGND.t898 36.0005
R3676 VGND.n721 VGND.t1561 36.0005
R3677 VGND.n721 VGND.t1563 36.0005
R3678 VGND.n682 VGND.t1579 36.0005
R3679 VGND.n682 VGND.t1583 36.0005
R3680 VGND.n678 VGND.t892 36.0005
R3681 VGND.n678 VGND.t840 36.0005
R3682 VGND.n675 VGND.t2590 36.0005
R3683 VGND.n675 VGND.t2592 36.0005
R3684 VGND.n74 VGND.n72 34.6358
R3685 VGND.n1109 VGND.n1091 34.6358
R3686 VGND.n1105 VGND.n1091 34.6358
R3687 VGND.n1105 VGND.n1104 34.6358
R3688 VGND.n1104 VGND.n1103 34.6358
R3689 VGND.n1103 VGND.n1093 34.6358
R3690 VGND.n1087 VGND.n1061 34.6358
R3691 VGND.n1082 VGND.n1062 34.6358
R3692 VGND.n1078 VGND.n1062 34.6358
R3693 VGND.n1078 VGND.n1077 34.6358
R3694 VGND.n1077 VGND.n1076 34.6358
R3695 VGND.n1076 VGND.n1064 34.6358
R3696 VGND.n130 VGND.n125 34.6358
R3697 VGND.n135 VGND.n134 34.6358
R3698 VGND.n598 VGND.n593 34.6358
R3699 VGND.n603 VGND.n602 34.6358
R3700 VGND.n976 VGND.n975 34.6358
R3701 VGND.n984 VGND.n983 34.6358
R3702 VGND.n980 VGND.n979 34.6358
R3703 VGND.n1020 VGND.n1000 34.6358
R3704 VGND.n1016 VGND.n1000 34.6358
R3705 VGND.n1016 VGND.n1015 34.6358
R3706 VGND.n1015 VGND.n1014 34.6358
R3707 VGND.n1014 VGND.n1002 34.6358
R3708 VGND.n1056 VGND.n1030 34.6358
R3709 VGND.n1051 VGND.n1031 34.6358
R3710 VGND.n1047 VGND.n1031 34.6358
R3711 VGND.n1047 VGND.n1046 34.6358
R3712 VGND.n1046 VGND.n1045 34.6358
R3713 VGND.n1045 VGND.n1033 34.6358
R3714 VGND.n160 VGND.n155 34.6358
R3715 VGND.n165 VGND.n164 34.6358
R3716 VGND.n17 VGND.n16 34.6358
R3717 VGND.n19 VGND.n10 34.6358
R3718 VGND.n23 VGND.n10 34.6358
R3719 VGND.n24 VGND.n23 34.6358
R3720 VGND.n25 VGND.n24 34.6358
R3721 VGND.n25 VGND.n8 34.6358
R3722 VGND.n46 VGND.n45 34.6358
R3723 VGND.n48 VGND.n37 34.6358
R3724 VGND.n52 VGND.n37 34.6358
R3725 VGND.n53 VGND.n52 34.6358
R3726 VGND.n54 VGND.n53 34.6358
R3727 VGND.n54 VGND.n35 34.6358
R3728 VGND.n100 VGND.n99 34.6358
R3729 VGND.n104 VGND.n103 34.6358
R3730 VGND.n2844 VGND.n2843 34.6358
R3731 VGND.n2848 VGND.n2847 34.6358
R3732 VGND.n2876 VGND.n2875 34.6358
R3733 VGND.n2880 VGND.n2879 34.6358
R3734 VGND.n78 VGND.n77 34.6358
R3735 VGND.n2919 VGND.n2913 34.6358
R3736 VGND.n2922 VGND.n2921 34.6358
R3737 VGND.n2922 VGND.n2909 34.6358
R3738 VGND.n2926 VGND.n2909 34.6358
R3739 VGND.n2927 VGND.n2926 34.6358
R3740 VGND.n2928 VGND.n2927 34.6358
R3741 VGND.n2944 VGND.n58 34.6358
R3742 VGND.n2959 VGND.n2958 34.6358
R3743 VGND.n2961 VGND.n2950 34.6358
R3744 VGND.n2965 VGND.n2950 34.6358
R3745 VGND.n2966 VGND.n2965 34.6358
R3746 VGND.n2967 VGND.n2966 34.6358
R3747 VGND.n2967 VGND.n2948 34.6358
R3748 VGND.n2976 VGND.n2971 34.6358
R3749 VGND.n2 VGND.t1605 34.4422
R3750 VGND.n995 VGND.n898 33.1299
R3751 VGND.n2901 VGND.n2900 33.1299
R3752 VGND.n80 VGND.n62 32.377
R3753 VGND.n986 VGND.n985 32.377
R3754 VGND.n106 VGND.n105 32.377
R3755 VGND.n2850 VGND.n2849 32.377
R3756 VGND.n2882 VGND.n2881 32.377
R3757 VGND.n80 VGND.n79 32.377
R3758 VGND.n986 VGND.n964 32.0005
R3759 VGND.n141 VGND.n138 30.4946
R3760 VGND.n609 VGND.n606 30.4946
R3761 VGND.n171 VGND.n168 30.4946
R3762 VGND.n109 VGND.n86 29.8709
R3763 VGND.n1099 VGND.n1098 28.9887
R3764 VGND.n1072 VGND.n1071 28.9887
R3765 VGND.n1010 VGND.n1009 28.9887
R3766 VGND.n1041 VGND.n1040 28.9887
R3767 VGND.n18 VGND.n17 27.8593
R3768 VGND.n47 VGND.n46 27.8593
R3769 VGND.n2920 VGND.n2919 27.8593
R3770 VGND.n2960 VGND.n2959 27.8593
R3771 VGND.n119 VGND.n118 27.0003
R3772 VGND.n2855 VGND.n2854 26.8591
R3773 VGND.n983 VGND.n968 26.3534
R3774 VGND.n103 VGND.n92 26.3534
R3775 VGND.n2847 VGND.n2836 26.3534
R3776 VGND.n2879 VGND.n2868 26.3534
R3777 VGND.n77 VGND.n67 26.3534
R3778 VGND.n142 VGND.n141 25.977
R3779 VGND.n610 VGND.n609 25.977
R3780 VGND.n585 VGND.n582 25.977
R3781 VGND.n172 VGND.n171 25.977
R3782 VGND.n2887 VGND.n2862 25.977
R3783 VGND.n1095 VGND.t255 24.9236
R3784 VGND.n1095 VGND.t267 24.9236
R3785 VGND.n1097 VGND.t2373 24.9236
R3786 VGND.n1097 VGND.t2313 24.9236
R3787 VGND.n1067 VGND.t179 24.9236
R3788 VGND.n1067 VGND.t180 24.9236
R3789 VGND.n1066 VGND.t257 24.9236
R3790 VGND.n1066 VGND.t269 24.9236
R3791 VGND.n1070 VGND.t181 24.9236
R3792 VGND.n1070 VGND.t2377 24.9236
R3793 VGND.n1069 VGND.t2374 24.9236
R3794 VGND.n1069 VGND.t2314 24.9236
R3795 VGND.n132 VGND.t2376 24.9236
R3796 VGND.n132 VGND.t408 24.9236
R3797 VGND.n131 VGND.t2366 24.9236
R3798 VGND.n131 VGND.t2514 24.9236
R3799 VGND.n122 VGND.t192 24.9236
R3800 VGND.n122 VGND.t2371 24.9236
R3801 VGND.n121 VGND.t2614 24.9236
R3802 VGND.n121 VGND.t263 24.9236
R3803 VGND.n140 VGND.t190 24.9236
R3804 VGND.n140 VGND.t191 24.9236
R3805 VGND.n139 VGND.t1081 24.9236
R3806 VGND.n139 VGND.t1082 24.9236
R3807 VGND.n600 VGND.t15 24.9236
R3808 VGND.n600 VGND.t1080 24.9236
R3809 VGND.n599 VGND.t5 24.9236
R3810 VGND.n599 VGND.t1074 24.9236
R3811 VGND.n590 VGND.t479 24.9236
R3812 VGND.n590 VGND.t14 24.9236
R3813 VGND.n589 VGND.t1683 24.9236
R3814 VGND.n589 VGND.t407 24.9236
R3815 VGND.n608 VGND.t481 24.9236
R3816 VGND.n608 VGND.t480 24.9236
R3817 VGND.n607 VGND.t1685 24.9236
R3818 VGND.n607 VGND.t1684 24.9236
R3819 VGND.n966 VGND.t265 24.9236
R3820 VGND.n966 VGND.t2511 24.9236
R3821 VGND.n967 VGND.t52 24.9236
R3822 VGND.n967 VGND.t2368 24.9236
R3823 VGND.n965 VGND.t56 24.9236
R3824 VGND.n965 VGND.t54 24.9236
R3825 VGND.n970 VGND.t2370 24.9236
R3826 VGND.n970 VGND.t2311 24.9236
R3827 VGND.n1005 VGND.t259 24.9236
R3828 VGND.n1005 VGND.t270 24.9236
R3829 VGND.n1004 VGND.t1075 24.9236
R3830 VGND.n1004 VGND.t1078 24.9236
R3831 VGND.n1008 VGND.t2375 24.9236
R3832 VGND.n1008 VGND.t2315 24.9236
R3833 VGND.n1007 VGND.t268 24.9236
R3834 VGND.n1007 VGND.t2512 24.9236
R3835 VGND.n1036 VGND.t2623 24.9236
R3836 VGND.n1036 VGND.t2624 24.9236
R3837 VGND.n1035 VGND.t2513 24.9236
R3838 VGND.n1035 VGND.t2515 24.9236
R3839 VGND.n1039 VGND.t2509 24.9236
R3840 VGND.n1039 VGND.t177 24.9236
R3841 VGND.n1038 VGND.t3 24.9236
R3842 VGND.n1038 VGND.t182 24.9236
R3843 VGND.n162 VGND.t175 24.9236
R3844 VGND.n162 VGND.t261 24.9236
R3845 VGND.n161 VGND.t12 24.9236
R3846 VGND.n161 VGND.t1077 24.9236
R3847 VGND.n152 VGND.t470 24.9236
R3848 VGND.n152 VGND.t17 24.9236
R3849 VGND.n151 VGND.t234 24.9236
R3850 VGND.n151 VGND.t11 24.9236
R3851 VGND.n170 VGND.t468 24.9236
R3852 VGND.n170 VGND.t469 24.9236
R3853 VGND.n169 VGND.t237 24.9236
R3854 VGND.n169 VGND.t235 24.9236
R3855 VGND.n13 VGND.t2497 24.9236
R3856 VGND.n13 VGND.t2416 24.9236
R3857 VGND.n12 VGND.t2426 24.9236
R3858 VGND.n12 VGND.t2434 24.9236
R3859 VGND.n42 VGND.t2476 24.9236
R3860 VGND.n42 VGND.t2508 24.9236
R3861 VGND.n41 VGND.t2432 24.9236
R3862 VGND.n41 VGND.t2471 24.9236
R3863 VGND.n40 VGND.t2482 24.9236
R3864 VGND.n40 VGND.t2450 24.9236
R3865 VGND.n39 VGND.t2442 24.9236
R3866 VGND.n39 VGND.t2500 24.9236
R3867 VGND.n95 VGND.t2422 24.9236
R3868 VGND.n95 VGND.t2463 24.9236
R3869 VGND.n94 VGND.t2480 24.9236
R3870 VGND.n94 VGND.t2420 24.9236
R3871 VGND.n91 VGND.t2430 24.9236
R3872 VGND.n91 VGND.t2251 24.9236
R3873 VGND.n90 VGND.t2486 24.9236
R3874 VGND.n90 VGND.t753 24.9236
R3875 VGND.n89 VGND.t2250 24.9236
R3876 VGND.n89 VGND.t2252 24.9236
R3877 VGND.n88 VGND.t1277 24.9236
R3878 VGND.n88 VGND.t459 24.9236
R3879 VGND.n2839 VGND.t2454 24.9236
R3880 VGND.n2839 VGND.t2487 24.9236
R3881 VGND.n2838 VGND.t2502 24.9236
R3882 VGND.n2838 VGND.t2452 24.9236
R3883 VGND.n2835 VGND.t2459 24.9236
R3884 VGND.n2835 VGND.t2238 24.9236
R3885 VGND.n2834 VGND.t2414 24.9236
R3886 VGND.n2834 VGND.t2680 24.9236
R3887 VGND.n2833 VGND.t715 24.9236
R3888 VGND.n2833 VGND.t720 24.9236
R3889 VGND.n2832 VGND.t1292 24.9236
R3890 VGND.n2832 VGND.t1905 24.9236
R3891 VGND.n2871 VGND.t2458 24.9236
R3892 VGND.n2871 VGND.t2492 24.9236
R3893 VGND.n2870 VGND.t2438 24.9236
R3894 VGND.n2870 VGND.t2479 24.9236
R3895 VGND.n2867 VGND.t2462 24.9236
R3896 VGND.n2867 VGND.t2668 24.9236
R3897 VGND.n2866 VGND.t2447 24.9236
R3898 VGND.n2866 VGND.t1323 24.9236
R3899 VGND.n2865 VGND.t2667 24.9236
R3900 VGND.n2865 VGND.t2665 24.9236
R3901 VGND.n2864 VGND.t1319 24.9236
R3902 VGND.n2864 VGND.t1313 24.9236
R3903 VGND.n65 VGND.t2469 24.9236
R3904 VGND.n65 VGND.t2506 24.9236
R3905 VGND.n66 VGND.t2473 24.9236
R3906 VGND.n66 VGND.t141 24.9236
R3907 VGND.n64 VGND.t137 24.9236
R3908 VGND.n64 VGND.t131 24.9236
R3909 VGND.n69 VGND.t2465 24.9236
R3910 VGND.n69 VGND.t2499 24.9236
R3911 VGND.n2915 VGND.t2448 24.9236
R3912 VGND.n2915 VGND.t2485 24.9236
R3913 VGND.n2914 VGND.t2436 24.9236
R3914 VGND.n2914 VGND.t2475 24.9236
R3915 VGND.n2912 VGND.t2457 24.9236
R3916 VGND.n2912 VGND.t2418 24.9236
R3917 VGND.n2911 VGND.t2444 24.9236
R3918 VGND.n2911 VGND.t2501 24.9236
R3919 VGND.n2955 VGND.t2493 24.9236
R3920 VGND.n2955 VGND.t2445 24.9236
R3921 VGND.n2954 VGND.t2484 24.9236
R3922 VGND.n2954 VGND.t2428 24.9236
R3923 VGND.n2953 VGND.t2504 24.9236
R3924 VGND.n2953 VGND.t2477 24.9236
R3925 VGND.n2952 VGND.t2489 24.9236
R3926 VGND.n2952 VGND.t2461 24.9236
R3927 VGND.n142 VGND.n116 24.4711
R3928 VGND.n610 VGND.n581 24.4711
R3929 VGND.n585 VGND.n584 24.4711
R3930 VGND.n996 VGND.n995 24.4711
R3931 VGND.n1025 VGND.n999 24.4711
R3932 VGND.n172 VGND.n148 24.4711
R3933 VGND.n106 VGND.n85 24.4711
R3934 VGND.n2850 VGND.n2829 24.4711
R3935 VGND.n2882 VGND.n2861 24.4711
R3936 VGND.n2887 VGND.n2886 24.4711
R3937 VGND.n2902 VGND.n2901 24.4711
R3938 VGND.n2933 VGND.n2932 24.4711
R3939 VGND.n2858 VGND.n2830 23.7181
R3940 VGND.n1111 VGND.n1109 23.7181
R3941 VGND.n1083 VGND.n1061 23.7181
R3942 VGND.n1083 VGND.n1082 23.7181
R3943 VGND.n146 VGND.n115 23.7181
R3944 VGND.n990 VGND.n899 23.7181
R3945 VGND.n1021 VGND.n1020 23.7181
R3946 VGND.n1052 VGND.n1030 23.7181
R3947 VGND.n1052 VGND.n1051 23.7181
R3948 VGND.n2992 VGND.n8 23.7181
R3949 VGND.n2945 VGND.n35 23.7181
R3950 VGND.n2928 VGND.n2907 23.7181
R3951 VGND.n2945 VGND.n2944 23.7181
R3952 VGND.n2977 VGND.n2948 23.7181
R3953 VGND.n2977 VGND.n2976 23.7181
R3954 VGND.n991 VGND.n990 23.3417
R3955 VGND.n2896 VGND.n84 23.3417
R3956 VGND.n2896 VGND.n61 23.3417
R3957 VGND.n1099 VGND.n1096 21.4593
R3958 VGND.n1072 VGND.n1068 21.4593
R3959 VGND.n1010 VGND.n1006 21.4593
R3960 VGND.n1041 VGND.n1037 21.4593
R3961 VGND.n98 VGND.n97 21.0905
R3962 VGND.n2842 VGND.n2841 21.0905
R3963 VGND.n2874 VGND.n2873 21.0905
R3964 VGND.n71 VGND.n70 21.0905
R3965 VGND.n99 VGND.n98 20.3299
R3966 VGND.n2843 VGND.n2842 20.3299
R3967 VGND.n2875 VGND.n2874 20.3299
R3968 VGND.n72 VGND.n71 20.3299
R3969 VGND.n138 VGND.n123 19.9534
R3970 VGND.n606 VGND.n591 19.9534
R3971 VGND.n168 VGND.n153 19.9534
R3972 VGND.n1026 VGND.n1025 19.2005
R3973 VGND.n1057 VGND.n1056 19.2005
R3974 VGND.n2934 VGND.n2933 19.2005
R3975 VGND.n2939 VGND.n58 19.2005
R3976 VGND.t2526 VGND.t226 16.8587
R3977 VGND.t1795 VGND.t224 16.8587
R3978 VGND.t1221 VGND.t708 16.8587
R3979 VGND.t2032 VGND.t710 16.8587
R3980 VGND.n1089 VGND.n1088 16.077
R3981 VGND.n2973 VGND.n2972 16.077
R3982 VGND.n1027 VGND.n1026 15.4358
R3983 VGND.n2935 VGND.n2934 15.4358
R3984 VGND.n118 VGND.n117 14.6829
R3985 VGND.n1058 VGND.n1057 14.6829
R3986 VGND.n2854 VGND.n2853 14.6829
R3987 VGND.n2940 VGND.n2939 14.6829
R3988 VGND.n127 VGND.n126 14.5711
R3989 VGND.n595 VGND.n594 14.5711
R3990 VGND.n974 VGND.n973 14.5711
R3991 VGND.n157 VGND.n156 14.5711
R3992 VGND.n614 VGND.n582 14.3064
R3993 VGND.n2891 VGND.n2862 14.3064
R3994 VGND.n134 VGND.n133 13.9299
R3995 VGND.n602 VGND.n601 13.9299
R3996 VGND.n979 VGND.n971 13.9299
R3997 VGND.n164 VGND.n163 13.9299
R3998 VGND.n1021 VGND.n999 13.5534
R3999 VGND.n2932 VGND.n2907 13.5534
R4000 VGND.n146 VGND.n116 13.177
R4001 VGND.n614 VGND.n581 13.177
R4002 VGND.n176 VGND.n148 13.177
R4003 VGND.n112 VGND.n85 13.177
R4004 VGND.n2858 VGND.n2829 13.177
R4005 VGND.n2891 VGND.n2861 13.177
R4006 VGND.n176 VGND.n149 12.8005
R4007 VGND.n112 VGND.n86 12.8005
R4008 VGND.n3006 VGND.t2697 12.5645
R4009 VGND.n1088 VGND.n1087 10.5417
R4010 VGND.n2972 VGND.n2971 10.5417
R4011 VGND.n1059 VGND.n1058 10.0534
R4012 VGND.n2941 VGND.n2940 10.0534
R4013 VGND.n1100 VGND.n1099 9.3005
R4014 VGND.n1101 VGND.n1093 9.3005
R4015 VGND.n1103 VGND.n1102 9.3005
R4016 VGND.n1104 VGND.n1092 9.3005
R4017 VGND.n1106 VGND.n1105 9.3005
R4018 VGND.n1107 VGND.n1091 9.3005
R4019 VGND.n1109 VGND.n1108 9.3005
R4020 VGND.n1112 VGND.n1111 9.3005
R4021 VGND.n1073 VGND.n1072 9.3005
R4022 VGND.n1074 VGND.n1064 9.3005
R4023 VGND.n1076 VGND.n1075 9.3005
R4024 VGND.n1077 VGND.n1063 9.3005
R4025 VGND.n1079 VGND.n1078 9.3005
R4026 VGND.n1080 VGND.n1062 9.3005
R4027 VGND.n1082 VGND.n1081 9.3005
R4028 VGND.n1085 VGND.n1061 9.3005
R4029 VGND.n1087 VGND.n1086 9.3005
R4030 VGND.n1084 VGND.n1083 9.3005
R4031 VGND.n144 VGND.n116 9.3005
R4032 VGND.n128 VGND.n125 9.3005
R4033 VGND.n130 VGND.n129 9.3005
R4034 VGND.n134 VGND.n124 9.3005
R4035 VGND.n136 VGND.n135 9.3005
R4036 VGND.n138 VGND.n137 9.3005
R4037 VGND.n141 VGND.n120 9.3005
R4038 VGND.n143 VGND.n142 9.3005
R4039 VGND.n119 VGND.n115 9.3005
R4040 VGND.n146 VGND.n145 9.3005
R4041 VGND.n584 VGND.n583 9.3005
R4042 VGND.n587 VGND.n582 9.3005
R4043 VGND.n612 VGND.n581 9.3005
R4044 VGND.n596 VGND.n593 9.3005
R4045 VGND.n598 VGND.n597 9.3005
R4046 VGND.n602 VGND.n592 9.3005
R4047 VGND.n604 VGND.n603 9.3005
R4048 VGND.n606 VGND.n605 9.3005
R4049 VGND.n609 VGND.n588 9.3005
R4050 VGND.n611 VGND.n610 9.3005
R4051 VGND.n586 VGND.n585 9.3005
R4052 VGND.n614 VGND.n613 9.3005
R4053 VGND.n997 VGND.n996 9.3005
R4054 VGND.n988 VGND.n899 9.3005
R4055 VGND.n975 VGND.n972 9.3005
R4056 VGND.n977 VGND.n976 9.3005
R4057 VGND.n979 VGND.n978 9.3005
R4058 VGND.n981 VGND.n980 9.3005
R4059 VGND.n983 VGND.n982 9.3005
R4060 VGND.n984 VGND.n963 9.3005
R4061 VGND.n987 VGND.n986 9.3005
R4062 VGND.n993 VGND.n992 9.3005
R4063 VGND.n995 VGND.n994 9.3005
R4064 VGND.n990 VGND.n989 9.3005
R4065 VGND.n1011 VGND.n1010 9.3005
R4066 VGND.n1012 VGND.n1002 9.3005
R4067 VGND.n1014 VGND.n1013 9.3005
R4068 VGND.n1015 VGND.n1001 9.3005
R4069 VGND.n1017 VGND.n1016 9.3005
R4070 VGND.n1018 VGND.n1000 9.3005
R4071 VGND.n1020 VGND.n1019 9.3005
R4072 VGND.n1023 VGND.n999 9.3005
R4073 VGND.n1025 VGND.n1024 9.3005
R4074 VGND.n1028 VGND.n1027 9.3005
R4075 VGND.n1022 VGND.n1021 9.3005
R4076 VGND.n1042 VGND.n1041 9.3005
R4077 VGND.n1043 VGND.n1033 9.3005
R4078 VGND.n1045 VGND.n1044 9.3005
R4079 VGND.n1046 VGND.n1032 9.3005
R4080 VGND.n1048 VGND.n1047 9.3005
R4081 VGND.n1049 VGND.n1031 9.3005
R4082 VGND.n1051 VGND.n1050 9.3005
R4083 VGND.n1054 VGND.n1030 9.3005
R4084 VGND.n1056 VGND.n1055 9.3005
R4085 VGND.n1053 VGND.n1052 9.3005
R4086 VGND.n174 VGND.n148 9.3005
R4087 VGND.n158 VGND.n155 9.3005
R4088 VGND.n160 VGND.n159 9.3005
R4089 VGND.n164 VGND.n154 9.3005
R4090 VGND.n166 VGND.n165 9.3005
R4091 VGND.n168 VGND.n167 9.3005
R4092 VGND.n171 VGND.n150 9.3005
R4093 VGND.n173 VGND.n172 9.3005
R4094 VGND.n176 VGND.n175 9.3005
R4095 VGND.n2992 VGND.n2991 9.3005
R4096 VGND.n16 VGND.n15 9.3005
R4097 VGND.n17 VGND.n11 9.3005
R4098 VGND.n20 VGND.n19 9.3005
R4099 VGND.n21 VGND.n10 9.3005
R4100 VGND.n23 VGND.n22 9.3005
R4101 VGND.n24 VGND.n9 9.3005
R4102 VGND.n26 VGND.n25 9.3005
R4103 VGND.n27 VGND.n8 9.3005
R4104 VGND.n110 VGND.n86 9.3005
R4105 VGND.n99 VGND.n93 9.3005
R4106 VGND.n101 VGND.n100 9.3005
R4107 VGND.n103 VGND.n102 9.3005
R4108 VGND.n104 VGND.n87 9.3005
R4109 VGND.n107 VGND.n106 9.3005
R4110 VGND.n108 VGND.n85 9.3005
R4111 VGND.n112 VGND.n111 9.3005
R4112 VGND.n2856 VGND.n2830 9.3005
R4113 VGND.n2843 VGND.n2837 9.3005
R4114 VGND.n2845 VGND.n2844 9.3005
R4115 VGND.n2847 VGND.n2846 9.3005
R4116 VGND.n2848 VGND.n2831 9.3005
R4117 VGND.n2851 VGND.n2850 9.3005
R4118 VGND.n2852 VGND.n2829 9.3005
R4119 VGND.n2858 VGND.n2857 9.3005
R4120 VGND.n2886 VGND.n2885 9.3005
R4121 VGND.n2875 VGND.n2869 9.3005
R4122 VGND.n2877 VGND.n2876 9.3005
R4123 VGND.n2879 VGND.n2878 9.3005
R4124 VGND.n2880 VGND.n2863 9.3005
R4125 VGND.n2883 VGND.n2882 9.3005
R4126 VGND.n2884 VGND.n2861 9.3005
R4127 VGND.n2889 VGND.n2862 9.3005
R4128 VGND.n2888 VGND.n2887 9.3005
R4129 VGND.n2891 VGND.n2890 9.3005
R4130 VGND.n2903 VGND.n2902 9.3005
R4131 VGND.n72 VGND.n68 9.3005
R4132 VGND.n75 VGND.n74 9.3005
R4133 VGND.n77 VGND.n76 9.3005
R4134 VGND.n78 VGND.n63 9.3005
R4135 VGND.n81 VGND.n80 9.3005
R4136 VGND.n83 VGND.n82 9.3005
R4137 VGND.n2899 VGND.n2898 9.3005
R4138 VGND.n2901 VGND.n60 9.3005
R4139 VGND.n2897 VGND.n2896 9.3005
R4140 VGND.n2936 VGND.n2935 9.3005
R4141 VGND.n2917 VGND.n2913 9.3005
R4142 VGND.n2919 VGND.n2918 9.3005
R4143 VGND.n2921 VGND.n2910 9.3005
R4144 VGND.n2923 VGND.n2922 9.3005
R4145 VGND.n2924 VGND.n2909 9.3005
R4146 VGND.n2926 VGND.n2925 9.3005
R4147 VGND.n2927 VGND.n2908 9.3005
R4148 VGND.n2929 VGND.n2928 9.3005
R4149 VGND.n2932 VGND.n2931 9.3005
R4150 VGND.n2933 VGND.n2905 9.3005
R4151 VGND.n2930 VGND.n2907 9.3005
R4152 VGND.n45 VGND.n44 9.3005
R4153 VGND.n46 VGND.n38 9.3005
R4154 VGND.n49 VGND.n48 9.3005
R4155 VGND.n50 VGND.n37 9.3005
R4156 VGND.n52 VGND.n51 9.3005
R4157 VGND.n53 VGND.n36 9.3005
R4158 VGND.n55 VGND.n54 9.3005
R4159 VGND.n56 VGND.n35 9.3005
R4160 VGND.n2945 VGND.n57 9.3005
R4161 VGND.n2944 VGND.n2943 9.3005
R4162 VGND.n2942 VGND.n58 9.3005
R4163 VGND.n2958 VGND.n2957 9.3005
R4164 VGND.n2959 VGND.n2951 9.3005
R4165 VGND.n2962 VGND.n2961 9.3005
R4166 VGND.n2963 VGND.n2950 9.3005
R4167 VGND.n2965 VGND.n2964 9.3005
R4168 VGND.n2966 VGND.n2949 9.3005
R4169 VGND.n2968 VGND.n2967 9.3005
R4170 VGND.n2969 VGND.n2948 9.3005
R4171 VGND.n2977 VGND.n2970 9.3005
R4172 VGND.n2976 VGND.n2975 9.3005
R4173 VGND.n2974 VGND.n2971 9.3005
R4174 VGND.n100 VGND.n92 8.28285
R4175 VGND.n2844 VGND.n2836 8.28285
R4176 VGND.n2876 VGND.n2868 8.28285
R4177 VGND.n2697 VGND.n235 7.9105
R4178 VGND.n2699 VGND.n2698 7.9105
R4179 VGND.n2804 VGND.n189 7.9105
R4180 VGND.n2803 VGND.n190 7.9105
R4181 VGND.n2798 VGND.n195 7.9105
R4182 VGND.n2797 VGND.n196 7.9105
R4183 VGND.n2792 VGND.n201 7.9105
R4184 VGND.n2791 VGND.n202 7.9105
R4185 VGND.n2786 VGND.n207 7.9105
R4186 VGND.n2785 VGND.n208 7.9105
R4187 VGND.n2780 VGND.n213 7.9105
R4188 VGND.n2779 VGND.n214 7.9105
R4189 VGND.n2774 VGND.n219 7.9105
R4190 VGND.n2773 VGND.n220 7.9105
R4191 VGND.n2768 VGND.n2767 7.9105
R4192 VGND.n2986 VGND.n2985 7.9105
R4193 VGND.n2517 VGND.n2516 7.9105
R4194 VGND.n2808 VGND.n185 7.9105
R4195 VGND.n2807 VGND.n186 7.9105
R4196 VGND.n2504 VGND.n2503 7.9105
R4197 VGND.n2502 VGND.n248 7.9105
R4198 VGND.n2501 VGND.n249 7.9105
R4199 VGND.n2500 VGND.n250 7.9105
R4200 VGND.n2499 VGND.n251 7.9105
R4201 VGND.n2498 VGND.n252 7.9105
R4202 VGND.n2497 VGND.n253 7.9105
R4203 VGND.n2496 VGND.n254 7.9105
R4204 VGND.n2495 VGND.n255 7.9105
R4205 VGND.n2494 VGND.n256 7.9105
R4206 VGND.n2493 VGND.n257 7.9105
R4207 VGND.n2492 VGND.n258 7.9105
R4208 VGND.n2491 VGND.n2490 7.9105
R4209 VGND.n639 VGND.n180 7.9105
R4210 VGND.n2812 VGND.n2811 7.9105
R4211 VGND.n375 VGND.n374 7.9105
R4212 VGND.n2166 VGND.n2165 7.9105
R4213 VGND.n2175 VGND.n2174 7.9105
R4214 VGND.n2192 VGND.n2191 7.9105
R4215 VGND.n2201 VGND.n2200 7.9105
R4216 VGND.n2218 VGND.n2217 7.9105
R4217 VGND.n2227 VGND.n2226 7.9105
R4218 VGND.n2244 VGND.n2243 7.9105
R4219 VGND.n2253 VGND.n2252 7.9105
R4220 VGND.n2275 VGND.n2274 7.9105
R4221 VGND.n2297 VGND.n328 7.9105
R4222 VGND.n2296 VGND.n329 7.9105
R4223 VGND.n2294 VGND.n2293 7.9105
R4224 VGND.n2430 VGND.n2429 7.9105
R4225 VGND.n1433 VGND.n1420 7.9105
R4226 VGND.n1432 VGND.n1431 7.9105
R4227 VGND.n2153 VGND.n2152 7.9105
R4228 VGND.n2162 VGND.n2161 7.9105
R4229 VGND.n2179 VGND.n2178 7.9105
R4230 VGND.n2188 VGND.n2187 7.9105
R4231 VGND.n2205 VGND.n2204 7.9105
R4232 VGND.n2214 VGND.n2213 7.9105
R4233 VGND.n2231 VGND.n2230 7.9105
R4234 VGND.n2240 VGND.n2239 7.9105
R4235 VGND.n2257 VGND.n2256 7.9105
R4236 VGND.n2271 VGND.n2270 7.9105
R4237 VGND.n2300 VGND.n327 7.9105
R4238 VGND.n2302 VGND.n2301 7.9105
R4239 VGND.n2314 VGND.n324 7.9105
R4240 VGND.n2313 VGND.n2312 7.9105
R4241 VGND.n1437 VGND.n1436 7.9105
R4242 VGND.n1496 VGND.n1495 7.9105
R4243 VGND.n2149 VGND.n381 7.9105
R4244 VGND.n2148 VGND.n382 7.9105
R4245 VGND.n2147 VGND.n383 7.9105
R4246 VGND.n2146 VGND.n384 7.9105
R4247 VGND.n2145 VGND.n385 7.9105
R4248 VGND.n2144 VGND.n386 7.9105
R4249 VGND.n2143 VGND.n387 7.9105
R4250 VGND.n2142 VGND.n388 7.9105
R4251 VGND.n2141 VGND.n389 7.9105
R4252 VGND.n2140 VGND.n390 7.9105
R4253 VGND.n2139 VGND.n2138 7.9105
R4254 VGND.n2318 VGND.n321 7.9105
R4255 VGND.n2317 VGND.n322 7.9105
R4256 VGND.n2126 VGND.n2125 7.9105
R4257 VGND.n1414 VGND.n617 7.9105
R4258 VGND.n1500 VGND.n1499 7.9105
R4259 VGND.n630 VGND.n629 7.9105
R4260 VGND.n1992 VGND.n1991 7.9105
R4261 VGND.n2001 VGND.n2000 7.9105
R4262 VGND.n2018 VGND.n2017 7.9105
R4263 VGND.n2027 VGND.n2026 7.9105
R4264 VGND.n2044 VGND.n2043 7.9105
R4265 VGND.n2053 VGND.n2052 7.9105
R4266 VGND.n2070 VGND.n2069 7.9105
R4267 VGND.n2079 VGND.n2078 7.9105
R4268 VGND.n2101 VGND.n2100 7.9105
R4269 VGND.n2322 VGND.n318 7.9105
R4270 VGND.n2321 VGND.n319 7.9105
R4271 VGND.n399 VGND.n398 7.9105
R4272 VGND.n2122 VGND.n2121 7.9105
R4273 VGND.n1412 VGND.n644 7.9105
R4274 VGND.n656 VGND.n655 7.9105
R4275 VGND.n1979 VGND.n1978 7.9105
R4276 VGND.n1988 VGND.n1987 7.9105
R4277 VGND.n2005 VGND.n2004 7.9105
R4278 VGND.n2014 VGND.n2013 7.9105
R4279 VGND.n2031 VGND.n2030 7.9105
R4280 VGND.n2040 VGND.n2039 7.9105
R4281 VGND.n2057 VGND.n2056 7.9105
R4282 VGND.n2066 VGND.n2065 7.9105
R4283 VGND.n2083 VGND.n2082 7.9105
R4284 VGND.n2097 VGND.n2096 7.9105
R4285 VGND.n2325 VGND.n316 7.9105
R4286 VGND.n2327 VGND.n2326 7.9105
R4287 VGND.n2339 VGND.n312 7.9105
R4288 VGND.n2338 VGND.n2337 7.9105
R4289 VGND.n1409 VGND.n660 7.9105
R4290 VGND.n1408 VGND.n661 7.9105
R4291 VGND.n1975 VGND.n437 7.9105
R4292 VGND.n1974 VGND.n438 7.9105
R4293 VGND.n1973 VGND.n439 7.9105
R4294 VGND.n1972 VGND.n440 7.9105
R4295 VGND.n1971 VGND.n441 7.9105
R4296 VGND.n1970 VGND.n442 7.9105
R4297 VGND.n1969 VGND.n443 7.9105
R4298 VGND.n1968 VGND.n444 7.9105
R4299 VGND.n1967 VGND.n445 7.9105
R4300 VGND.n1966 VGND.n446 7.9105
R4301 VGND.n1965 VGND.n1964 7.9105
R4302 VGND.n2343 VGND.n309 7.9105
R4303 VGND.n2342 VGND.n310 7.9105
R4304 VGND.n1952 VGND.n1951 7.9105
R4305 VGND.n1390 VGND.n1389 7.9105
R4306 VGND.n1405 VGND.n663 7.9105
R4307 VGND.n1404 VGND.n1403 7.9105
R4308 VGND.n1818 VGND.n1817 7.9105
R4309 VGND.n1827 VGND.n1826 7.9105
R4310 VGND.n1844 VGND.n1843 7.9105
R4311 VGND.n1853 VGND.n1852 7.9105
R4312 VGND.n1870 VGND.n1869 7.9105
R4313 VGND.n1879 VGND.n1878 7.9105
R4314 VGND.n1896 VGND.n1895 7.9105
R4315 VGND.n1905 VGND.n1904 7.9105
R4316 VGND.n1927 VGND.n1926 7.9105
R4317 VGND.n2347 VGND.n306 7.9105
R4318 VGND.n2346 VGND.n307 7.9105
R4319 VGND.n455 VGND.n454 7.9105
R4320 VGND.n1948 VGND.n1947 7.9105
R4321 VGND.n1386 VGND.n1372 7.9105
R4322 VGND.n1384 VGND.n1383 7.9105
R4323 VGND.n1805 VGND.n1804 7.9105
R4324 VGND.n1814 VGND.n1813 7.9105
R4325 VGND.n1831 VGND.n1830 7.9105
R4326 VGND.n1840 VGND.n1839 7.9105
R4327 VGND.n1857 VGND.n1856 7.9105
R4328 VGND.n1866 VGND.n1865 7.9105
R4329 VGND.n1883 VGND.n1882 7.9105
R4330 VGND.n1892 VGND.n1891 7.9105
R4331 VGND.n1909 VGND.n1908 7.9105
R4332 VGND.n1923 VGND.n1922 7.9105
R4333 VGND.n2350 VGND.n304 7.9105
R4334 VGND.n2352 VGND.n2351 7.9105
R4335 VGND.n2364 VGND.n300 7.9105
R4336 VGND.n2363 VGND.n2362 7.9105
R4337 VGND.n1368 VGND.n1304 7.9105
R4338 VGND.n1367 VGND.n1365 7.9105
R4339 VGND.n1801 VGND.n493 7.9105
R4340 VGND.n1800 VGND.n494 7.9105
R4341 VGND.n1799 VGND.n495 7.9105
R4342 VGND.n1798 VGND.n496 7.9105
R4343 VGND.n1797 VGND.n497 7.9105
R4344 VGND.n1796 VGND.n498 7.9105
R4345 VGND.n1795 VGND.n499 7.9105
R4346 VGND.n1794 VGND.n500 7.9105
R4347 VGND.n1793 VGND.n501 7.9105
R4348 VGND.n1792 VGND.n502 7.9105
R4349 VGND.n1791 VGND.n1790 7.9105
R4350 VGND.n2368 VGND.n297 7.9105
R4351 VGND.n2367 VGND.n298 7.9105
R4352 VGND.n1778 VGND.n1777 7.9105
R4353 VGND.n1528 VGND.n573 7.9105
R4354 VGND.n1527 VGND.n574 7.9105
R4355 VGND.n1526 VGND.n1525 7.9105
R4356 VGND.n1644 VGND.n1643 7.9105
R4357 VGND.n1653 VGND.n1652 7.9105
R4358 VGND.n1670 VGND.n1669 7.9105
R4359 VGND.n1679 VGND.n1678 7.9105
R4360 VGND.n1696 VGND.n1695 7.9105
R4361 VGND.n1705 VGND.n1704 7.9105
R4362 VGND.n1722 VGND.n1721 7.9105
R4363 VGND.n1731 VGND.n1730 7.9105
R4364 VGND.n1753 VGND.n1752 7.9105
R4365 VGND.n2372 VGND.n294 7.9105
R4366 VGND.n2371 VGND.n295 7.9105
R4367 VGND.n511 VGND.n510 7.9105
R4368 VGND.n1774 VGND.n1773 7.9105
R4369 VGND.n1532 VGND.n1531 7.9105
R4370 VGND.n1541 VGND.n1540 7.9105
R4371 VGND.n1631 VGND.n1630 7.9105
R4372 VGND.n1640 VGND.n1639 7.9105
R4373 VGND.n1657 VGND.n1656 7.9105
R4374 VGND.n1666 VGND.n1665 7.9105
R4375 VGND.n1683 VGND.n1682 7.9105
R4376 VGND.n1692 VGND.n1691 7.9105
R4377 VGND.n1709 VGND.n1708 7.9105
R4378 VGND.n1718 VGND.n1717 7.9105
R4379 VGND.n1735 VGND.n1734 7.9105
R4380 VGND.n1749 VGND.n1748 7.9105
R4381 VGND.n2375 VGND.n291 7.9105
R4382 VGND.n2377 VGND.n2376 7.9105
R4383 VGND.n2389 VGND.n287 7.9105
R4384 VGND.n2388 VGND.n2387 7.9105
R4385 VGND.n1298 VGND.n1297 7.9105
R4386 VGND.n1545 VGND.n1544 7.9105
R4387 VGND.n1627 VGND.n549 7.9105
R4388 VGND.n1626 VGND.n550 7.9105
R4389 VGND.n1625 VGND.n551 7.9105
R4390 VGND.n1624 VGND.n552 7.9105
R4391 VGND.n1623 VGND.n553 7.9105
R4392 VGND.n1622 VGND.n554 7.9105
R4393 VGND.n1621 VGND.n555 7.9105
R4394 VGND.n1620 VGND.n556 7.9105
R4395 VGND.n1619 VGND.n557 7.9105
R4396 VGND.n1618 VGND.n558 7.9105
R4397 VGND.n1617 VGND.n1616 7.9105
R4398 VGND.n2393 VGND.n282 7.9105
R4399 VGND.n2392 VGND.n283 7.9105
R4400 VGND.n1604 VGND.n1603 7.9105
R4401 VGND.n896 VGND.n826 7.9105
R4402 VGND.n895 VGND.n827 7.9105
R4403 VGND.n894 VGND.n893 7.9105
R4404 VGND.n1275 VGND.n688 7.9105
R4405 VGND.n1274 VGND.n689 7.9105
R4406 VGND.n1267 VGND.n694 7.9105
R4407 VGND.n1266 VGND.n695 7.9105
R4408 VGND.n1259 VGND.n700 7.9105
R4409 VGND.n1258 VGND.n701 7.9105
R4410 VGND.n1251 VGND.n706 7.9105
R4411 VGND.n1250 VGND.n707 7.9105
R4412 VGND.n1243 VGND.n712 7.9105
R4413 VGND.n1242 VGND.n713 7.9105
R4414 VGND.n2397 VGND.n2396 7.9105
R4415 VGND.n284 VGND.n279 7.9105
R4416 VGND.n2408 VGND.n2407 7.9105
R4417 VGND.n1117 VGND.n677 7.9105
R4418 VGND.n1285 VGND.n1284 7.9105
R4419 VGND.n1279 VGND.n685 7.9105
R4420 VGND.n1278 VGND.n686 7.9105
R4421 VGND.n1271 VGND.n691 7.9105
R4422 VGND.n1270 VGND.n692 7.9105
R4423 VGND.n1263 VGND.n697 7.9105
R4424 VGND.n1262 VGND.n698 7.9105
R4425 VGND.n1255 VGND.n703 7.9105
R4426 VGND.n1254 VGND.n704 7.9105
R4427 VGND.n1247 VGND.n709 7.9105
R4428 VGND.n1246 VGND.n710 7.9105
R4429 VGND.n1239 VGND.n715 7.9105
R4430 VGND.n1238 VGND.n716 7.9105
R4431 VGND.n1237 VGND.n783 7.9105
R4432 VGND.n2412 VGND.n2411 7.9105
R4433 VGND.n133 VGND.n130 7.90638
R4434 VGND.n126 VGND.n125 7.90638
R4435 VGND.n601 VGND.n598 7.90638
R4436 VGND.n594 VGND.n593 7.90638
R4437 VGND.n976 VGND.n971 7.90638
R4438 VGND.n975 VGND.n974 7.90638
R4439 VGND.n163 VGND.n160 7.90638
R4440 VGND.n156 VGND.n155 7.90638
R4441 VGND.n1098 VGND.n1094 7.4049
R4442 VGND.n1071 VGND.n1065 7.4049
R4443 VGND.n1009 VGND.n1003 7.4049
R4444 VGND.n1040 VGND.n1034 7.4049
R4445 VGND VGND.n149 7.12482
R4446 VGND.n97 VGND.n96 6.85473
R4447 VGND.n2841 VGND.n2840 6.85473
R4448 VGND.n2873 VGND.n2872 6.85473
R4449 VGND.n19 VGND.n18 6.77697
R4450 VGND.n48 VGND.n47 6.77697
R4451 VGND.n2921 VGND.n2920 6.77697
R4452 VGND.n2961 VGND.n2960 6.77697
R4453 VGND.n3005 VGND.n3004 6.4005
R4454 VGND.n969 VGND.n968 5.27109
R4455 VGND.n73 VGND.n67 5.27109
R4456 VGND.n2582 VGND.n2581 4.5005
R4457 VGND.n2640 VGND.n223 4.5005
R4458 VGND.n2585 VGND.n2584 4.5005
R4459 VGND.n2649 VGND.n222 4.5005
R4460 VGND.n2588 VGND.n2587 4.5005
R4461 VGND.n2637 VGND.n217 4.5005
R4462 VGND.n2591 VGND.n2590 4.5005
R4463 VGND.n2656 VGND.n216 4.5005
R4464 VGND.n2594 VGND.n2593 4.5005
R4465 VGND.n2634 VGND.n211 4.5005
R4466 VGND.n2597 VGND.n2596 4.5005
R4467 VGND.n2663 VGND.n210 4.5005
R4468 VGND.n2600 VGND.n2599 4.5005
R4469 VGND.n2631 VGND.n205 4.5005
R4470 VGND.n2603 VGND.n2602 4.5005
R4471 VGND.n2670 VGND.n204 4.5005
R4472 VGND.n2606 VGND.n2605 4.5005
R4473 VGND.n2628 VGND.n199 4.5005
R4474 VGND.n2609 VGND.n2608 4.5005
R4475 VGND.n2677 VGND.n198 4.5005
R4476 VGND.n2612 VGND.n2611 4.5005
R4477 VGND.n2625 VGND.n193 4.5005
R4478 VGND.n2615 VGND.n2614 4.5005
R4479 VGND.n2684 VGND.n192 4.5005
R4480 VGND.n2618 VGND.n2575 4.5005
R4481 VGND.n2622 VGND.n2619 4.5005
R4482 VGND.n2569 VGND.n2568 4.5005
R4483 VGND.n2693 VGND.n2692 4.5005
R4484 VGND.n2523 VGND.n2522 4.5005
R4485 VGND.n2526 VGND.n2525 4.5005
R4486 VGND.n2529 VGND.n2528 4.5005
R4487 VGND.n2532 VGND.n2531 4.5005
R4488 VGND.n2535 VGND.n2534 4.5005
R4489 VGND.n2538 VGND.n2537 4.5005
R4490 VGND.n2541 VGND.n2540 4.5005
R4491 VGND.n2544 VGND.n2543 4.5005
R4492 VGND.n2547 VGND.n2546 4.5005
R4493 VGND.n2550 VGND.n2549 4.5005
R4494 VGND.n2553 VGND.n2552 4.5005
R4495 VGND.n2556 VGND.n2555 4.5005
R4496 VGND.n2559 VGND.n2558 4.5005
R4497 VGND.n2562 VGND.n2561 4.5005
R4498 VGND.n2565 VGND.n2564 4.5005
R4499 VGND.n2574 VGND.n2567 4.5005
R4500 VGND.n2577 VGND.n2576 4.5005
R4501 VGND.n2580 VGND.n2579 4.5005
R4502 VGND.n2642 VGND.n30 4.5005
R4503 VGND.n820 VGND.n819 4.5005
R4504 VGND.n817 VGND.n816 4.5005
R4505 VGND.n1137 VGND.n1136 4.5005
R4506 VGND.n1149 VGND.n807 4.5005
R4507 VGND.n1156 VGND.n805 4.5005
R4508 VGND.n1153 VGND.n1151 4.5005
R4509 VGND.n1169 VGND.n1168 4.5005
R4510 VGND.n1181 VGND.n799 4.5005
R4511 VGND.n1188 VGND.n797 4.5005
R4512 VGND.n1185 VGND.n1183 4.5005
R4513 VGND.n1201 VGND.n1200 4.5005
R4514 VGND.n1213 VGND.n791 4.5005
R4515 VGND.n1219 VGND.n789 4.5005
R4516 VGND.n1216 VGND.n1215 4.5005
R4517 VGND.n786 VGND.n785 4.5005
R4518 VGND.n823 VGND.n822 4.5005
R4519 VGND.n1121 VGND.n1120 4.5005
R4520 VGND.n1126 VGND.n680 4.5005
R4521 VGND.n812 VGND.n681 4.5005
R4522 VGND.n1139 VGND.n1138 4.5005
R4523 VGND.n1148 VGND.n1147 4.5005
R4524 VGND.n1158 VGND.n1157 4.5005
R4525 VGND.n1152 VGND.n804 4.5005
R4526 VGND.n1171 VGND.n1170 4.5005
R4527 VGND.n1180 VGND.n1179 4.5005
R4528 VGND.n1190 VGND.n1189 4.5005
R4529 VGND.n1184 VGND.n796 4.5005
R4530 VGND.n1203 VGND.n1202 4.5005
R4531 VGND.n1212 VGND.n1211 4.5005
R4532 VGND.n1222 VGND.n1221 4.5005
R4533 VGND.n788 VGND.n784 4.5005
R4534 VGND.n1233 VGND.n1232 4.5005
R4535 VGND.n1113 VGND.n1112 4.41365
R4536 VGND VGND.n2990 4.35375
R4537 VGND.n1090 VGND.n1089 4.05427
R4538 VGND.n583 VGND.n0 4.05427
R4539 VGND.n998 VGND.n997 4.05427
R4540 VGND.n1029 VGND.n1028 4.05427
R4541 VGND.n1060 VGND.n1059 4.05427
R4542 VGND VGND.n59 3.99438
R4543 VGND.n2904 VGND 3.99438
R4544 VGND.n2937 VGND 3.99438
R4545 VGND VGND.n2938 3.99437
R4546 VGND VGND.n28 3.99437
R4547 VGND.n1234 VGND.n274 3.77268
R4548 VGND.n2988 VGND.n2987 3.77268
R4549 VGND.n1119 VGND.n1118 3.77268
R4550 VGND.n2696 VGND.n2695 3.77268
R4551 VGND.n1281 VGND.n1280 3.77268
R4552 VGND.n2805 VGND.n188 3.77268
R4553 VGND.n1277 VGND.n687 3.77268
R4554 VGND.n2802 VGND.n2801 3.77268
R4555 VGND.n1272 VGND.n690 3.77268
R4556 VGND.n2800 VGND.n2799 3.77268
R4557 VGND.n1269 VGND.n693 3.77268
R4558 VGND.n2796 VGND.n2795 3.77268
R4559 VGND.n1264 VGND.n696 3.77268
R4560 VGND.n2794 VGND.n2793 3.77268
R4561 VGND.n1261 VGND.n699 3.77268
R4562 VGND.n2790 VGND.n2789 3.77268
R4563 VGND.n1256 VGND.n702 3.77268
R4564 VGND.n2788 VGND.n2787 3.77268
R4565 VGND.n1253 VGND.n705 3.77268
R4566 VGND.n2784 VGND.n2783 3.77268
R4567 VGND.n1248 VGND.n708 3.77268
R4568 VGND.n2782 VGND.n2781 3.77268
R4569 VGND.n1245 VGND.n711 3.77268
R4570 VGND.n2778 VGND.n2777 3.77268
R4571 VGND.n1240 VGND.n714 3.77268
R4572 VGND.n2776 VGND.n2775 3.77268
R4573 VGND.n1220 VGND.n280 3.77268
R4574 VGND.n2772 VGND.n2771 3.77268
R4575 VGND.n1236 VGND.n1235 3.77268
R4576 VGND.n2770 VGND.n2769 3.77268
R4577 VGND.n1283 VGND.n1282 3.77268
R4578 VGND.n2694 VGND.n184 3.77268
R4579 VGND.n2578 VGND.n2577 3.75914
R4580 VGND.n2583 VGND.n2580 3.75914
R4581 VGND.n1217 VGND.n786 3.75914
R4582 VGND.n823 VGND.n821 3.75914
R4583 VGND.n2578 VGND.n2569 3.4105
R4584 VGND.n2618 VGND.n2617 3.4105
R4585 VGND.n2616 VGND.n2615 3.4105
R4586 VGND.n2613 VGND.n2612 3.4105
R4587 VGND.n2610 VGND.n2609 3.4105
R4588 VGND.n2607 VGND.n2606 3.4105
R4589 VGND.n2604 VGND.n2603 3.4105
R4590 VGND.n2601 VGND.n2600 3.4105
R4591 VGND.n2598 VGND.n2597 3.4105
R4592 VGND.n2595 VGND.n2594 3.4105
R4593 VGND.n2592 VGND.n2591 3.4105
R4594 VGND.n2589 VGND.n2588 3.4105
R4595 VGND.n2586 VGND.n2585 3.4105
R4596 VGND.n2583 VGND.n2582 3.4105
R4597 VGND.n2988 VGND.n30 3.4105
R4598 VGND.n2770 VGND.n223 3.4105
R4599 VGND.n2771 VGND.n222 3.4105
R4600 VGND.n2776 VGND.n217 3.4105
R4601 VGND.n2777 VGND.n216 3.4105
R4602 VGND.n2782 VGND.n211 3.4105
R4603 VGND.n2783 VGND.n210 3.4105
R4604 VGND.n2788 VGND.n205 3.4105
R4605 VGND.n2789 VGND.n204 3.4105
R4606 VGND.n2794 VGND.n199 3.4105
R4607 VGND.n2795 VGND.n198 3.4105
R4608 VGND.n2800 VGND.n193 3.4105
R4609 VGND.n2801 VGND.n192 3.4105
R4610 VGND.n2619 VGND.n188 3.4105
R4611 VGND.n2694 VGND.n2693 3.4105
R4612 VGND.n2695 VGND.n2567 3.4105
R4613 VGND.n2987 VGND.n2986 3.4105
R4614 VGND.n2697 VGND.n2696 3.4105
R4615 VGND.n2517 VGND.n236 3.4105
R4616 VGND.n2491 VGND.n31 3.4105
R4617 VGND.n2807 VGND.n2806 3.4105
R4618 VGND.n2805 VGND.n2804 3.4105
R4619 VGND.n375 VGND.n187 3.4105
R4620 VGND.n640 VGND.n639 3.4105
R4621 VGND.n2430 VGND.n260 3.4105
R4622 VGND.n2165 VGND.n2164 3.4105
R4623 VGND.n2503 VGND.n191 3.4105
R4624 VGND.n2803 VGND.n2802 3.4105
R4625 VGND.n2163 VGND.n2162 3.4105
R4626 VGND.n2152 VGND.n2151 3.4105
R4627 VGND.n1434 VGND.n1433 3.4105
R4628 VGND.n2313 VGND.n325 3.4105
R4629 VGND.n2178 VGND.n2177 3.4105
R4630 VGND.n2176 VGND.n2175 3.4105
R4631 VGND.n2502 VGND.n194 3.4105
R4632 VGND.n2799 VGND.n2798 3.4105
R4633 VGND.n2147 VGND.n361 3.4105
R4634 VGND.n2148 VGND.n376 3.4105
R4635 VGND.n2150 VGND.n2149 3.4105
R4636 VGND.n1436 VGND.n1435 3.4105
R4637 VGND.n2125 VGND.n395 3.4105
R4638 VGND.n2146 VGND.n357 3.4105
R4639 VGND.n2189 VGND.n2188 3.4105
R4640 VGND.n2191 VGND.n2190 3.4105
R4641 VGND.n2501 VGND.n197 3.4105
R4642 VGND.n2797 VGND.n2796 3.4105
R4643 VGND.n2017 VGND.n2016 3.4105
R4644 VGND.n2002 VGND.n2001 3.4105
R4645 VGND.n1991 VGND.n1990 3.4105
R4646 VGND.n630 VGND.n380 3.4105
R4647 VGND.n1414 VGND.n638 3.4105
R4648 VGND.n2122 VGND.n396 3.4105
R4649 VGND.n2028 VGND.n2027 3.4105
R4650 VGND.n2145 VGND.n353 3.4105
R4651 VGND.n2204 VGND.n2203 3.4105
R4652 VGND.n2202 VGND.n2201 3.4105
R4653 VGND.n2500 VGND.n200 3.4105
R4654 VGND.n2793 VGND.n2792 3.4105
R4655 VGND.n2030 VGND.n2029 3.4105
R4656 VGND.n2015 VGND.n2014 3.4105
R4657 VGND.n2004 VGND.n2003 3.4105
R4658 VGND.n1989 VGND.n1988 3.4105
R4659 VGND.n1978 VGND.n1977 3.4105
R4660 VGND.n1412 VGND.n1411 3.4105
R4661 VGND.n2338 VGND.n313 3.4105
R4662 VGND.n2041 VGND.n2040 3.4105
R4663 VGND.n2043 VGND.n2042 3.4105
R4664 VGND.n2144 VGND.n349 3.4105
R4665 VGND.n2215 VGND.n2214 3.4105
R4666 VGND.n2217 VGND.n2216 3.4105
R4667 VGND.n2499 VGND.n203 3.4105
R4668 VGND.n2791 VGND.n2790 3.4105
R4669 VGND.n1970 VGND.n416 3.4105
R4670 VGND.n1971 VGND.n420 3.4105
R4671 VGND.n1972 VGND.n424 3.4105
R4672 VGND.n1973 VGND.n428 3.4105
R4673 VGND.n1974 VGND.n432 3.4105
R4674 VGND.n1976 VGND.n1975 3.4105
R4675 VGND.n1410 VGND.n1409 3.4105
R4676 VGND.n1951 VGND.n451 3.4105
R4677 VGND.n1969 VGND.n412 3.4105
R4678 VGND.n2056 VGND.n2055 3.4105
R4679 VGND.n2054 VGND.n2053 3.4105
R4680 VGND.n2143 VGND.n345 3.4105
R4681 VGND.n2230 VGND.n2229 3.4105
R4682 VGND.n2228 VGND.n2227 3.4105
R4683 VGND.n2498 VGND.n206 3.4105
R4684 VGND.n2787 VGND.n2786 3.4105
R4685 VGND.n1880 VGND.n1879 3.4105
R4686 VGND.n1869 VGND.n1868 3.4105
R4687 VGND.n1854 VGND.n1853 3.4105
R4688 VGND.n1843 VGND.n1842 3.4105
R4689 VGND.n1828 VGND.n1827 3.4105
R4690 VGND.n1817 VGND.n1816 3.4105
R4691 VGND.n1404 VGND.n436 3.4105
R4692 VGND.n1389 VGND.n657 3.4105
R4693 VGND.n1948 VGND.n452 3.4105
R4694 VGND.n1895 VGND.n1894 3.4105
R4695 VGND.n1968 VGND.n408 3.4105
R4696 VGND.n2067 VGND.n2066 3.4105
R4697 VGND.n2069 VGND.n2068 3.4105
R4698 VGND.n2142 VGND.n341 3.4105
R4699 VGND.n2241 VGND.n2240 3.4105
R4700 VGND.n2243 VGND.n2242 3.4105
R4701 VGND.n2497 VGND.n209 3.4105
R4702 VGND.n2785 VGND.n2784 3.4105
R4703 VGND.n1893 VGND.n1892 3.4105
R4704 VGND.n1882 VGND.n1881 3.4105
R4705 VGND.n1867 VGND.n1866 3.4105
R4706 VGND.n1856 VGND.n1855 3.4105
R4707 VGND.n1841 VGND.n1840 3.4105
R4708 VGND.n1830 VGND.n1829 3.4105
R4709 VGND.n1815 VGND.n1814 3.4105
R4710 VGND.n1804 VGND.n1803 3.4105
R4711 VGND.n1386 VGND.n1385 3.4105
R4712 VGND.n2363 VGND.n301 3.4105
R4713 VGND.n1908 VGND.n1907 3.4105
R4714 VGND.n1906 VGND.n1905 3.4105
R4715 VGND.n1967 VGND.n404 3.4105
R4716 VGND.n2082 VGND.n2081 3.4105
R4717 VGND.n2080 VGND.n2079 3.4105
R4718 VGND.n2141 VGND.n337 3.4105
R4719 VGND.n2256 VGND.n2255 3.4105
R4720 VGND.n2254 VGND.n2253 3.4105
R4721 VGND.n2496 VGND.n212 3.4105
R4722 VGND.n2781 VGND.n2780 3.4105
R4723 VGND.n1793 VGND.n460 3.4105
R4724 VGND.n1794 VGND.n464 3.4105
R4725 VGND.n1795 VGND.n468 3.4105
R4726 VGND.n1796 VGND.n472 3.4105
R4727 VGND.n1797 VGND.n476 3.4105
R4728 VGND.n1798 VGND.n480 3.4105
R4729 VGND.n1799 VGND.n484 3.4105
R4730 VGND.n1800 VGND.n488 3.4105
R4731 VGND.n1802 VGND.n1801 3.4105
R4732 VGND.n1368 VGND.n570 3.4105
R4733 VGND.n1777 VGND.n507 3.4105
R4734 VGND.n1792 VGND.n456 3.4105
R4735 VGND.n1924 VGND.n1923 3.4105
R4736 VGND.n1926 VGND.n1925 3.4105
R4737 VGND.n1966 VGND.n400 3.4105
R4738 VGND.n2098 VGND.n2097 3.4105
R4739 VGND.n2100 VGND.n2099 3.4105
R4740 VGND.n2140 VGND.n333 3.4105
R4741 VGND.n2272 VGND.n2271 3.4105
R4742 VGND.n2274 VGND.n2273 3.4105
R4743 VGND.n2495 VGND.n215 3.4105
R4744 VGND.n2779 VGND.n2778 3.4105
R4745 VGND.n1752 VGND.n1751 3.4105
R4746 VGND.n1732 VGND.n1731 3.4105
R4747 VGND.n1721 VGND.n1720 3.4105
R4748 VGND.n1706 VGND.n1705 3.4105
R4749 VGND.n1695 VGND.n1694 3.4105
R4750 VGND.n1680 VGND.n1679 3.4105
R4751 VGND.n1669 VGND.n1668 3.4105
R4752 VGND.n1654 VGND.n1653 3.4105
R4753 VGND.n1643 VGND.n1642 3.4105
R4754 VGND.n1526 VGND.n492 3.4105
R4755 VGND.n1529 VGND.n1528 3.4105
R4756 VGND.n1774 VGND.n508 3.4105
R4757 VGND.n2373 VGND.n2372 3.4105
R4758 VGND.n1791 VGND.n293 3.4105
R4759 VGND.n2350 VGND.n2349 3.4105
R4760 VGND.n2348 VGND.n2347 3.4105
R4761 VGND.n1965 VGND.n305 3.4105
R4762 VGND.n2325 VGND.n2324 3.4105
R4763 VGND.n2323 VGND.n2322 3.4105
R4764 VGND.n2139 VGND.n317 3.4105
R4765 VGND.n2300 VGND.n2299 3.4105
R4766 VGND.n2298 VGND.n2297 3.4105
R4767 VGND.n2494 VGND.n218 3.4105
R4768 VGND.n2775 VGND.n2774 3.4105
R4769 VGND.n2375 VGND.n2374 3.4105
R4770 VGND.n1750 VGND.n1749 3.4105
R4771 VGND.n1734 VGND.n1733 3.4105
R4772 VGND.n1719 VGND.n1718 3.4105
R4773 VGND.n1708 VGND.n1707 3.4105
R4774 VGND.n1693 VGND.n1692 3.4105
R4775 VGND.n1682 VGND.n1681 3.4105
R4776 VGND.n1667 VGND.n1666 3.4105
R4777 VGND.n1656 VGND.n1655 3.4105
R4778 VGND.n1641 VGND.n1640 3.4105
R4779 VGND.n1630 VGND.n1629 3.4105
R4780 VGND.n1531 VGND.n1530 3.4105
R4781 VGND.n2388 VGND.n288 3.4105
R4782 VGND.n2376 VGND.n281 3.4105
R4783 VGND.n2371 VGND.n2370 3.4105
R4784 VGND.n2369 VGND.n2368 3.4105
R4785 VGND.n2351 VGND.n296 3.4105
R4786 VGND.n2346 VGND.n2345 3.4105
R4787 VGND.n2344 VGND.n2343 3.4105
R4788 VGND.n2326 VGND.n308 3.4105
R4789 VGND.n2321 VGND.n2320 3.4105
R4790 VGND.n2319 VGND.n2318 3.4105
R4791 VGND.n2301 VGND.n320 3.4105
R4792 VGND.n2296 VGND.n2295 3.4105
R4793 VGND.n2493 VGND.n221 3.4105
R4794 VGND.n2773 VGND.n2772 3.4105
R4795 VGND.n2394 VGND.n2393 3.4105
R4796 VGND.n1617 VGND.n292 3.4105
R4797 VGND.n1618 VGND.n512 3.4105
R4798 VGND.n1619 VGND.n516 3.4105
R4799 VGND.n1620 VGND.n520 3.4105
R4800 VGND.n1621 VGND.n524 3.4105
R4801 VGND.n1622 VGND.n528 3.4105
R4802 VGND.n1623 VGND.n532 3.4105
R4803 VGND.n1624 VGND.n536 3.4105
R4804 VGND.n1625 VGND.n540 3.4105
R4805 VGND.n1626 VGND.n544 3.4105
R4806 VGND.n1628 VGND.n1627 3.4105
R4807 VGND.n1298 VGND.n569 3.4105
R4808 VGND.n1603 VGND.n1602 3.4105
R4809 VGND.n2392 VGND.n2391 3.4105
R4810 VGND.n2390 VGND.n2389 3.4105
R4811 VGND.n510 VGND.n286 3.4105
R4812 VGND.n2367 VGND.n2366 3.4105
R4813 VGND.n2365 VGND.n2364 3.4105
R4814 VGND.n454 VGND.n299 3.4105
R4815 VGND.n2342 VGND.n2341 3.4105
R4816 VGND.n2340 VGND.n2339 3.4105
R4817 VGND.n398 VGND.n311 3.4105
R4818 VGND.n2317 VGND.n2316 3.4105
R4819 VGND.n2315 VGND.n2314 3.4105
R4820 VGND.n2294 VGND.n323 3.4105
R4821 VGND.n2492 VGND.n224 3.4105
R4822 VGND.n2769 VGND.n2768 3.4105
R4823 VGND.n285 VGND.n284 3.4105
R4824 VGND.n2396 VGND.n2395 3.4105
R4825 VGND.n1242 VGND.n1241 3.4105
R4826 VGND.n1244 VGND.n1243 3.4105
R4827 VGND.n1250 VGND.n1249 3.4105
R4828 VGND.n1252 VGND.n1251 3.4105
R4829 VGND.n1258 VGND.n1257 3.4105
R4830 VGND.n1260 VGND.n1259 3.4105
R4831 VGND.n1266 VGND.n1265 3.4105
R4832 VGND.n1268 VGND.n1267 3.4105
R4833 VGND.n1274 VGND.n1273 3.4105
R4834 VGND.n1276 VGND.n1275 3.4105
R4835 VGND.n894 VGND.n548 3.4105
R4836 VGND.n897 VGND.n896 3.4105
R4837 VGND.n2408 VGND.n277 3.4105
R4838 VGND.n895 VGND.n562 3.4105
R4839 VGND.n1544 VGND.n1543 3.4105
R4840 VGND.n1542 VGND.n1541 3.4105
R4841 VGND.n1527 VGND.n563 3.4105
R4842 VGND.n1367 VGND.n1366 3.4105
R4843 VGND.n1384 VGND.n662 3.4105
R4844 VGND.n1406 VGND.n1405 3.4105
R4845 VGND.n1408 VGND.n1407 3.4105
R4846 VGND.n656 VGND.n631 3.4105
R4847 VGND.n1499 VGND.n1498 3.4105
R4848 VGND.n1497 VGND.n1496 3.4105
R4849 VGND.n1432 VGND.n183 3.4105
R4850 VGND.n2811 VGND.n2810 3.4105
R4851 VGND.n2809 VGND.n2808 3.4105
R4852 VGND.n2698 VGND.n184 3.4105
R4853 VGND.n1235 VGND.n784 3.4105
R4854 VGND.n1221 VGND.n1220 3.4105
R4855 VGND.n1212 VGND.n714 3.4105
R4856 VGND.n1202 VGND.n711 3.4105
R4857 VGND.n1184 VGND.n708 3.4105
R4858 VGND.n1189 VGND.n705 3.4105
R4859 VGND.n1180 VGND.n702 3.4105
R4860 VGND.n1170 VGND.n699 3.4105
R4861 VGND.n1152 VGND.n696 3.4105
R4862 VGND.n1157 VGND.n693 3.4105
R4863 VGND.n1148 VGND.n690 3.4105
R4864 VGND.n1138 VGND.n687 3.4105
R4865 VGND.n1281 VGND.n681 3.4105
R4866 VGND.n1282 VGND.n680 3.4105
R4867 VGND.n1234 VGND.n1233 3.4105
R4868 VGND.n1217 VGND.n1216 3.4105
R4869 VGND.n1219 VGND.n1218 3.4105
R4870 VGND.n1214 VGND.n1213 3.4105
R4871 VGND.n1201 VGND.n790 3.4105
R4872 VGND.n1186 VGND.n1185 3.4105
R4873 VGND.n1188 VGND.n1187 3.4105
R4874 VGND.n1182 VGND.n1181 3.4105
R4875 VGND.n1169 VGND.n798 3.4105
R4876 VGND.n1154 VGND.n1153 3.4105
R4877 VGND.n1156 VGND.n1155 3.4105
R4878 VGND.n1150 VGND.n1149 3.4105
R4879 VGND.n1137 VGND.n806 3.4105
R4880 VGND.n818 VGND.n817 3.4105
R4881 VGND.n821 VGND.n820 3.4105
R4882 VGND.n1120 VGND.n1119 3.4105
R4883 VGND.n1237 VGND.n1236 3.4105
R4884 VGND.n1238 VGND.n280 3.4105
R4885 VGND.n1240 VGND.n1239 3.4105
R4886 VGND.n1246 VGND.n1245 3.4105
R4887 VGND.n1248 VGND.n1247 3.4105
R4888 VGND.n1254 VGND.n1253 3.4105
R4889 VGND.n1256 VGND.n1255 3.4105
R4890 VGND.n1262 VGND.n1261 3.4105
R4891 VGND.n1264 VGND.n1263 3.4105
R4892 VGND.n1270 VGND.n1269 3.4105
R4893 VGND.n1272 VGND.n1271 3.4105
R4894 VGND.n1278 VGND.n1277 3.4105
R4895 VGND.n1280 VGND.n1279 3.4105
R4896 VGND.n1284 VGND.n1283 3.4105
R4897 VGND.n1118 VGND.n1117 3.4105
R4898 VGND.n2411 VGND.n274 3.4105
R4899 VGND.n980 VGND.n969 3.01226
R4900 VGND.n74 VGND.n73 3.01226
R4901 VGND.n964 VGND.n899 2.63579
R4902 VGND.n2523 VGND 2.51836
R4903 VGND.n2526 VGND 2.51836
R4904 VGND.n2529 VGND 2.51836
R4905 VGND.n2532 VGND 2.51836
R4906 VGND.n2535 VGND 2.51836
R4907 VGND.n2538 VGND 2.51836
R4908 VGND.n2541 VGND 2.51836
R4909 VGND.n2544 VGND 2.51836
R4910 VGND.n2547 VGND 2.51836
R4911 VGND.n2550 VGND 2.51836
R4912 VGND.n2553 VGND 2.51836
R4913 VGND.n2556 VGND 2.51836
R4914 VGND.n2559 VGND 2.51836
R4915 VGND.n2562 VGND 2.51836
R4916 VGND.n2565 VGND 2.51836
R4917 VGND.n985 VGND.n984 2.25932
R4918 VGND.n105 VGND.n104 2.25932
R4919 VGND.n2849 VGND.n2848 2.25932
R4920 VGND.n2881 VGND.n2880 2.25932
R4921 VGND.n83 VGND.n62 2.25932
R4922 VGND.n79 VGND.n78 2.25932
R4923 VGND.n135 VGND.n123 1.88285
R4924 VGND.n603 VGND.n591 1.88285
R4925 VGND.n165 VGND.n153 1.88285
R4926 VGND.n2566 VGND 1.79514
R4927 VGND.n1114 VGND.n275 1.75987
R4928 VGND.n2566 VGND 1.57193
R4929 VGND.n2989 VGND.n2988 1.54254
R4930 VGND.n2986 VGND.n29 1.54254
R4931 VGND.n2491 VGND.n2432 1.54254
R4932 VGND.n2431 VGND.n2430 1.54254
R4933 VGND.n2313 VGND.n259 1.54254
R4934 VGND.n2125 VGND.n2124 1.54254
R4935 VGND.n2123 VGND.n2122 1.54254
R4936 VGND.n2338 VGND.n314 1.54254
R4937 VGND.n1951 VGND.n1950 1.54254
R4938 VGND.n1949 VGND.n1948 1.54254
R4939 VGND.n2363 VGND.n302 1.54254
R4940 VGND.n1777 VGND.n1776 1.54254
R4941 VGND.n1775 VGND.n1774 1.54254
R4942 VGND.n2388 VGND.n289 1.54254
R4943 VGND.n1603 VGND.n276 1.54254
R4944 VGND.n2409 VGND.n2408 1.54254
R4945 VGND.n1234 VGND.n275 1.54254
R4946 VGND.n2411 VGND.n2410 1.54254
R4947 VGND.n992 VGND.n898 1.50638
R4948 VGND.n2900 VGND.n2899 1.50638
R4949 VGND VGND.n2520 1.3946
R4950 VGND.n2519 VGND 1.3946
R4951 VGND.n2518 VGND 1.3946
R4952 VGND VGND.n237 1.3946
R4953 VGND VGND.n1417 1.3946
R4954 VGND.n1416 VGND 1.3946
R4955 VGND.n1415 VGND 1.3946
R4956 VGND.n1413 VGND 1.3946
R4957 VGND VGND.n641 1.3946
R4958 VGND VGND.n1388 1.3946
R4959 VGND.n1387 VGND 1.3946
R4960 VGND.n1369 VGND 1.3946
R4961 VGND.n1301 VGND 1.3946
R4962 VGND.n1300 VGND 1.3946
R4963 VGND.n1299 VGND 1.3946
R4964 VGND VGND.n669 1.3946
R4965 VGND.n1115 VGND 1.3946
R4966 VGND VGND.n1116 1.3946
R4967 VGND.n1114 VGND.n1113 1.04507
R4968 VGND.n2582 VGND.n223 1.00149
R4969 VGND.n2585 VGND.n222 1.00149
R4970 VGND.n2588 VGND.n217 1.00149
R4971 VGND.n2591 VGND.n216 1.00149
R4972 VGND.n2594 VGND.n211 1.00149
R4973 VGND.n2597 VGND.n210 1.00149
R4974 VGND.n2600 VGND.n205 1.00149
R4975 VGND.n2603 VGND.n204 1.00149
R4976 VGND.n2606 VGND.n199 1.00149
R4977 VGND.n2609 VGND.n198 1.00149
R4978 VGND.n2612 VGND.n193 1.00149
R4979 VGND.n2615 VGND.n192 1.00149
R4980 VGND.n2619 VGND.n2618 1.00149
R4981 VGND.n2693 VGND.n2569 1.00149
R4982 VGND.n2580 VGND.n30 1.00149
R4983 VGND.n820 VGND.n680 1.00149
R4984 VGND.n817 VGND.n681 1.00149
R4985 VGND.n1138 VGND.n1137 1.00149
R4986 VGND.n1149 VGND.n1148 1.00149
R4987 VGND.n1157 VGND.n1156 1.00149
R4988 VGND.n1153 VGND.n1152 1.00149
R4989 VGND.n1170 VGND.n1169 1.00149
R4990 VGND.n1181 VGND.n1180 1.00149
R4991 VGND.n1189 VGND.n1188 1.00149
R4992 VGND.n1185 VGND.n1184 1.00149
R4993 VGND.n1202 VGND.n1201 1.00149
R4994 VGND.n1213 VGND.n1212 1.00149
R4995 VGND.n1221 VGND.n1219 1.00149
R4996 VGND.n1216 VGND.n784 1.00149
R4997 VGND.n1233 VGND.n786 1.00149
R4998 VGND.n1120 VGND.n823 1.00149
R4999 VGND.n2577 VGND.n2567 0.973133
R5000 VGND.n2819 VGND.n2 0.9305
R5001 VGND.n97 VGND.n93 0.929432
R5002 VGND.n2841 VGND.n2837 0.929432
R5003 VGND.n2873 VGND.n2869 0.929432
R5004 VGND.n70 VGND.n68 0.929432
R5005 VGND.n59 VGND.n1 0.916608
R5006 VGND VGND.n2523 0.848714
R5007 VGND VGND.n2526 0.848714
R5008 VGND VGND.n2529 0.848714
R5009 VGND VGND.n2532 0.848714
R5010 VGND VGND.n2535 0.848714
R5011 VGND VGND.n2538 0.848714
R5012 VGND VGND.n2541 0.848714
R5013 VGND VGND.n2544 0.848714
R5014 VGND VGND.n2547 0.848714
R5015 VGND VGND.n2550 0.848714
R5016 VGND VGND.n2553 0.848714
R5017 VGND VGND.n2556 0.848714
R5018 VGND VGND.n2559 0.848714
R5019 VGND VGND.n2562 0.848714
R5020 VGND VGND.n2565 0.848714
R5021 VGND.n3006 VGND.n3005 0.7755
R5022 VGND.n3007 VGND.n3006 0.774207
R5023 VGND.n117 VGND.n115 0.753441
R5024 VGND.n16 VGND.n14 0.753441
R5025 VGND.n45 VGND.n43 0.753441
R5026 VGND.n2853 VGND.n2830 0.753441
R5027 VGND.n2916 VGND.n2913 0.753441
R5028 VGND.n2958 VGND.n2956 0.753441
R5029 VGND.n3009 VGND.n3008 0.573119
R5030 VGND VGND.n0 0.542567
R5031 VGND.n3009 VGND.n1 0.507317
R5032 VGND.n2990 VGND.n2989 0.404308
R5033 VGND.n1096 VGND.n1093 0.376971
R5034 VGND.n1068 VGND.n1064 0.376971
R5035 VGND.n992 VGND.n991 0.376971
R5036 VGND.n1006 VGND.n1002 0.376971
R5037 VGND.n1037 VGND.n1033 0.376971
R5038 VGND.n84 VGND.n83 0.376971
R5039 VGND.n2899 VGND.n61 0.376971
R5040 VGND VGND.n3009 0.37415
R5041 VGND.n277 VGND.n274 0.362676
R5042 VGND.n1602 VGND.n277 0.362676
R5043 VGND.n1602 VGND.n288 0.362676
R5044 VGND.n508 VGND.n288 0.362676
R5045 VGND.n508 VGND.n507 0.362676
R5046 VGND.n507 VGND.n301 0.362676
R5047 VGND.n452 VGND.n301 0.362676
R5048 VGND.n452 VGND.n451 0.362676
R5049 VGND.n451 VGND.n313 0.362676
R5050 VGND.n396 VGND.n313 0.362676
R5051 VGND.n396 VGND.n395 0.362676
R5052 VGND.n395 VGND.n325 0.362676
R5053 VGND.n325 VGND.n260 0.362676
R5054 VGND.n260 VGND.n31 0.362676
R5055 VGND.n2987 VGND.n31 0.362676
R5056 VGND.n1118 VGND.n897 0.362676
R5057 VGND.n897 VGND.n569 0.362676
R5058 VGND.n1530 VGND.n569 0.362676
R5059 VGND.n1530 VGND.n1529 0.362676
R5060 VGND.n1529 VGND.n570 0.362676
R5061 VGND.n1385 VGND.n570 0.362676
R5062 VGND.n1385 VGND.n657 0.362676
R5063 VGND.n1410 VGND.n657 0.362676
R5064 VGND.n1411 VGND.n1410 0.362676
R5065 VGND.n1411 VGND.n638 0.362676
R5066 VGND.n1435 VGND.n638 0.362676
R5067 VGND.n1435 VGND.n1434 0.362676
R5068 VGND.n1434 VGND.n640 0.362676
R5069 VGND.n640 VGND.n236 0.362676
R5070 VGND.n2696 VGND.n236 0.362676
R5071 VGND.n1280 VGND.n548 0.362676
R5072 VGND.n1628 VGND.n548 0.362676
R5073 VGND.n1629 VGND.n1628 0.362676
R5074 VGND.n1629 VGND.n492 0.362676
R5075 VGND.n1802 VGND.n492 0.362676
R5076 VGND.n1803 VGND.n1802 0.362676
R5077 VGND.n1803 VGND.n436 0.362676
R5078 VGND.n1976 VGND.n436 0.362676
R5079 VGND.n1977 VGND.n1976 0.362676
R5080 VGND.n1977 VGND.n380 0.362676
R5081 VGND.n2150 VGND.n380 0.362676
R5082 VGND.n2151 VGND.n2150 0.362676
R5083 VGND.n2151 VGND.n187 0.362676
R5084 VGND.n2806 VGND.n187 0.362676
R5085 VGND.n2806 VGND.n2805 0.362676
R5086 VGND.n1277 VGND.n1276 0.362676
R5087 VGND.n1276 VGND.n544 0.362676
R5088 VGND.n1641 VGND.n544 0.362676
R5089 VGND.n1642 VGND.n1641 0.362676
R5090 VGND.n1642 VGND.n488 0.362676
R5091 VGND.n1815 VGND.n488 0.362676
R5092 VGND.n1816 VGND.n1815 0.362676
R5093 VGND.n1816 VGND.n432 0.362676
R5094 VGND.n1989 VGND.n432 0.362676
R5095 VGND.n1990 VGND.n1989 0.362676
R5096 VGND.n1990 VGND.n376 0.362676
R5097 VGND.n2163 VGND.n376 0.362676
R5098 VGND.n2164 VGND.n2163 0.362676
R5099 VGND.n2164 VGND.n191 0.362676
R5100 VGND.n2802 VGND.n191 0.362676
R5101 VGND.n1273 VGND.n1272 0.362676
R5102 VGND.n1273 VGND.n540 0.362676
R5103 VGND.n1655 VGND.n540 0.362676
R5104 VGND.n1655 VGND.n1654 0.362676
R5105 VGND.n1654 VGND.n484 0.362676
R5106 VGND.n1829 VGND.n484 0.362676
R5107 VGND.n1829 VGND.n1828 0.362676
R5108 VGND.n1828 VGND.n428 0.362676
R5109 VGND.n2003 VGND.n428 0.362676
R5110 VGND.n2003 VGND.n2002 0.362676
R5111 VGND.n2002 VGND.n361 0.362676
R5112 VGND.n2177 VGND.n361 0.362676
R5113 VGND.n2177 VGND.n2176 0.362676
R5114 VGND.n2176 VGND.n194 0.362676
R5115 VGND.n2799 VGND.n194 0.362676
R5116 VGND.n1269 VGND.n1268 0.362676
R5117 VGND.n1268 VGND.n536 0.362676
R5118 VGND.n1667 VGND.n536 0.362676
R5119 VGND.n1668 VGND.n1667 0.362676
R5120 VGND.n1668 VGND.n480 0.362676
R5121 VGND.n1841 VGND.n480 0.362676
R5122 VGND.n1842 VGND.n1841 0.362676
R5123 VGND.n1842 VGND.n424 0.362676
R5124 VGND.n2015 VGND.n424 0.362676
R5125 VGND.n2016 VGND.n2015 0.362676
R5126 VGND.n2016 VGND.n357 0.362676
R5127 VGND.n2189 VGND.n357 0.362676
R5128 VGND.n2190 VGND.n2189 0.362676
R5129 VGND.n2190 VGND.n197 0.362676
R5130 VGND.n2796 VGND.n197 0.362676
R5131 VGND.n1265 VGND.n1264 0.362676
R5132 VGND.n1265 VGND.n532 0.362676
R5133 VGND.n1681 VGND.n532 0.362676
R5134 VGND.n1681 VGND.n1680 0.362676
R5135 VGND.n1680 VGND.n476 0.362676
R5136 VGND.n1855 VGND.n476 0.362676
R5137 VGND.n1855 VGND.n1854 0.362676
R5138 VGND.n1854 VGND.n420 0.362676
R5139 VGND.n2029 VGND.n420 0.362676
R5140 VGND.n2029 VGND.n2028 0.362676
R5141 VGND.n2028 VGND.n353 0.362676
R5142 VGND.n2203 VGND.n353 0.362676
R5143 VGND.n2203 VGND.n2202 0.362676
R5144 VGND.n2202 VGND.n200 0.362676
R5145 VGND.n2793 VGND.n200 0.362676
R5146 VGND.n1261 VGND.n1260 0.362676
R5147 VGND.n1260 VGND.n528 0.362676
R5148 VGND.n1693 VGND.n528 0.362676
R5149 VGND.n1694 VGND.n1693 0.362676
R5150 VGND.n1694 VGND.n472 0.362676
R5151 VGND.n1867 VGND.n472 0.362676
R5152 VGND.n1868 VGND.n1867 0.362676
R5153 VGND.n1868 VGND.n416 0.362676
R5154 VGND.n2041 VGND.n416 0.362676
R5155 VGND.n2042 VGND.n2041 0.362676
R5156 VGND.n2042 VGND.n349 0.362676
R5157 VGND.n2215 VGND.n349 0.362676
R5158 VGND.n2216 VGND.n2215 0.362676
R5159 VGND.n2216 VGND.n203 0.362676
R5160 VGND.n2790 VGND.n203 0.362676
R5161 VGND.n1257 VGND.n1256 0.362676
R5162 VGND.n1257 VGND.n524 0.362676
R5163 VGND.n1707 VGND.n524 0.362676
R5164 VGND.n1707 VGND.n1706 0.362676
R5165 VGND.n1706 VGND.n468 0.362676
R5166 VGND.n1881 VGND.n468 0.362676
R5167 VGND.n1881 VGND.n1880 0.362676
R5168 VGND.n1880 VGND.n412 0.362676
R5169 VGND.n2055 VGND.n412 0.362676
R5170 VGND.n2055 VGND.n2054 0.362676
R5171 VGND.n2054 VGND.n345 0.362676
R5172 VGND.n2229 VGND.n345 0.362676
R5173 VGND.n2229 VGND.n2228 0.362676
R5174 VGND.n2228 VGND.n206 0.362676
R5175 VGND.n2787 VGND.n206 0.362676
R5176 VGND.n1253 VGND.n1252 0.362676
R5177 VGND.n1252 VGND.n520 0.362676
R5178 VGND.n1719 VGND.n520 0.362676
R5179 VGND.n1720 VGND.n1719 0.362676
R5180 VGND.n1720 VGND.n464 0.362676
R5181 VGND.n1893 VGND.n464 0.362676
R5182 VGND.n1894 VGND.n1893 0.362676
R5183 VGND.n1894 VGND.n408 0.362676
R5184 VGND.n2067 VGND.n408 0.362676
R5185 VGND.n2068 VGND.n2067 0.362676
R5186 VGND.n2068 VGND.n341 0.362676
R5187 VGND.n2241 VGND.n341 0.362676
R5188 VGND.n2242 VGND.n2241 0.362676
R5189 VGND.n2242 VGND.n209 0.362676
R5190 VGND.n2784 VGND.n209 0.362676
R5191 VGND.n1249 VGND.n1248 0.362676
R5192 VGND.n1249 VGND.n516 0.362676
R5193 VGND.n1733 VGND.n516 0.362676
R5194 VGND.n1733 VGND.n1732 0.362676
R5195 VGND.n1732 VGND.n460 0.362676
R5196 VGND.n1907 VGND.n460 0.362676
R5197 VGND.n1907 VGND.n1906 0.362676
R5198 VGND.n1906 VGND.n404 0.362676
R5199 VGND.n2081 VGND.n404 0.362676
R5200 VGND.n2081 VGND.n2080 0.362676
R5201 VGND.n2080 VGND.n337 0.362676
R5202 VGND.n2255 VGND.n337 0.362676
R5203 VGND.n2255 VGND.n2254 0.362676
R5204 VGND.n2254 VGND.n212 0.362676
R5205 VGND.n2781 VGND.n212 0.362676
R5206 VGND.n1245 VGND.n1244 0.362676
R5207 VGND.n1244 VGND.n512 0.362676
R5208 VGND.n1750 VGND.n512 0.362676
R5209 VGND.n1751 VGND.n1750 0.362676
R5210 VGND.n1751 VGND.n456 0.362676
R5211 VGND.n1924 VGND.n456 0.362676
R5212 VGND.n1925 VGND.n1924 0.362676
R5213 VGND.n1925 VGND.n400 0.362676
R5214 VGND.n2098 VGND.n400 0.362676
R5215 VGND.n2099 VGND.n2098 0.362676
R5216 VGND.n2099 VGND.n333 0.362676
R5217 VGND.n2272 VGND.n333 0.362676
R5218 VGND.n2273 VGND.n2272 0.362676
R5219 VGND.n2273 VGND.n215 0.362676
R5220 VGND.n2778 VGND.n215 0.362676
R5221 VGND.n1241 VGND.n1240 0.362676
R5222 VGND.n1241 VGND.n292 0.362676
R5223 VGND.n2374 VGND.n292 0.362676
R5224 VGND.n2374 VGND.n2373 0.362676
R5225 VGND.n2373 VGND.n293 0.362676
R5226 VGND.n2349 VGND.n293 0.362676
R5227 VGND.n2349 VGND.n2348 0.362676
R5228 VGND.n2348 VGND.n305 0.362676
R5229 VGND.n2324 VGND.n305 0.362676
R5230 VGND.n2324 VGND.n2323 0.362676
R5231 VGND.n2323 VGND.n317 0.362676
R5232 VGND.n2299 VGND.n317 0.362676
R5233 VGND.n2299 VGND.n2298 0.362676
R5234 VGND.n2298 VGND.n218 0.362676
R5235 VGND.n2775 VGND.n218 0.362676
R5236 VGND.n2395 VGND.n280 0.362676
R5237 VGND.n2395 VGND.n2394 0.362676
R5238 VGND.n2394 VGND.n281 0.362676
R5239 VGND.n2370 VGND.n281 0.362676
R5240 VGND.n2370 VGND.n2369 0.362676
R5241 VGND.n2369 VGND.n296 0.362676
R5242 VGND.n2345 VGND.n296 0.362676
R5243 VGND.n2345 VGND.n2344 0.362676
R5244 VGND.n2344 VGND.n308 0.362676
R5245 VGND.n2320 VGND.n308 0.362676
R5246 VGND.n2320 VGND.n2319 0.362676
R5247 VGND.n2319 VGND.n320 0.362676
R5248 VGND.n2295 VGND.n320 0.362676
R5249 VGND.n2295 VGND.n221 0.362676
R5250 VGND.n2772 VGND.n221 0.362676
R5251 VGND.n1236 VGND.n285 0.362676
R5252 VGND.n2391 VGND.n285 0.362676
R5253 VGND.n2391 VGND.n2390 0.362676
R5254 VGND.n2390 VGND.n286 0.362676
R5255 VGND.n2366 VGND.n286 0.362676
R5256 VGND.n2366 VGND.n2365 0.362676
R5257 VGND.n2365 VGND.n299 0.362676
R5258 VGND.n2341 VGND.n299 0.362676
R5259 VGND.n2341 VGND.n2340 0.362676
R5260 VGND.n2340 VGND.n311 0.362676
R5261 VGND.n2316 VGND.n311 0.362676
R5262 VGND.n2316 VGND.n2315 0.362676
R5263 VGND.n2315 VGND.n323 0.362676
R5264 VGND.n323 VGND.n224 0.362676
R5265 VGND.n2769 VGND.n224 0.362676
R5266 VGND.n1283 VGND.n562 0.362676
R5267 VGND.n1543 VGND.n562 0.362676
R5268 VGND.n1543 VGND.n1542 0.362676
R5269 VGND.n1542 VGND.n563 0.362676
R5270 VGND.n1366 VGND.n563 0.362676
R5271 VGND.n1366 VGND.n662 0.362676
R5272 VGND.n1406 VGND.n662 0.362676
R5273 VGND.n1407 VGND.n1406 0.362676
R5274 VGND.n1407 VGND.n631 0.362676
R5275 VGND.n1498 VGND.n631 0.362676
R5276 VGND.n1498 VGND.n1497 0.362676
R5277 VGND.n1497 VGND.n183 0.362676
R5278 VGND.n2810 VGND.n183 0.362676
R5279 VGND.n2810 VGND.n2809 0.362676
R5280 VGND.n2809 VGND.n184 0.362676
R5281 VGND.n2617 VGND.n2578 0.349144
R5282 VGND.n2617 VGND.n2616 0.349144
R5283 VGND.n2616 VGND.n2613 0.349144
R5284 VGND.n2613 VGND.n2610 0.349144
R5285 VGND.n2610 VGND.n2607 0.349144
R5286 VGND.n2607 VGND.n2604 0.349144
R5287 VGND.n2604 VGND.n2601 0.349144
R5288 VGND.n2601 VGND.n2598 0.349144
R5289 VGND.n2598 VGND.n2595 0.349144
R5290 VGND.n2595 VGND.n2592 0.349144
R5291 VGND.n2592 VGND.n2589 0.349144
R5292 VGND.n2589 VGND.n2586 0.349144
R5293 VGND.n2586 VGND.n2583 0.349144
R5294 VGND.n1218 VGND.n1217 0.349144
R5295 VGND.n1218 VGND.n1214 0.349144
R5296 VGND.n1214 VGND.n790 0.349144
R5297 VGND.n1186 VGND.n790 0.349144
R5298 VGND.n1187 VGND.n1186 0.349144
R5299 VGND.n1187 VGND.n1182 0.349144
R5300 VGND.n1182 VGND.n798 0.349144
R5301 VGND.n1154 VGND.n798 0.349144
R5302 VGND.n1155 VGND.n1154 0.349144
R5303 VGND.n1155 VGND.n1150 0.349144
R5304 VGND.n1150 VGND.n806 0.349144
R5305 VGND.n818 VGND.n806 0.349144
R5306 VGND.n821 VGND.n818 0.349144
R5307 VGND.n2690 VGND.n2574 0.347091
R5308 VGND.n235 VGND.n234 0.347091
R5309 VGND.n2703 VGND.n2699 0.347091
R5310 VGND.n2708 VGND.n189 0.347091
R5311 VGND.n2713 VGND.n190 0.347091
R5312 VGND.n2718 VGND.n195 0.347091
R5313 VGND.n2723 VGND.n196 0.347091
R5314 VGND.n2728 VGND.n201 0.347091
R5315 VGND.n2733 VGND.n202 0.347091
R5316 VGND.n2738 VGND.n207 0.347091
R5317 VGND.n2743 VGND.n208 0.347091
R5318 VGND.n2748 VGND.n213 0.347091
R5319 VGND.n2753 VGND.n214 0.347091
R5320 VGND.n2758 VGND.n219 0.347091
R5321 VGND.n2763 VGND.n220 0.347091
R5322 VGND.n2767 VGND.n2766 0.347091
R5323 VGND.n2516 VGND.n2515 0.347091
R5324 VGND.n2512 VGND.n185 0.347091
R5325 VGND.n2507 VGND.n186 0.347091
R5326 VGND.n2504 VGND.n244 0.347091
R5327 VGND.n2437 VGND.n248 0.347091
R5328 VGND.n2442 VGND.n249 0.347091
R5329 VGND.n2447 VGND.n250 0.347091
R5330 VGND.n2452 VGND.n251 0.347091
R5331 VGND.n2457 VGND.n252 0.347091
R5332 VGND.n2462 VGND.n253 0.347091
R5333 VGND.n2467 VGND.n254 0.347091
R5334 VGND.n2472 VGND.n255 0.347091
R5335 VGND.n2477 VGND.n256 0.347091
R5336 VGND.n2482 VGND.n257 0.347091
R5337 VGND.n2487 VGND.n258 0.347091
R5338 VGND.n2815 VGND.n180 0.347091
R5339 VGND.n2812 VGND.n182 0.347091
R5340 VGND.n374 VGND.n373 0.347091
R5341 VGND.n2170 VGND.n2166 0.347091
R5342 VGND.n2174 VGND.n2173 0.347091
R5343 VGND.n2196 VGND.n2192 0.347091
R5344 VGND.n2200 VGND.n2199 0.347091
R5345 VGND.n2222 VGND.n2218 0.347091
R5346 VGND.n2226 VGND.n2225 0.347091
R5347 VGND.n2248 VGND.n2244 0.347091
R5348 VGND.n2252 VGND.n2251 0.347091
R5349 VGND.n2279 VGND.n2275 0.347091
R5350 VGND.n2284 VGND.n328 0.347091
R5351 VGND.n2289 VGND.n329 0.347091
R5352 VGND.n2293 VGND.n2292 0.347091
R5353 VGND.n1427 VGND.n1420 0.347091
R5354 VGND.n1431 VGND.n1430 0.347091
R5355 VGND.n2157 VGND.n2153 0.347091
R5356 VGND.n2161 VGND.n2160 0.347091
R5357 VGND.n2183 VGND.n2179 0.347091
R5358 VGND.n2187 VGND.n2186 0.347091
R5359 VGND.n2209 VGND.n2205 0.347091
R5360 VGND.n2213 VGND.n2212 0.347091
R5361 VGND.n2235 VGND.n2231 0.347091
R5362 VGND.n2239 VGND.n2238 0.347091
R5363 VGND.n2261 VGND.n2257 0.347091
R5364 VGND.n2270 VGND.n2269 0.347091
R5365 VGND.n2266 VGND.n327 0.347091
R5366 VGND.n2306 VGND.n2302 0.347091
R5367 VGND.n2309 VGND.n324 0.347091
R5368 VGND.n1441 VGND.n1437 0.347091
R5369 VGND.n1495 VGND.n1494 0.347091
R5370 VGND.n1491 VGND.n381 0.347091
R5371 VGND.n1486 VGND.n382 0.347091
R5372 VGND.n1481 VGND.n383 0.347091
R5373 VGND.n1476 VGND.n384 0.347091
R5374 VGND.n1471 VGND.n385 0.347091
R5375 VGND.n1466 VGND.n386 0.347091
R5376 VGND.n1461 VGND.n387 0.347091
R5377 VGND.n1456 VGND.n388 0.347091
R5378 VGND.n1451 VGND.n389 0.347091
R5379 VGND.n1446 VGND.n390 0.347091
R5380 VGND.n2138 VGND.n2137 0.347091
R5381 VGND.n2134 VGND.n321 0.347091
R5382 VGND.n2129 VGND.n322 0.347091
R5383 VGND.n1503 VGND.n617 0.347091
R5384 VGND.n1500 VGND.n619 0.347091
R5385 VGND.n629 VGND.n628 0.347091
R5386 VGND.n1996 VGND.n1992 0.347091
R5387 VGND.n2000 VGND.n1999 0.347091
R5388 VGND.n2022 VGND.n2018 0.347091
R5389 VGND.n2026 VGND.n2025 0.347091
R5390 VGND.n2048 VGND.n2044 0.347091
R5391 VGND.n2052 VGND.n2051 0.347091
R5392 VGND.n2074 VGND.n2070 0.347091
R5393 VGND.n2078 VGND.n2077 0.347091
R5394 VGND.n2105 VGND.n2101 0.347091
R5395 VGND.n2110 VGND.n318 0.347091
R5396 VGND.n2115 VGND.n319 0.347091
R5397 VGND.n2118 VGND.n399 0.347091
R5398 VGND.n651 VGND.n644 0.347091
R5399 VGND.n655 VGND.n654 0.347091
R5400 VGND.n1983 VGND.n1979 0.347091
R5401 VGND.n1987 VGND.n1986 0.347091
R5402 VGND.n2009 VGND.n2005 0.347091
R5403 VGND.n2013 VGND.n2012 0.347091
R5404 VGND.n2035 VGND.n2031 0.347091
R5405 VGND.n2039 VGND.n2038 0.347091
R5406 VGND.n2061 VGND.n2057 0.347091
R5407 VGND.n2065 VGND.n2064 0.347091
R5408 VGND.n2087 VGND.n2083 0.347091
R5409 VGND.n2096 VGND.n2095 0.347091
R5410 VGND.n2092 VGND.n316 0.347091
R5411 VGND.n2331 VGND.n2327 0.347091
R5412 VGND.n2334 VGND.n312 0.347091
R5413 VGND.n958 VGND.n660 0.347091
R5414 VGND.n953 VGND.n661 0.347091
R5415 VGND.n948 VGND.n437 0.347091
R5416 VGND.n943 VGND.n438 0.347091
R5417 VGND.n938 VGND.n439 0.347091
R5418 VGND.n933 VGND.n440 0.347091
R5419 VGND.n928 VGND.n441 0.347091
R5420 VGND.n923 VGND.n442 0.347091
R5421 VGND.n918 VGND.n443 0.347091
R5422 VGND.n913 VGND.n444 0.347091
R5423 VGND.n908 VGND.n445 0.347091
R5424 VGND.n903 VGND.n446 0.347091
R5425 VGND.n1964 VGND.n1963 0.347091
R5426 VGND.n1960 VGND.n309 0.347091
R5427 VGND.n1955 VGND.n310 0.347091
R5428 VGND.n1394 VGND.n1390 0.347091
R5429 VGND.n1399 VGND.n663 0.347091
R5430 VGND.n1403 VGND.n1402 0.347091
R5431 VGND.n1822 VGND.n1818 0.347091
R5432 VGND.n1826 VGND.n1825 0.347091
R5433 VGND.n1848 VGND.n1844 0.347091
R5434 VGND.n1852 VGND.n1851 0.347091
R5435 VGND.n1874 VGND.n1870 0.347091
R5436 VGND.n1878 VGND.n1877 0.347091
R5437 VGND.n1900 VGND.n1896 0.347091
R5438 VGND.n1904 VGND.n1903 0.347091
R5439 VGND.n1931 VGND.n1927 0.347091
R5440 VGND.n1936 VGND.n306 0.347091
R5441 VGND.n1941 VGND.n307 0.347091
R5442 VGND.n1944 VGND.n455 0.347091
R5443 VGND.n1379 VGND.n1372 0.347091
R5444 VGND.n1383 VGND.n1382 0.347091
R5445 VGND.n1809 VGND.n1805 0.347091
R5446 VGND.n1813 VGND.n1812 0.347091
R5447 VGND.n1835 VGND.n1831 0.347091
R5448 VGND.n1839 VGND.n1838 0.347091
R5449 VGND.n1861 VGND.n1857 0.347091
R5450 VGND.n1865 VGND.n1864 0.347091
R5451 VGND.n1887 VGND.n1883 0.347091
R5452 VGND.n1891 VGND.n1890 0.347091
R5453 VGND.n1913 VGND.n1909 0.347091
R5454 VGND.n1922 VGND.n1921 0.347091
R5455 VGND.n1918 VGND.n304 0.347091
R5456 VGND.n2356 VGND.n2352 0.347091
R5457 VGND.n2359 VGND.n300 0.347091
R5458 VGND.n1311 VGND.n1304 0.347091
R5459 VGND.n1365 VGND.n1364 0.347091
R5460 VGND.n1361 VGND.n493 0.347091
R5461 VGND.n1356 VGND.n494 0.347091
R5462 VGND.n1351 VGND.n495 0.347091
R5463 VGND.n1346 VGND.n496 0.347091
R5464 VGND.n1341 VGND.n497 0.347091
R5465 VGND.n1336 VGND.n498 0.347091
R5466 VGND.n1331 VGND.n499 0.347091
R5467 VGND.n1326 VGND.n500 0.347091
R5468 VGND.n1321 VGND.n501 0.347091
R5469 VGND.n1316 VGND.n502 0.347091
R5470 VGND.n1790 VGND.n1789 0.347091
R5471 VGND.n1786 VGND.n297 0.347091
R5472 VGND.n1781 VGND.n298 0.347091
R5473 VGND.n1516 VGND.n573 0.347091
R5474 VGND.n1521 VGND.n574 0.347091
R5475 VGND.n1525 VGND.n1524 0.347091
R5476 VGND.n1648 VGND.n1644 0.347091
R5477 VGND.n1652 VGND.n1651 0.347091
R5478 VGND.n1674 VGND.n1670 0.347091
R5479 VGND.n1678 VGND.n1677 0.347091
R5480 VGND.n1700 VGND.n1696 0.347091
R5481 VGND.n1704 VGND.n1703 0.347091
R5482 VGND.n1726 VGND.n1722 0.347091
R5483 VGND.n1730 VGND.n1729 0.347091
R5484 VGND.n1757 VGND.n1753 0.347091
R5485 VGND.n1762 VGND.n294 0.347091
R5486 VGND.n1767 VGND.n295 0.347091
R5487 VGND.n1770 VGND.n511 0.347091
R5488 VGND.n1536 VGND.n1532 0.347091
R5489 VGND.n1540 VGND.n1539 0.347091
R5490 VGND.n1635 VGND.n1631 0.347091
R5491 VGND.n1639 VGND.n1638 0.347091
R5492 VGND.n1661 VGND.n1657 0.347091
R5493 VGND.n1665 VGND.n1664 0.347091
R5494 VGND.n1687 VGND.n1683 0.347091
R5495 VGND.n1691 VGND.n1690 0.347091
R5496 VGND.n1713 VGND.n1709 0.347091
R5497 VGND.n1717 VGND.n1716 0.347091
R5498 VGND.n1739 VGND.n1735 0.347091
R5499 VGND.n1748 VGND.n1747 0.347091
R5500 VGND.n1744 VGND.n291 0.347091
R5501 VGND.n2381 VGND.n2377 0.347091
R5502 VGND.n2384 VGND.n287 0.347091
R5503 VGND.n1297 VGND.n1296 0.347091
R5504 VGND.n1549 VGND.n1545 0.347091
R5505 VGND.n1554 VGND.n549 0.347091
R5506 VGND.n1559 VGND.n550 0.347091
R5507 VGND.n1564 VGND.n551 0.347091
R5508 VGND.n1569 VGND.n552 0.347091
R5509 VGND.n1574 VGND.n553 0.347091
R5510 VGND.n1579 VGND.n554 0.347091
R5511 VGND.n1584 VGND.n555 0.347091
R5512 VGND.n1589 VGND.n556 0.347091
R5513 VGND.n1594 VGND.n557 0.347091
R5514 VGND.n1599 VGND.n558 0.347091
R5515 VGND.n1616 VGND.n1615 0.347091
R5516 VGND.n1612 VGND.n282 0.347091
R5517 VGND.n1607 VGND.n283 0.347091
R5518 VGND.n834 VGND.n826 0.347091
R5519 VGND.n839 VGND.n827 0.347091
R5520 VGND.n893 VGND.n892 0.347091
R5521 VGND.n889 VGND.n688 0.347091
R5522 VGND.n884 VGND.n689 0.347091
R5523 VGND.n879 VGND.n694 0.347091
R5524 VGND.n874 VGND.n695 0.347091
R5525 VGND.n869 VGND.n700 0.347091
R5526 VGND.n864 VGND.n701 0.347091
R5527 VGND.n859 VGND.n706 0.347091
R5528 VGND.n854 VGND.n707 0.347091
R5529 VGND.n849 VGND.n712 0.347091
R5530 VGND.n844 VGND.n713 0.347091
R5531 VGND.n2401 VGND.n2397 0.347091
R5532 VGND.n2404 VGND.n279 0.347091
R5533 VGND.n1123 VGND.n1121 0.347091
R5534 VGND.n1130 VGND.n1126 0.347091
R5535 VGND.n1133 VGND.n812 0.347091
R5536 VGND.n1143 VGND.n1139 0.347091
R5537 VGND.n1147 VGND.n1146 0.347091
R5538 VGND.n1162 VGND.n1158 0.347091
R5539 VGND.n1165 VGND.n804 0.347091
R5540 VGND.n1175 VGND.n1171 0.347091
R5541 VGND.n1179 VGND.n1178 0.347091
R5542 VGND.n1194 VGND.n1190 0.347091
R5543 VGND.n1197 VGND.n796 0.347091
R5544 VGND.n1207 VGND.n1203 0.347091
R5545 VGND.n1211 VGND.n1210 0.347091
R5546 VGND.n1226 VGND.n1222 0.347091
R5547 VGND.n1229 VGND.n788 0.347091
R5548 VGND.n1288 VGND.n677 0.347091
R5549 VGND.n1285 VGND.n679 0.347091
R5550 VGND.n724 VGND.n685 0.347091
R5551 VGND.n729 VGND.n686 0.347091
R5552 VGND.n734 VGND.n691 0.347091
R5553 VGND.n739 VGND.n692 0.347091
R5554 VGND.n744 VGND.n697 0.347091
R5555 VGND.n749 VGND.n698 0.347091
R5556 VGND.n754 VGND.n703 0.347091
R5557 VGND.n759 VGND.n704 0.347091
R5558 VGND.n764 VGND.n709 0.347091
R5559 VGND.n769 VGND.n710 0.347091
R5560 VGND.n774 VGND.n715 0.347091
R5561 VGND.n779 VGND.n716 0.347091
R5562 VGND.n783 VGND.n782 0.347091
R5563 VGND.n2644 VGND.n2640 0.34283
R5564 VGND.n2649 VGND.n2647 0.34283
R5565 VGND.n2651 VGND.n2637 0.34283
R5566 VGND.n2656 VGND.n2654 0.34283
R5567 VGND.n2658 VGND.n2634 0.34283
R5568 VGND.n2663 VGND.n2661 0.34283
R5569 VGND.n2665 VGND.n2631 0.34283
R5570 VGND.n2670 VGND.n2668 0.34283
R5571 VGND.n2672 VGND.n2628 0.34283
R5572 VGND.n2677 VGND.n2675 0.34283
R5573 VGND.n2679 VGND.n2625 0.34283
R5574 VGND.n2684 VGND.n2682 0.34283
R5575 VGND.n2686 VGND.n2622 0.34283
R5576 VGND.n2692 VGND.n2570 0.34283
R5577 VGND.n3008 VGND.n2 0.247202
R5578 VGND.n2904 VGND.n59 0.213567
R5579 VGND.n2937 VGND.n2904 0.213567
R5580 VGND.n2938 VGND.n2937 0.213567
R5581 VGND.n2938 VGND.n28 0.213567
R5582 VGND.n1113 VGND.n1090 0.213567
R5583 VGND.n1090 VGND.n1060 0.213567
R5584 VGND.n1060 VGND.n1029 0.213567
R5585 VGND.n1029 VGND.n998 0.213567
R5586 VGND.n998 VGND.n0 0.213567
R5587 VGND.n2990 VGND.n28 0.2073
R5588 VGND.n1115 VGND.n1114 0.17205
R5589 VGND.n2695 VGND 0.169807
R5590 VGND.n2694 VGND 0.169807
R5591 VGND VGND.n188 0.169807
R5592 VGND.n2801 VGND 0.169807
R5593 VGND.n2800 VGND 0.169807
R5594 VGND.n2795 VGND 0.169807
R5595 VGND.n2794 VGND 0.169807
R5596 VGND.n2789 VGND 0.169807
R5597 VGND.n2788 VGND 0.169807
R5598 VGND.n2783 VGND 0.169807
R5599 VGND.n2782 VGND 0.169807
R5600 VGND.n2777 VGND 0.169807
R5601 VGND.n2776 VGND 0.169807
R5602 VGND.n2771 VGND 0.169807
R5603 VGND.n2770 VGND 0.169807
R5604 VGND VGND.n2697 0.169807
R5605 VGND.n2698 VGND 0.169807
R5606 VGND.n2804 VGND 0.169807
R5607 VGND.n2803 VGND 0.169807
R5608 VGND.n2798 VGND 0.169807
R5609 VGND.n2797 VGND 0.169807
R5610 VGND.n2792 VGND 0.169807
R5611 VGND.n2791 VGND 0.169807
R5612 VGND.n2786 VGND 0.169807
R5613 VGND.n2785 VGND 0.169807
R5614 VGND.n2780 VGND 0.169807
R5615 VGND.n2779 VGND 0.169807
R5616 VGND.n2774 VGND 0.169807
R5617 VGND.n2773 VGND 0.169807
R5618 VGND.n2768 VGND 0.169807
R5619 VGND.n2517 VGND 0.169807
R5620 VGND.n2808 VGND 0.169807
R5621 VGND.n2807 VGND 0.169807
R5622 VGND.n2503 VGND 0.169807
R5623 VGND.n2502 VGND 0.169807
R5624 VGND.n2501 VGND 0.169807
R5625 VGND.n2500 VGND 0.169807
R5626 VGND.n2499 VGND 0.169807
R5627 VGND.n2498 VGND 0.169807
R5628 VGND.n2497 VGND 0.169807
R5629 VGND.n2496 VGND 0.169807
R5630 VGND.n2495 VGND 0.169807
R5631 VGND.n2494 VGND 0.169807
R5632 VGND.n2493 VGND 0.169807
R5633 VGND.n2492 VGND 0.169807
R5634 VGND.n639 VGND 0.169807
R5635 VGND.n2811 VGND 0.169807
R5636 VGND VGND.n375 0.169807
R5637 VGND.n2165 VGND 0.169807
R5638 VGND.n2175 VGND 0.169807
R5639 VGND.n2191 VGND 0.169807
R5640 VGND.n2201 VGND 0.169807
R5641 VGND.n2217 VGND 0.169807
R5642 VGND.n2227 VGND 0.169807
R5643 VGND.n2243 VGND 0.169807
R5644 VGND.n2253 VGND 0.169807
R5645 VGND.n2274 VGND 0.169807
R5646 VGND.n2297 VGND 0.169807
R5647 VGND.n2296 VGND 0.169807
R5648 VGND.n2294 VGND 0.169807
R5649 VGND.n1433 VGND 0.169807
R5650 VGND.n1432 VGND 0.169807
R5651 VGND.n2152 VGND 0.169807
R5652 VGND.n2162 VGND 0.169807
R5653 VGND.n2178 VGND 0.169807
R5654 VGND.n2188 VGND 0.169807
R5655 VGND.n2204 VGND 0.169807
R5656 VGND.n2214 VGND 0.169807
R5657 VGND.n2230 VGND 0.169807
R5658 VGND.n2240 VGND 0.169807
R5659 VGND.n2256 VGND 0.169807
R5660 VGND.n2271 VGND 0.169807
R5661 VGND VGND.n2300 0.169807
R5662 VGND.n2301 VGND 0.169807
R5663 VGND.n2314 VGND 0.169807
R5664 VGND.n1436 VGND 0.169807
R5665 VGND.n1496 VGND 0.169807
R5666 VGND.n2149 VGND 0.169807
R5667 VGND.n2148 VGND 0.169807
R5668 VGND.n2147 VGND 0.169807
R5669 VGND.n2146 VGND 0.169807
R5670 VGND.n2145 VGND 0.169807
R5671 VGND.n2144 VGND 0.169807
R5672 VGND.n2143 VGND 0.169807
R5673 VGND.n2142 VGND 0.169807
R5674 VGND.n2141 VGND 0.169807
R5675 VGND.n2140 VGND 0.169807
R5676 VGND.n2139 VGND 0.169807
R5677 VGND.n2318 VGND 0.169807
R5678 VGND.n2317 VGND 0.169807
R5679 VGND.n1414 VGND 0.169807
R5680 VGND.n1499 VGND 0.169807
R5681 VGND.n630 VGND 0.169807
R5682 VGND.n1991 VGND 0.169807
R5683 VGND.n2001 VGND 0.169807
R5684 VGND.n2017 VGND 0.169807
R5685 VGND.n2027 VGND 0.169807
R5686 VGND.n2043 VGND 0.169807
R5687 VGND.n2053 VGND 0.169807
R5688 VGND.n2069 VGND 0.169807
R5689 VGND.n2079 VGND 0.169807
R5690 VGND.n2100 VGND 0.169807
R5691 VGND.n2322 VGND 0.169807
R5692 VGND.n2321 VGND 0.169807
R5693 VGND.n398 VGND 0.169807
R5694 VGND.n1412 VGND 0.169807
R5695 VGND.n656 VGND 0.169807
R5696 VGND.n1978 VGND 0.169807
R5697 VGND.n1988 VGND 0.169807
R5698 VGND.n2004 VGND 0.169807
R5699 VGND.n2014 VGND 0.169807
R5700 VGND.n2030 VGND 0.169807
R5701 VGND.n2040 VGND 0.169807
R5702 VGND.n2056 VGND 0.169807
R5703 VGND.n2066 VGND 0.169807
R5704 VGND.n2082 VGND 0.169807
R5705 VGND.n2097 VGND 0.169807
R5706 VGND VGND.n2325 0.169807
R5707 VGND.n2326 VGND 0.169807
R5708 VGND.n2339 VGND 0.169807
R5709 VGND.n1409 VGND 0.169807
R5710 VGND.n1408 VGND 0.169807
R5711 VGND.n1975 VGND 0.169807
R5712 VGND.n1974 VGND 0.169807
R5713 VGND.n1973 VGND 0.169807
R5714 VGND.n1972 VGND 0.169807
R5715 VGND.n1971 VGND 0.169807
R5716 VGND.n1970 VGND 0.169807
R5717 VGND.n1969 VGND 0.169807
R5718 VGND.n1968 VGND 0.169807
R5719 VGND.n1967 VGND 0.169807
R5720 VGND.n1966 VGND 0.169807
R5721 VGND.n1965 VGND 0.169807
R5722 VGND.n2343 VGND 0.169807
R5723 VGND.n2342 VGND 0.169807
R5724 VGND.n1389 VGND 0.169807
R5725 VGND.n1405 VGND 0.169807
R5726 VGND.n1404 VGND 0.169807
R5727 VGND.n1817 VGND 0.169807
R5728 VGND.n1827 VGND 0.169807
R5729 VGND.n1843 VGND 0.169807
R5730 VGND.n1853 VGND 0.169807
R5731 VGND.n1869 VGND 0.169807
R5732 VGND.n1879 VGND 0.169807
R5733 VGND.n1895 VGND 0.169807
R5734 VGND.n1905 VGND 0.169807
R5735 VGND.n1926 VGND 0.169807
R5736 VGND.n2347 VGND 0.169807
R5737 VGND.n2346 VGND 0.169807
R5738 VGND.n454 VGND 0.169807
R5739 VGND.n1386 VGND 0.169807
R5740 VGND.n1384 VGND 0.169807
R5741 VGND.n1804 VGND 0.169807
R5742 VGND.n1814 VGND 0.169807
R5743 VGND.n1830 VGND 0.169807
R5744 VGND.n1840 VGND 0.169807
R5745 VGND.n1856 VGND 0.169807
R5746 VGND.n1866 VGND 0.169807
R5747 VGND.n1882 VGND 0.169807
R5748 VGND.n1892 VGND 0.169807
R5749 VGND.n1908 VGND 0.169807
R5750 VGND.n1923 VGND 0.169807
R5751 VGND VGND.n2350 0.169807
R5752 VGND.n2351 VGND 0.169807
R5753 VGND.n2364 VGND 0.169807
R5754 VGND.n1368 VGND 0.169807
R5755 VGND.n1367 VGND 0.169807
R5756 VGND.n1801 VGND 0.169807
R5757 VGND.n1800 VGND 0.169807
R5758 VGND.n1799 VGND 0.169807
R5759 VGND.n1798 VGND 0.169807
R5760 VGND.n1797 VGND 0.169807
R5761 VGND.n1796 VGND 0.169807
R5762 VGND.n1795 VGND 0.169807
R5763 VGND.n1794 VGND 0.169807
R5764 VGND.n1793 VGND 0.169807
R5765 VGND.n1792 VGND 0.169807
R5766 VGND.n1791 VGND 0.169807
R5767 VGND.n2368 VGND 0.169807
R5768 VGND.n2367 VGND 0.169807
R5769 VGND.n1528 VGND 0.169807
R5770 VGND.n1527 VGND 0.169807
R5771 VGND.n1526 VGND 0.169807
R5772 VGND.n1643 VGND 0.169807
R5773 VGND.n1653 VGND 0.169807
R5774 VGND.n1669 VGND 0.169807
R5775 VGND.n1679 VGND 0.169807
R5776 VGND.n1695 VGND 0.169807
R5777 VGND.n1705 VGND 0.169807
R5778 VGND.n1721 VGND 0.169807
R5779 VGND.n1731 VGND 0.169807
R5780 VGND.n1752 VGND 0.169807
R5781 VGND.n2372 VGND 0.169807
R5782 VGND.n2371 VGND 0.169807
R5783 VGND.n510 VGND 0.169807
R5784 VGND.n1531 VGND 0.169807
R5785 VGND.n1541 VGND 0.169807
R5786 VGND.n1630 VGND 0.169807
R5787 VGND.n1640 VGND 0.169807
R5788 VGND.n1656 VGND 0.169807
R5789 VGND.n1666 VGND 0.169807
R5790 VGND.n1682 VGND 0.169807
R5791 VGND.n1692 VGND 0.169807
R5792 VGND.n1708 VGND 0.169807
R5793 VGND.n1718 VGND 0.169807
R5794 VGND.n1734 VGND 0.169807
R5795 VGND.n1749 VGND 0.169807
R5796 VGND VGND.n2375 0.169807
R5797 VGND.n2376 VGND 0.169807
R5798 VGND.n2389 VGND 0.169807
R5799 VGND.n1298 VGND 0.169807
R5800 VGND.n1544 VGND 0.169807
R5801 VGND.n1627 VGND 0.169807
R5802 VGND.n1626 VGND 0.169807
R5803 VGND.n1625 VGND 0.169807
R5804 VGND.n1624 VGND 0.169807
R5805 VGND.n1623 VGND 0.169807
R5806 VGND.n1622 VGND 0.169807
R5807 VGND.n1621 VGND 0.169807
R5808 VGND.n1620 VGND 0.169807
R5809 VGND.n1619 VGND 0.169807
R5810 VGND.n1618 VGND 0.169807
R5811 VGND.n1617 VGND 0.169807
R5812 VGND.n2393 VGND 0.169807
R5813 VGND.n2392 VGND 0.169807
R5814 VGND.n896 VGND 0.169807
R5815 VGND.n895 VGND 0.169807
R5816 VGND.n894 VGND 0.169807
R5817 VGND.n1275 VGND 0.169807
R5818 VGND.n1274 VGND 0.169807
R5819 VGND.n1267 VGND 0.169807
R5820 VGND.n1266 VGND 0.169807
R5821 VGND.n1259 VGND 0.169807
R5822 VGND.n1258 VGND 0.169807
R5823 VGND.n1251 VGND 0.169807
R5824 VGND.n1250 VGND 0.169807
R5825 VGND.n1243 VGND 0.169807
R5826 VGND.n1242 VGND 0.169807
R5827 VGND.n2396 VGND 0.169807
R5828 VGND.n284 VGND 0.169807
R5829 VGND.n1119 VGND 0.169807
R5830 VGND.n1282 VGND 0.169807
R5831 VGND.n1281 VGND 0.169807
R5832 VGND VGND.n687 0.169807
R5833 VGND VGND.n690 0.169807
R5834 VGND VGND.n693 0.169807
R5835 VGND VGND.n696 0.169807
R5836 VGND VGND.n699 0.169807
R5837 VGND VGND.n702 0.169807
R5838 VGND VGND.n705 0.169807
R5839 VGND VGND.n708 0.169807
R5840 VGND VGND.n711 0.169807
R5841 VGND VGND.n714 0.169807
R5842 VGND.n1220 VGND 0.169807
R5843 VGND.n1235 VGND 0.169807
R5844 VGND.n1117 VGND 0.169807
R5845 VGND.n1284 VGND 0.169807
R5846 VGND.n1279 VGND 0.169807
R5847 VGND.n1278 VGND 0.169807
R5848 VGND.n1271 VGND 0.169807
R5849 VGND.n1270 VGND 0.169807
R5850 VGND.n1263 VGND 0.169807
R5851 VGND.n1262 VGND 0.169807
R5852 VGND.n1255 VGND 0.169807
R5853 VGND.n1254 VGND 0.169807
R5854 VGND.n1247 VGND 0.169807
R5855 VGND.n1246 VGND 0.169807
R5856 VGND.n1239 VGND 0.169807
R5857 VGND.n1238 VGND 0.169807
R5858 VGND.n1237 VGND 0.169807
R5859 VGND.n109 VGND 0.159538
R5860 VGND.n2855 VGND 0.159538
R5861 VGND.n2410 VGND.n275 0.154425
R5862 VGND.n2410 VGND.n2409 0.154425
R5863 VGND.n2409 VGND.n276 0.154425
R5864 VGND.n289 VGND.n276 0.154425
R5865 VGND.n1775 VGND.n289 0.154425
R5866 VGND.n1776 VGND.n1775 0.154425
R5867 VGND.n1776 VGND.n302 0.154425
R5868 VGND.n1949 VGND.n302 0.154425
R5869 VGND.n1950 VGND.n1949 0.154425
R5870 VGND.n1950 VGND.n314 0.154425
R5871 VGND.n2123 VGND.n314 0.154425
R5872 VGND.n2124 VGND.n2123 0.154425
R5873 VGND.n2124 VGND.n259 0.154425
R5874 VGND.n2431 VGND.n259 0.154425
R5875 VGND.n2432 VGND.n2431 0.154425
R5876 VGND.n2432 VGND.n29 0.154425
R5877 VGND.n2989 VGND.n29 0.154425
R5878 VGND.n1116 VGND.n1115 0.154425
R5879 VGND.n1116 VGND.n669 0.154425
R5880 VGND.n1299 VGND.n669 0.154425
R5881 VGND.n1300 VGND.n1299 0.154425
R5882 VGND.n1301 VGND.n1300 0.154425
R5883 VGND.n1369 VGND.n1301 0.154425
R5884 VGND.n1387 VGND.n1369 0.154425
R5885 VGND.n1388 VGND.n1387 0.154425
R5886 VGND.n1388 VGND.n641 0.154425
R5887 VGND.n1413 VGND.n641 0.154425
R5888 VGND.n1415 VGND.n1413 0.154425
R5889 VGND.n1416 VGND.n1415 0.154425
R5890 VGND.n1417 VGND.n1416 0.154425
R5891 VGND.n1417 VGND.n237 0.154425
R5892 VGND.n2518 VGND.n237 0.154425
R5893 VGND.n2519 VGND.n2518 0.154425
R5894 VGND.n2520 VGND.n2519 0.154425
R5895 VGND.n2644 VGND.n2643 0.145386
R5896 VGND.n2647 VGND.n2638 0.145386
R5897 VGND.n2651 VGND.n2650 0.145386
R5898 VGND.n2654 VGND.n2635 0.145386
R5899 VGND.n2658 VGND.n2657 0.145386
R5900 VGND.n2661 VGND.n2632 0.145386
R5901 VGND.n2665 VGND.n2664 0.145386
R5902 VGND.n2668 VGND.n2629 0.145386
R5903 VGND.n2672 VGND.n2671 0.145386
R5904 VGND.n2675 VGND.n2626 0.145386
R5905 VGND.n2679 VGND.n2678 0.145386
R5906 VGND.n2682 VGND.n2623 0.145386
R5907 VGND.n2686 VGND.n2685 0.145386
R5908 VGND.n2621 VGND.n2570 0.145386
R5909 VGND.n2691 VGND.n2690 0.145386
R5910 VGND.n234 VGND.n232 0.145386
R5911 VGND.n2703 VGND.n2702 0.145386
R5912 VGND.n2708 VGND.n2707 0.145386
R5913 VGND.n2713 VGND.n2712 0.145386
R5914 VGND.n2718 VGND.n2717 0.145386
R5915 VGND.n2723 VGND.n2722 0.145386
R5916 VGND.n2728 VGND.n2727 0.145386
R5917 VGND.n2733 VGND.n2732 0.145386
R5918 VGND.n2738 VGND.n2737 0.145386
R5919 VGND.n2743 VGND.n2742 0.145386
R5920 VGND.n2748 VGND.n2747 0.145386
R5921 VGND.n2753 VGND.n2752 0.145386
R5922 VGND.n2758 VGND.n2757 0.145386
R5923 VGND.n2763 VGND.n2762 0.145386
R5924 VGND.n2766 VGND.n227 0.145386
R5925 VGND.n2515 VGND.n242 0.145386
R5926 VGND.n2512 VGND.n2511 0.145386
R5927 VGND.n2507 VGND.n2506 0.145386
R5928 VGND.n246 VGND.n244 0.145386
R5929 VGND.n2437 VGND.n2436 0.145386
R5930 VGND.n2442 VGND.n2441 0.145386
R5931 VGND.n2447 VGND.n2446 0.145386
R5932 VGND.n2452 VGND.n2451 0.145386
R5933 VGND.n2457 VGND.n2456 0.145386
R5934 VGND.n2462 VGND.n2461 0.145386
R5935 VGND.n2467 VGND.n2466 0.145386
R5936 VGND.n2472 VGND.n2471 0.145386
R5937 VGND.n2477 VGND.n2476 0.145386
R5938 VGND.n2482 VGND.n2481 0.145386
R5939 VGND.n2487 VGND.n2486 0.145386
R5940 VGND.n2815 VGND.n2814 0.145386
R5941 VGND.n366 VGND.n182 0.145386
R5942 VGND.n373 VGND.n370 0.145386
R5943 VGND.n2170 VGND.n2169 0.145386
R5944 VGND.n2173 VGND.n364 0.145386
R5945 VGND.n2196 VGND.n2195 0.145386
R5946 VGND.n2199 VGND.n356 0.145386
R5947 VGND.n2222 VGND.n2221 0.145386
R5948 VGND.n2225 VGND.n348 0.145386
R5949 VGND.n2248 VGND.n2247 0.145386
R5950 VGND.n2251 VGND.n340 0.145386
R5951 VGND.n2279 VGND.n2278 0.145386
R5952 VGND.n2284 VGND.n2283 0.145386
R5953 VGND.n2289 VGND.n2288 0.145386
R5954 VGND.n2292 VGND.n332 0.145386
R5955 VGND.n1427 VGND.n1426 0.145386
R5956 VGND.n1430 VGND.n1423 0.145386
R5957 VGND.n2157 VGND.n2156 0.145386
R5958 VGND.n2160 VGND.n379 0.145386
R5959 VGND.n2183 VGND.n2182 0.145386
R5960 VGND.n2186 VGND.n360 0.145386
R5961 VGND.n2209 VGND.n2208 0.145386
R5962 VGND.n2212 VGND.n352 0.145386
R5963 VGND.n2235 VGND.n2234 0.145386
R5964 VGND.n2238 VGND.n344 0.145386
R5965 VGND.n2261 VGND.n2260 0.145386
R5966 VGND.n2269 VGND.n336 0.145386
R5967 VGND.n2266 VGND.n2265 0.145386
R5968 VGND.n2306 VGND.n2305 0.145386
R5969 VGND.n2310 VGND.n2309 0.145386
R5970 VGND.n1441 VGND.n1440 0.145386
R5971 VGND.n1494 VGND.n634 0.145386
R5972 VGND.n1491 VGND.n1490 0.145386
R5973 VGND.n1486 VGND.n1485 0.145386
R5974 VGND.n1481 VGND.n1480 0.145386
R5975 VGND.n1476 VGND.n1475 0.145386
R5976 VGND.n1471 VGND.n1470 0.145386
R5977 VGND.n1466 VGND.n1465 0.145386
R5978 VGND.n1461 VGND.n1460 0.145386
R5979 VGND.n1456 VGND.n1455 0.145386
R5980 VGND.n1451 VGND.n1450 0.145386
R5981 VGND.n1446 VGND.n1445 0.145386
R5982 VGND.n2137 VGND.n393 0.145386
R5983 VGND.n2134 VGND.n2133 0.145386
R5984 VGND.n2129 VGND.n2128 0.145386
R5985 VGND.n1503 VGND.n1502 0.145386
R5986 VGND.n621 VGND.n619 0.145386
R5987 VGND.n628 VGND.n625 0.145386
R5988 VGND.n1996 VGND.n1995 0.145386
R5989 VGND.n1999 VGND.n431 0.145386
R5990 VGND.n2022 VGND.n2021 0.145386
R5991 VGND.n2025 VGND.n423 0.145386
R5992 VGND.n2048 VGND.n2047 0.145386
R5993 VGND.n2051 VGND.n415 0.145386
R5994 VGND.n2074 VGND.n2073 0.145386
R5995 VGND.n2077 VGND.n407 0.145386
R5996 VGND.n2105 VGND.n2104 0.145386
R5997 VGND.n2110 VGND.n2109 0.145386
R5998 VGND.n2115 VGND.n2114 0.145386
R5999 VGND.n2119 VGND.n2118 0.145386
R6000 VGND.n651 VGND.n650 0.145386
R6001 VGND.n654 VGND.n647 0.145386
R6002 VGND.n1983 VGND.n1982 0.145386
R6003 VGND.n1986 VGND.n435 0.145386
R6004 VGND.n2009 VGND.n2008 0.145386
R6005 VGND.n2012 VGND.n427 0.145386
R6006 VGND.n2035 VGND.n2034 0.145386
R6007 VGND.n2038 VGND.n419 0.145386
R6008 VGND.n2061 VGND.n2060 0.145386
R6009 VGND.n2064 VGND.n411 0.145386
R6010 VGND.n2087 VGND.n2086 0.145386
R6011 VGND.n2095 VGND.n403 0.145386
R6012 VGND.n2092 VGND.n2091 0.145386
R6013 VGND.n2331 VGND.n2330 0.145386
R6014 VGND.n2335 VGND.n2334 0.145386
R6015 VGND.n958 VGND.n957 0.145386
R6016 VGND.n953 VGND.n952 0.145386
R6017 VGND.n948 VGND.n947 0.145386
R6018 VGND.n943 VGND.n942 0.145386
R6019 VGND.n938 VGND.n937 0.145386
R6020 VGND.n933 VGND.n932 0.145386
R6021 VGND.n928 VGND.n927 0.145386
R6022 VGND.n923 VGND.n922 0.145386
R6023 VGND.n918 VGND.n917 0.145386
R6024 VGND.n913 VGND.n912 0.145386
R6025 VGND.n908 VGND.n907 0.145386
R6026 VGND.n903 VGND.n902 0.145386
R6027 VGND.n1963 VGND.n449 0.145386
R6028 VGND.n1960 VGND.n1959 0.145386
R6029 VGND.n1955 VGND.n1954 0.145386
R6030 VGND.n1394 VGND.n1393 0.145386
R6031 VGND.n1399 VGND.n1398 0.145386
R6032 VGND.n1402 VGND.n666 0.145386
R6033 VGND.n1822 VGND.n1821 0.145386
R6034 VGND.n1825 VGND.n487 0.145386
R6035 VGND.n1848 VGND.n1847 0.145386
R6036 VGND.n1851 VGND.n479 0.145386
R6037 VGND.n1874 VGND.n1873 0.145386
R6038 VGND.n1877 VGND.n471 0.145386
R6039 VGND.n1900 VGND.n1899 0.145386
R6040 VGND.n1903 VGND.n463 0.145386
R6041 VGND.n1931 VGND.n1930 0.145386
R6042 VGND.n1936 VGND.n1935 0.145386
R6043 VGND.n1941 VGND.n1940 0.145386
R6044 VGND.n1945 VGND.n1944 0.145386
R6045 VGND.n1379 VGND.n1378 0.145386
R6046 VGND.n1382 VGND.n1375 0.145386
R6047 VGND.n1809 VGND.n1808 0.145386
R6048 VGND.n1812 VGND.n491 0.145386
R6049 VGND.n1835 VGND.n1834 0.145386
R6050 VGND.n1838 VGND.n483 0.145386
R6051 VGND.n1861 VGND.n1860 0.145386
R6052 VGND.n1864 VGND.n475 0.145386
R6053 VGND.n1887 VGND.n1886 0.145386
R6054 VGND.n1890 VGND.n467 0.145386
R6055 VGND.n1913 VGND.n1912 0.145386
R6056 VGND.n1921 VGND.n459 0.145386
R6057 VGND.n1918 VGND.n1917 0.145386
R6058 VGND.n2356 VGND.n2355 0.145386
R6059 VGND.n2360 VGND.n2359 0.145386
R6060 VGND.n1311 VGND.n1310 0.145386
R6061 VGND.n1364 VGND.n1307 0.145386
R6062 VGND.n1361 VGND.n1360 0.145386
R6063 VGND.n1356 VGND.n1355 0.145386
R6064 VGND.n1351 VGND.n1350 0.145386
R6065 VGND.n1346 VGND.n1345 0.145386
R6066 VGND.n1341 VGND.n1340 0.145386
R6067 VGND.n1336 VGND.n1335 0.145386
R6068 VGND.n1331 VGND.n1330 0.145386
R6069 VGND.n1326 VGND.n1325 0.145386
R6070 VGND.n1321 VGND.n1320 0.145386
R6071 VGND.n1316 VGND.n1315 0.145386
R6072 VGND.n1789 VGND.n505 0.145386
R6073 VGND.n1786 VGND.n1785 0.145386
R6074 VGND.n1781 VGND.n1780 0.145386
R6075 VGND.n1516 VGND.n1515 0.145386
R6076 VGND.n1521 VGND.n1520 0.145386
R6077 VGND.n1524 VGND.n577 0.145386
R6078 VGND.n1648 VGND.n1647 0.145386
R6079 VGND.n1651 VGND.n543 0.145386
R6080 VGND.n1674 VGND.n1673 0.145386
R6081 VGND.n1677 VGND.n535 0.145386
R6082 VGND.n1700 VGND.n1699 0.145386
R6083 VGND.n1703 VGND.n527 0.145386
R6084 VGND.n1726 VGND.n1725 0.145386
R6085 VGND.n1729 VGND.n519 0.145386
R6086 VGND.n1757 VGND.n1756 0.145386
R6087 VGND.n1762 VGND.n1761 0.145386
R6088 VGND.n1767 VGND.n1766 0.145386
R6089 VGND.n1771 VGND.n1770 0.145386
R6090 VGND.n1536 VGND.n1535 0.145386
R6091 VGND.n1539 VGND.n566 0.145386
R6092 VGND.n1635 VGND.n1634 0.145386
R6093 VGND.n1638 VGND.n547 0.145386
R6094 VGND.n1661 VGND.n1660 0.145386
R6095 VGND.n1664 VGND.n539 0.145386
R6096 VGND.n1687 VGND.n1686 0.145386
R6097 VGND.n1690 VGND.n531 0.145386
R6098 VGND.n1713 VGND.n1712 0.145386
R6099 VGND.n1716 VGND.n523 0.145386
R6100 VGND.n1739 VGND.n1738 0.145386
R6101 VGND.n1747 VGND.n515 0.145386
R6102 VGND.n1744 VGND.n1743 0.145386
R6103 VGND.n2381 VGND.n2380 0.145386
R6104 VGND.n2385 VGND.n2384 0.145386
R6105 VGND.n1296 VGND.n674 0.145386
R6106 VGND.n1549 VGND.n1548 0.145386
R6107 VGND.n1554 VGND.n1553 0.145386
R6108 VGND.n1559 VGND.n1558 0.145386
R6109 VGND.n1564 VGND.n1563 0.145386
R6110 VGND.n1569 VGND.n1568 0.145386
R6111 VGND.n1574 VGND.n1573 0.145386
R6112 VGND.n1579 VGND.n1578 0.145386
R6113 VGND.n1584 VGND.n1583 0.145386
R6114 VGND.n1589 VGND.n1588 0.145386
R6115 VGND.n1594 VGND.n1593 0.145386
R6116 VGND.n1599 VGND.n1598 0.145386
R6117 VGND.n1615 VGND.n561 0.145386
R6118 VGND.n1612 VGND.n1611 0.145386
R6119 VGND.n1607 VGND.n1606 0.145386
R6120 VGND.n834 VGND.n833 0.145386
R6121 VGND.n839 VGND.n838 0.145386
R6122 VGND.n892 VGND.n830 0.145386
R6123 VGND.n889 VGND.n888 0.145386
R6124 VGND.n884 VGND.n883 0.145386
R6125 VGND.n879 VGND.n878 0.145386
R6126 VGND.n874 VGND.n873 0.145386
R6127 VGND.n869 VGND.n868 0.145386
R6128 VGND.n864 VGND.n863 0.145386
R6129 VGND.n859 VGND.n858 0.145386
R6130 VGND.n854 VGND.n853 0.145386
R6131 VGND.n849 VGND.n848 0.145386
R6132 VGND.n844 VGND.n843 0.145386
R6133 VGND.n2401 VGND.n2400 0.145386
R6134 VGND.n2405 VGND.n2404 0.145386
R6135 VGND.n1124 VGND.n1123 0.145386
R6136 VGND.n1130 VGND.n1129 0.145386
R6137 VGND.n1134 VGND.n1133 0.145386
R6138 VGND.n1143 VGND.n1142 0.145386
R6139 VGND.n1146 VGND.n810 0.145386
R6140 VGND.n1162 VGND.n1161 0.145386
R6141 VGND.n1166 VGND.n1165 0.145386
R6142 VGND.n1175 VGND.n1174 0.145386
R6143 VGND.n1178 VGND.n802 0.145386
R6144 VGND.n1194 VGND.n1193 0.145386
R6145 VGND.n1198 VGND.n1197 0.145386
R6146 VGND.n1207 VGND.n1206 0.145386
R6147 VGND.n1210 VGND.n794 0.145386
R6148 VGND.n1226 VGND.n1225 0.145386
R6149 VGND.n1230 VGND.n1229 0.145386
R6150 VGND.n1288 VGND.n1287 0.145386
R6151 VGND.n683 VGND.n679 0.145386
R6152 VGND.n724 VGND.n723 0.145386
R6153 VGND.n729 VGND.n728 0.145386
R6154 VGND.n734 VGND.n733 0.145386
R6155 VGND.n739 VGND.n738 0.145386
R6156 VGND.n744 VGND.n743 0.145386
R6157 VGND.n749 VGND.n748 0.145386
R6158 VGND.n754 VGND.n753 0.145386
R6159 VGND.n759 VGND.n758 0.145386
R6160 VGND.n764 VGND.n763 0.145386
R6161 VGND.n769 VGND.n768 0.145386
R6162 VGND.n774 VGND.n773 0.145386
R6163 VGND.n779 VGND.n778 0.145386
R6164 VGND.n782 VGND.n719 0.145386
R6165 VGND.n1100 VGND.n1094 0.144904
R6166 VGND.n1073 VGND.n1065 0.144904
R6167 VGND.n1011 VGND.n1003 0.144904
R6168 VGND.n1042 VGND.n1034 0.144904
R6169 VGND.n2567 VGND.n2566 0.138284
R6170 VGND.n232 VGND.n231 0.122659
R6171 VGND.n2702 VGND.n2701 0.122659
R6172 VGND.n2707 VGND.n2706 0.122659
R6173 VGND.n2712 VGND.n2711 0.122659
R6174 VGND.n2717 VGND.n2716 0.122659
R6175 VGND.n2722 VGND.n2721 0.122659
R6176 VGND.n2727 VGND.n2726 0.122659
R6177 VGND.n2732 VGND.n2731 0.122659
R6178 VGND.n2737 VGND.n2736 0.122659
R6179 VGND.n2742 VGND.n2741 0.122659
R6180 VGND.n2747 VGND.n2746 0.122659
R6181 VGND.n2752 VGND.n2751 0.122659
R6182 VGND.n2757 VGND.n2756 0.122659
R6183 VGND.n2762 VGND.n2761 0.122659
R6184 VGND.n227 VGND.n226 0.122659
R6185 VGND.n242 VGND.n241 0.122659
R6186 VGND.n2511 VGND.n2510 0.122659
R6187 VGND.n2506 VGND.n2505 0.122659
R6188 VGND.n247 VGND.n246 0.122659
R6189 VGND.n2436 VGND.n2435 0.122659
R6190 VGND.n2441 VGND.n2440 0.122659
R6191 VGND.n2446 VGND.n2445 0.122659
R6192 VGND.n2451 VGND.n2450 0.122659
R6193 VGND.n2456 VGND.n2455 0.122659
R6194 VGND.n2461 VGND.n2460 0.122659
R6195 VGND.n2466 VGND.n2465 0.122659
R6196 VGND.n2471 VGND.n2470 0.122659
R6197 VGND.n2476 VGND.n2475 0.122659
R6198 VGND.n2481 VGND.n2480 0.122659
R6199 VGND.n2486 VGND.n2485 0.122659
R6200 VGND.n2814 VGND.n2813 0.122659
R6201 VGND.n367 VGND.n366 0.122659
R6202 VGND.n370 VGND.n369 0.122659
R6203 VGND.n2169 VGND.n2168 0.122659
R6204 VGND.n364 VGND.n363 0.122659
R6205 VGND.n2195 VGND.n2194 0.122659
R6206 VGND.n356 VGND.n355 0.122659
R6207 VGND.n2221 VGND.n2220 0.122659
R6208 VGND.n348 VGND.n347 0.122659
R6209 VGND.n2247 VGND.n2246 0.122659
R6210 VGND.n340 VGND.n339 0.122659
R6211 VGND.n2278 VGND.n2277 0.122659
R6212 VGND.n2283 VGND.n2282 0.122659
R6213 VGND.n2288 VGND.n2287 0.122659
R6214 VGND.n332 VGND.n331 0.122659
R6215 VGND.n1426 VGND.n1425 0.122659
R6216 VGND.n1423 VGND.n1422 0.122659
R6217 VGND.n2156 VGND.n2155 0.122659
R6218 VGND.n379 VGND.n378 0.122659
R6219 VGND.n2182 VGND.n2181 0.122659
R6220 VGND.n360 VGND.n359 0.122659
R6221 VGND.n2208 VGND.n2207 0.122659
R6222 VGND.n352 VGND.n351 0.122659
R6223 VGND.n2234 VGND.n2233 0.122659
R6224 VGND.n344 VGND.n343 0.122659
R6225 VGND.n2260 VGND.n2259 0.122659
R6226 VGND.n336 VGND.n335 0.122659
R6227 VGND.n2265 VGND.n2264 0.122659
R6228 VGND.n2305 VGND.n2304 0.122659
R6229 VGND.n2311 VGND.n2310 0.122659
R6230 VGND.n1440 VGND.n1439 0.122659
R6231 VGND.n634 VGND.n633 0.122659
R6232 VGND.n1490 VGND.n1489 0.122659
R6233 VGND.n1485 VGND.n1484 0.122659
R6234 VGND.n1480 VGND.n1479 0.122659
R6235 VGND.n1475 VGND.n1474 0.122659
R6236 VGND.n1470 VGND.n1469 0.122659
R6237 VGND.n1465 VGND.n1464 0.122659
R6238 VGND.n1460 VGND.n1459 0.122659
R6239 VGND.n1455 VGND.n1454 0.122659
R6240 VGND.n1450 VGND.n1449 0.122659
R6241 VGND.n1445 VGND.n1444 0.122659
R6242 VGND.n393 VGND.n392 0.122659
R6243 VGND.n2133 VGND.n2132 0.122659
R6244 VGND.n2128 VGND.n2127 0.122659
R6245 VGND.n1502 VGND.n1501 0.122659
R6246 VGND.n622 VGND.n621 0.122659
R6247 VGND.n625 VGND.n624 0.122659
R6248 VGND.n1995 VGND.n1994 0.122659
R6249 VGND.n431 VGND.n430 0.122659
R6250 VGND.n2021 VGND.n2020 0.122659
R6251 VGND.n423 VGND.n422 0.122659
R6252 VGND.n2047 VGND.n2046 0.122659
R6253 VGND.n415 VGND.n414 0.122659
R6254 VGND.n2073 VGND.n2072 0.122659
R6255 VGND.n407 VGND.n406 0.122659
R6256 VGND.n2104 VGND.n2103 0.122659
R6257 VGND.n2109 VGND.n2108 0.122659
R6258 VGND.n2114 VGND.n2113 0.122659
R6259 VGND.n2120 VGND.n2119 0.122659
R6260 VGND.n650 VGND.n649 0.122659
R6261 VGND.n647 VGND.n646 0.122659
R6262 VGND.n1982 VGND.n1981 0.122659
R6263 VGND.n435 VGND.n434 0.122659
R6264 VGND.n2008 VGND.n2007 0.122659
R6265 VGND.n427 VGND.n426 0.122659
R6266 VGND.n2034 VGND.n2033 0.122659
R6267 VGND.n419 VGND.n418 0.122659
R6268 VGND.n2060 VGND.n2059 0.122659
R6269 VGND.n411 VGND.n410 0.122659
R6270 VGND.n2086 VGND.n2085 0.122659
R6271 VGND.n403 VGND.n402 0.122659
R6272 VGND.n2091 VGND.n2090 0.122659
R6273 VGND.n2330 VGND.n2329 0.122659
R6274 VGND.n2336 VGND.n2335 0.122659
R6275 VGND.n957 VGND.n956 0.122659
R6276 VGND.n952 VGND.n951 0.122659
R6277 VGND.n947 VGND.n946 0.122659
R6278 VGND.n942 VGND.n941 0.122659
R6279 VGND.n937 VGND.n936 0.122659
R6280 VGND.n932 VGND.n931 0.122659
R6281 VGND.n927 VGND.n926 0.122659
R6282 VGND.n922 VGND.n921 0.122659
R6283 VGND.n917 VGND.n916 0.122659
R6284 VGND.n912 VGND.n911 0.122659
R6285 VGND.n907 VGND.n906 0.122659
R6286 VGND.n902 VGND.n901 0.122659
R6287 VGND.n449 VGND.n448 0.122659
R6288 VGND.n1959 VGND.n1958 0.122659
R6289 VGND.n1954 VGND.n1953 0.122659
R6290 VGND.n1393 VGND.n1392 0.122659
R6291 VGND.n1398 VGND.n1397 0.122659
R6292 VGND.n666 VGND.n665 0.122659
R6293 VGND.n1821 VGND.n1820 0.122659
R6294 VGND.n487 VGND.n486 0.122659
R6295 VGND.n1847 VGND.n1846 0.122659
R6296 VGND.n479 VGND.n478 0.122659
R6297 VGND.n1873 VGND.n1872 0.122659
R6298 VGND.n471 VGND.n470 0.122659
R6299 VGND.n1899 VGND.n1898 0.122659
R6300 VGND.n463 VGND.n462 0.122659
R6301 VGND.n1930 VGND.n1929 0.122659
R6302 VGND.n1935 VGND.n1934 0.122659
R6303 VGND.n1940 VGND.n1939 0.122659
R6304 VGND.n1946 VGND.n1945 0.122659
R6305 VGND.n1378 VGND.n1377 0.122659
R6306 VGND.n1375 VGND.n1374 0.122659
R6307 VGND.n1808 VGND.n1807 0.122659
R6308 VGND.n491 VGND.n490 0.122659
R6309 VGND.n1834 VGND.n1833 0.122659
R6310 VGND.n483 VGND.n482 0.122659
R6311 VGND.n1860 VGND.n1859 0.122659
R6312 VGND.n475 VGND.n474 0.122659
R6313 VGND.n1886 VGND.n1885 0.122659
R6314 VGND.n467 VGND.n466 0.122659
R6315 VGND.n1912 VGND.n1911 0.122659
R6316 VGND.n459 VGND.n458 0.122659
R6317 VGND.n1917 VGND.n1916 0.122659
R6318 VGND.n2355 VGND.n2354 0.122659
R6319 VGND.n2361 VGND.n2360 0.122659
R6320 VGND.n1310 VGND.n1309 0.122659
R6321 VGND.n1307 VGND.n1306 0.122659
R6322 VGND.n1360 VGND.n1359 0.122659
R6323 VGND.n1355 VGND.n1354 0.122659
R6324 VGND.n1350 VGND.n1349 0.122659
R6325 VGND.n1345 VGND.n1344 0.122659
R6326 VGND.n1340 VGND.n1339 0.122659
R6327 VGND.n1335 VGND.n1334 0.122659
R6328 VGND.n1330 VGND.n1329 0.122659
R6329 VGND.n1325 VGND.n1324 0.122659
R6330 VGND.n1320 VGND.n1319 0.122659
R6331 VGND.n1315 VGND.n1314 0.122659
R6332 VGND.n505 VGND.n504 0.122659
R6333 VGND.n1785 VGND.n1784 0.122659
R6334 VGND.n1780 VGND.n1779 0.122659
R6335 VGND.n1515 VGND.n1514 0.122659
R6336 VGND.n1520 VGND.n1519 0.122659
R6337 VGND.n577 VGND.n576 0.122659
R6338 VGND.n1647 VGND.n1646 0.122659
R6339 VGND.n543 VGND.n542 0.122659
R6340 VGND.n1673 VGND.n1672 0.122659
R6341 VGND.n535 VGND.n534 0.122659
R6342 VGND.n1699 VGND.n1698 0.122659
R6343 VGND.n527 VGND.n526 0.122659
R6344 VGND.n1725 VGND.n1724 0.122659
R6345 VGND.n519 VGND.n518 0.122659
R6346 VGND.n1756 VGND.n1755 0.122659
R6347 VGND.n1761 VGND.n1760 0.122659
R6348 VGND.n1766 VGND.n1765 0.122659
R6349 VGND.n1772 VGND.n1771 0.122659
R6350 VGND.n1535 VGND.n1534 0.122659
R6351 VGND.n566 VGND.n565 0.122659
R6352 VGND.n1634 VGND.n1633 0.122659
R6353 VGND.n547 VGND.n546 0.122659
R6354 VGND.n1660 VGND.n1659 0.122659
R6355 VGND.n539 VGND.n538 0.122659
R6356 VGND.n1686 VGND.n1685 0.122659
R6357 VGND.n531 VGND.n530 0.122659
R6358 VGND.n1712 VGND.n1711 0.122659
R6359 VGND.n523 VGND.n522 0.122659
R6360 VGND.n1738 VGND.n1737 0.122659
R6361 VGND.n515 VGND.n514 0.122659
R6362 VGND.n1743 VGND.n1742 0.122659
R6363 VGND.n2380 VGND.n2379 0.122659
R6364 VGND.n2386 VGND.n2385 0.122659
R6365 VGND.n674 VGND.n673 0.122659
R6366 VGND.n1548 VGND.n1547 0.122659
R6367 VGND.n1553 VGND.n1552 0.122659
R6368 VGND.n1558 VGND.n1557 0.122659
R6369 VGND.n1563 VGND.n1562 0.122659
R6370 VGND.n1568 VGND.n1567 0.122659
R6371 VGND.n1573 VGND.n1572 0.122659
R6372 VGND.n1578 VGND.n1577 0.122659
R6373 VGND.n1583 VGND.n1582 0.122659
R6374 VGND.n1588 VGND.n1587 0.122659
R6375 VGND.n1593 VGND.n1592 0.122659
R6376 VGND.n1598 VGND.n1597 0.122659
R6377 VGND.n561 VGND.n560 0.122659
R6378 VGND.n1611 VGND.n1610 0.122659
R6379 VGND.n1606 VGND.n1605 0.122659
R6380 VGND.n833 VGND.n832 0.122659
R6381 VGND.n838 VGND.n837 0.122659
R6382 VGND.n830 VGND.n829 0.122659
R6383 VGND.n888 VGND.n887 0.122659
R6384 VGND.n883 VGND.n882 0.122659
R6385 VGND.n878 VGND.n877 0.122659
R6386 VGND.n873 VGND.n872 0.122659
R6387 VGND.n868 VGND.n867 0.122659
R6388 VGND.n863 VGND.n862 0.122659
R6389 VGND.n858 VGND.n857 0.122659
R6390 VGND.n853 VGND.n852 0.122659
R6391 VGND.n848 VGND.n847 0.122659
R6392 VGND.n843 VGND.n842 0.122659
R6393 VGND.n2400 VGND.n2399 0.122659
R6394 VGND.n2406 VGND.n2405 0.122659
R6395 VGND.n1125 VGND.n1124 0.122659
R6396 VGND.n1129 VGND.n1128 0.122659
R6397 VGND.n1135 VGND.n1134 0.122659
R6398 VGND.n1142 VGND.n1141 0.122659
R6399 VGND.n810 VGND.n809 0.122659
R6400 VGND.n1161 VGND.n1160 0.122659
R6401 VGND.n1167 VGND.n1166 0.122659
R6402 VGND.n1174 VGND.n1173 0.122659
R6403 VGND.n802 VGND.n801 0.122659
R6404 VGND.n1193 VGND.n1192 0.122659
R6405 VGND.n1199 VGND.n1198 0.122659
R6406 VGND.n1206 VGND.n1205 0.122659
R6407 VGND.n794 VGND.n793 0.122659
R6408 VGND.n1225 VGND.n1224 0.122659
R6409 VGND.n1231 VGND.n1230 0.122659
R6410 VGND.n1287 VGND.n1286 0.122659
R6411 VGND.n684 VGND.n683 0.122659
R6412 VGND.n723 VGND.n722 0.122659
R6413 VGND.n728 VGND.n727 0.122659
R6414 VGND.n733 VGND.n732 0.122659
R6415 VGND.n738 VGND.n737 0.122659
R6416 VGND.n743 VGND.n742 0.122659
R6417 VGND.n748 VGND.n747 0.122659
R6418 VGND.n753 VGND.n752 0.122659
R6419 VGND.n758 VGND.n757 0.122659
R6420 VGND.n763 VGND.n762 0.122659
R6421 VGND.n768 VGND.n767 0.122659
R6422 VGND.n773 VGND.n772 0.122659
R6423 VGND.n778 VGND.n777 0.122659
R6424 VGND.n719 VGND.n718 0.122659
R6425 VGND VGND.n109 0.120838
R6426 VGND.n1108 VGND.n1107 0.120292
R6427 VGND.n1107 VGND.n1106 0.120292
R6428 VGND.n1106 VGND.n1092 0.120292
R6429 VGND.n1102 VGND.n1092 0.120292
R6430 VGND.n1102 VGND.n1101 0.120292
R6431 VGND.n1101 VGND.n1100 0.120292
R6432 VGND.n1086 VGND.n1085 0.120292
R6433 VGND.n1081 VGND.n1080 0.120292
R6434 VGND.n1080 VGND.n1079 0.120292
R6435 VGND.n1079 VGND.n1063 0.120292
R6436 VGND.n1075 VGND.n1063 0.120292
R6437 VGND.n1075 VGND.n1074 0.120292
R6438 VGND.n1074 VGND.n1073 0.120292
R6439 VGND.n143 VGND.n120 0.120292
R6440 VGND.n137 VGND.n120 0.120292
R6441 VGND.n137 VGND.n136 0.120292
R6442 VGND.n136 VGND.n124 0.120292
R6443 VGND.n129 VGND.n124 0.120292
R6444 VGND.n129 VGND.n128 0.120292
R6445 VGND.n128 VGND.n127 0.120292
R6446 VGND.n586 VGND.n583 0.120292
R6447 VGND.n587 VGND.n586 0.120292
R6448 VGND.n611 VGND.n588 0.120292
R6449 VGND.n605 VGND.n588 0.120292
R6450 VGND.n605 VGND.n604 0.120292
R6451 VGND.n604 VGND.n592 0.120292
R6452 VGND.n597 VGND.n592 0.120292
R6453 VGND.n597 VGND.n596 0.120292
R6454 VGND.n596 VGND.n595 0.120292
R6455 VGND.n994 VGND.n993 0.120292
R6456 VGND.n987 VGND.n963 0.120292
R6457 VGND.n982 VGND.n963 0.120292
R6458 VGND.n982 VGND.n981 0.120292
R6459 VGND.n978 VGND.n977 0.120292
R6460 VGND.n977 VGND.n972 0.120292
R6461 VGND.n973 VGND.n972 0.120292
R6462 VGND.n1024 VGND.n1023 0.120292
R6463 VGND.n1019 VGND.n1018 0.120292
R6464 VGND.n1018 VGND.n1017 0.120292
R6465 VGND.n1017 VGND.n1001 0.120292
R6466 VGND.n1013 VGND.n1001 0.120292
R6467 VGND.n1013 VGND.n1012 0.120292
R6468 VGND.n1012 VGND.n1011 0.120292
R6469 VGND.n1055 VGND.n1054 0.120292
R6470 VGND.n1050 VGND.n1049 0.120292
R6471 VGND.n1049 VGND.n1048 0.120292
R6472 VGND.n1048 VGND.n1032 0.120292
R6473 VGND.n1044 VGND.n1032 0.120292
R6474 VGND.n1044 VGND.n1043 0.120292
R6475 VGND.n1043 VGND.n1042 0.120292
R6476 VGND.n173 VGND.n150 0.120292
R6477 VGND.n167 VGND.n150 0.120292
R6478 VGND.n167 VGND.n166 0.120292
R6479 VGND.n166 VGND.n154 0.120292
R6480 VGND.n159 VGND.n154 0.120292
R6481 VGND.n159 VGND.n158 0.120292
R6482 VGND.n158 VGND.n157 0.120292
R6483 VGND.n15 VGND.n11 0.120292
R6484 VGND.n20 VGND.n11 0.120292
R6485 VGND.n21 VGND.n20 0.120292
R6486 VGND.n22 VGND.n21 0.120292
R6487 VGND.n22 VGND.n9 0.120292
R6488 VGND.n26 VGND.n9 0.120292
R6489 VGND.n27 VGND.n26 0.120292
R6490 VGND.n101 VGND.n93 0.120292
R6491 VGND.n102 VGND.n101 0.120292
R6492 VGND.n102 VGND.n87 0.120292
R6493 VGND.n107 VGND.n87 0.120292
R6494 VGND.n108 VGND.n107 0.120292
R6495 VGND.n2845 VGND.n2837 0.120292
R6496 VGND.n2846 VGND.n2845 0.120292
R6497 VGND.n2846 VGND.n2831 0.120292
R6498 VGND.n2851 VGND.n2831 0.120292
R6499 VGND.n2852 VGND.n2851 0.120292
R6500 VGND.n2877 VGND.n2869 0.120292
R6501 VGND.n2878 VGND.n2877 0.120292
R6502 VGND.n2878 VGND.n2863 0.120292
R6503 VGND.n2883 VGND.n2863 0.120292
R6504 VGND.n2884 VGND.n2883 0.120292
R6505 VGND.n2888 VGND.n2885 0.120292
R6506 VGND.n75 VGND.n68 0.120292
R6507 VGND.n76 VGND.n75 0.120292
R6508 VGND.n76 VGND.n63 0.120292
R6509 VGND.n81 VGND.n63 0.120292
R6510 VGND.n82 VGND.n81 0.120292
R6511 VGND.n2903 VGND.n60 0.120292
R6512 VGND.n2918 VGND.n2917 0.120292
R6513 VGND.n2918 VGND.n2910 0.120292
R6514 VGND.n2923 VGND.n2910 0.120292
R6515 VGND.n2924 VGND.n2923 0.120292
R6516 VGND.n2925 VGND.n2924 0.120292
R6517 VGND.n2925 VGND.n2908 0.120292
R6518 VGND.n2929 VGND.n2908 0.120292
R6519 VGND.n2931 VGND.n2905 0.120292
R6520 VGND.n2936 VGND.n2905 0.120292
R6521 VGND.n44 VGND.n38 0.120292
R6522 VGND.n49 VGND.n38 0.120292
R6523 VGND.n50 VGND.n49 0.120292
R6524 VGND.n51 VGND.n50 0.120292
R6525 VGND.n51 VGND.n36 0.120292
R6526 VGND.n55 VGND.n36 0.120292
R6527 VGND.n56 VGND.n55 0.120292
R6528 VGND.n2943 VGND.n2942 0.120292
R6529 VGND.n2942 VGND.n2941 0.120292
R6530 VGND.n2957 VGND.n2951 0.120292
R6531 VGND.n2962 VGND.n2951 0.120292
R6532 VGND.n2963 VGND.n2962 0.120292
R6533 VGND.n2964 VGND.n2963 0.120292
R6534 VGND.n2964 VGND.n2949 0.120292
R6535 VGND.n2968 VGND.n2949 0.120292
R6536 VGND.n2969 VGND.n2968 0.120292
R6537 VGND.n2975 VGND.n2974 0.120292
R6538 VGND.n2974 VGND.n2973 0.120292
R6539 VGND VGND.n2855 0.119536
R6540 VGND.n1094 VGND 0.117202
R6541 VGND.n1065 VGND 0.117202
R6542 VGND.n1003 VGND 0.117202
R6543 VGND.n1034 VGND 0.117202
R6544 VGND.n1086 VGND 0.0981562
R6545 VGND.n994 VGND 0.0981562
R6546 VGND.n1055 VGND 0.0981562
R6547 VGND VGND.n143 0.0968542
R6548 VGND VGND.n611 0.0968542
R6549 VGND VGND.n987 0.0968542
R6550 VGND.n1024 VGND 0.0968542
R6551 VGND VGND.n173 0.0968542
R6552 VGND.n15 VGND 0.0968542
R6553 VGND VGND.n2888 0.0968542
R6554 VGND VGND.n60 0.0968542
R6555 VGND.n2917 VGND 0.0968542
R6556 VGND.n44 VGND 0.0968542
R6557 VGND.n2957 VGND 0.0968542
R6558 VGND.n2520 VGND 0.088625
R6559 VGND.n2695 VGND 0.0790114
R6560 VGND VGND.n2694 0.0790114
R6561 VGND VGND.n188 0.0790114
R6562 VGND.n2801 VGND 0.0790114
R6563 VGND VGND.n2800 0.0790114
R6564 VGND.n2795 VGND 0.0790114
R6565 VGND VGND.n2794 0.0790114
R6566 VGND.n2789 VGND 0.0790114
R6567 VGND VGND.n2788 0.0790114
R6568 VGND.n2783 VGND 0.0790114
R6569 VGND VGND.n2782 0.0790114
R6570 VGND.n2777 VGND 0.0790114
R6571 VGND VGND.n2776 0.0790114
R6572 VGND.n2771 VGND 0.0790114
R6573 VGND VGND.n2770 0.0790114
R6574 VGND.n2988 VGND 0.0790114
R6575 VGND.n2697 VGND 0.0790114
R6576 VGND.n2698 VGND 0.0790114
R6577 VGND.n2804 VGND 0.0790114
R6578 VGND VGND.n2803 0.0790114
R6579 VGND.n2798 VGND 0.0790114
R6580 VGND VGND.n2797 0.0790114
R6581 VGND.n2792 VGND 0.0790114
R6582 VGND VGND.n2791 0.0790114
R6583 VGND.n2786 VGND 0.0790114
R6584 VGND VGND.n2785 0.0790114
R6585 VGND.n2780 VGND 0.0790114
R6586 VGND VGND.n2779 0.0790114
R6587 VGND.n2774 VGND 0.0790114
R6588 VGND VGND.n2773 0.0790114
R6589 VGND.n2768 VGND 0.0790114
R6590 VGND.n2986 VGND 0.0790114
R6591 VGND VGND.n2517 0.0790114
R6592 VGND.n2808 VGND 0.0790114
R6593 VGND VGND.n2807 0.0790114
R6594 VGND.n2503 VGND 0.0790114
R6595 VGND VGND.n2502 0.0790114
R6596 VGND VGND.n2501 0.0790114
R6597 VGND VGND.n2500 0.0790114
R6598 VGND VGND.n2499 0.0790114
R6599 VGND VGND.n2498 0.0790114
R6600 VGND VGND.n2497 0.0790114
R6601 VGND VGND.n2496 0.0790114
R6602 VGND VGND.n2495 0.0790114
R6603 VGND VGND.n2494 0.0790114
R6604 VGND VGND.n2493 0.0790114
R6605 VGND VGND.n2492 0.0790114
R6606 VGND VGND.n2491 0.0790114
R6607 VGND.n639 VGND 0.0790114
R6608 VGND.n2811 VGND 0.0790114
R6609 VGND.n375 VGND 0.0790114
R6610 VGND.n2165 VGND 0.0790114
R6611 VGND.n2175 VGND 0.0790114
R6612 VGND.n2191 VGND 0.0790114
R6613 VGND.n2201 VGND 0.0790114
R6614 VGND.n2217 VGND 0.0790114
R6615 VGND.n2227 VGND 0.0790114
R6616 VGND.n2243 VGND 0.0790114
R6617 VGND.n2253 VGND 0.0790114
R6618 VGND.n2274 VGND 0.0790114
R6619 VGND.n2297 VGND 0.0790114
R6620 VGND VGND.n2296 0.0790114
R6621 VGND VGND.n2294 0.0790114
R6622 VGND.n2430 VGND 0.0790114
R6623 VGND.n1433 VGND 0.0790114
R6624 VGND VGND.n1432 0.0790114
R6625 VGND.n2152 VGND 0.0790114
R6626 VGND.n2162 VGND 0.0790114
R6627 VGND.n2178 VGND 0.0790114
R6628 VGND.n2188 VGND 0.0790114
R6629 VGND.n2204 VGND 0.0790114
R6630 VGND.n2214 VGND 0.0790114
R6631 VGND.n2230 VGND 0.0790114
R6632 VGND.n2240 VGND 0.0790114
R6633 VGND.n2256 VGND 0.0790114
R6634 VGND.n2271 VGND 0.0790114
R6635 VGND.n2300 VGND 0.0790114
R6636 VGND.n2301 VGND 0.0790114
R6637 VGND.n2314 VGND 0.0790114
R6638 VGND VGND.n2313 0.0790114
R6639 VGND.n1436 VGND 0.0790114
R6640 VGND.n1496 VGND 0.0790114
R6641 VGND.n2149 VGND 0.0790114
R6642 VGND VGND.n2148 0.0790114
R6643 VGND VGND.n2147 0.0790114
R6644 VGND VGND.n2146 0.0790114
R6645 VGND VGND.n2145 0.0790114
R6646 VGND VGND.n2144 0.0790114
R6647 VGND VGND.n2143 0.0790114
R6648 VGND VGND.n2142 0.0790114
R6649 VGND VGND.n2141 0.0790114
R6650 VGND VGND.n2140 0.0790114
R6651 VGND VGND.n2139 0.0790114
R6652 VGND.n2318 VGND 0.0790114
R6653 VGND VGND.n2317 0.0790114
R6654 VGND.n2125 VGND 0.0790114
R6655 VGND VGND.n1414 0.0790114
R6656 VGND.n1499 VGND 0.0790114
R6657 VGND VGND.n630 0.0790114
R6658 VGND.n1991 VGND 0.0790114
R6659 VGND.n2001 VGND 0.0790114
R6660 VGND.n2017 VGND 0.0790114
R6661 VGND.n2027 VGND 0.0790114
R6662 VGND.n2043 VGND 0.0790114
R6663 VGND.n2053 VGND 0.0790114
R6664 VGND.n2069 VGND 0.0790114
R6665 VGND.n2079 VGND 0.0790114
R6666 VGND.n2100 VGND 0.0790114
R6667 VGND.n2322 VGND 0.0790114
R6668 VGND VGND.n2321 0.0790114
R6669 VGND.n398 VGND 0.0790114
R6670 VGND.n2122 VGND 0.0790114
R6671 VGND VGND.n1412 0.0790114
R6672 VGND VGND.n656 0.0790114
R6673 VGND.n1978 VGND 0.0790114
R6674 VGND.n1988 VGND 0.0790114
R6675 VGND.n2004 VGND 0.0790114
R6676 VGND.n2014 VGND 0.0790114
R6677 VGND.n2030 VGND 0.0790114
R6678 VGND.n2040 VGND 0.0790114
R6679 VGND.n2056 VGND 0.0790114
R6680 VGND.n2066 VGND 0.0790114
R6681 VGND.n2082 VGND 0.0790114
R6682 VGND.n2097 VGND 0.0790114
R6683 VGND.n2325 VGND 0.0790114
R6684 VGND.n2326 VGND 0.0790114
R6685 VGND.n2339 VGND 0.0790114
R6686 VGND VGND.n2338 0.0790114
R6687 VGND.n1409 VGND 0.0790114
R6688 VGND VGND.n1408 0.0790114
R6689 VGND.n1975 VGND 0.0790114
R6690 VGND VGND.n1974 0.0790114
R6691 VGND VGND.n1973 0.0790114
R6692 VGND VGND.n1972 0.0790114
R6693 VGND VGND.n1971 0.0790114
R6694 VGND VGND.n1970 0.0790114
R6695 VGND VGND.n1969 0.0790114
R6696 VGND VGND.n1968 0.0790114
R6697 VGND VGND.n1967 0.0790114
R6698 VGND VGND.n1966 0.0790114
R6699 VGND VGND.n1965 0.0790114
R6700 VGND.n2343 VGND 0.0790114
R6701 VGND VGND.n2342 0.0790114
R6702 VGND.n1951 VGND 0.0790114
R6703 VGND.n1389 VGND 0.0790114
R6704 VGND.n1405 VGND 0.0790114
R6705 VGND VGND.n1404 0.0790114
R6706 VGND.n1817 VGND 0.0790114
R6707 VGND.n1827 VGND 0.0790114
R6708 VGND.n1843 VGND 0.0790114
R6709 VGND.n1853 VGND 0.0790114
R6710 VGND.n1869 VGND 0.0790114
R6711 VGND.n1879 VGND 0.0790114
R6712 VGND.n1895 VGND 0.0790114
R6713 VGND.n1905 VGND 0.0790114
R6714 VGND.n1926 VGND 0.0790114
R6715 VGND.n2347 VGND 0.0790114
R6716 VGND VGND.n2346 0.0790114
R6717 VGND.n454 VGND 0.0790114
R6718 VGND.n1948 VGND 0.0790114
R6719 VGND VGND.n1386 0.0790114
R6720 VGND VGND.n1384 0.0790114
R6721 VGND.n1804 VGND 0.0790114
R6722 VGND.n1814 VGND 0.0790114
R6723 VGND.n1830 VGND 0.0790114
R6724 VGND.n1840 VGND 0.0790114
R6725 VGND.n1856 VGND 0.0790114
R6726 VGND.n1866 VGND 0.0790114
R6727 VGND.n1882 VGND 0.0790114
R6728 VGND.n1892 VGND 0.0790114
R6729 VGND.n1908 VGND 0.0790114
R6730 VGND.n1923 VGND 0.0790114
R6731 VGND.n2350 VGND 0.0790114
R6732 VGND.n2351 VGND 0.0790114
R6733 VGND.n2364 VGND 0.0790114
R6734 VGND VGND.n2363 0.0790114
R6735 VGND VGND.n1368 0.0790114
R6736 VGND VGND.n1367 0.0790114
R6737 VGND.n1801 VGND 0.0790114
R6738 VGND VGND.n1800 0.0790114
R6739 VGND VGND.n1799 0.0790114
R6740 VGND VGND.n1798 0.0790114
R6741 VGND VGND.n1797 0.0790114
R6742 VGND VGND.n1796 0.0790114
R6743 VGND VGND.n1795 0.0790114
R6744 VGND VGND.n1794 0.0790114
R6745 VGND VGND.n1793 0.0790114
R6746 VGND VGND.n1792 0.0790114
R6747 VGND VGND.n1791 0.0790114
R6748 VGND.n2368 VGND 0.0790114
R6749 VGND VGND.n2367 0.0790114
R6750 VGND.n1777 VGND 0.0790114
R6751 VGND.n1528 VGND 0.0790114
R6752 VGND VGND.n1527 0.0790114
R6753 VGND VGND.n1526 0.0790114
R6754 VGND.n1643 VGND 0.0790114
R6755 VGND.n1653 VGND 0.0790114
R6756 VGND.n1669 VGND 0.0790114
R6757 VGND.n1679 VGND 0.0790114
R6758 VGND.n1695 VGND 0.0790114
R6759 VGND.n1705 VGND 0.0790114
R6760 VGND.n1721 VGND 0.0790114
R6761 VGND.n1731 VGND 0.0790114
R6762 VGND.n1752 VGND 0.0790114
R6763 VGND.n2372 VGND 0.0790114
R6764 VGND VGND.n2371 0.0790114
R6765 VGND.n510 VGND 0.0790114
R6766 VGND.n1774 VGND 0.0790114
R6767 VGND.n1531 VGND 0.0790114
R6768 VGND.n1541 VGND 0.0790114
R6769 VGND.n1630 VGND 0.0790114
R6770 VGND.n1640 VGND 0.0790114
R6771 VGND.n1656 VGND 0.0790114
R6772 VGND.n1666 VGND 0.0790114
R6773 VGND.n1682 VGND 0.0790114
R6774 VGND.n1692 VGND 0.0790114
R6775 VGND.n1708 VGND 0.0790114
R6776 VGND.n1718 VGND 0.0790114
R6777 VGND.n1734 VGND 0.0790114
R6778 VGND.n1749 VGND 0.0790114
R6779 VGND.n2375 VGND 0.0790114
R6780 VGND.n2376 VGND 0.0790114
R6781 VGND.n2389 VGND 0.0790114
R6782 VGND VGND.n2388 0.0790114
R6783 VGND VGND.n1298 0.0790114
R6784 VGND.n1544 VGND 0.0790114
R6785 VGND.n1627 VGND 0.0790114
R6786 VGND VGND.n1626 0.0790114
R6787 VGND VGND.n1625 0.0790114
R6788 VGND VGND.n1624 0.0790114
R6789 VGND VGND.n1623 0.0790114
R6790 VGND VGND.n1622 0.0790114
R6791 VGND VGND.n1621 0.0790114
R6792 VGND VGND.n1620 0.0790114
R6793 VGND VGND.n1619 0.0790114
R6794 VGND VGND.n1618 0.0790114
R6795 VGND VGND.n1617 0.0790114
R6796 VGND.n2393 VGND 0.0790114
R6797 VGND VGND.n2392 0.0790114
R6798 VGND.n1603 VGND 0.0790114
R6799 VGND.n896 VGND 0.0790114
R6800 VGND VGND.n895 0.0790114
R6801 VGND VGND.n894 0.0790114
R6802 VGND.n1275 VGND 0.0790114
R6803 VGND VGND.n1274 0.0790114
R6804 VGND.n1267 VGND 0.0790114
R6805 VGND VGND.n1266 0.0790114
R6806 VGND.n1259 VGND 0.0790114
R6807 VGND VGND.n1258 0.0790114
R6808 VGND.n1251 VGND 0.0790114
R6809 VGND VGND.n1250 0.0790114
R6810 VGND.n1243 VGND 0.0790114
R6811 VGND VGND.n1242 0.0790114
R6812 VGND.n2396 VGND 0.0790114
R6813 VGND.n284 VGND 0.0790114
R6814 VGND.n2408 VGND 0.0790114
R6815 VGND.n1119 VGND 0.0790114
R6816 VGND.n1282 VGND 0.0790114
R6817 VGND VGND.n1281 0.0790114
R6818 VGND.n687 VGND 0.0790114
R6819 VGND.n690 VGND 0.0790114
R6820 VGND.n693 VGND 0.0790114
R6821 VGND.n696 VGND 0.0790114
R6822 VGND.n699 VGND 0.0790114
R6823 VGND.n702 VGND 0.0790114
R6824 VGND.n705 VGND 0.0790114
R6825 VGND.n708 VGND 0.0790114
R6826 VGND.n711 VGND 0.0790114
R6827 VGND.n714 VGND 0.0790114
R6828 VGND.n1220 VGND 0.0790114
R6829 VGND.n1235 VGND 0.0790114
R6830 VGND VGND.n1234 0.0790114
R6831 VGND.n1117 VGND 0.0790114
R6832 VGND.n1284 VGND 0.0790114
R6833 VGND.n1279 VGND 0.0790114
R6834 VGND VGND.n1278 0.0790114
R6835 VGND.n1271 VGND 0.0790114
R6836 VGND VGND.n1270 0.0790114
R6837 VGND.n1263 VGND 0.0790114
R6838 VGND VGND.n1262 0.0790114
R6839 VGND.n1255 VGND 0.0790114
R6840 VGND VGND.n1254 0.0790114
R6841 VGND.n1247 VGND 0.0790114
R6842 VGND VGND.n1246 0.0790114
R6843 VGND.n1239 VGND 0.0790114
R6844 VGND VGND.n1238 0.0790114
R6845 VGND VGND.n1237 0.0790114
R6846 VGND.n2411 VGND 0.0790114
R6847 VGND.n3008 VGND.n3007 0.0732323
R6848 VGND.n2643 VGND.n2642 0.0729432
R6849 VGND.n2640 VGND.n2638 0.0729432
R6850 VGND.n2650 VGND.n2649 0.0729432
R6851 VGND.n2637 VGND.n2635 0.0729432
R6852 VGND.n2657 VGND.n2656 0.0729432
R6853 VGND.n2634 VGND.n2632 0.0729432
R6854 VGND.n2664 VGND.n2663 0.0729432
R6855 VGND.n2631 VGND.n2629 0.0729432
R6856 VGND.n2671 VGND.n2670 0.0729432
R6857 VGND.n2628 VGND.n2626 0.0729432
R6858 VGND.n2678 VGND.n2677 0.0729432
R6859 VGND.n2625 VGND.n2623 0.0729432
R6860 VGND.n2685 VGND.n2684 0.0729432
R6861 VGND.n2622 VGND.n2621 0.0729432
R6862 VGND.n2692 VGND.n2691 0.0729432
R6863 VGND.n2642 VGND 0.0612143
R6864 VGND.n2640 VGND 0.0612143
R6865 VGND.n2649 VGND 0.0612143
R6866 VGND.n2637 VGND 0.0612143
R6867 VGND.n2656 VGND 0.0612143
R6868 VGND.n2634 VGND 0.0612143
R6869 VGND.n2663 VGND 0.0612143
R6870 VGND.n2631 VGND 0.0612143
R6871 VGND.n2670 VGND 0.0612143
R6872 VGND.n2628 VGND 0.0612143
R6873 VGND.n2677 VGND 0.0612143
R6874 VGND.n2625 VGND 0.0612143
R6875 VGND.n2684 VGND 0.0612143
R6876 VGND.n2622 VGND 0.0612143
R6877 VGND.n2692 VGND 0.0612143
R6878 VGND.n2564 VGND 0.0608448
R6879 VGND.n2561 VGND 0.0608448
R6880 VGND.n2558 VGND 0.0608448
R6881 VGND.n2555 VGND 0.0608448
R6882 VGND.n2552 VGND 0.0608448
R6883 VGND.n2549 VGND 0.0608448
R6884 VGND.n2546 VGND 0.0608448
R6885 VGND.n2543 VGND 0.0608448
R6886 VGND.n2540 VGND 0.0608448
R6887 VGND.n2537 VGND 0.0608448
R6888 VGND.n2534 VGND 0.0608448
R6889 VGND.n2531 VGND 0.0608448
R6890 VGND.n2528 VGND 0.0608448
R6891 VGND.n2525 VGND 0.0608448
R6892 VGND.n2522 VGND 0.0608448
R6893 VGND.n1108 VGND 0.0603958
R6894 VGND.n1085 VGND 0.0603958
R6895 VGND VGND.n1084 0.0603958
R6896 VGND.n1081 VGND 0.0603958
R6897 VGND.n145 VGND 0.0603958
R6898 VGND VGND.n144 0.0603958
R6899 VGND.n127 VGND 0.0603958
R6900 VGND.n613 VGND 0.0603958
R6901 VGND VGND.n612 0.0603958
R6902 VGND.n595 VGND 0.0603958
R6903 VGND.n989 VGND 0.0603958
R6904 VGND VGND.n988 0.0603958
R6905 VGND.n981 VGND 0.0603958
R6906 VGND.n978 VGND 0.0603958
R6907 VGND.n973 VGND 0.0603958
R6908 VGND.n1023 VGND 0.0603958
R6909 VGND VGND.n1022 0.0603958
R6910 VGND.n1019 VGND 0.0603958
R6911 VGND.n1054 VGND 0.0603958
R6912 VGND VGND.n1053 0.0603958
R6913 VGND.n1050 VGND 0.0603958
R6914 VGND.n175 VGND 0.0603958
R6915 VGND VGND.n174 0.0603958
R6916 VGND.n157 VGND 0.0603958
R6917 VGND VGND.n27 0.0603958
R6918 VGND.n2991 VGND 0.0603958
R6919 VGND.n111 VGND 0.0603958
R6920 VGND VGND.n110 0.0603958
R6921 VGND.n2857 VGND 0.0603958
R6922 VGND VGND.n2856 0.0603958
R6923 VGND.n2890 VGND 0.0603958
R6924 VGND VGND.n2889 0.0603958
R6925 VGND.n2885 VGND 0.0603958
R6926 VGND.n2897 VGND 0.0603958
R6927 VGND.n2898 VGND 0.0603958
R6928 VGND VGND.n2929 0.0603958
R6929 VGND.n2930 VGND 0.0603958
R6930 VGND.n2931 VGND 0.0603958
R6931 VGND VGND.n56 0.0603958
R6932 VGND.n57 VGND 0.0603958
R6933 VGND.n2943 VGND 0.0603958
R6934 VGND VGND.n2969 0.0603958
R6935 VGND.n2970 VGND 0.0603958
R6936 VGND.n2975 VGND 0.0603958
R6937 VGND.n822 VGND 0.0489375
R6938 VGND.n785 VGND 0.0489375
R6939 VGND.n2579 VGND 0.0489375
R6940 VGND.n2576 VGND 0.0489375
R6941 VGND.n2581 VGND 0.0489375
R6942 VGND.n2584 VGND 0.0489375
R6943 VGND.n2587 VGND 0.0489375
R6944 VGND.n2590 VGND 0.0489375
R6945 VGND.n2593 VGND 0.0489375
R6946 VGND.n2596 VGND 0.0489375
R6947 VGND.n2599 VGND 0.0489375
R6948 VGND.n2602 VGND 0.0489375
R6949 VGND.n2605 VGND 0.0489375
R6950 VGND.n2608 VGND 0.0489375
R6951 VGND.n2611 VGND 0.0489375
R6952 VGND.n2614 VGND 0.0489375
R6953 VGND.n2575 VGND 0.0489375
R6954 VGND.n2568 VGND 0.0489375
R6955 VGND.n819 VGND 0.0489375
R6956 VGND.n816 VGND 0.0489375
R6957 VGND.n1136 VGND 0.0489375
R6958 VGND.n807 VGND 0.0489375
R6959 VGND.n805 VGND 0.0489375
R6960 VGND.n1151 VGND 0.0489375
R6961 VGND.n1168 VGND 0.0489375
R6962 VGND.n799 VGND 0.0489375
R6963 VGND.n797 VGND 0.0489375
R6964 VGND.n1183 VGND 0.0489375
R6965 VGND.n1200 VGND 0.0489375
R6966 VGND.n791 VGND 0.0489375
R6967 VGND.n789 VGND 0.0489375
R6968 VGND.n1215 VGND 0.0489375
R6969 VGND VGND.n2573 0.0360114
R6970 VGND VGND.n229 0.0360114
R6971 VGND.n231 VGND 0.0360114
R6972 VGND.n2701 VGND 0.0360114
R6973 VGND.n2706 VGND 0.0360114
R6974 VGND.n2711 VGND 0.0360114
R6975 VGND.n2716 VGND 0.0360114
R6976 VGND.n2721 VGND 0.0360114
R6977 VGND.n2726 VGND 0.0360114
R6978 VGND.n2731 VGND 0.0360114
R6979 VGND.n2736 VGND 0.0360114
R6980 VGND.n2741 VGND 0.0360114
R6981 VGND.n2746 VGND 0.0360114
R6982 VGND.n2751 VGND 0.0360114
R6983 VGND.n2756 VGND 0.0360114
R6984 VGND.n2761 VGND 0.0360114
R6985 VGND.n226 VGND 0.0360114
R6986 VGND VGND.n239 0.0360114
R6987 VGND.n241 VGND 0.0360114
R6988 VGND.n2510 VGND 0.0360114
R6989 VGND.n2505 VGND 0.0360114
R6990 VGND VGND.n247 0.0360114
R6991 VGND.n2435 VGND 0.0360114
R6992 VGND.n2440 VGND 0.0360114
R6993 VGND.n2445 VGND 0.0360114
R6994 VGND.n2450 VGND 0.0360114
R6995 VGND.n2455 VGND 0.0360114
R6996 VGND.n2460 VGND 0.0360114
R6997 VGND.n2465 VGND 0.0360114
R6998 VGND.n2470 VGND 0.0360114
R6999 VGND.n2475 VGND 0.0360114
R7000 VGND.n2480 VGND 0.0360114
R7001 VGND.n2485 VGND 0.0360114
R7002 VGND VGND.n179 0.0360114
R7003 VGND.n2813 VGND 0.0360114
R7004 VGND VGND.n367 0.0360114
R7005 VGND.n369 VGND 0.0360114
R7006 VGND.n2168 VGND 0.0360114
R7007 VGND.n363 VGND 0.0360114
R7008 VGND.n2194 VGND 0.0360114
R7009 VGND.n355 VGND 0.0360114
R7010 VGND.n2220 VGND 0.0360114
R7011 VGND.n347 VGND 0.0360114
R7012 VGND.n2246 VGND 0.0360114
R7013 VGND.n339 VGND 0.0360114
R7014 VGND.n2277 VGND 0.0360114
R7015 VGND.n2282 VGND 0.0360114
R7016 VGND.n2287 VGND 0.0360114
R7017 VGND.n331 VGND 0.0360114
R7018 VGND VGND.n1419 0.0360114
R7019 VGND.n1425 VGND 0.0360114
R7020 VGND.n1422 VGND 0.0360114
R7021 VGND.n2155 VGND 0.0360114
R7022 VGND.n378 VGND 0.0360114
R7023 VGND.n2181 VGND 0.0360114
R7024 VGND.n359 VGND 0.0360114
R7025 VGND.n2207 VGND 0.0360114
R7026 VGND.n351 VGND 0.0360114
R7027 VGND.n2233 VGND 0.0360114
R7028 VGND.n343 VGND 0.0360114
R7029 VGND.n2259 VGND 0.0360114
R7030 VGND.n335 VGND 0.0360114
R7031 VGND.n2264 VGND 0.0360114
R7032 VGND.n2304 VGND 0.0360114
R7033 VGND VGND.n2311 0.0360114
R7034 VGND VGND.n637 0.0360114
R7035 VGND.n1439 VGND 0.0360114
R7036 VGND.n633 VGND 0.0360114
R7037 VGND.n1489 VGND 0.0360114
R7038 VGND.n1484 VGND 0.0360114
R7039 VGND.n1479 VGND 0.0360114
R7040 VGND.n1474 VGND 0.0360114
R7041 VGND.n1469 VGND 0.0360114
R7042 VGND.n1464 VGND 0.0360114
R7043 VGND.n1459 VGND 0.0360114
R7044 VGND.n1454 VGND 0.0360114
R7045 VGND.n1449 VGND 0.0360114
R7046 VGND.n1444 VGND 0.0360114
R7047 VGND.n392 VGND 0.0360114
R7048 VGND.n2132 VGND 0.0360114
R7049 VGND.n2127 VGND 0.0360114
R7050 VGND VGND.n616 0.0360114
R7051 VGND.n1501 VGND 0.0360114
R7052 VGND VGND.n622 0.0360114
R7053 VGND.n624 VGND 0.0360114
R7054 VGND.n1994 VGND 0.0360114
R7055 VGND.n430 VGND 0.0360114
R7056 VGND.n2020 VGND 0.0360114
R7057 VGND.n422 VGND 0.0360114
R7058 VGND.n2046 VGND 0.0360114
R7059 VGND.n414 VGND 0.0360114
R7060 VGND.n2072 VGND 0.0360114
R7061 VGND.n406 VGND 0.0360114
R7062 VGND.n2103 VGND 0.0360114
R7063 VGND.n2108 VGND 0.0360114
R7064 VGND.n2113 VGND 0.0360114
R7065 VGND VGND.n2120 0.0360114
R7066 VGND VGND.n643 0.0360114
R7067 VGND.n649 VGND 0.0360114
R7068 VGND.n646 VGND 0.0360114
R7069 VGND.n1981 VGND 0.0360114
R7070 VGND.n434 VGND 0.0360114
R7071 VGND.n2007 VGND 0.0360114
R7072 VGND.n426 VGND 0.0360114
R7073 VGND.n2033 VGND 0.0360114
R7074 VGND.n418 VGND 0.0360114
R7075 VGND.n2059 VGND 0.0360114
R7076 VGND.n410 VGND 0.0360114
R7077 VGND.n2085 VGND 0.0360114
R7078 VGND.n402 VGND 0.0360114
R7079 VGND.n2090 VGND 0.0360114
R7080 VGND.n2329 VGND 0.0360114
R7081 VGND VGND.n2336 0.0360114
R7082 VGND VGND.n659 0.0360114
R7083 VGND.n956 VGND 0.0360114
R7084 VGND.n951 VGND 0.0360114
R7085 VGND.n946 VGND 0.0360114
R7086 VGND.n941 VGND 0.0360114
R7087 VGND.n936 VGND 0.0360114
R7088 VGND.n931 VGND 0.0360114
R7089 VGND.n926 VGND 0.0360114
R7090 VGND.n921 VGND 0.0360114
R7091 VGND.n916 VGND 0.0360114
R7092 VGND.n911 VGND 0.0360114
R7093 VGND.n906 VGND 0.0360114
R7094 VGND.n901 VGND 0.0360114
R7095 VGND.n448 VGND 0.0360114
R7096 VGND.n1958 VGND 0.0360114
R7097 VGND.n1953 VGND 0.0360114
R7098 VGND VGND.n668 0.0360114
R7099 VGND.n1392 VGND 0.0360114
R7100 VGND.n1397 VGND 0.0360114
R7101 VGND.n665 VGND 0.0360114
R7102 VGND.n1820 VGND 0.0360114
R7103 VGND.n486 VGND 0.0360114
R7104 VGND.n1846 VGND 0.0360114
R7105 VGND.n478 VGND 0.0360114
R7106 VGND.n1872 VGND 0.0360114
R7107 VGND.n470 VGND 0.0360114
R7108 VGND.n1898 VGND 0.0360114
R7109 VGND.n462 VGND 0.0360114
R7110 VGND.n1929 VGND 0.0360114
R7111 VGND.n1934 VGND 0.0360114
R7112 VGND.n1939 VGND 0.0360114
R7113 VGND VGND.n1946 0.0360114
R7114 VGND VGND.n1371 0.0360114
R7115 VGND.n1377 VGND 0.0360114
R7116 VGND.n1374 VGND 0.0360114
R7117 VGND.n1807 VGND 0.0360114
R7118 VGND.n490 VGND 0.0360114
R7119 VGND.n1833 VGND 0.0360114
R7120 VGND.n482 VGND 0.0360114
R7121 VGND.n1859 VGND 0.0360114
R7122 VGND.n474 VGND 0.0360114
R7123 VGND.n1885 VGND 0.0360114
R7124 VGND.n466 VGND 0.0360114
R7125 VGND.n1911 VGND 0.0360114
R7126 VGND.n458 VGND 0.0360114
R7127 VGND.n1916 VGND 0.0360114
R7128 VGND.n2354 VGND 0.0360114
R7129 VGND VGND.n2361 0.0360114
R7130 VGND VGND.n1303 0.0360114
R7131 VGND.n1309 VGND 0.0360114
R7132 VGND.n1306 VGND 0.0360114
R7133 VGND.n1359 VGND 0.0360114
R7134 VGND.n1354 VGND 0.0360114
R7135 VGND.n1349 VGND 0.0360114
R7136 VGND.n1344 VGND 0.0360114
R7137 VGND.n1339 VGND 0.0360114
R7138 VGND.n1334 VGND 0.0360114
R7139 VGND.n1329 VGND 0.0360114
R7140 VGND.n1324 VGND 0.0360114
R7141 VGND.n1319 VGND 0.0360114
R7142 VGND.n1314 VGND 0.0360114
R7143 VGND.n504 VGND 0.0360114
R7144 VGND.n1784 VGND 0.0360114
R7145 VGND.n1779 VGND 0.0360114
R7146 VGND VGND.n572 0.0360114
R7147 VGND.n1514 VGND 0.0360114
R7148 VGND.n1519 VGND 0.0360114
R7149 VGND.n576 VGND 0.0360114
R7150 VGND.n1646 VGND 0.0360114
R7151 VGND.n542 VGND 0.0360114
R7152 VGND.n1672 VGND 0.0360114
R7153 VGND.n534 VGND 0.0360114
R7154 VGND.n1698 VGND 0.0360114
R7155 VGND.n526 VGND 0.0360114
R7156 VGND.n1724 VGND 0.0360114
R7157 VGND.n518 VGND 0.0360114
R7158 VGND.n1755 VGND 0.0360114
R7159 VGND.n1760 VGND 0.0360114
R7160 VGND.n1765 VGND 0.0360114
R7161 VGND VGND.n1772 0.0360114
R7162 VGND VGND.n568 0.0360114
R7163 VGND.n1534 VGND 0.0360114
R7164 VGND.n565 VGND 0.0360114
R7165 VGND.n1633 VGND 0.0360114
R7166 VGND.n546 VGND 0.0360114
R7167 VGND.n1659 VGND 0.0360114
R7168 VGND.n538 VGND 0.0360114
R7169 VGND.n1685 VGND 0.0360114
R7170 VGND.n530 VGND 0.0360114
R7171 VGND.n1711 VGND 0.0360114
R7172 VGND.n522 VGND 0.0360114
R7173 VGND.n1737 VGND 0.0360114
R7174 VGND.n514 VGND 0.0360114
R7175 VGND.n1742 VGND 0.0360114
R7176 VGND.n2379 VGND 0.0360114
R7177 VGND VGND.n2386 0.0360114
R7178 VGND VGND.n671 0.0360114
R7179 VGND.n673 VGND 0.0360114
R7180 VGND.n1547 VGND 0.0360114
R7181 VGND.n1552 VGND 0.0360114
R7182 VGND.n1557 VGND 0.0360114
R7183 VGND.n1562 VGND 0.0360114
R7184 VGND.n1567 VGND 0.0360114
R7185 VGND.n1572 VGND 0.0360114
R7186 VGND.n1577 VGND 0.0360114
R7187 VGND.n1582 VGND 0.0360114
R7188 VGND.n1587 VGND 0.0360114
R7189 VGND.n1592 VGND 0.0360114
R7190 VGND.n1597 VGND 0.0360114
R7191 VGND.n560 VGND 0.0360114
R7192 VGND.n1610 VGND 0.0360114
R7193 VGND.n1605 VGND 0.0360114
R7194 VGND VGND.n825 0.0360114
R7195 VGND.n832 VGND 0.0360114
R7196 VGND.n837 VGND 0.0360114
R7197 VGND.n829 VGND 0.0360114
R7198 VGND.n887 VGND 0.0360114
R7199 VGND.n882 VGND 0.0360114
R7200 VGND.n877 VGND 0.0360114
R7201 VGND.n872 VGND 0.0360114
R7202 VGND.n867 VGND 0.0360114
R7203 VGND.n862 VGND 0.0360114
R7204 VGND.n857 VGND 0.0360114
R7205 VGND.n852 VGND 0.0360114
R7206 VGND.n847 VGND 0.0360114
R7207 VGND.n842 VGND 0.0360114
R7208 VGND.n2399 VGND 0.0360114
R7209 VGND VGND.n2406 0.0360114
R7210 VGND VGND.n815 0.0360114
R7211 VGND VGND.n1125 0.0360114
R7212 VGND.n1128 VGND 0.0360114
R7213 VGND VGND.n1135 0.0360114
R7214 VGND.n1141 VGND 0.0360114
R7215 VGND.n809 VGND 0.0360114
R7216 VGND.n1160 VGND 0.0360114
R7217 VGND VGND.n1167 0.0360114
R7218 VGND.n1173 VGND 0.0360114
R7219 VGND.n801 VGND 0.0360114
R7220 VGND.n1192 VGND 0.0360114
R7221 VGND VGND.n1199 0.0360114
R7222 VGND.n1205 VGND 0.0360114
R7223 VGND.n793 VGND 0.0360114
R7224 VGND.n1224 VGND 0.0360114
R7225 VGND VGND.n1231 0.0360114
R7226 VGND VGND.n676 0.0360114
R7227 VGND.n1286 VGND 0.0360114
R7228 VGND VGND.n684 0.0360114
R7229 VGND.n722 VGND 0.0360114
R7230 VGND.n727 VGND 0.0360114
R7231 VGND.n732 VGND 0.0360114
R7232 VGND.n737 VGND 0.0360114
R7233 VGND.n742 VGND 0.0360114
R7234 VGND.n747 VGND 0.0360114
R7235 VGND.n752 VGND 0.0360114
R7236 VGND.n757 VGND 0.0360114
R7237 VGND.n762 VGND 0.0360114
R7238 VGND.n767 VGND 0.0360114
R7239 VGND.n772 VGND 0.0360114
R7240 VGND.n777 VGND 0.0360114
R7241 VGND.n718 VGND 0.0360114
R7242 VGND.n1112 VGND 0.0343542
R7243 VGND.n1084 VGND 0.0343542
R7244 VGND.n145 VGND 0.0343542
R7245 VGND.n613 VGND 0.0343542
R7246 VGND.n989 VGND 0.0343542
R7247 VGND.n1022 VGND 0.0343542
R7248 VGND.n1053 VGND 0.0343542
R7249 VGND.n175 VGND 0.0343542
R7250 VGND.n2991 VGND 0.0330521
R7251 VGND.n111 VGND 0.0330521
R7252 VGND.n2857 VGND 0.0330521
R7253 VGND.n2890 VGND 0.0330521
R7254 VGND VGND.n2897 0.0330521
R7255 VGND VGND.n2930 0.0330521
R7256 VGND VGND.n57 0.0330521
R7257 VGND VGND.n2970 0.0330521
R7258 VGND.n2990 VGND 0.024
R7259 VGND.n1 VGND 0.024
R7260 VGND.n144 VGND 0.0239375
R7261 VGND.n612 VGND 0.0239375
R7262 VGND.n174 VGND 0.0239375
R7263 VGND.n2889 VGND 0.0239375
R7264 VGND.n2898 VGND 0.0239375
R7265 VGND.n1089 VGND 0.0226354
R7266 VGND VGND.n119 0.0226354
R7267 VGND.n997 VGND 0.0226354
R7268 VGND.n988 VGND 0.0226354
R7269 VGND.n1028 VGND 0.0226354
R7270 VGND VGND.n2903 0.0226354
R7271 VGND.n2941 VGND 0.0226354
R7272 VGND.n2973 VGND 0.0226354
R7273 VGND VGND.n587 0.0213333
R7274 VGND.n993 VGND 0.0213333
R7275 VGND.n1059 VGND 0.0213333
R7276 VGND VGND.n108 0.0213333
R7277 VGND.n110 VGND 0.0213333
R7278 VGND VGND.n2852 0.0213333
R7279 VGND.n2856 VGND 0.0213333
R7280 VGND VGND.n2884 0.0213333
R7281 VGND.n82 VGND 0.0213333
R7282 VGND VGND.n2936 0.0213333
R7283 VGND.n2990 VGND 0.0161667
R7284 VGND.n2574 VGND 0.0104432
R7285 VGND.n235 VGND 0.0104432
R7286 VGND.n2699 VGND 0.0104432
R7287 VGND VGND.n189 0.0104432
R7288 VGND VGND.n190 0.0104432
R7289 VGND VGND.n195 0.0104432
R7290 VGND VGND.n196 0.0104432
R7291 VGND VGND.n201 0.0104432
R7292 VGND VGND.n202 0.0104432
R7293 VGND VGND.n207 0.0104432
R7294 VGND VGND.n208 0.0104432
R7295 VGND VGND.n213 0.0104432
R7296 VGND VGND.n214 0.0104432
R7297 VGND VGND.n219 0.0104432
R7298 VGND VGND.n220 0.0104432
R7299 VGND.n2767 VGND 0.0104432
R7300 VGND.n2985 VGND 0.0104432
R7301 VGND.n2516 VGND 0.0104432
R7302 VGND VGND.n185 0.0104432
R7303 VGND VGND.n186 0.0104432
R7304 VGND VGND.n2504 0.0104432
R7305 VGND.n248 VGND 0.0104432
R7306 VGND VGND.n249 0.0104432
R7307 VGND VGND.n250 0.0104432
R7308 VGND VGND.n251 0.0104432
R7309 VGND VGND.n252 0.0104432
R7310 VGND VGND.n253 0.0104432
R7311 VGND VGND.n254 0.0104432
R7312 VGND VGND.n255 0.0104432
R7313 VGND VGND.n256 0.0104432
R7314 VGND VGND.n257 0.0104432
R7315 VGND VGND.n258 0.0104432
R7316 VGND.n2490 VGND 0.0104432
R7317 VGND.n180 VGND 0.0104432
R7318 VGND VGND.n2812 0.0104432
R7319 VGND.n374 VGND 0.0104432
R7320 VGND.n2166 VGND 0.0104432
R7321 VGND.n2174 VGND 0.0104432
R7322 VGND.n2192 VGND 0.0104432
R7323 VGND.n2200 VGND 0.0104432
R7324 VGND.n2218 VGND 0.0104432
R7325 VGND.n2226 VGND 0.0104432
R7326 VGND.n2244 VGND 0.0104432
R7327 VGND.n2252 VGND 0.0104432
R7328 VGND.n2275 VGND 0.0104432
R7329 VGND VGND.n328 0.0104432
R7330 VGND VGND.n329 0.0104432
R7331 VGND.n2293 VGND 0.0104432
R7332 VGND.n2429 VGND 0.0104432
R7333 VGND.n1420 VGND 0.0104432
R7334 VGND.n1431 VGND 0.0104432
R7335 VGND.n2153 VGND 0.0104432
R7336 VGND.n2161 VGND 0.0104432
R7337 VGND.n2179 VGND 0.0104432
R7338 VGND.n2187 VGND 0.0104432
R7339 VGND.n2205 VGND 0.0104432
R7340 VGND.n2213 VGND 0.0104432
R7341 VGND.n2231 VGND 0.0104432
R7342 VGND.n2239 VGND 0.0104432
R7343 VGND.n2257 VGND 0.0104432
R7344 VGND.n2270 VGND 0.0104432
R7345 VGND VGND.n327 0.0104432
R7346 VGND.n2302 VGND 0.0104432
R7347 VGND VGND.n324 0.0104432
R7348 VGND.n2312 VGND 0.0104432
R7349 VGND.n1437 VGND 0.0104432
R7350 VGND.n1495 VGND 0.0104432
R7351 VGND VGND.n381 0.0104432
R7352 VGND VGND.n382 0.0104432
R7353 VGND VGND.n383 0.0104432
R7354 VGND VGND.n384 0.0104432
R7355 VGND VGND.n385 0.0104432
R7356 VGND VGND.n386 0.0104432
R7357 VGND VGND.n387 0.0104432
R7358 VGND VGND.n388 0.0104432
R7359 VGND VGND.n389 0.0104432
R7360 VGND VGND.n390 0.0104432
R7361 VGND.n2138 VGND 0.0104432
R7362 VGND VGND.n321 0.0104432
R7363 VGND VGND.n322 0.0104432
R7364 VGND VGND.n2126 0.0104432
R7365 VGND.n617 VGND 0.0104432
R7366 VGND VGND.n1500 0.0104432
R7367 VGND.n629 VGND 0.0104432
R7368 VGND.n1992 VGND 0.0104432
R7369 VGND.n2000 VGND 0.0104432
R7370 VGND.n2018 VGND 0.0104432
R7371 VGND.n2026 VGND 0.0104432
R7372 VGND.n2044 VGND 0.0104432
R7373 VGND.n2052 VGND 0.0104432
R7374 VGND.n2070 VGND 0.0104432
R7375 VGND.n2078 VGND 0.0104432
R7376 VGND.n2101 VGND 0.0104432
R7377 VGND VGND.n318 0.0104432
R7378 VGND VGND.n319 0.0104432
R7379 VGND VGND.n399 0.0104432
R7380 VGND.n2121 VGND 0.0104432
R7381 VGND.n644 VGND 0.0104432
R7382 VGND.n655 VGND 0.0104432
R7383 VGND.n1979 VGND 0.0104432
R7384 VGND.n1987 VGND 0.0104432
R7385 VGND.n2005 VGND 0.0104432
R7386 VGND.n2013 VGND 0.0104432
R7387 VGND.n2031 VGND 0.0104432
R7388 VGND.n2039 VGND 0.0104432
R7389 VGND.n2057 VGND 0.0104432
R7390 VGND.n2065 VGND 0.0104432
R7391 VGND.n2083 VGND 0.0104432
R7392 VGND.n2096 VGND 0.0104432
R7393 VGND VGND.n316 0.0104432
R7394 VGND.n2327 VGND 0.0104432
R7395 VGND VGND.n312 0.0104432
R7396 VGND.n2337 VGND 0.0104432
R7397 VGND.n660 VGND 0.0104432
R7398 VGND VGND.n661 0.0104432
R7399 VGND VGND.n437 0.0104432
R7400 VGND VGND.n438 0.0104432
R7401 VGND VGND.n439 0.0104432
R7402 VGND VGND.n440 0.0104432
R7403 VGND VGND.n441 0.0104432
R7404 VGND VGND.n442 0.0104432
R7405 VGND VGND.n443 0.0104432
R7406 VGND VGND.n444 0.0104432
R7407 VGND VGND.n445 0.0104432
R7408 VGND VGND.n446 0.0104432
R7409 VGND.n1964 VGND 0.0104432
R7410 VGND VGND.n309 0.0104432
R7411 VGND VGND.n310 0.0104432
R7412 VGND VGND.n1952 0.0104432
R7413 VGND.n1390 VGND 0.0104432
R7414 VGND VGND.n663 0.0104432
R7415 VGND.n1403 VGND 0.0104432
R7416 VGND.n1818 VGND 0.0104432
R7417 VGND.n1826 VGND 0.0104432
R7418 VGND.n1844 VGND 0.0104432
R7419 VGND.n1852 VGND 0.0104432
R7420 VGND.n1870 VGND 0.0104432
R7421 VGND.n1878 VGND 0.0104432
R7422 VGND.n1896 VGND 0.0104432
R7423 VGND.n1904 VGND 0.0104432
R7424 VGND.n1927 VGND 0.0104432
R7425 VGND VGND.n306 0.0104432
R7426 VGND VGND.n307 0.0104432
R7427 VGND VGND.n455 0.0104432
R7428 VGND.n1947 VGND 0.0104432
R7429 VGND.n1372 VGND 0.0104432
R7430 VGND.n1383 VGND 0.0104432
R7431 VGND.n1805 VGND 0.0104432
R7432 VGND.n1813 VGND 0.0104432
R7433 VGND.n1831 VGND 0.0104432
R7434 VGND.n1839 VGND 0.0104432
R7435 VGND.n1857 VGND 0.0104432
R7436 VGND.n1865 VGND 0.0104432
R7437 VGND.n1883 VGND 0.0104432
R7438 VGND.n1891 VGND 0.0104432
R7439 VGND.n1909 VGND 0.0104432
R7440 VGND.n1922 VGND 0.0104432
R7441 VGND VGND.n304 0.0104432
R7442 VGND.n2352 VGND 0.0104432
R7443 VGND VGND.n300 0.0104432
R7444 VGND.n2362 VGND 0.0104432
R7445 VGND.n1304 VGND 0.0104432
R7446 VGND.n1365 VGND 0.0104432
R7447 VGND VGND.n493 0.0104432
R7448 VGND VGND.n494 0.0104432
R7449 VGND VGND.n495 0.0104432
R7450 VGND VGND.n496 0.0104432
R7451 VGND VGND.n497 0.0104432
R7452 VGND VGND.n498 0.0104432
R7453 VGND VGND.n499 0.0104432
R7454 VGND VGND.n500 0.0104432
R7455 VGND VGND.n501 0.0104432
R7456 VGND VGND.n502 0.0104432
R7457 VGND.n1790 VGND 0.0104432
R7458 VGND VGND.n297 0.0104432
R7459 VGND VGND.n298 0.0104432
R7460 VGND VGND.n1778 0.0104432
R7461 VGND.n573 VGND 0.0104432
R7462 VGND VGND.n574 0.0104432
R7463 VGND.n1525 VGND 0.0104432
R7464 VGND.n1644 VGND 0.0104432
R7465 VGND.n1652 VGND 0.0104432
R7466 VGND.n1670 VGND 0.0104432
R7467 VGND.n1678 VGND 0.0104432
R7468 VGND.n1696 VGND 0.0104432
R7469 VGND.n1704 VGND 0.0104432
R7470 VGND.n1722 VGND 0.0104432
R7471 VGND.n1730 VGND 0.0104432
R7472 VGND.n1753 VGND 0.0104432
R7473 VGND VGND.n294 0.0104432
R7474 VGND VGND.n295 0.0104432
R7475 VGND VGND.n511 0.0104432
R7476 VGND.n1773 VGND 0.0104432
R7477 VGND.n1532 VGND 0.0104432
R7478 VGND.n1540 VGND 0.0104432
R7479 VGND.n1631 VGND 0.0104432
R7480 VGND.n1639 VGND 0.0104432
R7481 VGND.n1657 VGND 0.0104432
R7482 VGND.n1665 VGND 0.0104432
R7483 VGND.n1683 VGND 0.0104432
R7484 VGND.n1691 VGND 0.0104432
R7485 VGND.n1709 VGND 0.0104432
R7486 VGND.n1717 VGND 0.0104432
R7487 VGND.n1735 VGND 0.0104432
R7488 VGND.n1748 VGND 0.0104432
R7489 VGND VGND.n291 0.0104432
R7490 VGND.n2377 VGND 0.0104432
R7491 VGND VGND.n287 0.0104432
R7492 VGND.n2387 VGND 0.0104432
R7493 VGND.n1297 VGND 0.0104432
R7494 VGND.n1545 VGND 0.0104432
R7495 VGND VGND.n549 0.0104432
R7496 VGND VGND.n550 0.0104432
R7497 VGND VGND.n551 0.0104432
R7498 VGND VGND.n552 0.0104432
R7499 VGND VGND.n553 0.0104432
R7500 VGND VGND.n554 0.0104432
R7501 VGND VGND.n555 0.0104432
R7502 VGND VGND.n556 0.0104432
R7503 VGND VGND.n557 0.0104432
R7504 VGND VGND.n558 0.0104432
R7505 VGND.n1616 VGND 0.0104432
R7506 VGND VGND.n282 0.0104432
R7507 VGND VGND.n283 0.0104432
R7508 VGND VGND.n1604 0.0104432
R7509 VGND.n826 VGND 0.0104432
R7510 VGND VGND.n827 0.0104432
R7511 VGND.n893 VGND 0.0104432
R7512 VGND VGND.n688 0.0104432
R7513 VGND VGND.n689 0.0104432
R7514 VGND VGND.n694 0.0104432
R7515 VGND VGND.n695 0.0104432
R7516 VGND VGND.n700 0.0104432
R7517 VGND VGND.n701 0.0104432
R7518 VGND VGND.n706 0.0104432
R7519 VGND VGND.n707 0.0104432
R7520 VGND VGND.n712 0.0104432
R7521 VGND VGND.n713 0.0104432
R7522 VGND.n2397 VGND 0.0104432
R7523 VGND VGND.n279 0.0104432
R7524 VGND.n2407 VGND 0.0104432
R7525 VGND.n1121 VGND 0.0104432
R7526 VGND.n1126 VGND 0.0104432
R7527 VGND VGND.n812 0.0104432
R7528 VGND.n1139 VGND 0.0104432
R7529 VGND.n1147 VGND 0.0104432
R7530 VGND.n1158 VGND 0.0104432
R7531 VGND VGND.n804 0.0104432
R7532 VGND.n1171 VGND 0.0104432
R7533 VGND.n1179 VGND 0.0104432
R7534 VGND.n1190 VGND 0.0104432
R7535 VGND VGND.n796 0.0104432
R7536 VGND.n1203 VGND 0.0104432
R7537 VGND.n1211 VGND 0.0104432
R7538 VGND.n1222 VGND 0.0104432
R7539 VGND VGND.n788 0.0104432
R7540 VGND.n1232 VGND 0.0104432
R7541 VGND.n677 VGND 0.0104432
R7542 VGND VGND.n1285 0.0104432
R7543 VGND.n685 VGND 0.0104432
R7544 VGND VGND.n686 0.0104432
R7545 VGND VGND.n691 0.0104432
R7546 VGND VGND.n692 0.0104432
R7547 VGND VGND.n697 0.0104432
R7548 VGND VGND.n698 0.0104432
R7549 VGND VGND.n703 0.0104432
R7550 VGND VGND.n704 0.0104432
R7551 VGND VGND.n709 0.0104432
R7552 VGND VGND.n710 0.0104432
R7553 VGND VGND.n715 0.0104432
R7554 VGND VGND.n716 0.0104432
R7555 VGND.n783 VGND 0.0104432
R7556 VGND.n2412 VGND 0.0104432
R7557 VGND.n3007 VGND 0.00851991
R7558 Iout.n1020 Iout.t116 239.927
R7559 Iout.n509 Iout.t201 239.927
R7560 Iout.n513 Iout.t158 239.927
R7561 Iout.n507 Iout.t124 239.927
R7562 Iout.n504 Iout.t7 239.927
R7563 Iout.n500 Iout.t142 239.927
R7564 Iout.n192 Iout.t155 239.927
R7565 Iout.n195 Iout.t0 239.927
R7566 Iout.n199 Iout.t75 239.927
R7567 Iout.n202 Iout.t8 239.927
R7568 Iout.n206 Iout.t98 239.927
R7569 Iout.n210 Iout.t94 239.927
R7570 Iout.n214 Iout.t4 239.927
R7571 Iout.n218 Iout.t50 239.927
R7572 Iout.n222 Iout.t114 239.927
R7573 Iout.n226 Iout.t126 239.927
R7574 Iout.n232 Iout.t40 239.927
R7575 Iout.n235 Iout.t66 239.927
R7576 Iout.n238 Iout.t205 239.927
R7577 Iout.n241 Iout.t131 239.927
R7578 Iout.n244 Iout.t6 239.927
R7579 Iout.n247 Iout.t174 239.927
R7580 Iout.n250 Iout.t105 239.927
R7581 Iout.n255 Iout.t111 239.927
R7582 Iout.n252 Iout.t198 239.927
R7583 Iout.n489 Iout.t81 239.927
R7584 Iout.n494 Iout.t178 239.927
R7585 Iout.n491 Iout.t129 239.927
R7586 Iout.n519 Iout.t139 239.927
R7587 Iout.n149 Iout.t157 239.927
R7588 Iout.n146 Iout.t255 239.927
R7589 Iout.n1010 Iout.t147 239.927
R7590 Iout.n1007 Iout.t247 239.927
R7591 Iout.n140 Iout.t53 239.927
R7592 Iout.n143 Iout.t171 239.927
R7593 Iout.n525 Iout.t231 239.927
R7594 Iout.n480 Iout.t196 239.927
R7595 Iout.n483 Iout.t58 239.927
R7596 Iout.n478 Iout.t65 239.927
R7597 Iout.n259 Iout.t32 239.927
R7598 Iout.n186 Iout.t172 239.927
R7599 Iout.n271 Iout.t37 239.927
R7600 Iout.n180 Iout.t59 239.927
R7601 Iout.n283 Iout.t237 239.927
R7602 Iout.n174 Iout.t242 239.927
R7603 Iout.n168 Iout.t195 239.927
R7604 Iout.n301 Iout.t189 239.927
R7605 Iout.n289 Iout.t228 239.927
R7606 Iout.n177 Iout.t103 239.927
R7607 Iout.n277 Iout.t70 239.927
R7608 Iout.n183 Iout.t39 239.927
R7609 Iout.n265 Iout.t92 239.927
R7610 Iout.n189 Iout.t216 239.927
R7611 Iout.n472 Iout.t177 239.927
R7612 Iout.n469 Iout.t9 239.927
R7613 Iout.n156 Iout.t165 239.927
R7614 Iout.n531 Iout.t10 239.927
R7615 Iout.n534 Iout.t213 239.927
R7616 Iout.n536 Iout.t69 239.927
R7617 Iout.n133 Iout.t123 239.927
R7618 Iout.n136 Iout.t248 239.927
R7619 Iout.n542 Iout.t31 239.927
R7620 Iout.n460 Iout.t29 239.927
R7621 Iout.n463 Iout.t221 239.927
R7622 Iout.n458 Iout.t160 239.927
R7623 Iout.n305 Iout.t26 239.927
R7624 Iout.n308 Iout.t80 239.927
R7625 Iout.n311 Iout.t226 239.927
R7626 Iout.n314 Iout.t83 239.927
R7627 Iout.n317 Iout.t113 239.927
R7628 Iout.n320 Iout.t67 239.927
R7629 Iout.n392 Iout.t253 239.927
R7630 Iout.n378 Iout.t112 239.927
R7631 Iout.n376 Iout.t183 239.927
R7632 Iout.n394 Iout.t73 239.927
R7633 Iout.n408 Iout.t199 239.927
R7634 Iout.n410 Iout.t91 239.927
R7635 Iout.n424 Iout.t246 239.927
R7636 Iout.n426 Iout.t206 239.927
R7637 Iout.n447 Iout.t176 239.927
R7638 Iout.n452 Iout.t186 239.927
R7639 Iout.n449 Iout.t164 239.927
R7640 Iout.n548 Iout.t191 239.927
R7641 Iout.n130 Iout.t203 239.927
R7642 Iout.n559 Iout.t169 239.927
R7643 Iout.n557 Iout.t34 239.927
R7644 Iout.n554 Iout.t25 239.927
R7645 Iout.n434 Iout.t78 239.927
R7646 Iout.n438 Iout.t104 239.927
R7647 Iout.n441 Iout.t41 239.927
R7648 Iout.n432 Iout.t20 239.927
R7649 Iout.n418 Iout.t85 239.927
R7650 Iout.n416 Iout.t49 239.927
R7651 Iout.n402 Iout.t99 239.927
R7652 Iout.n357 Iout.t115 239.927
R7653 Iout.n360 Iout.t76 239.927
R7654 Iout.n363 Iout.t251 239.927
R7655 Iout.n366 Iout.t187 239.927
R7656 Iout.n354 Iout.t145 239.927
R7657 Iout.n351 Iout.t207 239.927
R7658 Iout.n348 Iout.t149 239.927
R7659 Iout.n345 Iout.t192 239.927
R7660 Iout.n342 Iout.t219 239.927
R7661 Iout.n339 Iout.t225 239.927
R7662 Iout.n336 Iout.t209 239.927
R7663 Iout.n333 Iout.t182 239.927
R7664 Iout.n117 Iout.t240 239.927
R7665 Iout.n582 Iout.t222 239.927
R7666 Iout.n111 Iout.t55 239.927
R7667 Iout.n594 Iout.t128 239.927
R7668 Iout.n105 Iout.t13 239.927
R7669 Iout.n606 Iout.t151 239.927
R7670 Iout.n99 Iout.t179 239.927
R7671 Iout.n618 Iout.t72 239.927
R7672 Iout.n624 Iout.t143 239.927
R7673 Iout.n90 Iout.t197 239.927
R7674 Iout.n636 Iout.t12 239.927
R7675 Iout.n81 Iout.t90 239.927
R7676 Iout.n648 Iout.t63 239.927
R7677 Iout.n96 Iout.t214 239.927
R7678 Iout.n612 Iout.t33 239.927
R7679 Iout.n102 Iout.t56 239.927
R7680 Iout.n600 Iout.t134 239.927
R7681 Iout.n108 Iout.t79 239.927
R7682 Iout.n588 Iout.t235 239.927
R7683 Iout.n687 Iout.t156 239.927
R7684 Iout.n684 Iout.t193 239.927
R7685 Iout.n681 Iout.t100 239.927
R7686 Iout.n678 Iout.t249 239.927
R7687 Iout.n675 Iout.t215 239.927
R7688 Iout.n672 Iout.t84 239.927
R7689 Iout.n747 Iout.t250 239.927
R7690 Iout.n50 Iout.t229 239.927
R7691 Iout.n759 Iout.t95 239.927
R7692 Iout.n44 Iout.t61 239.927
R7693 Iout.n771 Iout.t220 239.927
R7694 Iout.n42 Iout.t45 239.927
R7695 Iout.n56 Iout.t254 239.927
R7696 Iout.n735 Iout.t77 239.927
R7697 Iout.n62 Iout.t184 239.927
R7698 Iout.n723 Iout.t217 239.927
R7699 Iout.n717 Iout.t152 239.927
R7700 Iout.n65 Iout.t146 239.927
R7701 Iout.n729 Iout.t3 239.927
R7702 Iout.n59 Iout.t15 239.927
R7703 Iout.n805 Iout.t96 239.927
R7704 Iout.n808 Iout.t162 239.927
R7705 Iout.n811 Iout.t62 239.927
R7706 Iout.n814 Iout.t87 239.927
R7707 Iout.n817 Iout.t2 239.927
R7708 Iout.n820 Iout.t64 239.927
R7709 Iout.n823 Iout.t52 239.927
R7710 Iout.n802 Iout.t210 239.927
R7711 Iout.n799 Iout.t185 239.927
R7712 Iout.n890 Iout.t107 239.927
R7713 Iout.n888 Iout.t245 239.927
R7714 Iout.n881 Iout.t42 239.927
R7715 Iout.n869 Iout.t110 239.927
R7716 Iout.n867 Iout.t130 239.927
R7717 Iout.n855 Iout.t16 239.927
R7718 Iout.n853 Iout.t148 239.927
R7719 Iout.n841 Iout.t230 239.927
R7720 Iout.n839 Iout.t68 239.927
R7721 Iout.n827 Iout.t5 239.927
R7722 Iout.n883 Iout.t57 239.927
R7723 Iout.n895 Iout.t54 239.927
R7724 Iout.n897 Iout.t218 239.927
R7725 Iout.n909 Iout.t108 239.927
R7726 Iout.n911 Iout.t121 239.927
R7727 Iout.n923 Iout.t47 239.927
R7728 Iout.n926 Iout.t163 239.927
R7729 Iout.n22 Iout.t168 239.927
R7730 Iout.n876 Iout.t102 239.927
R7731 Iout.n874 Iout.t232 239.927
R7732 Iout.n862 Iout.t11 239.927
R7733 Iout.n860 Iout.t167 239.927
R7734 Iout.n848 Iout.t136 239.927
R7735 Iout.n846 Iout.t97 239.927
R7736 Iout.n834 Iout.t224 239.927
R7737 Iout.n832 Iout.t51 239.927
R7738 Iout.n902 Iout.t30 239.927
R7739 Iout.n904 Iout.t236 239.927
R7740 Iout.n916 Iout.t227 239.927
R7741 Iout.n918 Iout.t27 239.927
R7742 Iout.n931 Iout.t19 239.927
R7743 Iout.n934 Iout.t1 239.927
R7744 Iout.n796 Iout.t43 239.927
R7745 Iout.n793 Iout.t166 239.927
R7746 Iout.n790 Iout.t38 239.927
R7747 Iout.n787 Iout.t252 239.927
R7748 Iout.n784 Iout.t140 239.927
R7749 Iout.n781 Iout.t241 239.927
R7750 Iout.n938 Iout.t159 239.927
R7751 Iout.n741 Iout.t35 239.927
R7752 Iout.n53 Iout.t133 239.927
R7753 Iout.n753 Iout.t122 239.927
R7754 Iout.n47 Iout.t204 239.927
R7755 Iout.n765 Iout.t101 239.927
R7756 Iout.n38 Iout.t212 239.927
R7757 Iout.n777 Iout.t44 239.927
R7758 Iout.n71 Iout.t60 239.927
R7759 Iout.n705 Iout.t181 239.927
R7760 Iout.n77 Iout.t154 239.927
R7761 Iout.n944 Iout.t137 239.927
R7762 Iout.n19 Iout.t89 239.927
R7763 Iout.n68 Iout.t22 239.927
R7764 Iout.n711 Iout.t71 239.927
R7765 Iout.n74 Iout.t170 239.927
R7766 Iout.n699 Iout.t127 239.927
R7767 Iout.n950 Iout.t141 239.927
R7768 Iout.n953 Iout.t239 239.927
R7769 Iout.n669 Iout.t23 239.927
R7770 Iout.n666 Iout.t161 239.927
R7771 Iout.n663 Iout.t17 239.927
R7772 Iout.n660 Iout.t223 239.927
R7773 Iout.n657 Iout.t175 239.927
R7774 Iout.n654 Iout.t138 239.927
R7775 Iout.n690 Iout.t202 239.927
R7776 Iout.n695 Iout.t109 239.927
R7777 Iout.n692 Iout.t36 239.927
R7778 Iout.n957 Iout.t200 239.927
R7779 Iout.n114 Iout.t117 239.927
R7780 Iout.n576 Iout.t233 239.927
R7781 Iout.n573 Iout.t82 239.927
R7782 Iout.n963 Iout.t238 239.927
R7783 Iout.n14 Iout.t119 239.927
R7784 Iout.n93 Iout.t173 239.927
R7785 Iout.n630 Iout.t180 239.927
R7786 Iout.n87 Iout.t21 239.927
R7787 Iout.n642 Iout.t234 239.927
R7788 Iout.n85 Iout.t106 239.927
R7789 Iout.n563 Iout.t125 239.927
R7790 Iout.n969 Iout.t135 239.927
R7791 Iout.n972 Iout.t93 239.927
R7792 Iout.n569 Iout.t48 239.927
R7793 Iout.n123 Iout.t14 239.927
R7794 Iout.n120 Iout.t118 239.927
R7795 Iout.n976 Iout.t208 239.927
R7796 Iout.n400 Iout.t132 239.927
R7797 Iout.n386 Iout.t194 239.927
R7798 Iout.n384 Iout.t243 239.927
R7799 Iout.n370 Iout.t190 239.927
R7800 Iout.n982 Iout.t120 239.927
R7801 Iout.n9 Iout.t28 239.927
R7802 Iout.n127 Iout.t188 239.927
R7803 Iout.n988 Iout.t74 239.927
R7804 Iout.n991 Iout.t144 239.927
R7805 Iout.n323 Iout.t18 239.927
R7806 Iout.n326 Iout.t46 239.927
R7807 Iout.n329 Iout.t150 239.927
R7808 Iout.n995 Iout.t86 239.927
R7809 Iout.n1001 Iout.t153 239.927
R7810 Iout.n4 Iout.t244 239.927
R7811 Iout.n295 Iout.t24 239.927
R7812 Iout.n172 Iout.t211 239.927
R7813 Iout.n1014 Iout.t88 239.927
R7814 Iout.n1021 Iout.n1020 7.9105
R7815 Iout.n510 Iout.n509 7.9105
R7816 Iout.n514 Iout.n513 7.9105
R7817 Iout.n508 Iout.n507 7.9105
R7818 Iout.n505 Iout.n504 7.9105
R7819 Iout.n501 Iout.n500 7.9105
R7820 Iout.n193 Iout.n192 7.9105
R7821 Iout.n196 Iout.n195 7.9105
R7822 Iout.n200 Iout.n199 7.9105
R7823 Iout.n203 Iout.n202 7.9105
R7824 Iout.n207 Iout.n206 7.9105
R7825 Iout.n211 Iout.n210 7.9105
R7826 Iout.n215 Iout.n214 7.9105
R7827 Iout.n219 Iout.n218 7.9105
R7828 Iout.n223 Iout.n222 7.9105
R7829 Iout.n227 Iout.n226 7.9105
R7830 Iout.n233 Iout.n232 7.9105
R7831 Iout.n236 Iout.n235 7.9105
R7832 Iout.n239 Iout.n238 7.9105
R7833 Iout.n242 Iout.n241 7.9105
R7834 Iout.n245 Iout.n244 7.9105
R7835 Iout.n248 Iout.n247 7.9105
R7836 Iout.n251 Iout.n250 7.9105
R7837 Iout.n256 Iout.n255 7.9105
R7838 Iout.n253 Iout.n252 7.9105
R7839 Iout.n490 Iout.n489 7.9105
R7840 Iout.n495 Iout.n494 7.9105
R7841 Iout.n492 Iout.n491 7.9105
R7842 Iout.n520 Iout.n519 7.9105
R7843 Iout.n150 Iout.n149 7.9105
R7844 Iout.n147 Iout.n146 7.9105
R7845 Iout.n1011 Iout.n1010 7.9105
R7846 Iout.n1008 Iout.n1007 7.9105
R7847 Iout.n141 Iout.n140 7.9105
R7848 Iout.n144 Iout.n143 7.9105
R7849 Iout.n526 Iout.n525 7.9105
R7850 Iout.n481 Iout.n480 7.9105
R7851 Iout.n484 Iout.n483 7.9105
R7852 Iout.n479 Iout.n478 7.9105
R7853 Iout.n260 Iout.n259 7.9105
R7854 Iout.n187 Iout.n186 7.9105
R7855 Iout.n272 Iout.n271 7.9105
R7856 Iout.n181 Iout.n180 7.9105
R7857 Iout.n284 Iout.n283 7.9105
R7858 Iout.n175 Iout.n174 7.9105
R7859 Iout.n169 Iout.n168 7.9105
R7860 Iout.n302 Iout.n301 7.9105
R7861 Iout.n290 Iout.n289 7.9105
R7862 Iout.n178 Iout.n177 7.9105
R7863 Iout.n278 Iout.n277 7.9105
R7864 Iout.n184 Iout.n183 7.9105
R7865 Iout.n266 Iout.n265 7.9105
R7866 Iout.n190 Iout.n189 7.9105
R7867 Iout.n473 Iout.n472 7.9105
R7868 Iout.n470 Iout.n469 7.9105
R7869 Iout.n157 Iout.n156 7.9105
R7870 Iout.n532 Iout.n531 7.9105
R7871 Iout.n535 Iout.n534 7.9105
R7872 Iout.n537 Iout.n536 7.9105
R7873 Iout.n134 Iout.n133 7.9105
R7874 Iout.n137 Iout.n136 7.9105
R7875 Iout.n543 Iout.n542 7.9105
R7876 Iout.n461 Iout.n460 7.9105
R7877 Iout.n464 Iout.n463 7.9105
R7878 Iout.n459 Iout.n458 7.9105
R7879 Iout.n306 Iout.n305 7.9105
R7880 Iout.n309 Iout.n308 7.9105
R7881 Iout.n312 Iout.n311 7.9105
R7882 Iout.n315 Iout.n314 7.9105
R7883 Iout.n318 Iout.n317 7.9105
R7884 Iout.n321 Iout.n320 7.9105
R7885 Iout.n393 Iout.n392 7.9105
R7886 Iout.n379 Iout.n378 7.9105
R7887 Iout.n377 Iout.n376 7.9105
R7888 Iout.n395 Iout.n394 7.9105
R7889 Iout.n409 Iout.n408 7.9105
R7890 Iout.n411 Iout.n410 7.9105
R7891 Iout.n425 Iout.n424 7.9105
R7892 Iout.n427 Iout.n426 7.9105
R7893 Iout.n448 Iout.n447 7.9105
R7894 Iout.n453 Iout.n452 7.9105
R7895 Iout.n450 Iout.n449 7.9105
R7896 Iout.n549 Iout.n548 7.9105
R7897 Iout.n131 Iout.n130 7.9105
R7898 Iout.n560 Iout.n559 7.9105
R7899 Iout.n558 Iout.n557 7.9105
R7900 Iout.n555 Iout.n554 7.9105
R7901 Iout.n435 Iout.n434 7.9105
R7902 Iout.n439 Iout.n438 7.9105
R7903 Iout.n442 Iout.n441 7.9105
R7904 Iout.n433 Iout.n432 7.9105
R7905 Iout.n419 Iout.n418 7.9105
R7906 Iout.n417 Iout.n416 7.9105
R7907 Iout.n403 Iout.n402 7.9105
R7908 Iout.n358 Iout.n357 7.9105
R7909 Iout.n361 Iout.n360 7.9105
R7910 Iout.n364 Iout.n363 7.9105
R7911 Iout.n367 Iout.n366 7.9105
R7912 Iout.n355 Iout.n354 7.9105
R7913 Iout.n352 Iout.n351 7.9105
R7914 Iout.n349 Iout.n348 7.9105
R7915 Iout.n346 Iout.n345 7.9105
R7916 Iout.n343 Iout.n342 7.9105
R7917 Iout.n340 Iout.n339 7.9105
R7918 Iout.n337 Iout.n336 7.9105
R7919 Iout.n334 Iout.n333 7.9105
R7920 Iout.n118 Iout.n117 7.9105
R7921 Iout.n583 Iout.n582 7.9105
R7922 Iout.n112 Iout.n111 7.9105
R7923 Iout.n595 Iout.n594 7.9105
R7924 Iout.n106 Iout.n105 7.9105
R7925 Iout.n607 Iout.n606 7.9105
R7926 Iout.n100 Iout.n99 7.9105
R7927 Iout.n619 Iout.n618 7.9105
R7928 Iout.n625 Iout.n624 7.9105
R7929 Iout.n91 Iout.n90 7.9105
R7930 Iout.n637 Iout.n636 7.9105
R7931 Iout.n82 Iout.n81 7.9105
R7932 Iout.n649 Iout.n648 7.9105
R7933 Iout.n97 Iout.n96 7.9105
R7934 Iout.n613 Iout.n612 7.9105
R7935 Iout.n103 Iout.n102 7.9105
R7936 Iout.n601 Iout.n600 7.9105
R7937 Iout.n109 Iout.n108 7.9105
R7938 Iout.n589 Iout.n588 7.9105
R7939 Iout.n688 Iout.n687 7.9105
R7940 Iout.n685 Iout.n684 7.9105
R7941 Iout.n682 Iout.n681 7.9105
R7942 Iout.n679 Iout.n678 7.9105
R7943 Iout.n676 Iout.n675 7.9105
R7944 Iout.n673 Iout.n672 7.9105
R7945 Iout.n748 Iout.n747 7.9105
R7946 Iout.n51 Iout.n50 7.9105
R7947 Iout.n760 Iout.n759 7.9105
R7948 Iout.n45 Iout.n44 7.9105
R7949 Iout.n772 Iout.n771 7.9105
R7950 Iout.n43 Iout.n42 7.9105
R7951 Iout.n57 Iout.n56 7.9105
R7952 Iout.n736 Iout.n735 7.9105
R7953 Iout.n63 Iout.n62 7.9105
R7954 Iout.n724 Iout.n723 7.9105
R7955 Iout.n718 Iout.n717 7.9105
R7956 Iout.n66 Iout.n65 7.9105
R7957 Iout.n730 Iout.n729 7.9105
R7958 Iout.n60 Iout.n59 7.9105
R7959 Iout.n806 Iout.n805 7.9105
R7960 Iout.n809 Iout.n808 7.9105
R7961 Iout.n812 Iout.n811 7.9105
R7962 Iout.n815 Iout.n814 7.9105
R7963 Iout.n818 Iout.n817 7.9105
R7964 Iout.n821 Iout.n820 7.9105
R7965 Iout.n824 Iout.n823 7.9105
R7966 Iout.n803 Iout.n802 7.9105
R7967 Iout.n800 Iout.n799 7.9105
R7968 Iout.n891 Iout.n890 7.9105
R7969 Iout.n889 Iout.n888 7.9105
R7970 Iout.n882 Iout.n881 7.9105
R7971 Iout.n870 Iout.n869 7.9105
R7972 Iout.n868 Iout.n867 7.9105
R7973 Iout.n856 Iout.n855 7.9105
R7974 Iout.n854 Iout.n853 7.9105
R7975 Iout.n842 Iout.n841 7.9105
R7976 Iout.n840 Iout.n839 7.9105
R7977 Iout.n828 Iout.n827 7.9105
R7978 Iout.n884 Iout.n883 7.9105
R7979 Iout.n896 Iout.n895 7.9105
R7980 Iout.n898 Iout.n897 7.9105
R7981 Iout.n910 Iout.n909 7.9105
R7982 Iout.n912 Iout.n911 7.9105
R7983 Iout.n924 Iout.n923 7.9105
R7984 Iout.n927 Iout.n926 7.9105
R7985 Iout.n23 Iout.n22 7.9105
R7986 Iout.n877 Iout.n876 7.9105
R7987 Iout.n875 Iout.n874 7.9105
R7988 Iout.n863 Iout.n862 7.9105
R7989 Iout.n861 Iout.n860 7.9105
R7990 Iout.n849 Iout.n848 7.9105
R7991 Iout.n847 Iout.n846 7.9105
R7992 Iout.n835 Iout.n834 7.9105
R7993 Iout.n833 Iout.n832 7.9105
R7994 Iout.n903 Iout.n902 7.9105
R7995 Iout.n905 Iout.n904 7.9105
R7996 Iout.n917 Iout.n916 7.9105
R7997 Iout.n919 Iout.n918 7.9105
R7998 Iout.n932 Iout.n931 7.9105
R7999 Iout.n935 Iout.n934 7.9105
R8000 Iout.n797 Iout.n796 7.9105
R8001 Iout.n794 Iout.n793 7.9105
R8002 Iout.n791 Iout.n790 7.9105
R8003 Iout.n788 Iout.n787 7.9105
R8004 Iout.n785 Iout.n784 7.9105
R8005 Iout.n782 Iout.n781 7.9105
R8006 Iout.n939 Iout.n938 7.9105
R8007 Iout.n742 Iout.n741 7.9105
R8008 Iout.n54 Iout.n53 7.9105
R8009 Iout.n754 Iout.n753 7.9105
R8010 Iout.n48 Iout.n47 7.9105
R8011 Iout.n766 Iout.n765 7.9105
R8012 Iout.n39 Iout.n38 7.9105
R8013 Iout.n778 Iout.n777 7.9105
R8014 Iout.n72 Iout.n71 7.9105
R8015 Iout.n706 Iout.n705 7.9105
R8016 Iout.n78 Iout.n77 7.9105
R8017 Iout.n945 Iout.n944 7.9105
R8018 Iout.n20 Iout.n19 7.9105
R8019 Iout.n69 Iout.n68 7.9105
R8020 Iout.n712 Iout.n711 7.9105
R8021 Iout.n75 Iout.n74 7.9105
R8022 Iout.n700 Iout.n699 7.9105
R8023 Iout.n951 Iout.n950 7.9105
R8024 Iout.n954 Iout.n953 7.9105
R8025 Iout.n670 Iout.n669 7.9105
R8026 Iout.n667 Iout.n666 7.9105
R8027 Iout.n664 Iout.n663 7.9105
R8028 Iout.n661 Iout.n660 7.9105
R8029 Iout.n658 Iout.n657 7.9105
R8030 Iout.n655 Iout.n654 7.9105
R8031 Iout.n691 Iout.n690 7.9105
R8032 Iout.n696 Iout.n695 7.9105
R8033 Iout.n693 Iout.n692 7.9105
R8034 Iout.n958 Iout.n957 7.9105
R8035 Iout.n115 Iout.n114 7.9105
R8036 Iout.n577 Iout.n576 7.9105
R8037 Iout.n574 Iout.n573 7.9105
R8038 Iout.n964 Iout.n963 7.9105
R8039 Iout.n15 Iout.n14 7.9105
R8040 Iout.n94 Iout.n93 7.9105
R8041 Iout.n631 Iout.n630 7.9105
R8042 Iout.n88 Iout.n87 7.9105
R8043 Iout.n643 Iout.n642 7.9105
R8044 Iout.n86 Iout.n85 7.9105
R8045 Iout.n564 Iout.n563 7.9105
R8046 Iout.n970 Iout.n969 7.9105
R8047 Iout.n973 Iout.n972 7.9105
R8048 Iout.n570 Iout.n569 7.9105
R8049 Iout.n124 Iout.n123 7.9105
R8050 Iout.n121 Iout.n120 7.9105
R8051 Iout.n977 Iout.n976 7.9105
R8052 Iout.n401 Iout.n400 7.9105
R8053 Iout.n387 Iout.n386 7.9105
R8054 Iout.n385 Iout.n384 7.9105
R8055 Iout.n371 Iout.n370 7.9105
R8056 Iout.n983 Iout.n982 7.9105
R8057 Iout.n10 Iout.n9 7.9105
R8058 Iout.n128 Iout.n127 7.9105
R8059 Iout.n989 Iout.n988 7.9105
R8060 Iout.n992 Iout.n991 7.9105
R8061 Iout.n324 Iout.n323 7.9105
R8062 Iout.n327 Iout.n326 7.9105
R8063 Iout.n330 Iout.n329 7.9105
R8064 Iout.n996 Iout.n995 7.9105
R8065 Iout.n1002 Iout.n1001 7.9105
R8066 Iout.n5 Iout.n4 7.9105
R8067 Iout.n296 Iout.n295 7.9105
R8068 Iout.n173 Iout.n172 7.9105
R8069 Iout.n1015 Iout.n1014 7.9105
R8070 Iout.n886 Iout.n885 3.86101
R8071 Iout.n880 Iout.n879 3.86101
R8072 Iout.n894 Iout.n893 3.86101
R8073 Iout.n872 Iout.n871 3.86101
R8074 Iout.n900 Iout.n899 3.86101
R8075 Iout.n866 Iout.n865 3.86101
R8076 Iout.n908 Iout.n907 3.86101
R8077 Iout.n858 Iout.n857 3.86101
R8078 Iout.n914 Iout.n913 3.86101
R8079 Iout.n852 Iout.n851 3.86101
R8080 Iout.n922 Iout.n921 3.86101
R8081 Iout.n844 Iout.n843 3.86101
R8082 Iout.n929 Iout.n928 3.86101
R8083 Iout.n838 Iout.n837 3.86101
R8084 Iout.n925 Iout.n21 3.86101
R8085 Iout.n830 Iout.n829 3.86101
R8086 Iout.n879 Iout.n878 3.4105
R8087 Iout.n887 Iout.n886 3.4105
R8088 Iout.n893 Iout.n892 3.4105
R8089 Iout.n798 Iout.n28 3.4105
R8090 Iout.n801 Iout.n29 3.4105
R8091 Iout.n804 Iout.n30 3.4105
R8092 Iout.n807 Iout.n31 3.4105
R8093 Iout.n873 Iout.n872 3.4105
R8094 Iout.n744 Iout.n743 3.4105
R8095 Iout.n740 Iout.n739 3.4105
R8096 Iout.n732 Iout.n731 3.4105
R8097 Iout.n728 Iout.n727 3.4105
R8098 Iout.n720 Iout.n719 3.4105
R8099 Iout.n795 Iout.n27 3.4105
R8100 Iout.n901 Iout.n900 3.4105
R8101 Iout.n722 Iout.n721 3.4105
R8102 Iout.n726 Iout.n725 3.4105
R8103 Iout.n734 Iout.n733 3.4105
R8104 Iout.n738 Iout.n737 3.4105
R8105 Iout.n746 Iout.n745 3.4105
R8106 Iout.n750 Iout.n749 3.4105
R8107 Iout.n752 Iout.n751 3.4105
R8108 Iout.n810 Iout.n32 3.4105
R8109 Iout.n865 Iout.n864 3.4105
R8110 Iout.n668 Iout.n55 3.4105
R8111 Iout.n671 Iout.n58 3.4105
R8112 Iout.n674 Iout.n61 3.4105
R8113 Iout.n677 Iout.n64 3.4105
R8114 Iout.n680 Iout.n67 3.4105
R8115 Iout.n683 Iout.n70 3.4105
R8116 Iout.n686 Iout.n73 3.4105
R8117 Iout.n714 Iout.n713 3.4105
R8118 Iout.n716 Iout.n715 3.4105
R8119 Iout.n792 Iout.n26 3.4105
R8120 Iout.n907 Iout.n906 3.4105
R8121 Iout.n587 Iout.n586 3.4105
R8122 Iout.n591 Iout.n590 3.4105
R8123 Iout.n599 Iout.n598 3.4105
R8124 Iout.n603 Iout.n602 3.4105
R8125 Iout.n611 Iout.n610 3.4105
R8126 Iout.n615 Iout.n614 3.4105
R8127 Iout.n623 Iout.n622 3.4105
R8128 Iout.n627 Iout.n626 3.4105
R8129 Iout.n665 Iout.n52 3.4105
R8130 Iout.n758 Iout.n757 3.4105
R8131 Iout.n756 Iout.n755 3.4105
R8132 Iout.n813 Iout.n33 3.4105
R8133 Iout.n859 Iout.n858 3.4105
R8134 Iout.n629 Iout.n628 3.4105
R8135 Iout.n621 Iout.n620 3.4105
R8136 Iout.n617 Iout.n616 3.4105
R8137 Iout.n609 Iout.n608 3.4105
R8138 Iout.n605 Iout.n604 3.4105
R8139 Iout.n597 Iout.n596 3.4105
R8140 Iout.n593 Iout.n592 3.4105
R8141 Iout.n585 Iout.n584 3.4105
R8142 Iout.n581 Iout.n580 3.4105
R8143 Iout.n579 Iout.n578 3.4105
R8144 Iout.n689 Iout.n76 3.4105
R8145 Iout.n710 Iout.n709 3.4105
R8146 Iout.n708 Iout.n707 3.4105
R8147 Iout.n789 Iout.n25 3.4105
R8148 Iout.n915 Iout.n914 3.4105
R8149 Iout.n572 Iout.n571 3.4105
R8150 Iout.n335 Iout.n116 3.4105
R8151 Iout.n338 Iout.n113 3.4105
R8152 Iout.n341 Iout.n110 3.4105
R8153 Iout.n344 Iout.n107 3.4105
R8154 Iout.n347 Iout.n104 3.4105
R8155 Iout.n350 Iout.n101 3.4105
R8156 Iout.n353 Iout.n98 3.4105
R8157 Iout.n356 Iout.n95 3.4105
R8158 Iout.n359 Iout.n92 3.4105
R8159 Iout.n633 Iout.n632 3.4105
R8160 Iout.n635 Iout.n634 3.4105
R8161 Iout.n662 Iout.n49 3.4105
R8162 Iout.n762 Iout.n761 3.4105
R8163 Iout.n764 Iout.n763 3.4105
R8164 Iout.n816 Iout.n34 3.4105
R8165 Iout.n851 Iout.n850 3.4105
R8166 Iout.n399 Iout.n398 3.4105
R8167 Iout.n405 Iout.n404 3.4105
R8168 Iout.n415 Iout.n414 3.4105
R8169 Iout.n421 Iout.n420 3.4105
R8170 Iout.n431 Iout.n430 3.4105
R8171 Iout.n444 Iout.n443 3.4105
R8172 Iout.n440 Iout.n159 3.4105
R8173 Iout.n437 Iout.n436 3.4105
R8174 Iout.n553 Iout.n552 3.4105
R8175 Iout.n556 Iout.n119 3.4105
R8176 Iout.n562 Iout.n561 3.4105
R8177 Iout.n568 Iout.n567 3.4105
R8178 Iout.n566 Iout.n565 3.4105
R8179 Iout.n575 Iout.n79 3.4105
R8180 Iout.n698 Iout.n697 3.4105
R8181 Iout.n702 Iout.n701 3.4105
R8182 Iout.n704 Iout.n703 3.4105
R8183 Iout.n786 Iout.n24 3.4105
R8184 Iout.n921 Iout.n920 3.4105
R8185 Iout.n129 Iout.n125 3.4105
R8186 Iout.n547 Iout.n546 3.4105
R8187 Iout.n551 Iout.n550 3.4105
R8188 Iout.n451 Iout.n158 3.4105
R8189 Iout.n455 Iout.n454 3.4105
R8190 Iout.n446 Iout.n445 3.4105
R8191 Iout.n429 Iout.n428 3.4105
R8192 Iout.n423 Iout.n422 3.4105
R8193 Iout.n413 Iout.n412 3.4105
R8194 Iout.n407 Iout.n406 3.4105
R8195 Iout.n397 Iout.n396 3.4105
R8196 Iout.n391 Iout.n390 3.4105
R8197 Iout.n389 Iout.n388 3.4105
R8198 Iout.n362 Iout.n89 3.4105
R8199 Iout.n641 Iout.n640 3.4105
R8200 Iout.n639 Iout.n638 3.4105
R8201 Iout.n659 Iout.n46 3.4105
R8202 Iout.n770 Iout.n769 3.4105
R8203 Iout.n768 Iout.n767 3.4105
R8204 Iout.n819 Iout.n35 3.4105
R8205 Iout.n845 Iout.n844 3.4105
R8206 Iout.n325 Iout.n165 3.4105
R8207 Iout.n322 Iout.n164 3.4105
R8208 Iout.n319 Iout.n163 3.4105
R8209 Iout.n316 Iout.n162 3.4105
R8210 Iout.n313 Iout.n161 3.4105
R8211 Iout.n310 Iout.n160 3.4105
R8212 Iout.n307 Iout.n155 3.4105
R8213 Iout.n457 Iout.n456 3.4105
R8214 Iout.n466 Iout.n465 3.4105
R8215 Iout.n462 Iout.n126 3.4105
R8216 Iout.n545 Iout.n544 3.4105
R8217 Iout.n541 Iout.n540 3.4105
R8218 Iout.n135 Iout.n3 3.4105
R8219 Iout.n987 Iout.n986 3.4105
R8220 Iout.n985 Iout.n984 3.4105
R8221 Iout.n122 Iout.n8 3.4105
R8222 Iout.n968 Iout.n967 3.4105
R8223 Iout.n966 Iout.n965 3.4105
R8224 Iout.n694 Iout.n13 3.4105
R8225 Iout.n949 Iout.n948 3.4105
R8226 Iout.n947 Iout.n946 3.4105
R8227 Iout.n783 Iout.n18 3.4105
R8228 Iout.n930 Iout.n929 3.4105
R8229 Iout.n1004 Iout.n1003 3.4105
R8230 Iout.n539 Iout.n538 3.4105
R8231 Iout.n533 Iout.n132 3.4105
R8232 Iout.n530 Iout.n529 3.4105
R8233 Iout.n468 Iout.n467 3.4105
R8234 Iout.n471 Iout.n153 3.4105
R8235 Iout.n475 Iout.n474 3.4105
R8236 Iout.n264 Iout.n263 3.4105
R8237 Iout.n268 Iout.n267 3.4105
R8238 Iout.n276 Iout.n275 3.4105
R8239 Iout.n280 Iout.n279 3.4105
R8240 Iout.n288 Iout.n287 3.4105
R8241 Iout.n292 Iout.n291 3.4105
R8242 Iout.n300 Iout.n299 3.4105
R8243 Iout.n328 Iout.n166 3.4105
R8244 Iout.n381 Iout.n380 3.4105
R8245 Iout.n383 Iout.n382 3.4105
R8246 Iout.n365 Iout.n83 3.4105
R8247 Iout.n645 Iout.n644 3.4105
R8248 Iout.n647 Iout.n646 3.4105
R8249 Iout.n656 Iout.n40 3.4105
R8250 Iout.n774 Iout.n773 3.4105
R8251 Iout.n776 Iout.n775 3.4105
R8252 Iout.n822 Iout.n36 3.4105
R8253 Iout.n837 Iout.n836 3.4105
R8254 Iout.n298 Iout.n297 3.4105
R8255 Iout.n294 Iout.n293 3.4105
R8256 Iout.n286 Iout.n285 3.4105
R8257 Iout.n282 Iout.n281 3.4105
R8258 Iout.n274 Iout.n273 3.4105
R8259 Iout.n270 Iout.n269 3.4105
R8260 Iout.n262 Iout.n261 3.4105
R8261 Iout.n477 Iout.n476 3.4105
R8262 Iout.n486 Iout.n485 3.4105
R8263 Iout.n482 Iout.n151 3.4105
R8264 Iout.n528 Iout.n527 3.4105
R8265 Iout.n524 Iout.n523 3.4105
R8266 Iout.n142 Iout.n138 3.4105
R8267 Iout.n1006 Iout.n1005 3.4105
R8268 Iout.n1009 Iout.n0 3.4105
R8269 Iout.n1000 Iout.n999 3.4105
R8270 Iout.n998 Iout.n997 3.4105
R8271 Iout.n990 Iout.n6 3.4105
R8272 Iout.n981 Iout.n980 3.4105
R8273 Iout.n979 Iout.n978 3.4105
R8274 Iout.n971 Iout.n11 3.4105
R8275 Iout.n962 Iout.n961 3.4105
R8276 Iout.n960 Iout.n959 3.4105
R8277 Iout.n952 Iout.n16 3.4105
R8278 Iout.n943 Iout.n942 3.4105
R8279 Iout.n941 Iout.n940 3.4105
R8280 Iout.n933 Iout.n21 3.4105
R8281 Iout.n1017 Iout.n1016 3.4105
R8282 Iout.n148 Iout.n2 3.4105
R8283 Iout.n518 Iout.n517 3.4105
R8284 Iout.n522 Iout.n521 3.4105
R8285 Iout.n493 Iout.n139 3.4105
R8286 Iout.n497 Iout.n496 3.4105
R8287 Iout.n488 Iout.n487 3.4105
R8288 Iout.n254 Iout.n154 3.4105
R8289 Iout.n258 Iout.n257 3.4105
R8290 Iout.n249 Iout.n188 3.4105
R8291 Iout.n246 Iout.n185 3.4105
R8292 Iout.n243 Iout.n182 3.4105
R8293 Iout.n240 Iout.n179 3.4105
R8294 Iout.n237 Iout.n176 3.4105
R8295 Iout.n234 Iout.n170 3.4105
R8296 Iout.n231 Iout.n230 3.4105
R8297 Iout.n171 Iout.n167 3.4105
R8298 Iout.n304 Iout.n303 3.4105
R8299 Iout.n332 Iout.n331 3.4105
R8300 Iout.n375 Iout.n374 3.4105
R8301 Iout.n373 Iout.n372 3.4105
R8302 Iout.n369 Iout.n368 3.4105
R8303 Iout.n84 Iout.n80 3.4105
R8304 Iout.n651 Iout.n650 3.4105
R8305 Iout.n653 Iout.n652 3.4105
R8306 Iout.n41 Iout.n37 3.4105
R8307 Iout.n780 Iout.n779 3.4105
R8308 Iout.n826 Iout.n825 3.4105
R8309 Iout.n831 Iout.n830 3.4105
R8310 Iout.n229 Iout.n228 3.4105
R8311 Iout.n225 Iout.n224 3.4105
R8312 Iout.n221 Iout.n220 3.4105
R8313 Iout.n217 Iout.n216 3.4105
R8314 Iout.n213 Iout.n212 3.4105
R8315 Iout.n209 Iout.n208 3.4105
R8316 Iout.n205 Iout.n204 3.4105
R8317 Iout.n201 Iout.n191 3.4105
R8318 Iout.n198 Iout.n197 3.4105
R8319 Iout.n194 Iout.n152 3.4105
R8320 Iout.n499 Iout.n498 3.4105
R8321 Iout.n503 Iout.n502 3.4105
R8322 Iout.n506 Iout.n145 3.4105
R8323 Iout.n516 Iout.n515 3.4105
R8324 Iout.n512 Iout.n511 3.4105
R8325 Iout.n1019 Iout.n1018 3.4105
R8326 Iout.n936 Iout.n23 1.43848
R8327 Iout.n936 Iout.n935 1.34612
R8328 Iout.n939 Iout.n937 1.34612
R8329 Iout.n20 Iout.n17 1.34612
R8330 Iout.n955 Iout.n954 1.34612
R8331 Iout.n958 Iout.n956 1.34612
R8332 Iout.n15 Iout.n12 1.34612
R8333 Iout.n974 Iout.n973 1.34612
R8334 Iout.n977 Iout.n975 1.34612
R8335 Iout.n10 Iout.n7 1.34612
R8336 Iout.n993 Iout.n992 1.34612
R8337 Iout.n996 Iout.n994 1.34612
R8338 Iout.n5 Iout.n1 1.34612
R8339 Iout.n1012 Iout.n1011 1.34612
R8340 Iout.n1015 Iout.n1013 1.34612
R8341 Iout.n1022 Iout.n1021 1.34612
R8342 Iout.n197 Iout.n154 0.451012
R8343 Iout.n476 Iout.n154 0.451012
R8344 Iout.n476 Iout.n475 0.451012
R8345 Iout.n475 Iout.n155 0.451012
R8346 Iout.n445 Iout.n155 0.451012
R8347 Iout.n445 Iout.n444 0.451012
R8348 Iout.n444 Iout.n107 0.451012
R8349 Iout.n604 Iout.n107 0.451012
R8350 Iout.n604 Iout.n603 0.451012
R8351 Iout.n603 Iout.n64 0.451012
R8352 Iout.n733 Iout.n64 0.451012
R8353 Iout.n733 Iout.n732 0.451012
R8354 Iout.n732 Iout.n29 0.451012
R8355 Iout.n886 Iout.n29 0.451012
R8356 Iout.n258 Iout.n191 0.451012
R8357 Iout.n262 Iout.n258 0.451012
R8358 Iout.n263 Iout.n262 0.451012
R8359 Iout.n263 Iout.n160 0.451012
R8360 Iout.n429 Iout.n160 0.451012
R8361 Iout.n430 Iout.n429 0.451012
R8362 Iout.n430 Iout.n104 0.451012
R8363 Iout.n609 Iout.n104 0.451012
R8364 Iout.n610 Iout.n609 0.451012
R8365 Iout.n610 Iout.n61 0.451012
R8366 Iout.n738 Iout.n61 0.451012
R8367 Iout.n739 Iout.n738 0.451012
R8368 Iout.n739 Iout.n30 0.451012
R8369 Iout.n879 Iout.n30 0.451012
R8370 Iout.n487 Iout.n152 0.451012
R8371 Iout.n487 Iout.n486 0.451012
R8372 Iout.n486 Iout.n153 0.451012
R8373 Iout.n456 Iout.n153 0.451012
R8374 Iout.n456 Iout.n455 0.451012
R8375 Iout.n455 Iout.n159 0.451012
R8376 Iout.n159 Iout.n110 0.451012
R8377 Iout.n597 Iout.n110 0.451012
R8378 Iout.n598 Iout.n597 0.451012
R8379 Iout.n598 Iout.n67 0.451012
R8380 Iout.n726 Iout.n67 0.451012
R8381 Iout.n727 Iout.n726 0.451012
R8382 Iout.n727 Iout.n28 0.451012
R8383 Iout.n893 Iout.n28 0.451012
R8384 Iout.n204 Iout.n188 0.451012
R8385 Iout.n269 Iout.n188 0.451012
R8386 Iout.n269 Iout.n268 0.451012
R8387 Iout.n268 Iout.n161 0.451012
R8388 Iout.n422 Iout.n161 0.451012
R8389 Iout.n422 Iout.n421 0.451012
R8390 Iout.n421 Iout.n101 0.451012
R8391 Iout.n616 Iout.n101 0.451012
R8392 Iout.n616 Iout.n615 0.451012
R8393 Iout.n615 Iout.n58 0.451012
R8394 Iout.n745 Iout.n58 0.451012
R8395 Iout.n745 Iout.n744 0.451012
R8396 Iout.n744 Iout.n31 0.451012
R8397 Iout.n872 Iout.n31 0.451012
R8398 Iout.n498 Iout.n497 0.451012
R8399 Iout.n497 Iout.n151 0.451012
R8400 Iout.n467 Iout.n151 0.451012
R8401 Iout.n467 Iout.n466 0.451012
R8402 Iout.n466 Iout.n158 0.451012
R8403 Iout.n436 Iout.n158 0.451012
R8404 Iout.n436 Iout.n113 0.451012
R8405 Iout.n592 Iout.n113 0.451012
R8406 Iout.n592 Iout.n591 0.451012
R8407 Iout.n591 Iout.n70 0.451012
R8408 Iout.n721 Iout.n70 0.451012
R8409 Iout.n721 Iout.n720 0.451012
R8410 Iout.n720 Iout.n27 0.451012
R8411 Iout.n900 Iout.n27 0.451012
R8412 Iout.n208 Iout.n185 0.451012
R8413 Iout.n274 Iout.n185 0.451012
R8414 Iout.n275 Iout.n274 0.451012
R8415 Iout.n275 Iout.n162 0.451012
R8416 Iout.n413 Iout.n162 0.451012
R8417 Iout.n414 Iout.n413 0.451012
R8418 Iout.n414 Iout.n98 0.451012
R8419 Iout.n621 Iout.n98 0.451012
R8420 Iout.n622 Iout.n621 0.451012
R8421 Iout.n622 Iout.n55 0.451012
R8422 Iout.n750 Iout.n55 0.451012
R8423 Iout.n751 Iout.n750 0.451012
R8424 Iout.n751 Iout.n32 0.451012
R8425 Iout.n865 Iout.n32 0.451012
R8426 Iout.n502 Iout.n139 0.451012
R8427 Iout.n528 Iout.n139 0.451012
R8428 Iout.n529 Iout.n528 0.451012
R8429 Iout.n529 Iout.n126 0.451012
R8430 Iout.n551 Iout.n126 0.451012
R8431 Iout.n552 Iout.n551 0.451012
R8432 Iout.n552 Iout.n116 0.451012
R8433 Iout.n585 Iout.n116 0.451012
R8434 Iout.n586 Iout.n585 0.451012
R8435 Iout.n586 Iout.n73 0.451012
R8436 Iout.n714 Iout.n73 0.451012
R8437 Iout.n715 Iout.n714 0.451012
R8438 Iout.n715 Iout.n26 0.451012
R8439 Iout.n907 Iout.n26 0.451012
R8440 Iout.n212 Iout.n182 0.451012
R8441 Iout.n281 Iout.n182 0.451012
R8442 Iout.n281 Iout.n280 0.451012
R8443 Iout.n280 Iout.n163 0.451012
R8444 Iout.n406 Iout.n163 0.451012
R8445 Iout.n406 Iout.n405 0.451012
R8446 Iout.n405 Iout.n95 0.451012
R8447 Iout.n628 Iout.n95 0.451012
R8448 Iout.n628 Iout.n627 0.451012
R8449 Iout.n627 Iout.n52 0.451012
R8450 Iout.n757 Iout.n52 0.451012
R8451 Iout.n757 Iout.n756 0.451012
R8452 Iout.n756 Iout.n33 0.451012
R8453 Iout.n858 Iout.n33 0.451012
R8454 Iout.n522 Iout.n145 0.451012
R8455 Iout.n523 Iout.n522 0.451012
R8456 Iout.n523 Iout.n132 0.451012
R8457 Iout.n545 Iout.n132 0.451012
R8458 Iout.n546 Iout.n545 0.451012
R8459 Iout.n546 Iout.n119 0.451012
R8460 Iout.n572 Iout.n119 0.451012
R8461 Iout.n580 Iout.n572 0.451012
R8462 Iout.n580 Iout.n579 0.451012
R8463 Iout.n579 Iout.n76 0.451012
R8464 Iout.n709 Iout.n76 0.451012
R8465 Iout.n709 Iout.n708 0.451012
R8466 Iout.n708 Iout.n25 0.451012
R8467 Iout.n914 Iout.n25 0.451012
R8468 Iout.n216 Iout.n179 0.451012
R8469 Iout.n286 Iout.n179 0.451012
R8470 Iout.n287 Iout.n286 0.451012
R8471 Iout.n287 Iout.n164 0.451012
R8472 Iout.n397 Iout.n164 0.451012
R8473 Iout.n398 Iout.n397 0.451012
R8474 Iout.n398 Iout.n92 0.451012
R8475 Iout.n633 Iout.n92 0.451012
R8476 Iout.n634 Iout.n633 0.451012
R8477 Iout.n634 Iout.n49 0.451012
R8478 Iout.n762 Iout.n49 0.451012
R8479 Iout.n763 Iout.n762 0.451012
R8480 Iout.n763 Iout.n34 0.451012
R8481 Iout.n851 Iout.n34 0.451012
R8482 Iout.n517 Iout.n516 0.451012
R8483 Iout.n517 Iout.n138 0.451012
R8484 Iout.n539 Iout.n138 0.451012
R8485 Iout.n540 Iout.n539 0.451012
R8486 Iout.n540 Iout.n125 0.451012
R8487 Iout.n562 Iout.n125 0.451012
R8488 Iout.n567 Iout.n562 0.451012
R8489 Iout.n567 Iout.n566 0.451012
R8490 Iout.n566 Iout.n79 0.451012
R8491 Iout.n698 Iout.n79 0.451012
R8492 Iout.n702 Iout.n698 0.451012
R8493 Iout.n703 Iout.n702 0.451012
R8494 Iout.n703 Iout.n24 0.451012
R8495 Iout.n921 Iout.n24 0.451012
R8496 Iout.n220 Iout.n176 0.451012
R8497 Iout.n293 Iout.n176 0.451012
R8498 Iout.n293 Iout.n292 0.451012
R8499 Iout.n292 Iout.n165 0.451012
R8500 Iout.n390 Iout.n165 0.451012
R8501 Iout.n390 Iout.n389 0.451012
R8502 Iout.n389 Iout.n89 0.451012
R8503 Iout.n640 Iout.n89 0.451012
R8504 Iout.n640 Iout.n639 0.451012
R8505 Iout.n639 Iout.n46 0.451012
R8506 Iout.n769 Iout.n46 0.451012
R8507 Iout.n769 Iout.n768 0.451012
R8508 Iout.n768 Iout.n35 0.451012
R8509 Iout.n844 Iout.n35 0.451012
R8510 Iout.n511 Iout.n2 0.451012
R8511 Iout.n1005 Iout.n2 0.451012
R8512 Iout.n1005 Iout.n1004 0.451012
R8513 Iout.n1004 Iout.n3 0.451012
R8514 Iout.n986 Iout.n3 0.451012
R8515 Iout.n986 Iout.n985 0.451012
R8516 Iout.n985 Iout.n8 0.451012
R8517 Iout.n967 Iout.n8 0.451012
R8518 Iout.n967 Iout.n966 0.451012
R8519 Iout.n966 Iout.n13 0.451012
R8520 Iout.n948 Iout.n13 0.451012
R8521 Iout.n948 Iout.n947 0.451012
R8522 Iout.n947 Iout.n18 0.451012
R8523 Iout.n929 Iout.n18 0.451012
R8524 Iout.n224 Iout.n170 0.451012
R8525 Iout.n298 Iout.n170 0.451012
R8526 Iout.n299 Iout.n298 0.451012
R8527 Iout.n299 Iout.n166 0.451012
R8528 Iout.n381 Iout.n166 0.451012
R8529 Iout.n382 Iout.n381 0.451012
R8530 Iout.n382 Iout.n83 0.451012
R8531 Iout.n645 Iout.n83 0.451012
R8532 Iout.n646 Iout.n645 0.451012
R8533 Iout.n646 Iout.n40 0.451012
R8534 Iout.n774 Iout.n40 0.451012
R8535 Iout.n775 Iout.n774 0.451012
R8536 Iout.n775 Iout.n36 0.451012
R8537 Iout.n837 Iout.n36 0.451012
R8538 Iout.n1018 Iout.n1017 0.451012
R8539 Iout.n1017 Iout.n0 0.451012
R8540 Iout.n999 Iout.n0 0.451012
R8541 Iout.n999 Iout.n998 0.451012
R8542 Iout.n998 Iout.n6 0.451012
R8543 Iout.n980 Iout.n6 0.451012
R8544 Iout.n980 Iout.n979 0.451012
R8545 Iout.n979 Iout.n11 0.451012
R8546 Iout.n961 Iout.n11 0.451012
R8547 Iout.n961 Iout.n960 0.451012
R8548 Iout.n960 Iout.n16 0.451012
R8549 Iout.n942 Iout.n16 0.451012
R8550 Iout.n942 Iout.n941 0.451012
R8551 Iout.n941 Iout.n21 0.451012
R8552 Iout.n230 Iout.n229 0.451012
R8553 Iout.n230 Iout.n167 0.451012
R8554 Iout.n304 Iout.n167 0.451012
R8555 Iout.n332 Iout.n304 0.451012
R8556 Iout.n374 Iout.n332 0.451012
R8557 Iout.n374 Iout.n373 0.451012
R8558 Iout.n373 Iout.n369 0.451012
R8559 Iout.n369 Iout.n80 0.451012
R8560 Iout.n651 Iout.n80 0.451012
R8561 Iout.n652 Iout.n651 0.451012
R8562 Iout.n652 Iout.n37 0.451012
R8563 Iout.n780 Iout.n37 0.451012
R8564 Iout.n826 Iout.n780 0.451012
R8565 Iout.n830 Iout.n826 0.451012
R8566 Iout.n231 Iout 0.2919
R8567 Iout.n303 Iout 0.2919
R8568 Iout Iout.n300 0.2919
R8569 Iout.n375 Iout 0.2919
R8570 Iout.n380 Iout 0.2919
R8571 Iout.n391 Iout 0.2919
R8572 Iout.n368 Iout 0.2919
R8573 Iout Iout.n365 0.2919
R8574 Iout Iout.n362 0.2919
R8575 Iout Iout.n359 0.2919
R8576 Iout.n650 Iout 0.2919
R8577 Iout Iout.n647 0.2919
R8578 Iout.n638 Iout 0.2919
R8579 Iout Iout.n635 0.2919
R8580 Iout.n626 Iout 0.2919
R8581 Iout.n41 Iout 0.2919
R8582 Iout.n773 Iout 0.2919
R8583 Iout Iout.n770 0.2919
R8584 Iout.n761 Iout 0.2919
R8585 Iout Iout.n758 0.2919
R8586 Iout.n749 Iout 0.2919
R8587 Iout.n825 Iout 0.2919
R8588 Iout Iout.n822 0.2919
R8589 Iout Iout.n819 0.2919
R8590 Iout Iout.n816 0.2919
R8591 Iout Iout.n813 0.2919
R8592 Iout Iout.n810 0.2919
R8593 Iout Iout.n807 0.2919
R8594 Iout.n829 Iout 0.2919
R8595 Iout.n838 Iout 0.2919
R8596 Iout.n843 Iout 0.2919
R8597 Iout.n852 Iout 0.2919
R8598 Iout.n857 Iout 0.2919
R8599 Iout.n866 Iout 0.2919
R8600 Iout.n871 Iout 0.2919
R8601 Iout.n880 Iout 0.2919
R8602 Iout Iout.n925 0.2919
R8603 Iout.n928 Iout 0.2919
R8604 Iout.n922 Iout 0.2919
R8605 Iout.n913 Iout 0.2919
R8606 Iout.n908 Iout 0.2919
R8607 Iout.n899 Iout 0.2919
R8608 Iout.n894 Iout 0.2919
R8609 Iout.n885 Iout 0.2919
R8610 Iout.n831 Iout 0.2919
R8611 Iout.n836 Iout 0.2919
R8612 Iout.n845 Iout 0.2919
R8613 Iout.n850 Iout 0.2919
R8614 Iout.n859 Iout 0.2919
R8615 Iout.n864 Iout 0.2919
R8616 Iout.n873 Iout 0.2919
R8617 Iout.n878 Iout 0.2919
R8618 Iout.n887 Iout 0.2919
R8619 Iout.n892 Iout 0.2919
R8620 Iout.n933 Iout 0.2919
R8621 Iout.n930 Iout 0.2919
R8622 Iout.n920 Iout 0.2919
R8623 Iout.n915 Iout 0.2919
R8624 Iout.n906 Iout 0.2919
R8625 Iout.n901 Iout 0.2919
R8626 Iout.n940 Iout 0.2919
R8627 Iout Iout.n783 0.2919
R8628 Iout Iout.n786 0.2919
R8629 Iout Iout.n789 0.2919
R8630 Iout Iout.n792 0.2919
R8631 Iout Iout.n795 0.2919
R8632 Iout Iout.n798 0.2919
R8633 Iout Iout.n801 0.2919
R8634 Iout Iout.n804 0.2919
R8635 Iout.n779 Iout 0.2919
R8636 Iout Iout.n776 0.2919
R8637 Iout.n767 Iout 0.2919
R8638 Iout Iout.n764 0.2919
R8639 Iout.n755 Iout 0.2919
R8640 Iout Iout.n752 0.2919
R8641 Iout.n743 Iout 0.2919
R8642 Iout Iout.n740 0.2919
R8643 Iout.n731 Iout 0.2919
R8644 Iout Iout.n728 0.2919
R8645 Iout.n719 Iout 0.2919
R8646 Iout Iout.n943 0.2919
R8647 Iout.n946 Iout 0.2919
R8648 Iout Iout.n704 0.2919
R8649 Iout.n707 Iout 0.2919
R8650 Iout Iout.n716 0.2919
R8651 Iout.n952 Iout 0.2919
R8652 Iout.n949 Iout 0.2919
R8653 Iout.n701 Iout 0.2919
R8654 Iout Iout.n710 0.2919
R8655 Iout.n713 Iout 0.2919
R8656 Iout Iout.n722 0.2919
R8657 Iout.n725 Iout 0.2919
R8658 Iout Iout.n734 0.2919
R8659 Iout.n737 Iout 0.2919
R8660 Iout Iout.n746 0.2919
R8661 Iout.n653 Iout 0.2919
R8662 Iout.n656 Iout 0.2919
R8663 Iout.n659 Iout 0.2919
R8664 Iout.n662 Iout 0.2919
R8665 Iout.n665 Iout 0.2919
R8666 Iout.n668 Iout 0.2919
R8667 Iout.n671 Iout 0.2919
R8668 Iout.n674 Iout 0.2919
R8669 Iout.n677 Iout 0.2919
R8670 Iout.n680 Iout 0.2919
R8671 Iout.n683 Iout 0.2919
R8672 Iout.n686 Iout 0.2919
R8673 Iout.n959 Iout 0.2919
R8674 Iout Iout.n694 0.2919
R8675 Iout.n697 Iout 0.2919
R8676 Iout.n689 Iout 0.2919
R8677 Iout Iout.n962 0.2919
R8678 Iout.n965 Iout 0.2919
R8679 Iout Iout.n575 0.2919
R8680 Iout.n578 Iout 0.2919
R8681 Iout Iout.n587 0.2919
R8682 Iout.n590 Iout 0.2919
R8683 Iout Iout.n599 0.2919
R8684 Iout.n602 Iout 0.2919
R8685 Iout Iout.n611 0.2919
R8686 Iout.n614 Iout 0.2919
R8687 Iout Iout.n623 0.2919
R8688 Iout.n84 Iout 0.2919
R8689 Iout.n644 Iout 0.2919
R8690 Iout Iout.n641 0.2919
R8691 Iout.n632 Iout 0.2919
R8692 Iout Iout.n629 0.2919
R8693 Iout.n620 Iout 0.2919
R8694 Iout Iout.n617 0.2919
R8695 Iout.n608 Iout 0.2919
R8696 Iout Iout.n605 0.2919
R8697 Iout.n596 Iout 0.2919
R8698 Iout Iout.n593 0.2919
R8699 Iout.n584 Iout 0.2919
R8700 Iout Iout.n581 0.2919
R8701 Iout.n971 Iout 0.2919
R8702 Iout.n968 Iout 0.2919
R8703 Iout.n565 Iout 0.2919
R8704 Iout.n978 Iout 0.2919
R8705 Iout Iout.n122 0.2919
R8706 Iout Iout.n568 0.2919
R8707 Iout.n571 Iout 0.2919
R8708 Iout Iout.n335 0.2919
R8709 Iout Iout.n338 0.2919
R8710 Iout Iout.n341 0.2919
R8711 Iout Iout.n344 0.2919
R8712 Iout Iout.n347 0.2919
R8713 Iout Iout.n350 0.2919
R8714 Iout Iout.n353 0.2919
R8715 Iout Iout.n356 0.2919
R8716 Iout.n372 Iout 0.2919
R8717 Iout.n383 Iout 0.2919
R8718 Iout.n388 Iout 0.2919
R8719 Iout.n399 Iout 0.2919
R8720 Iout.n404 Iout 0.2919
R8721 Iout.n415 Iout 0.2919
R8722 Iout.n420 Iout 0.2919
R8723 Iout.n431 Iout 0.2919
R8724 Iout.n443 Iout 0.2919
R8725 Iout Iout.n440 0.2919
R8726 Iout Iout.n437 0.2919
R8727 Iout.n553 Iout 0.2919
R8728 Iout.n556 Iout 0.2919
R8729 Iout.n561 Iout 0.2919
R8730 Iout Iout.n981 0.2919
R8731 Iout.n984 Iout 0.2919
R8732 Iout.n990 Iout 0.2919
R8733 Iout.n987 Iout 0.2919
R8734 Iout Iout.n129 0.2919
R8735 Iout Iout.n547 0.2919
R8736 Iout.n550 Iout 0.2919
R8737 Iout Iout.n451 0.2919
R8738 Iout.n454 Iout 0.2919
R8739 Iout.n446 Iout 0.2919
R8740 Iout.n428 Iout 0.2919
R8741 Iout.n423 Iout 0.2919
R8742 Iout.n412 Iout 0.2919
R8743 Iout.n407 Iout 0.2919
R8744 Iout.n396 Iout 0.2919
R8745 Iout.n331 Iout 0.2919
R8746 Iout Iout.n328 0.2919
R8747 Iout Iout.n325 0.2919
R8748 Iout Iout.n322 0.2919
R8749 Iout Iout.n319 0.2919
R8750 Iout Iout.n316 0.2919
R8751 Iout Iout.n313 0.2919
R8752 Iout Iout.n310 0.2919
R8753 Iout Iout.n307 0.2919
R8754 Iout.n457 Iout 0.2919
R8755 Iout.n465 Iout 0.2919
R8756 Iout Iout.n462 0.2919
R8757 Iout.n544 Iout 0.2919
R8758 Iout Iout.n541 0.2919
R8759 Iout Iout.n135 0.2919
R8760 Iout.n997 Iout 0.2919
R8761 Iout Iout.n1000 0.2919
R8762 Iout.n1003 Iout 0.2919
R8763 Iout.n538 Iout 0.2919
R8764 Iout.n533 Iout 0.2919
R8765 Iout.n530 Iout 0.2919
R8766 Iout Iout.n468 0.2919
R8767 Iout Iout.n471 0.2919
R8768 Iout.n474 Iout 0.2919
R8769 Iout Iout.n264 0.2919
R8770 Iout.n267 Iout 0.2919
R8771 Iout Iout.n276 0.2919
R8772 Iout.n279 Iout 0.2919
R8773 Iout Iout.n288 0.2919
R8774 Iout.n291 Iout 0.2919
R8775 Iout.n171 Iout 0.2919
R8776 Iout.n297 Iout 0.2919
R8777 Iout Iout.n294 0.2919
R8778 Iout.n285 Iout 0.2919
R8779 Iout Iout.n282 0.2919
R8780 Iout.n273 Iout 0.2919
R8781 Iout Iout.n270 0.2919
R8782 Iout.n261 Iout 0.2919
R8783 Iout.n477 Iout 0.2919
R8784 Iout.n485 Iout 0.2919
R8785 Iout Iout.n482 0.2919
R8786 Iout.n527 Iout 0.2919
R8787 Iout Iout.n524 0.2919
R8788 Iout Iout.n142 0.2919
R8789 Iout.n1006 Iout 0.2919
R8790 Iout.n1009 Iout 0.2919
R8791 Iout.n1016 Iout 0.2919
R8792 Iout Iout.n148 0.2919
R8793 Iout Iout.n518 0.2919
R8794 Iout.n521 Iout 0.2919
R8795 Iout Iout.n493 0.2919
R8796 Iout.n496 Iout 0.2919
R8797 Iout.n488 Iout 0.2919
R8798 Iout Iout.n254 0.2919
R8799 Iout.n257 Iout 0.2919
R8800 Iout.n249 Iout 0.2919
R8801 Iout.n246 Iout 0.2919
R8802 Iout.n243 Iout 0.2919
R8803 Iout.n240 Iout 0.2919
R8804 Iout.n237 Iout 0.2919
R8805 Iout.n234 Iout 0.2919
R8806 Iout.n228 Iout 0.2919
R8807 Iout Iout.n225 0.2919
R8808 Iout Iout.n221 0.2919
R8809 Iout Iout.n217 0.2919
R8810 Iout Iout.n213 0.2919
R8811 Iout Iout.n209 0.2919
R8812 Iout Iout.n205 0.2919
R8813 Iout Iout.n201 0.2919
R8814 Iout Iout.n198 0.2919
R8815 Iout Iout.n194 0.2919
R8816 Iout.n499 Iout 0.2919
R8817 Iout.n503 Iout 0.2919
R8818 Iout.n506 Iout 0.2919
R8819 Iout.n515 Iout 0.2919
R8820 Iout Iout.n512 0.2919
R8821 Iout.n1019 Iout 0.2919
R8822 Iout.n1013 Iout.n1012 0.092855
R8823 Iout.n1012 Iout.n1 0.092855
R8824 Iout.n994 Iout.n1 0.092855
R8825 Iout.n994 Iout.n993 0.092855
R8826 Iout.n993 Iout.n7 0.092855
R8827 Iout.n975 Iout.n7 0.092855
R8828 Iout.n975 Iout.n974 0.092855
R8829 Iout.n974 Iout.n12 0.092855
R8830 Iout.n956 Iout.n12 0.092855
R8831 Iout.n956 Iout.n955 0.092855
R8832 Iout.n955 Iout.n17 0.092855
R8833 Iout.n937 Iout.n17 0.092855
R8834 Iout.n937 Iout.n936 0.092855
R8835 Iout.n197 Iout 0.0818902
R8836 Iout.n191 Iout 0.0818902
R8837 Iout.n152 Iout 0.0818902
R8838 Iout.n204 Iout 0.0818902
R8839 Iout.n498 Iout 0.0818902
R8840 Iout.n208 Iout 0.0818902
R8841 Iout.n502 Iout 0.0818902
R8842 Iout.n212 Iout 0.0818902
R8843 Iout.n145 Iout 0.0818902
R8844 Iout.n216 Iout 0.0818902
R8845 Iout.n516 Iout 0.0818902
R8846 Iout.n220 Iout 0.0818902
R8847 Iout.n511 Iout 0.0818902
R8848 Iout.n224 Iout 0.0818902
R8849 Iout.n1018 Iout 0.0818902
R8850 Iout.n229 Iout 0.0818902
R8851 Iout.n1013 Iout 0.072645
R8852 Iout.n302 Iout 0.0532071
R8853 Iout Iout.n377 0.0532071
R8854 Iout.n379 Iout 0.0532071
R8855 Iout.n367 Iout 0.0532071
R8856 Iout.n364 Iout 0.0532071
R8857 Iout.n361 Iout 0.0532071
R8858 Iout.n649 Iout 0.0532071
R8859 Iout Iout.n82 0.0532071
R8860 Iout.n637 Iout 0.0532071
R8861 Iout Iout.n91 0.0532071
R8862 Iout Iout.n43 0.0532071
R8863 Iout.n772 Iout 0.0532071
R8864 Iout Iout.n45 0.0532071
R8865 Iout.n760 Iout 0.0532071
R8866 Iout Iout.n51 0.0532071
R8867 Iout.n824 Iout 0.0532071
R8868 Iout.n821 Iout 0.0532071
R8869 Iout.n818 Iout 0.0532071
R8870 Iout.n815 Iout 0.0532071
R8871 Iout.n812 Iout 0.0532071
R8872 Iout.n809 Iout 0.0532071
R8873 Iout.n828 Iout 0.0532071
R8874 Iout Iout.n840 0.0532071
R8875 Iout.n842 Iout 0.0532071
R8876 Iout Iout.n854 0.0532071
R8877 Iout.n856 Iout 0.0532071
R8878 Iout Iout.n868 0.0532071
R8879 Iout.n870 Iout 0.0532071
R8880 Iout.n927 Iout 0.0532071
R8881 Iout Iout.n924 0.0532071
R8882 Iout.n912 Iout 0.0532071
R8883 Iout Iout.n910 0.0532071
R8884 Iout.n898 Iout 0.0532071
R8885 Iout Iout.n896 0.0532071
R8886 Iout.n884 Iout 0.0532071
R8887 Iout Iout.n882 0.0532071
R8888 Iout Iout.n833 0.0532071
R8889 Iout.n835 Iout 0.0532071
R8890 Iout Iout.n847 0.0532071
R8891 Iout.n849 Iout 0.0532071
R8892 Iout Iout.n861 0.0532071
R8893 Iout.n863 Iout 0.0532071
R8894 Iout Iout.n875 0.0532071
R8895 Iout.n877 Iout 0.0532071
R8896 Iout Iout.n889 0.0532071
R8897 Iout Iout.n932 0.0532071
R8898 Iout.n919 Iout 0.0532071
R8899 Iout Iout.n917 0.0532071
R8900 Iout.n905 Iout 0.0532071
R8901 Iout Iout.n903 0.0532071
R8902 Iout.n891 Iout 0.0532071
R8903 Iout.n782 Iout 0.0532071
R8904 Iout.n785 Iout 0.0532071
R8905 Iout.n788 Iout 0.0532071
R8906 Iout.n791 Iout 0.0532071
R8907 Iout.n794 Iout 0.0532071
R8908 Iout.n797 Iout 0.0532071
R8909 Iout.n800 Iout 0.0532071
R8910 Iout.n803 Iout 0.0532071
R8911 Iout.n806 Iout 0.0532071
R8912 Iout.n778 Iout 0.0532071
R8913 Iout Iout.n39 0.0532071
R8914 Iout.n766 Iout 0.0532071
R8915 Iout Iout.n48 0.0532071
R8916 Iout.n754 Iout 0.0532071
R8917 Iout Iout.n54 0.0532071
R8918 Iout.n742 Iout 0.0532071
R8919 Iout Iout.n60 0.0532071
R8920 Iout.n730 Iout 0.0532071
R8921 Iout Iout.n66 0.0532071
R8922 Iout.n945 Iout 0.0532071
R8923 Iout.n78 Iout 0.0532071
R8924 Iout.n706 Iout 0.0532071
R8925 Iout Iout.n72 0.0532071
R8926 Iout.n718 Iout 0.0532071
R8927 Iout Iout.n951 0.0532071
R8928 Iout.n700 Iout 0.0532071
R8929 Iout Iout.n75 0.0532071
R8930 Iout.n712 Iout 0.0532071
R8931 Iout Iout.n69 0.0532071
R8932 Iout.n724 Iout 0.0532071
R8933 Iout Iout.n63 0.0532071
R8934 Iout.n736 Iout 0.0532071
R8935 Iout Iout.n57 0.0532071
R8936 Iout.n748 Iout 0.0532071
R8937 Iout Iout.n655 0.0532071
R8938 Iout Iout.n658 0.0532071
R8939 Iout Iout.n661 0.0532071
R8940 Iout Iout.n664 0.0532071
R8941 Iout Iout.n667 0.0532071
R8942 Iout Iout.n670 0.0532071
R8943 Iout Iout.n673 0.0532071
R8944 Iout Iout.n676 0.0532071
R8945 Iout Iout.n679 0.0532071
R8946 Iout Iout.n682 0.0532071
R8947 Iout Iout.n685 0.0532071
R8948 Iout.n693 Iout 0.0532071
R8949 Iout.n696 Iout 0.0532071
R8950 Iout Iout.n691 0.0532071
R8951 Iout Iout.n688 0.0532071
R8952 Iout.n964 Iout 0.0532071
R8953 Iout.n574 Iout 0.0532071
R8954 Iout.n577 Iout 0.0532071
R8955 Iout Iout.n115 0.0532071
R8956 Iout.n589 Iout 0.0532071
R8957 Iout Iout.n109 0.0532071
R8958 Iout.n601 Iout 0.0532071
R8959 Iout Iout.n103 0.0532071
R8960 Iout.n613 Iout 0.0532071
R8961 Iout Iout.n97 0.0532071
R8962 Iout.n625 Iout 0.0532071
R8963 Iout Iout.n86 0.0532071
R8964 Iout.n643 Iout 0.0532071
R8965 Iout Iout.n88 0.0532071
R8966 Iout.n631 Iout 0.0532071
R8967 Iout Iout.n94 0.0532071
R8968 Iout.n619 Iout 0.0532071
R8969 Iout Iout.n100 0.0532071
R8970 Iout.n607 Iout 0.0532071
R8971 Iout Iout.n106 0.0532071
R8972 Iout.n595 Iout 0.0532071
R8973 Iout Iout.n112 0.0532071
R8974 Iout.n583 Iout 0.0532071
R8975 Iout Iout.n970 0.0532071
R8976 Iout.n564 Iout 0.0532071
R8977 Iout Iout.n118 0.0532071
R8978 Iout.n121 Iout 0.0532071
R8979 Iout.n124 Iout 0.0532071
R8980 Iout.n570 Iout 0.0532071
R8981 Iout.n334 Iout 0.0532071
R8982 Iout.n337 Iout 0.0532071
R8983 Iout.n340 Iout 0.0532071
R8984 Iout.n343 Iout 0.0532071
R8985 Iout.n346 Iout 0.0532071
R8986 Iout.n349 Iout 0.0532071
R8987 Iout.n352 Iout 0.0532071
R8988 Iout.n355 Iout 0.0532071
R8989 Iout.n358 Iout 0.0532071
R8990 Iout.n371 Iout 0.0532071
R8991 Iout Iout.n385 0.0532071
R8992 Iout.n387 Iout 0.0532071
R8993 Iout Iout.n401 0.0532071
R8994 Iout.n403 Iout 0.0532071
R8995 Iout Iout.n417 0.0532071
R8996 Iout.n419 Iout 0.0532071
R8997 Iout Iout.n433 0.0532071
R8998 Iout.n442 Iout 0.0532071
R8999 Iout.n439 Iout 0.0532071
R9000 Iout.n435 Iout 0.0532071
R9001 Iout Iout.n555 0.0532071
R9002 Iout Iout.n558 0.0532071
R9003 Iout.n983 Iout 0.0532071
R9004 Iout.n560 Iout 0.0532071
R9005 Iout Iout.n989 0.0532071
R9006 Iout.n128 Iout 0.0532071
R9007 Iout.n131 Iout 0.0532071
R9008 Iout.n549 Iout 0.0532071
R9009 Iout.n450 Iout 0.0532071
R9010 Iout.n453 Iout 0.0532071
R9011 Iout Iout.n448 0.0532071
R9012 Iout.n427 Iout 0.0532071
R9013 Iout Iout.n425 0.0532071
R9014 Iout.n411 Iout 0.0532071
R9015 Iout Iout.n409 0.0532071
R9016 Iout.n395 Iout 0.0532071
R9017 Iout Iout.n393 0.0532071
R9018 Iout.n330 Iout 0.0532071
R9019 Iout.n327 Iout 0.0532071
R9020 Iout.n324 Iout 0.0532071
R9021 Iout.n321 Iout 0.0532071
R9022 Iout.n318 Iout 0.0532071
R9023 Iout.n315 Iout 0.0532071
R9024 Iout.n312 Iout 0.0532071
R9025 Iout.n309 Iout 0.0532071
R9026 Iout.n306 Iout 0.0532071
R9027 Iout Iout.n459 0.0532071
R9028 Iout.n464 Iout 0.0532071
R9029 Iout.n461 Iout 0.0532071
R9030 Iout.n543 Iout 0.0532071
R9031 Iout.n137 Iout 0.0532071
R9032 Iout.n134 Iout 0.0532071
R9033 Iout.n1002 Iout 0.0532071
R9034 Iout.n537 Iout 0.0532071
R9035 Iout Iout.n535 0.0532071
R9036 Iout Iout.n532 0.0532071
R9037 Iout.n157 Iout 0.0532071
R9038 Iout.n470 Iout 0.0532071
R9039 Iout.n473 Iout 0.0532071
R9040 Iout.n190 Iout 0.0532071
R9041 Iout.n266 Iout 0.0532071
R9042 Iout Iout.n184 0.0532071
R9043 Iout.n278 Iout 0.0532071
R9044 Iout Iout.n178 0.0532071
R9045 Iout.n290 Iout 0.0532071
R9046 Iout Iout.n169 0.0532071
R9047 Iout Iout.n173 0.0532071
R9048 Iout.n296 Iout 0.0532071
R9049 Iout Iout.n175 0.0532071
R9050 Iout.n284 Iout 0.0532071
R9051 Iout Iout.n181 0.0532071
R9052 Iout.n272 Iout 0.0532071
R9053 Iout Iout.n187 0.0532071
R9054 Iout.n260 Iout 0.0532071
R9055 Iout Iout.n479 0.0532071
R9056 Iout.n484 Iout 0.0532071
R9057 Iout.n481 Iout 0.0532071
R9058 Iout.n526 Iout 0.0532071
R9059 Iout.n144 Iout 0.0532071
R9060 Iout.n141 Iout 0.0532071
R9061 Iout Iout.n1008 0.0532071
R9062 Iout.n147 Iout 0.0532071
R9063 Iout.n150 Iout 0.0532071
R9064 Iout.n520 Iout 0.0532071
R9065 Iout.n492 Iout 0.0532071
R9066 Iout.n495 Iout 0.0532071
R9067 Iout Iout.n490 0.0532071
R9068 Iout.n253 Iout 0.0532071
R9069 Iout.n256 Iout 0.0532071
R9070 Iout Iout.n251 0.0532071
R9071 Iout Iout.n248 0.0532071
R9072 Iout Iout.n245 0.0532071
R9073 Iout Iout.n242 0.0532071
R9074 Iout Iout.n239 0.0532071
R9075 Iout Iout.n236 0.0532071
R9076 Iout Iout.n233 0.0532071
R9077 Iout.n227 Iout 0.0532071
R9078 Iout.n223 Iout 0.0532071
R9079 Iout.n219 Iout 0.0532071
R9080 Iout.n215 Iout 0.0532071
R9081 Iout.n211 Iout 0.0532071
R9082 Iout.n207 Iout 0.0532071
R9083 Iout.n203 Iout 0.0532071
R9084 Iout.n200 Iout 0.0532071
R9085 Iout.n196 Iout 0.0532071
R9086 Iout.n193 Iout 0.0532071
R9087 Iout Iout.n501 0.0532071
R9088 Iout Iout.n505 0.0532071
R9089 Iout Iout.n508 0.0532071
R9090 Iout.n514 Iout 0.0532071
R9091 Iout.n510 Iout 0.0532071
R9092 Iout.n1020 Iout 0.03925
R9093 Iout.n509 Iout 0.03925
R9094 Iout.n513 Iout 0.03925
R9095 Iout.n507 Iout 0.03925
R9096 Iout.n504 Iout 0.03925
R9097 Iout.n500 Iout 0.03925
R9098 Iout.n192 Iout 0.03925
R9099 Iout.n195 Iout 0.03925
R9100 Iout.n199 Iout 0.03925
R9101 Iout.n202 Iout 0.03925
R9102 Iout.n206 Iout 0.03925
R9103 Iout.n210 Iout 0.03925
R9104 Iout.n214 Iout 0.03925
R9105 Iout.n218 Iout 0.03925
R9106 Iout.n222 Iout 0.03925
R9107 Iout.n226 Iout 0.03925
R9108 Iout.n232 Iout 0.03925
R9109 Iout.n235 Iout 0.03925
R9110 Iout.n238 Iout 0.03925
R9111 Iout.n241 Iout 0.03925
R9112 Iout.n244 Iout 0.03925
R9113 Iout.n247 Iout 0.03925
R9114 Iout.n250 Iout 0.03925
R9115 Iout.n255 Iout 0.03925
R9116 Iout.n252 Iout 0.03925
R9117 Iout.n489 Iout 0.03925
R9118 Iout.n494 Iout 0.03925
R9119 Iout.n491 Iout 0.03925
R9120 Iout.n519 Iout 0.03925
R9121 Iout.n149 Iout 0.03925
R9122 Iout.n146 Iout 0.03925
R9123 Iout.n1010 Iout 0.03925
R9124 Iout.n1007 Iout 0.03925
R9125 Iout.n140 Iout 0.03925
R9126 Iout.n143 Iout 0.03925
R9127 Iout.n525 Iout 0.03925
R9128 Iout.n480 Iout 0.03925
R9129 Iout.n483 Iout 0.03925
R9130 Iout.n478 Iout 0.03925
R9131 Iout.n259 Iout 0.03925
R9132 Iout.n186 Iout 0.03925
R9133 Iout.n271 Iout 0.03925
R9134 Iout.n180 Iout 0.03925
R9135 Iout.n283 Iout 0.03925
R9136 Iout.n174 Iout 0.03925
R9137 Iout.n168 Iout 0.03925
R9138 Iout.n301 Iout 0.03925
R9139 Iout.n289 Iout 0.03925
R9140 Iout.n177 Iout 0.03925
R9141 Iout.n277 Iout 0.03925
R9142 Iout.n183 Iout 0.03925
R9143 Iout.n265 Iout 0.03925
R9144 Iout.n189 Iout 0.03925
R9145 Iout.n472 Iout 0.03925
R9146 Iout.n469 Iout 0.03925
R9147 Iout.n156 Iout 0.03925
R9148 Iout.n531 Iout 0.03925
R9149 Iout.n534 Iout 0.03925
R9150 Iout.n536 Iout 0.03925
R9151 Iout.n133 Iout 0.03925
R9152 Iout.n136 Iout 0.03925
R9153 Iout.n542 Iout 0.03925
R9154 Iout.n460 Iout 0.03925
R9155 Iout.n463 Iout 0.03925
R9156 Iout.n458 Iout 0.03925
R9157 Iout.n305 Iout 0.03925
R9158 Iout.n308 Iout 0.03925
R9159 Iout.n311 Iout 0.03925
R9160 Iout.n314 Iout 0.03925
R9161 Iout.n317 Iout 0.03925
R9162 Iout.n320 Iout 0.03925
R9163 Iout.n392 Iout 0.03925
R9164 Iout.n378 Iout 0.03925
R9165 Iout.n376 Iout 0.03925
R9166 Iout.n394 Iout 0.03925
R9167 Iout.n408 Iout 0.03925
R9168 Iout.n410 Iout 0.03925
R9169 Iout.n424 Iout 0.03925
R9170 Iout.n426 Iout 0.03925
R9171 Iout.n447 Iout 0.03925
R9172 Iout.n452 Iout 0.03925
R9173 Iout.n449 Iout 0.03925
R9174 Iout.n548 Iout 0.03925
R9175 Iout.n130 Iout 0.03925
R9176 Iout.n559 Iout 0.03925
R9177 Iout.n557 Iout 0.03925
R9178 Iout.n554 Iout 0.03925
R9179 Iout.n434 Iout 0.03925
R9180 Iout.n438 Iout 0.03925
R9181 Iout.n441 Iout 0.03925
R9182 Iout.n432 Iout 0.03925
R9183 Iout.n418 Iout 0.03925
R9184 Iout.n416 Iout 0.03925
R9185 Iout.n402 Iout 0.03925
R9186 Iout.n357 Iout 0.03925
R9187 Iout.n360 Iout 0.03925
R9188 Iout.n363 Iout 0.03925
R9189 Iout.n366 Iout 0.03925
R9190 Iout.n354 Iout 0.03925
R9191 Iout.n351 Iout 0.03925
R9192 Iout.n348 Iout 0.03925
R9193 Iout.n345 Iout 0.03925
R9194 Iout.n342 Iout 0.03925
R9195 Iout.n339 Iout 0.03925
R9196 Iout.n336 Iout 0.03925
R9197 Iout.n333 Iout 0.03925
R9198 Iout.n117 Iout 0.03925
R9199 Iout.n582 Iout 0.03925
R9200 Iout.n111 Iout 0.03925
R9201 Iout.n594 Iout 0.03925
R9202 Iout.n105 Iout 0.03925
R9203 Iout.n606 Iout 0.03925
R9204 Iout.n99 Iout 0.03925
R9205 Iout.n618 Iout 0.03925
R9206 Iout.n624 Iout 0.03925
R9207 Iout.n90 Iout 0.03925
R9208 Iout.n636 Iout 0.03925
R9209 Iout.n81 Iout 0.03925
R9210 Iout.n648 Iout 0.03925
R9211 Iout.n96 Iout 0.03925
R9212 Iout.n612 Iout 0.03925
R9213 Iout.n102 Iout 0.03925
R9214 Iout.n600 Iout 0.03925
R9215 Iout.n108 Iout 0.03925
R9216 Iout.n588 Iout 0.03925
R9217 Iout.n687 Iout 0.03925
R9218 Iout.n684 Iout 0.03925
R9219 Iout.n681 Iout 0.03925
R9220 Iout.n678 Iout 0.03925
R9221 Iout.n675 Iout 0.03925
R9222 Iout.n672 Iout 0.03925
R9223 Iout.n747 Iout 0.03925
R9224 Iout.n50 Iout 0.03925
R9225 Iout.n759 Iout 0.03925
R9226 Iout.n44 Iout 0.03925
R9227 Iout.n771 Iout 0.03925
R9228 Iout.n42 Iout 0.03925
R9229 Iout.n56 Iout 0.03925
R9230 Iout.n735 Iout 0.03925
R9231 Iout.n62 Iout 0.03925
R9232 Iout.n723 Iout 0.03925
R9233 Iout.n717 Iout 0.03925
R9234 Iout.n65 Iout 0.03925
R9235 Iout.n729 Iout 0.03925
R9236 Iout.n59 Iout 0.03925
R9237 Iout.n805 Iout 0.03925
R9238 Iout.n808 Iout 0.03925
R9239 Iout.n811 Iout 0.03925
R9240 Iout.n814 Iout 0.03925
R9241 Iout.n817 Iout 0.03925
R9242 Iout.n820 Iout 0.03925
R9243 Iout.n823 Iout 0.03925
R9244 Iout.n802 Iout 0.03925
R9245 Iout.n799 Iout 0.03925
R9246 Iout.n890 Iout 0.03925
R9247 Iout.n888 Iout 0.03925
R9248 Iout.n881 Iout 0.03925
R9249 Iout.n869 Iout 0.03925
R9250 Iout.n867 Iout 0.03925
R9251 Iout.n855 Iout 0.03925
R9252 Iout.n853 Iout 0.03925
R9253 Iout.n841 Iout 0.03925
R9254 Iout.n839 Iout 0.03925
R9255 Iout.n827 Iout 0.03925
R9256 Iout.n883 Iout 0.03925
R9257 Iout.n895 Iout 0.03925
R9258 Iout.n897 Iout 0.03925
R9259 Iout.n909 Iout 0.03925
R9260 Iout.n911 Iout 0.03925
R9261 Iout.n923 Iout 0.03925
R9262 Iout.n926 Iout 0.03925
R9263 Iout.n22 Iout 0.03925
R9264 Iout.n876 Iout 0.03925
R9265 Iout.n874 Iout 0.03925
R9266 Iout.n862 Iout 0.03925
R9267 Iout.n860 Iout 0.03925
R9268 Iout.n848 Iout 0.03925
R9269 Iout.n846 Iout 0.03925
R9270 Iout.n834 Iout 0.03925
R9271 Iout.n832 Iout 0.03925
R9272 Iout.n902 Iout 0.03925
R9273 Iout.n904 Iout 0.03925
R9274 Iout.n916 Iout 0.03925
R9275 Iout.n918 Iout 0.03925
R9276 Iout.n931 Iout 0.03925
R9277 Iout.n934 Iout 0.03925
R9278 Iout.n796 Iout 0.03925
R9279 Iout.n793 Iout 0.03925
R9280 Iout.n790 Iout 0.03925
R9281 Iout.n787 Iout 0.03925
R9282 Iout.n784 Iout 0.03925
R9283 Iout.n781 Iout 0.03925
R9284 Iout.n938 Iout 0.03925
R9285 Iout.n741 Iout 0.03925
R9286 Iout.n53 Iout 0.03925
R9287 Iout.n753 Iout 0.03925
R9288 Iout.n47 Iout 0.03925
R9289 Iout.n765 Iout 0.03925
R9290 Iout.n38 Iout 0.03925
R9291 Iout.n777 Iout 0.03925
R9292 Iout.n71 Iout 0.03925
R9293 Iout.n705 Iout 0.03925
R9294 Iout.n77 Iout 0.03925
R9295 Iout.n944 Iout 0.03925
R9296 Iout.n19 Iout 0.03925
R9297 Iout.n68 Iout 0.03925
R9298 Iout.n711 Iout 0.03925
R9299 Iout.n74 Iout 0.03925
R9300 Iout.n699 Iout 0.03925
R9301 Iout.n950 Iout 0.03925
R9302 Iout.n953 Iout 0.03925
R9303 Iout.n669 Iout 0.03925
R9304 Iout.n666 Iout 0.03925
R9305 Iout.n663 Iout 0.03925
R9306 Iout.n660 Iout 0.03925
R9307 Iout.n657 Iout 0.03925
R9308 Iout.n654 Iout 0.03925
R9309 Iout.n690 Iout 0.03925
R9310 Iout.n695 Iout 0.03925
R9311 Iout.n692 Iout 0.03925
R9312 Iout.n957 Iout 0.03925
R9313 Iout.n114 Iout 0.03925
R9314 Iout.n576 Iout 0.03925
R9315 Iout.n573 Iout 0.03925
R9316 Iout.n963 Iout 0.03925
R9317 Iout.n14 Iout 0.03925
R9318 Iout.n93 Iout 0.03925
R9319 Iout.n630 Iout 0.03925
R9320 Iout.n87 Iout 0.03925
R9321 Iout.n642 Iout 0.03925
R9322 Iout.n85 Iout 0.03925
R9323 Iout.n563 Iout 0.03925
R9324 Iout.n969 Iout 0.03925
R9325 Iout.n972 Iout 0.03925
R9326 Iout.n569 Iout 0.03925
R9327 Iout.n123 Iout 0.03925
R9328 Iout.n120 Iout 0.03925
R9329 Iout.n976 Iout 0.03925
R9330 Iout.n400 Iout 0.03925
R9331 Iout.n386 Iout 0.03925
R9332 Iout.n384 Iout 0.03925
R9333 Iout.n370 Iout 0.03925
R9334 Iout.n982 Iout 0.03925
R9335 Iout.n9 Iout 0.03925
R9336 Iout.n127 Iout 0.03925
R9337 Iout.n988 Iout 0.03925
R9338 Iout.n991 Iout 0.03925
R9339 Iout.n323 Iout 0.03925
R9340 Iout.n326 Iout 0.03925
R9341 Iout.n329 Iout 0.03925
R9342 Iout.n995 Iout 0.03925
R9343 Iout.n1001 Iout 0.03925
R9344 Iout.n4 Iout 0.03925
R9345 Iout.n295 Iout 0.03925
R9346 Iout.n172 Iout 0.03925
R9347 Iout.n1014 Iout 0.03925
R9348 Iout.n1022 Iout 0.02071
R9349 Iout Iout.n1022 0.00379
R9350 Iout.n303 Iout.n302 0.00105952
R9351 Iout.n377 Iout.n375 0.00105952
R9352 Iout.n380 Iout.n379 0.00105952
R9353 Iout.n368 Iout.n367 0.00105952
R9354 Iout.n365 Iout.n364 0.00105952
R9355 Iout.n362 Iout.n361 0.00105952
R9356 Iout.n650 Iout.n649 0.00105952
R9357 Iout.n647 Iout.n82 0.00105952
R9358 Iout.n638 Iout.n637 0.00105952
R9359 Iout.n635 Iout.n91 0.00105952
R9360 Iout.n43 Iout.n41 0.00105952
R9361 Iout.n773 Iout.n772 0.00105952
R9362 Iout.n770 Iout.n45 0.00105952
R9363 Iout.n761 Iout.n760 0.00105952
R9364 Iout.n758 Iout.n51 0.00105952
R9365 Iout.n825 Iout.n824 0.00105952
R9366 Iout.n822 Iout.n821 0.00105952
R9367 Iout.n819 Iout.n818 0.00105952
R9368 Iout.n816 Iout.n815 0.00105952
R9369 Iout.n813 Iout.n812 0.00105952
R9370 Iout.n810 Iout.n809 0.00105952
R9371 Iout.n829 Iout.n828 0.00105952
R9372 Iout.n840 Iout.n838 0.00105952
R9373 Iout.n843 Iout.n842 0.00105952
R9374 Iout.n854 Iout.n852 0.00105952
R9375 Iout.n857 Iout.n856 0.00105952
R9376 Iout.n868 Iout.n866 0.00105952
R9377 Iout.n871 Iout.n870 0.00105952
R9378 Iout.n925 Iout.n23 0.00105952
R9379 Iout.n928 Iout.n927 0.00105952
R9380 Iout.n924 Iout.n922 0.00105952
R9381 Iout.n913 Iout.n912 0.00105952
R9382 Iout.n910 Iout.n908 0.00105952
R9383 Iout.n899 Iout.n898 0.00105952
R9384 Iout.n896 Iout.n894 0.00105952
R9385 Iout.n885 Iout.n884 0.00105952
R9386 Iout.n882 Iout.n880 0.00105952
R9387 Iout.n833 Iout.n831 0.00105952
R9388 Iout.n836 Iout.n835 0.00105952
R9389 Iout.n847 Iout.n845 0.00105952
R9390 Iout.n850 Iout.n849 0.00105952
R9391 Iout.n861 Iout.n859 0.00105952
R9392 Iout.n864 Iout.n863 0.00105952
R9393 Iout.n875 Iout.n873 0.00105952
R9394 Iout.n878 Iout.n877 0.00105952
R9395 Iout.n889 Iout.n887 0.00105952
R9396 Iout.n935 Iout.n933 0.00105952
R9397 Iout.n932 Iout.n930 0.00105952
R9398 Iout.n920 Iout.n919 0.00105952
R9399 Iout.n917 Iout.n915 0.00105952
R9400 Iout.n906 Iout.n905 0.00105952
R9401 Iout.n903 Iout.n901 0.00105952
R9402 Iout.n892 Iout.n891 0.00105952
R9403 Iout.n940 Iout.n939 0.00105952
R9404 Iout.n783 Iout.n782 0.00105952
R9405 Iout.n786 Iout.n785 0.00105952
R9406 Iout.n789 Iout.n788 0.00105952
R9407 Iout.n792 Iout.n791 0.00105952
R9408 Iout.n795 Iout.n794 0.00105952
R9409 Iout.n798 Iout.n797 0.00105952
R9410 Iout.n801 Iout.n800 0.00105952
R9411 Iout.n804 Iout.n803 0.00105952
R9412 Iout.n807 Iout.n806 0.00105952
R9413 Iout.n779 Iout.n778 0.00105952
R9414 Iout.n776 Iout.n39 0.00105952
R9415 Iout.n767 Iout.n766 0.00105952
R9416 Iout.n764 Iout.n48 0.00105952
R9417 Iout.n755 Iout.n754 0.00105952
R9418 Iout.n752 Iout.n54 0.00105952
R9419 Iout.n743 Iout.n742 0.00105952
R9420 Iout.n740 Iout.n60 0.00105952
R9421 Iout.n731 Iout.n730 0.00105952
R9422 Iout.n728 Iout.n66 0.00105952
R9423 Iout.n943 Iout.n20 0.00105952
R9424 Iout.n946 Iout.n945 0.00105952
R9425 Iout.n704 Iout.n78 0.00105952
R9426 Iout.n707 Iout.n706 0.00105952
R9427 Iout.n716 Iout.n72 0.00105952
R9428 Iout.n719 Iout.n718 0.00105952
R9429 Iout.n954 Iout.n952 0.00105952
R9430 Iout.n951 Iout.n949 0.00105952
R9431 Iout.n701 Iout.n700 0.00105952
R9432 Iout.n710 Iout.n75 0.00105952
R9433 Iout.n713 Iout.n712 0.00105952
R9434 Iout.n722 Iout.n69 0.00105952
R9435 Iout.n725 Iout.n724 0.00105952
R9436 Iout.n734 Iout.n63 0.00105952
R9437 Iout.n737 Iout.n736 0.00105952
R9438 Iout.n746 Iout.n57 0.00105952
R9439 Iout.n749 Iout.n748 0.00105952
R9440 Iout.n655 Iout.n653 0.00105952
R9441 Iout.n658 Iout.n656 0.00105952
R9442 Iout.n661 Iout.n659 0.00105952
R9443 Iout.n664 Iout.n662 0.00105952
R9444 Iout.n667 Iout.n665 0.00105952
R9445 Iout.n670 Iout.n668 0.00105952
R9446 Iout.n673 Iout.n671 0.00105952
R9447 Iout.n676 Iout.n674 0.00105952
R9448 Iout.n679 Iout.n677 0.00105952
R9449 Iout.n682 Iout.n680 0.00105952
R9450 Iout.n685 Iout.n683 0.00105952
R9451 Iout.n959 Iout.n958 0.00105952
R9452 Iout.n694 Iout.n693 0.00105952
R9453 Iout.n697 Iout.n696 0.00105952
R9454 Iout.n691 Iout.n689 0.00105952
R9455 Iout.n688 Iout.n686 0.00105952
R9456 Iout.n962 Iout.n15 0.00105952
R9457 Iout.n965 Iout.n964 0.00105952
R9458 Iout.n575 Iout.n574 0.00105952
R9459 Iout.n578 Iout.n577 0.00105952
R9460 Iout.n587 Iout.n115 0.00105952
R9461 Iout.n590 Iout.n589 0.00105952
R9462 Iout.n599 Iout.n109 0.00105952
R9463 Iout.n602 Iout.n601 0.00105952
R9464 Iout.n611 Iout.n103 0.00105952
R9465 Iout.n614 Iout.n613 0.00105952
R9466 Iout.n623 Iout.n97 0.00105952
R9467 Iout.n626 Iout.n625 0.00105952
R9468 Iout.n86 Iout.n84 0.00105952
R9469 Iout.n644 Iout.n643 0.00105952
R9470 Iout.n641 Iout.n88 0.00105952
R9471 Iout.n632 Iout.n631 0.00105952
R9472 Iout.n629 Iout.n94 0.00105952
R9473 Iout.n620 Iout.n619 0.00105952
R9474 Iout.n617 Iout.n100 0.00105952
R9475 Iout.n608 Iout.n607 0.00105952
R9476 Iout.n605 Iout.n106 0.00105952
R9477 Iout.n596 Iout.n595 0.00105952
R9478 Iout.n593 Iout.n112 0.00105952
R9479 Iout.n584 Iout.n583 0.00105952
R9480 Iout.n973 Iout.n971 0.00105952
R9481 Iout.n970 Iout.n968 0.00105952
R9482 Iout.n565 Iout.n564 0.00105952
R9483 Iout.n581 Iout.n118 0.00105952
R9484 Iout.n978 Iout.n977 0.00105952
R9485 Iout.n122 Iout.n121 0.00105952
R9486 Iout.n568 Iout.n124 0.00105952
R9487 Iout.n571 Iout.n570 0.00105952
R9488 Iout.n335 Iout.n334 0.00105952
R9489 Iout.n338 Iout.n337 0.00105952
R9490 Iout.n341 Iout.n340 0.00105952
R9491 Iout.n344 Iout.n343 0.00105952
R9492 Iout.n347 Iout.n346 0.00105952
R9493 Iout.n350 Iout.n349 0.00105952
R9494 Iout.n353 Iout.n352 0.00105952
R9495 Iout.n356 Iout.n355 0.00105952
R9496 Iout.n359 Iout.n358 0.00105952
R9497 Iout.n372 Iout.n371 0.00105952
R9498 Iout.n385 Iout.n383 0.00105952
R9499 Iout.n388 Iout.n387 0.00105952
R9500 Iout.n401 Iout.n399 0.00105952
R9501 Iout.n404 Iout.n403 0.00105952
R9502 Iout.n417 Iout.n415 0.00105952
R9503 Iout.n420 Iout.n419 0.00105952
R9504 Iout.n433 Iout.n431 0.00105952
R9505 Iout.n443 Iout.n442 0.00105952
R9506 Iout.n440 Iout.n439 0.00105952
R9507 Iout.n437 Iout.n435 0.00105952
R9508 Iout.n555 Iout.n553 0.00105952
R9509 Iout.n558 Iout.n556 0.00105952
R9510 Iout.n981 Iout.n10 0.00105952
R9511 Iout.n984 Iout.n983 0.00105952
R9512 Iout.n561 Iout.n560 0.00105952
R9513 Iout.n992 Iout.n990 0.00105952
R9514 Iout.n989 Iout.n987 0.00105952
R9515 Iout.n129 Iout.n128 0.00105952
R9516 Iout.n547 Iout.n131 0.00105952
R9517 Iout.n550 Iout.n549 0.00105952
R9518 Iout.n451 Iout.n450 0.00105952
R9519 Iout.n454 Iout.n453 0.00105952
R9520 Iout.n448 Iout.n446 0.00105952
R9521 Iout.n428 Iout.n427 0.00105952
R9522 Iout.n425 Iout.n423 0.00105952
R9523 Iout.n412 Iout.n411 0.00105952
R9524 Iout.n409 Iout.n407 0.00105952
R9525 Iout.n396 Iout.n395 0.00105952
R9526 Iout.n393 Iout.n391 0.00105952
R9527 Iout.n331 Iout.n330 0.00105952
R9528 Iout.n328 Iout.n327 0.00105952
R9529 Iout.n325 Iout.n324 0.00105952
R9530 Iout.n322 Iout.n321 0.00105952
R9531 Iout.n319 Iout.n318 0.00105952
R9532 Iout.n316 Iout.n315 0.00105952
R9533 Iout.n313 Iout.n312 0.00105952
R9534 Iout.n310 Iout.n309 0.00105952
R9535 Iout.n307 Iout.n306 0.00105952
R9536 Iout.n459 Iout.n457 0.00105952
R9537 Iout.n465 Iout.n464 0.00105952
R9538 Iout.n462 Iout.n461 0.00105952
R9539 Iout.n544 Iout.n543 0.00105952
R9540 Iout.n541 Iout.n137 0.00105952
R9541 Iout.n997 Iout.n996 0.00105952
R9542 Iout.n135 Iout.n134 0.00105952
R9543 Iout.n1000 Iout.n5 0.00105952
R9544 Iout.n1003 Iout.n1002 0.00105952
R9545 Iout.n538 Iout.n537 0.00105952
R9546 Iout.n535 Iout.n533 0.00105952
R9547 Iout.n532 Iout.n530 0.00105952
R9548 Iout.n468 Iout.n157 0.00105952
R9549 Iout.n471 Iout.n470 0.00105952
R9550 Iout.n474 Iout.n473 0.00105952
R9551 Iout.n264 Iout.n190 0.00105952
R9552 Iout.n267 Iout.n266 0.00105952
R9553 Iout.n276 Iout.n184 0.00105952
R9554 Iout.n279 Iout.n278 0.00105952
R9555 Iout.n288 Iout.n178 0.00105952
R9556 Iout.n291 Iout.n290 0.00105952
R9557 Iout.n300 Iout.n169 0.00105952
R9558 Iout.n173 Iout.n171 0.00105952
R9559 Iout.n297 Iout.n296 0.00105952
R9560 Iout.n294 Iout.n175 0.00105952
R9561 Iout.n285 Iout.n284 0.00105952
R9562 Iout.n282 Iout.n181 0.00105952
R9563 Iout.n273 Iout.n272 0.00105952
R9564 Iout.n270 Iout.n187 0.00105952
R9565 Iout.n261 Iout.n260 0.00105952
R9566 Iout.n479 Iout.n477 0.00105952
R9567 Iout.n485 Iout.n484 0.00105952
R9568 Iout.n482 Iout.n481 0.00105952
R9569 Iout.n527 Iout.n526 0.00105952
R9570 Iout.n524 Iout.n144 0.00105952
R9571 Iout.n142 Iout.n141 0.00105952
R9572 Iout.n1008 Iout.n1006 0.00105952
R9573 Iout.n1011 Iout.n1009 0.00105952
R9574 Iout.n1016 Iout.n1015 0.00105952
R9575 Iout.n148 Iout.n147 0.00105952
R9576 Iout.n518 Iout.n150 0.00105952
R9577 Iout.n521 Iout.n520 0.00105952
R9578 Iout.n493 Iout.n492 0.00105952
R9579 Iout.n496 Iout.n495 0.00105952
R9580 Iout.n490 Iout.n488 0.00105952
R9581 Iout.n254 Iout.n253 0.00105952
R9582 Iout.n257 Iout.n256 0.00105952
R9583 Iout.n251 Iout.n249 0.00105952
R9584 Iout.n248 Iout.n246 0.00105952
R9585 Iout.n245 Iout.n243 0.00105952
R9586 Iout.n242 Iout.n240 0.00105952
R9587 Iout.n239 Iout.n237 0.00105952
R9588 Iout.n236 Iout.n234 0.00105952
R9589 Iout.n233 Iout.n231 0.00105952
R9590 Iout.n228 Iout.n227 0.00105952
R9591 Iout.n225 Iout.n223 0.00105952
R9592 Iout.n221 Iout.n219 0.00105952
R9593 Iout.n217 Iout.n215 0.00105952
R9594 Iout.n213 Iout.n211 0.00105952
R9595 Iout.n209 Iout.n207 0.00105952
R9596 Iout.n205 Iout.n203 0.00105952
R9597 Iout.n201 Iout.n200 0.00105952
R9598 Iout.n198 Iout.n196 0.00105952
R9599 Iout.n194 Iout.n193 0.00105952
R9600 Iout.n501 Iout.n499 0.00105952
R9601 Iout.n505 Iout.n503 0.00105952
R9602 Iout.n508 Iout.n506 0.00105952
R9603 Iout.n515 Iout.n514 0.00105952
R9604 Iout.n512 Iout.n510 0.00105952
R9605 Iout.n1021 Iout.n1019 0.00105952
R9606 VPWR.n2773 VPWR.n2759 2618.82
R9607 VPWR.n2771 VPWR.n2765 2618.82
R9608 VPWR.n2789 VPWR.n2759 1916.47
R9609 VPWR.n2764 VPWR.n2763 1916.47
R9610 VPWR.n2763 VPWR.n2757 1916.47
R9611 VPWR.n2765 VPWR.n2758 1916.47
R9612 VPWR.n2788 VPWR.n2760 1912.94
R9613 VPWR.n2785 VPWR.n2779 1560
R9614 VPWR.n2786 VPWR.n2760 1408.24
R9615 VPWR.n2789 VPWR.n2788 1210.59
R9616 VPWR.n2787 VPWR.n2757 1210.59
R9617 VPWR.n2316 VPWR.t766 1005.7
R9618 VPWR.t986 VPWR.n453 1005.7
R9619 VPWR.t820 VPWR.n2146 1005.7
R9620 VPWR.n607 VPWR.t938 1005.7
R9621 VPWR.n2120 VPWR.t673 1005.7
R9622 VPWR.t774 VPWR.n645 1005.7
R9623 VPWR.t734 VPWR.n1950 1005.7
R9624 VPWR.n799 VPWR.t836 1005.7
R9625 VPWR.n1924 VPWR.t670 1005.7
R9626 VPWR.t845 VPWR.n837 1005.7
R9627 VPWR.n415 VPWR.t664 1005.7
R9628 VPWR.t946 VPWR.n1754 1005.7
R9629 VPWR.t932 VPWR.n2342 1005.7
R9630 VPWR.n991 VPWR.t804 1005.7
R9631 VPWR.t978 VPWR.n261 1005.7
R9632 VPWR.n1728 VPWR.t915 1005.7
R9633 VPWR.n2527 VPWR.t839 1005.7
R9634 VPWR.n1029 VPWR.t737 1005.7
R9635 VPWR.t1846 VPWR.n2245 938.953
R9636 VPWR.n2246 VPWR.t1442 938.953
R9637 VPWR.t1887 VPWR.n2255 938.953
R9638 VPWR.n2256 VPWR.t1464 938.953
R9639 VPWR.t1710 VPWR.n2265 938.953
R9640 VPWR.n2266 VPWR.t220 938.953
R9641 VPWR.t1628 VPWR.n2275 938.953
R9642 VPWR.n2276 VPWR.t509 938.953
R9643 VPWR.t1909 VPWR.n2285 938.953
R9644 VPWR.n2286 VPWR.t1070 938.953
R9645 VPWR.t82 VPWR.n2295 938.953
R9646 VPWR.n2296 VPWR.t1494 938.953
R9647 VPWR.t1600 VPWR.n2305 938.953
R9648 VPWR.n2306 VPWR.t1478 938.953
R9649 VPWR.t451 VPWR.n2315 938.953
R9650 VPWR.n510 VPWR.t1242 938.953
R9651 VPWR.n509 VPWR.t1400 938.953
R9652 VPWR.n505 VPWR.t30 938.953
R9653 VPWR.n501 VPWR.t1285 938.953
R9654 VPWR.n497 VPWR.t1526 938.953
R9655 VPWR.n493 VPWR.t1558 938.953
R9656 VPWR.n489 VPWR.t425 938.953
R9657 VPWR.n485 VPWR.t1861 938.953
R9658 VPWR.n481 VPWR.t236 938.953
R9659 VPWR.n477 VPWR.t314 938.953
R9660 VPWR.n473 VPWR.t116 938.953
R9661 VPWR.n469 VPWR.t565 938.953
R9662 VPWR.n465 VPWR.t1112 938.953
R9663 VPWR.n461 VPWR.t1084 938.953
R9664 VPWR.n457 VPWR.t471 938.953
R9665 VPWR.n2217 VPWR.t1019 938.953
R9666 VPWR.n2216 VPWR.t1683 938.953
R9667 VPWR.n2207 VPWR.t997 938.953
R9668 VPWR.n2206 VPWR.t584 938.953
R9669 VPWR.n2197 VPWR.t1254 938.953
R9670 VPWR.n2196 VPWR.t1520 938.953
R9671 VPWR.n2187 VPWR.t270 938.953
R9672 VPWR.n2186 VPWR.t1424 938.953
R9673 VPWR.n2177 VPWR.t1895 938.953
R9674 VPWR.n2176 VPWR.t304 938.953
R9675 VPWR.n2167 VPWR.t84 938.953
R9676 VPWR.n2166 VPWR.t423 938.953
R9677 VPWR.n2157 VPWR.t1612 938.953
R9678 VPWR.n2156 VPWR.t1646 938.953
R9679 VPWR.n2147 VPWR.t441 938.953
R9680 VPWR.t1037 VPWR.n550 938.953
R9681 VPWR.t1798 VPWR.n554 938.953
R9682 VPWR.t16 VPWR.n558 938.953
R9683 VPWR.t1918 VPWR.n562 938.953
R9684 VPWR.t1584 VPWR.n566 938.953
R9685 VPWR.t1808 VPWR.n570 938.953
R9686 VPWR.t431 VPWR.n574 938.953
R9687 VPWR.t497 VPWR.n578 938.953
R9688 VPWR.t242 VPWR.n582 938.953
R9689 VPWR.t320 VPWR.n586 938.953
R9690 VPWR.t108 VPWR.n590 938.953
R9691 VPWR.t256 VPWR.n594 938.953
R9692 VPWR.t1122 VPWR.n598 938.953
R9693 VPWR.t601 VPWR.n602 938.953
R9694 VPWR.t457 VPWR.n606 938.953
R9695 VPWR.t336 VPWR.n2049 938.953
R9696 VPWR.n2050 VPWR.t1693 938.953
R9697 VPWR.t1269 VPWR.n2059 938.953
R9698 VPWR.n2060 VPWR.t140 938.953
R9699 VPWR.t1592 VPWR.n2069 938.953
R9700 VPWR.n2070 VPWR.t284 938.953
R9701 VPWR.t539 VPWR.n2079 938.953
R9702 VPWR.n2080 VPWR.t519 938.953
R9703 VPWR.t1178 VPWR.n2089 938.953
R9704 VPWR.n2090 VPWR.t349 938.953
R9705 VPWR.t70 VPWR.n2099 938.953
R9706 VPWR.n2100 VPWR.t1108 938.953
R9707 VPWR.t1411 VPWR.n2109 938.953
R9708 VPWR.n2110 VPWR.t1480 938.953
R9709 VPWR.t1375 VPWR.n2119 938.953
R9710 VPWR.n702 VPWR.t1844 938.953
R9711 VPWR.n701 VPWR.t1440 938.953
R9712 VPWR.n697 VPWR.t1883 938.953
R9713 VPWR.n693 VPWR.t1462 938.953
R9714 VPWR.n689 VPWR.t1708 938.953
R9715 VPWR.n685 VPWR.t218 938.953
R9716 VPWR.n681 VPWR.t1626 938.953
R9717 VPWR.n677 VPWR.t1436 938.953
R9718 VPWR.n673 VPWR.t1907 938.953
R9719 VPWR.n669 VPWR.t1066 938.953
R9720 VPWR.n665 VPWR.t80 938.953
R9721 VPWR.n661 VPWR.t1490 938.953
R9722 VPWR.n657 VPWR.t1363 938.953
R9723 VPWR.n653 VPWR.t1476 938.953
R9724 VPWR.n649 VPWR.t449 938.953
R9725 VPWR.n2021 VPWR.t1850 938.953
R9726 VPWR.n2020 VPWR.t178 938.953
R9727 VPWR.n2011 VPWR.t56 938.953
R9728 VPWR.n2010 VPWR.t1291 938.953
R9729 VPWR.n2001 VPWR.t1695 938.953
R9730 VPWR.n2000 VPWR.t46 938.953
R9731 VPWR.n1991 VPWR.t1090 938.953
R9732 VPWR.n1990 VPWR.t515 938.953
R9733 VPWR.n1981 VPWR.t1168 938.953
R9734 VPWR.n1980 VPWR.t342 938.953
R9735 VPWR.n1971 VPWR.t74 938.953
R9736 VPWR.n1970 VPWR.t1614 938.953
R9737 VPWR.n1961 VPWR.t1606 938.953
R9738 VPWR.n1960 VPWR.t1074 938.953
R9739 VPWR.n1951 VPWR.t1367 938.953
R9740 VPWR.t1017 VPWR.n742 938.953
R9741 VPWR.t1681 VPWR.n746 938.953
R9742 VPWR.t995 VPWR.n750 938.953
R9743 VPWR.t582 VPWR.n754 938.953
R9744 VPWR.t1252 VPWR.n758 938.953
R9745 VPWR.t1518 VPWR.n762 938.953
R9746 VPWR.t266 VPWR.n766 938.953
R9747 VPWR.t1422 VPWR.n770 938.953
R9748 VPWR.t1893 VPWR.n774 938.953
R9749 VPWR.t302 VPWR.n778 938.953
R9750 VPWR.t100 VPWR.n782 938.953
R9751 VPWR.t421 VPWR.n786 938.953
R9752 VPWR.t1610 VPWR.n790 938.953
R9753 VPWR.t1644 VPWR.n794 938.953
R9754 VPWR.t437 VPWR.n798 938.953
R9755 VPWR.t338 VPWR.n1853 938.953
R9756 VPWR.n1854 VPWR.t1540 938.953
R9757 VPWR.t1271 VPWR.n1863 938.953
R9758 VPWR.n1864 VPWR.t142 938.953
R9759 VPWR.t1594 VPWR.n1873 938.953
R9760 VPWR.n1874 VPWR.t286 938.953
R9761 VPWR.t543 VPWR.n1883 938.953
R9762 VPWR.n1884 VPWR.t1387 938.953
R9763 VPWR.t1180 VPWR.n1893 938.953
R9764 VPWR.n1894 VPWR.t351 938.953
R9765 VPWR.t72 VPWR.n1903 938.953
R9766 VPWR.n1904 VPWR.t1110 938.953
R9767 VPWR.t1413 VPWR.n1913 938.953
R9768 VPWR.n1914 VPWR.t1482 938.953
R9769 VPWR.t1379 VPWR.n1923 938.953
R9770 VPWR.n894 VPWR.t595 938.953
R9771 VPWR.n893 VPWR.t1417 938.953
R9772 VPWR.n889 VPWR.t993 938.953
R9773 VPWR.n885 VPWR.t580 938.953
R9774 VPWR.n881 VPWR.t1250 938.953
R9775 VPWR.n877 VPWR.t1514 938.953
R9776 VPWR.n873 VPWR.t1458 938.953
R9777 VPWR.n869 VPWR.t1420 938.953
R9778 VPWR.n865 VPWR.t1889 938.953
R9779 VPWR.n861 VPWR.t300 938.953
R9780 VPWR.n857 VPWR.t96 938.953
R9781 VPWR.n853 VPWR.t419 938.953
R9782 VPWR.n849 VPWR.t1608 938.953
R9783 VPWR.n845 VPWR.t1232 938.953
R9784 VPWR.n841 VPWR.t433 938.953
R9785 VPWR.t1234 VPWR.n358 938.953
R9786 VPWR.t1542 VPWR.n362 938.953
R9787 VPWR.t1273 VPWR.n366 938.953
R9788 VPWR.t576 VPWR.n370 938.953
R9789 VPWR.t1596 VPWR.n374 938.953
R9790 VPWR.t1550 VPWR.n378 938.953
R9791 VPWR.t545 VPWR.n382 938.953
R9792 VPWR.t1389 VPWR.n386 938.953
R9793 VPWR.t1182 VPWR.n390 938.953
R9794 VPWR.t353 VPWR.n394 938.953
R9795 VPWR.t58 VPWR.n398 938.953
R9796 VPWR.t246 VPWR.n402 938.953
R9797 VPWR.t1415 VPWR.n406 938.953
R9798 VPWR.t1484 VPWR.n410 938.953
R9799 VPWR.t1381 VPWR.n414 938.953
R9800 VPWR.n1825 VPWR.t1035 938.953
R9801 VPWR.n1824 VPWR.t1796 938.953
R9802 VPWR.n1815 VPWR.t14 938.953
R9803 VPWR.n1814 VPWR.t1916 938.953
R9804 VPWR.n1805 VPWR.t1582 938.953
R9805 VPWR.n1804 VPWR.t1806 938.953
R9806 VPWR.n1795 VPWR.t429 938.953
R9807 VPWR.n1794 VPWR.t495 938.953
R9808 VPWR.n1785 VPWR.t240 938.953
R9809 VPWR.n1784 VPWR.t318 938.953
R9810 VPWR.n1775 VPWR.t106 938.953
R9811 VPWR.n1774 VPWR.t254 938.953
R9812 VPWR.n1765 VPWR.t1120 938.953
R9813 VPWR.n1764 VPWR.t599 938.953
R9814 VPWR.n1755 VPWR.t455 938.953
R9815 VPWR.n2413 VPWR.t1039 938.953
R9816 VPWR.n2412 VPWR.t1800 938.953
R9817 VPWR.n2403 VPWR.t20 938.953
R9818 VPWR.n2402 VPWR.t1920 938.953
R9819 VPWR.n2393 VPWR.t1586 938.953
R9820 VPWR.n2392 VPWR.t1810 938.953
R9821 VPWR.n2383 VPWR.t1104 938.953
R9822 VPWR.n2382 VPWR.t499 938.953
R9823 VPWR.n2373 VPWR.t244 938.953
R9824 VPWR.n2372 VPWR.t185 938.953
R9825 VPWR.n2363 VPWR.t110 938.953
R9826 VPWR.n2362 VPWR.t260 938.953
R9827 VPWR.n2353 VPWR.t1124 938.953
R9828 VPWR.n2352 VPWR.t1140 938.953
R9829 VPWR.n2343 VPWR.t463 938.953
R9830 VPWR.t1025 VPWR.n934 938.953
R9831 VPWR.t1407 VPWR.n938 938.953
R9832 VPWR.t384 VPWR.n942 938.953
R9833 VPWR.t553 VPWR.n946 938.953
R9834 VPWR.t1704 VPWR.n950 938.953
R9835 VPWR.t212 VPWR.n954 938.953
R9836 VPWR.t1622 VPWR.n958 938.953
R9837 VPWR.t1432 VPWR.n962 938.953
R9838 VPWR.t1901 VPWR.n966 938.953
R9839 VPWR.t1058 VPWR.n970 938.953
R9840 VPWR.t90 VPWR.n974 938.953
R9841 VPWR.t559 VPWR.n978 938.953
R9842 VPWR.t1359 VPWR.n982 938.953
R9843 VPWR.t1652 VPWR.n986 938.953
R9844 VPWR.t445 VPWR.n990 938.953
R9845 VPWR.n318 VPWR.t1244 938.953
R9846 VPWR.n317 VPWR.t1402 938.953
R9847 VPWR.n313 VPWR.t12 938.953
R9848 VPWR.n309 VPWR.t1287 938.953
R9849 VPWR.n305 VPWR.t1528 938.953
R9850 VPWR.n301 VPWR.t1560 938.953
R9851 VPWR.n297 VPWR.t427 938.953
R9852 VPWR.n293 VPWR.t1863 938.953
R9853 VPWR.n289 VPWR.t238 938.953
R9854 VPWR.n285 VPWR.t316 938.953
R9855 VPWR.n281 VPWR.t118 938.953
R9856 VPWR.n277 VPWR.t567 938.953
R9857 VPWR.n273 VPWR.t1114 938.953
R9858 VPWR.n269 VPWR.t1086 938.953
R9859 VPWR.n265 VPWR.t473 938.953
R9860 VPWR.t613 VPWR.n1451 938.953
R9861 VPWR.t707 VPWR.n1457 938.953
R9862 VPWR.n1458 VPWR.t747 938.953
R9863 VPWR.t967 VPWR.n1470 938.953
R9864 VPWR.n1471 VPWR.t610 938.953
R9865 VPWR.t752 VPWR.n1484 938.953
R9866 VPWR.n1485 VPWR.t865 938.953
R9867 VPWR.t886 VPWR.n1498 938.953
R9868 VPWR.n1499 VPWR.t641 938.953
R9869 VPWR.n1514 VPWR.t771 938.953
R9870 VPWR.n1513 VPWR.t897 938.953
R9871 VPWR.n1697 VPWR.t889 938.953
R9872 VPWR.n1696 VPWR.t667 938.953
R9873 VPWR.n1685 VPWR.t809 938.953
R9874 VPWR.t923 VPWR.n1727 938.953
R9875 VPWR.t929 VPWR.n2442 938.953
R9876 VPWR.n2443 VPWR.t651 938.953
R9877 VPWR.t689 VPWR.n2454 938.953
R9878 VPWR.n2455 VPWR.t907 938.953
R9879 VPWR.t926 VPWR.n2466 938.953
R9880 VPWR.n2467 VPWR.t699 938.953
R9881 VPWR.t795 VPWR.n2478 938.953
R9882 VPWR.n2479 VPWR.t831 938.953
R9883 VPWR.t972 VPWR.n2490 938.953
R9884 VPWR.n2491 VPWR.t715 938.953
R9885 VPWR.t850 VPWR.n2502 938.953
R9886 VPWR.n2503 VPWR.t881 938.953
R9887 VPWR.t621 VPWR.n2514 938.953
R9888 VPWR.n2515 VPWR.t760 938.953
R9889 VPWR.t870 VPWR.n2526 938.953
R9890 VPWR.n1165 VPWR.t801 938.953
R9891 VPWR.n1164 VPWR.t918 938.953
R9892 VPWR.n1160 VPWR.t954 938.953
R9893 VPWR.n1156 VPWR.t790 938.953
R9894 VPWR.n1152 VPWR.t798 938.953
R9895 VPWR.n1148 VPWR.t962 938.953
R9896 VPWR.n1144 VPWR.t681 938.953
R9897 VPWR.n1140 VPWR.t723 938.953
R9898 VPWR.n1136 VPWR.t855 938.953
R9899 VPWR.n1132 VPWR.t991 938.953
R9900 VPWR.n1128 VPWR.t731 938.953
R9901 VPWR.n1124 VPWR.t763 938.953
R9902 VPWR.n1120 VPWR.t878 938.953
R9903 VPWR.n1676 VPWR.t631 938.953
R9904 VPWR.n1675 VPWR.t742 938.953
R9905 VPWR.n1247 VPWR.t348 877.144
R9906 VPWR.n2659 VPWR.t1755 877.144
R9907 VPWR.n2779 VPWR.n2758 857.648
R9908 VPWR.n1116 VPWR.t660 745.917
R9909 VPWR.n99 VPWR.t783 745.917
R9910 VPWR.n258 VPWR.t1221 745.917
R9911 VPWR.n68 VPWR.t851 745.917
R9912 VPWR.n314 VPWR.t1245 745.917
R9913 VPWR.n98 VPWR.t930 745.917
R9914 VPWR.n931 VPWR.t1205 745.917
R9915 VPWR.n324 VPWR.t1215 745.917
R9916 VPWR.n325 VPWR.t1040 745.917
R9917 VPWR.n286 VPWR.t1864 745.917
R9918 VPWR.n75 VPWR.t832 745.917
R9919 VPWR.n939 VPWR.t1408 745.917
R9920 VPWR.n337 VPWR.t1105 745.917
R9921 VPWR.n290 VPWR.t428 745.917
R9922 VPWR.n80 VPWR.t796 745.917
R9923 VPWR.n900 VPWR.t1219 745.917
R9924 VPWR.n901 VPWR.t1036 745.917
R9925 VPWR.n904 VPWR.t1797 745.917
R9926 VPWR.n355 VPWR.t1225 745.917
R9927 VPWR.n359 VPWR.t1235 745.917
R9928 VPWR.n363 VPWR.t1543 745.917
R9929 VPWR.n333 VPWR.t1587 745.917
R9930 VPWR.n298 VPWR.t1529 745.917
R9931 VPWR.n86 VPWR.t927 745.917
R9932 VPWR.n905 VPWR.t15 745.917
R9933 VPWR.n371 VPWR.t577 745.917
R9934 VPWR.n332 VPWR.t1921 745.917
R9935 VPWR.n302 VPWR.t1288 745.917
R9936 VPWR.n87 VPWR.t908 745.917
R9937 VPWR.n449 VPWR.t1201 745.917
R9938 VPWR.n448 VPWR.t1847 745.917
R9939 VPWR.n445 VPWR.t1443 745.917
R9940 VPWR.n444 VPWR.t1888 745.917
R9941 VPWR.n440 VPWR.t1711 745.917
R9942 VPWR.n437 VPWR.t221 745.917
R9943 VPWR.n436 VPWR.t1629 745.917
R9944 VPWR.n433 VPWR.t510 745.917
R9945 VPWR.n432 VPWR.t1910 745.917
R9946 VPWR.n429 VPWR.t1071 745.917
R9947 VPWR.n428 VPWR.t83 745.917
R9948 VPWR.n425 VPWR.t1495 745.917
R9949 VPWR.n424 VPWR.t1601 745.917
R9950 VPWR.n421 VPWR.t1479 745.917
R9951 VPWR.n420 VPWR.t452 745.917
R9952 VPWR.n441 VPWR.t1465 745.917
R9953 VPWR.n450 VPWR.t1223 745.917
R9954 VPWR.n506 VPWR.t1243 745.917
R9955 VPWR.n502 VPWR.t1401 745.917
R9956 VPWR.n498 VPWR.t31 745.917
R9957 VPWR.n490 VPWR.t1527 745.917
R9958 VPWR.n486 VPWR.t1559 745.917
R9959 VPWR.n482 VPWR.t426 745.917
R9960 VPWR.n478 VPWR.t1862 745.917
R9961 VPWR.n474 VPWR.t237 745.917
R9962 VPWR.n470 VPWR.t315 745.917
R9963 VPWR.n466 VPWR.t117 745.917
R9964 VPWR.n462 VPWR.t566 745.917
R9965 VPWR.n458 VPWR.t1113 745.917
R9966 VPWR.n454 VPWR.t1085 745.917
R9967 VPWR.n451 VPWR.t472 745.917
R9968 VPWR.n494 VPWR.t1286 745.917
R9969 VPWR.n516 VPWR.t1207 745.917
R9970 VPWR.n517 VPWR.t1020 745.917
R9971 VPWR.n520 VPWR.t1684 745.917
R9972 VPWR.n521 VPWR.t998 745.917
R9973 VPWR.n525 VPWR.t1255 745.917
R9974 VPWR.n528 VPWR.t1521 745.917
R9975 VPWR.n529 VPWR.t271 745.917
R9976 VPWR.n532 VPWR.t1425 745.917
R9977 VPWR.n533 VPWR.t1896 745.917
R9978 VPWR.n536 VPWR.t305 745.917
R9979 VPWR.n537 VPWR.t85 745.917
R9980 VPWR.n540 VPWR.t424 745.917
R9981 VPWR.n541 VPWR.t1613 745.917
R9982 VPWR.n544 VPWR.t1647 745.917
R9983 VPWR.n545 VPWR.t442 745.917
R9984 VPWR.n524 VPWR.t585 745.917
R9985 VPWR.n547 VPWR.t1217 745.917
R9986 VPWR.n551 VPWR.t1038 745.917
R9987 VPWR.n555 VPWR.t1799 745.917
R9988 VPWR.n559 VPWR.t17 745.917
R9989 VPWR.n567 VPWR.t1585 745.917
R9990 VPWR.n571 VPWR.t1809 745.917
R9991 VPWR.n575 VPWR.t432 745.917
R9992 VPWR.n579 VPWR.t498 745.917
R9993 VPWR.n583 VPWR.t243 745.917
R9994 VPWR.n587 VPWR.t321 745.917
R9995 VPWR.n591 VPWR.t109 745.917
R9996 VPWR.n595 VPWR.t257 745.917
R9997 VPWR.n599 VPWR.t1123 745.917
R9998 VPWR.n603 VPWR.t602 745.917
R9999 VPWR.n546 VPWR.t458 745.917
R10000 VPWR.n563 VPWR.t1919 745.917
R10001 VPWR.n641 VPWR.t1229 745.917
R10002 VPWR.n640 VPWR.t337 745.917
R10003 VPWR.n637 VPWR.t1694 745.917
R10004 VPWR.n636 VPWR.t1270 745.917
R10005 VPWR.n632 VPWR.t1593 745.917
R10006 VPWR.n629 VPWR.t285 745.917
R10007 VPWR.n628 VPWR.t540 745.917
R10008 VPWR.n625 VPWR.t520 745.917
R10009 VPWR.n624 VPWR.t1179 745.917
R10010 VPWR.n621 VPWR.t350 745.917
R10011 VPWR.n620 VPWR.t71 745.917
R10012 VPWR.n617 VPWR.t1109 745.917
R10013 VPWR.n616 VPWR.t1412 745.917
R10014 VPWR.n613 VPWR.t1481 745.917
R10015 VPWR.n612 VPWR.t1376 745.917
R10016 VPWR.n633 VPWR.t141 745.917
R10017 VPWR.n642 VPWR.t1203 745.917
R10018 VPWR.n698 VPWR.t1845 745.917
R10019 VPWR.n694 VPWR.t1441 745.917
R10020 VPWR.n690 VPWR.t1884 745.917
R10021 VPWR.n682 VPWR.t1709 745.917
R10022 VPWR.n678 VPWR.t219 745.917
R10023 VPWR.n674 VPWR.t1627 745.917
R10024 VPWR.n670 VPWR.t1437 745.917
R10025 VPWR.n666 VPWR.t1908 745.917
R10026 VPWR.n662 VPWR.t1067 745.917
R10027 VPWR.n658 VPWR.t81 745.917
R10028 VPWR.n654 VPWR.t1491 745.917
R10029 VPWR.n650 VPWR.t1364 745.917
R10030 VPWR.n646 VPWR.t1477 745.917
R10031 VPWR.n643 VPWR.t450 745.917
R10032 VPWR.n686 VPWR.t1463 745.917
R10033 VPWR.n708 VPWR.t1199 745.917
R10034 VPWR.n709 VPWR.t1851 745.917
R10035 VPWR.n712 VPWR.t179 745.917
R10036 VPWR.n713 VPWR.t57 745.917
R10037 VPWR.n717 VPWR.t1696 745.917
R10038 VPWR.n720 VPWR.t47 745.917
R10039 VPWR.n721 VPWR.t1091 745.917
R10040 VPWR.n724 VPWR.t516 745.917
R10041 VPWR.n725 VPWR.t1169 745.917
R10042 VPWR.n728 VPWR.t343 745.917
R10043 VPWR.n729 VPWR.t75 745.917
R10044 VPWR.n732 VPWR.t1615 745.917
R10045 VPWR.n733 VPWR.t1607 745.917
R10046 VPWR.n736 VPWR.t1075 745.917
R10047 VPWR.n737 VPWR.t1368 745.917
R10048 VPWR.n716 VPWR.t1292 745.917
R10049 VPWR.n739 VPWR.t1209 745.917
R10050 VPWR.n743 VPWR.t1018 745.917
R10051 VPWR.n747 VPWR.t1682 745.917
R10052 VPWR.n751 VPWR.t996 745.917
R10053 VPWR.n759 VPWR.t1253 745.917
R10054 VPWR.n763 VPWR.t1519 745.917
R10055 VPWR.n767 VPWR.t267 745.917
R10056 VPWR.n771 VPWR.t1423 745.917
R10057 VPWR.n775 VPWR.t1894 745.917
R10058 VPWR.n779 VPWR.t303 745.917
R10059 VPWR.n783 VPWR.t101 745.917
R10060 VPWR.n787 VPWR.t422 745.917
R10061 VPWR.n791 VPWR.t1611 745.917
R10062 VPWR.n795 VPWR.t1645 745.917
R10063 VPWR.n738 VPWR.t438 745.917
R10064 VPWR.n755 VPWR.t583 745.917
R10065 VPWR.n833 VPWR.t1227 745.917
R10066 VPWR.n832 VPWR.t339 745.917
R10067 VPWR.n829 VPWR.t1541 745.917
R10068 VPWR.n828 VPWR.t1272 745.917
R10069 VPWR.n824 VPWR.t1595 745.917
R10070 VPWR.n821 VPWR.t287 745.917
R10071 VPWR.n820 VPWR.t544 745.917
R10072 VPWR.n817 VPWR.t1388 745.917
R10073 VPWR.n816 VPWR.t1181 745.917
R10074 VPWR.n813 VPWR.t352 745.917
R10075 VPWR.n812 VPWR.t73 745.917
R10076 VPWR.n809 VPWR.t1111 745.917
R10077 VPWR.n808 VPWR.t1414 745.917
R10078 VPWR.n805 VPWR.t1483 745.917
R10079 VPWR.n804 VPWR.t1380 745.917
R10080 VPWR.n825 VPWR.t143 745.917
R10081 VPWR.n834 VPWR.t1213 745.917
R10082 VPWR.n890 VPWR.t596 745.917
R10083 VPWR.n886 VPWR.t1418 745.917
R10084 VPWR.n882 VPWR.t994 745.917
R10085 VPWR.n874 VPWR.t1251 745.917
R10086 VPWR.n870 VPWR.t1515 745.917
R10087 VPWR.n866 VPWR.t1459 745.917
R10088 VPWR.n862 VPWR.t1421 745.917
R10089 VPWR.n858 VPWR.t1890 745.917
R10090 VPWR.n854 VPWR.t301 745.917
R10091 VPWR.n850 VPWR.t97 745.917
R10092 VPWR.n846 VPWR.t420 745.917
R10093 VPWR.n842 VPWR.t1609 745.917
R10094 VPWR.n838 VPWR.t1233 745.917
R10095 VPWR.n835 VPWR.t434 745.917
R10096 VPWR.n878 VPWR.t581 745.917
R10097 VPWR.n908 VPWR.t1917 745.917
R10098 VPWR.n947 VPWR.t554 745.917
R10099 VPWR.n1149 VPWR.t791 745.917
R10100 VPWR.n367 VPWR.t1274 745.917
R10101 VPWR.n329 VPWR.t21 745.917
R10102 VPWR.n306 VPWR.t13 745.917
R10103 VPWR.n92 VPWR.t690 745.917
R10104 VPWR.n943 VPWR.t385 745.917
R10105 VPWR.n1153 VPWR.t955 745.917
R10106 VPWR.n909 VPWR.t1583 745.917
R10107 VPWR.n951 VPWR.t1705 745.917
R10108 VPWR.n1145 VPWR.t799 745.917
R10109 VPWR.n375 VPWR.t1597 745.917
R10110 VPWR.n383 VPWR.t546 745.917
R10111 VPWR.n387 VPWR.t1390 745.917
R10112 VPWR.n391 VPWR.t1183 745.917
R10113 VPWR.n395 VPWR.t354 745.917
R10114 VPWR.n399 VPWR.t59 745.917
R10115 VPWR.n403 VPWR.t247 745.917
R10116 VPWR.n407 VPWR.t1416 745.917
R10117 VPWR.n411 VPWR.t1485 745.917
R10118 VPWR.n354 VPWR.t1382 745.917
R10119 VPWR.n379 VPWR.t1551 745.917
R10120 VPWR.n336 VPWR.t1811 745.917
R10121 VPWR.n294 VPWR.t1561 745.917
R10122 VPWR.n81 VPWR.t700 745.917
R10123 VPWR.n955 VPWR.t213 745.917
R10124 VPWR.n1141 VPWR.t963 745.917
R10125 VPWR.n912 VPWR.t1807 745.917
R10126 VPWR.n916 VPWR.t496 745.917
R10127 VPWR.n917 VPWR.t241 745.917
R10128 VPWR.n920 VPWR.t319 745.917
R10129 VPWR.n921 VPWR.t107 745.917
R10130 VPWR.n924 VPWR.t255 745.917
R10131 VPWR.n925 VPWR.t1121 745.917
R10132 VPWR.n928 VPWR.t600 745.917
R10133 VPWR.n929 VPWR.t456 745.917
R10134 VPWR.n913 VPWR.t430 745.917
R10135 VPWR.n959 VPWR.t1623 745.917
R10136 VPWR.n1137 VPWR.t682 745.917
R10137 VPWR.n328 VPWR.t1801 745.917
R10138 VPWR.n310 VPWR.t1403 745.917
R10139 VPWR.n93 VPWR.t652 745.917
R10140 VPWR.n1157 VPWR.t919 745.917
R10141 VPWR.n963 VPWR.t1433 745.917
R10142 VPWR.n1133 VPWR.t724 745.917
R10143 VPWR.n340 VPWR.t500 745.917
R10144 VPWR.n344 VPWR.t186 745.917
R10145 VPWR.n345 VPWR.t111 745.917
R10146 VPWR.n348 VPWR.t261 745.917
R10147 VPWR.n349 VPWR.t1125 745.917
R10148 VPWR.n352 VPWR.t1141 745.917
R10149 VPWR.n353 VPWR.t464 745.917
R10150 VPWR.n341 VPWR.t245 745.917
R10151 VPWR.n282 VPWR.t239 745.917
R10152 VPWR.n74 VPWR.t973 745.917
R10153 VPWR.n1129 VPWR.t856 745.917
R10154 VPWR.n967 VPWR.t1902 745.917
R10155 VPWR.n971 VPWR.t1059 745.917
R10156 VPWR.n975 VPWR.t91 745.917
R10157 VPWR.n979 VPWR.t560 745.917
R10158 VPWR.n983 VPWR.t1360 745.917
R10159 VPWR.n987 VPWR.t1653 745.917
R10160 VPWR.n930 VPWR.t446 745.917
R10161 VPWR.n935 VPWR.t1026 745.917
R10162 VPWR.n1161 VPWR.t802 745.917
R10163 VPWR.n278 VPWR.t317 745.917
R10164 VPWR.n69 VPWR.t716 745.917
R10165 VPWR.n1125 VPWR.t992 745.917
R10166 VPWR.n1121 VPWR.t732 745.917
R10167 VPWR.n274 VPWR.t119 745.917
R10168 VPWR.n270 VPWR.t568 745.917
R10169 VPWR.n262 VPWR.t1087 745.917
R10170 VPWR.n259 VPWR.t474 745.917
R10171 VPWR.n266 VPWR.t1115 745.917
R10172 VPWR.n1026 VPWR.t879 745.917
R10173 VPWR.n1117 VPWR.t764 745.917
R10174 VPWR.n63 VPWR.t882 745.917
R10175 VPWR.n62 VPWR.t622 745.917
R10176 VPWR.n57 VPWR.t761 745.917
R10177 VPWR.n56 VPWR.t871 745.917
R10178 VPWR.n1027 VPWR.t632 745.917
R10179 VPWR.n1028 VPWR.t743 745.917
R10180 VPWR.n2792 VPWR.n2757 702.354
R10181 VPWR.n2792 VPWR.n2758 702.354
R10182 VPWR.n2790 VPWR.n2789 702.354
R10183 VPWR.n2790 VPWR.n2757 702.354
R10184 VPWR.n2773 VPWR.n2764 702.354
R10185 VPWR.n2786 VPWR.n2785 702.354
R10186 VPWR.n2771 VPWR.n2764 702.354
R10187 VPWR.n2751 VPWR.t400 651.634
R10188 VPWR.n2767 VPWR.t1211 651.505
R10189 VPWR.n2761 VPWR.t1911 651.505
R10190 VPWR.n2798 VPWR.t1860 651.431
R10191 VPWR.n1447 VPWR.t826 648.04
R10192 VPWR.n1415 VPWR.t772 648.04
R10193 VPWR.n1435 VPWR.t968 648.04
R10194 VPWR.n1439 VPWR.t748 648.04
R10195 VPWR.n1431 VPWR.t611 648.04
R10196 VPWR.n1427 VPWR.t753 648.04
R10197 VPWR.n1423 VPWR.t866 648.04
R10198 VPWR.n1443 VPWR.t708 648.04
R10199 VPWR.n1419 VPWR.t887 648.04
R10200 VPWR.n1411 VPWR.t642 648.04
R10201 VPWR.n1454 VPWR.t614 648.04
R10202 VPWR.n1016 VPWR.t898 648.04
R10203 VPWR.n1683 VPWR.t668 648.04
R10204 VPWR.n1003 VPWR.t810 648.04
R10205 VPWR.n999 VPWR.t924 648.04
R10206 VPWR.n1020 VPWR.t890 648.04
R10207 VPWR.n1028 VPWR.t738 646.071
R10208 VPWR.n1116 VPWR.t655 646.071
R10209 VPWR.n1027 VPWR.t627 646.071
R10210 VPWR.n56 VPWR.t840 646.071
R10211 VPWR.n62 VPWR.t617 646.071
R10212 VPWR.n99 VPWR.t778 646.071
R10213 VPWR.n1021 VPWR.t175 646.071
R10214 VPWR.n1448 VPWR.t1849 646.071
R10215 VPWR.n266 VPWR.t1651 646.071
R10216 VPWR.n258 VPWR.t1024 646.071
R10217 VPWR.n274 VPWR.t263 646.071
R10218 VPWR.n68 VPWR.t843 646.071
R10219 VPWR.n1416 VPWR.t79 646.071
R10220 VPWR.n314 VPWR.t1795 646.071
R10221 VPWR.n98 VPWR.t635 646.071
R10222 VPWR.n935 VPWR.t1439 646.071
R10223 VPWR.n931 VPWR.t1237 646.071
R10224 VPWR.n967 VPWR.t1069 646.071
R10225 VPWR.n341 VPWR.t194 646.071
R10226 VPWR.n324 VPWR.t1032 646.071
R10227 VPWR.n325 VPWR.t1537 646.071
R10228 VPWR.n340 VPWR.t1904 646.071
R10229 VPWR.n286 VPWR.t1892 646.071
R10230 VPWR.n75 VPWR.t829 646.071
R10231 VPWR.n939 VPWR.t1886 646.071
R10232 VPWR.n337 VPWR.t506 646.071
R10233 VPWR.n290 VPWR.t1868 646.071
R10234 VPWR.n80 VPWR.t813 646.071
R10235 VPWR.n913 VPWR.t502 646.071
R10236 VPWR.n900 VPWR.t1028 646.071
R10237 VPWR.n901 VPWR.t1803 646.071
R10238 VPWR.n904 VPWR.t25 646.071
R10239 VPWR.n912 VPWR.t265 646.071
R10240 VPWR.n379 VPWR.t1107 646.071
R10241 VPWR.n355 VPWR.t594 646.071
R10242 VPWR.n359 VPWR.t1549 646.071
R10243 VPWR.n363 VPWR.t29 646.071
R10244 VPWR.n375 VPWR.t1817 646.071
R10245 VPWR.n333 VPWR.t215 646.071
R10246 VPWR.n298 VPWR.t1517 646.071
R10247 VPWR.n86 VPWR.t942 646.071
R10248 VPWR.n905 VPWR.t1294 646.071
R10249 VPWR.n371 VPWR.t1525 646.071
R10250 VPWR.n332 VPWR.t1337 646.071
R10251 VPWR.n302 VPWR.t1581 646.071
R10252 VPWR.n87 VPWR.t903 646.071
R10253 VPWR.n441 VPWR.t1715 646.071
R10254 VPWR.n449 VPWR.t1241 646.071
R10255 VPWR.n448 VPWR.t177 646.071
R10256 VPWR.n445 VPWR.t39 646.071
R10257 VPWR.n444 VPWR.t1925 646.071
R10258 VPWR.n440 VPWR.t1555 646.071
R10259 VPWR.n437 VPWR.t1386 646.071
R10260 VPWR.n436 VPWR.t514 646.071
R10261 VPWR.n433 VPWR.t233 646.071
R10262 VPWR.n432 VPWR.t291 646.071
R10263 VPWR.n429 VPWR.t63 646.071
R10264 VPWR.n428 VPWR.t1499 646.071
R10265 VPWR.n425 VPWR.t1605 646.071
R10266 VPWR.n424 VPWR.t1083 646.071
R10267 VPWR.n421 VPWR.t1384 646.071
R10268 VPWR.n420 VPWR.t767 646.071
R10269 VPWR.n494 VPWR.t1579 646.071
R10270 VPWR.n450 VPWR.t1022 646.071
R10271 VPWR.n506 VPWR.t1793 646.071
R10272 VPWR.n502 VPWR.t19 646.071
R10273 VPWR.n498 VPWR.t1467 646.071
R10274 VPWR.n490 VPWR.t1513 646.071
R10275 VPWR.n486 VPWR.t1455 646.071
R10276 VPWR.n482 VPWR.t1866 646.071
R10277 VPWR.n478 VPWR.t1843 646.071
R10278 VPWR.n474 VPWR.t323 646.071
R10279 VPWR.n470 VPWR.t95 646.071
R10280 VPWR.n466 VPWR.t259 646.071
R10281 VPWR.n462 VPWR.t1117 646.071
R10282 VPWR.n458 VPWR.t1649 646.071
R10283 VPWR.n454 VPWR.t468 646.071
R10284 VPWR.n451 VPWR.t987 646.071
R10285 VPWR.n524 VPWR.t1703 646.071
R10286 VPWR.n516 VPWR.t335 646.071
R10287 VPWR.n517 VPWR.t1690 646.071
R10288 VPWR.n520 VPWR.t1882 646.071
R10289 VPWR.n521 VPWR.t1284 646.071
R10290 VPWR.n525 VPWR.t281 646.071
R10291 VPWR.n528 VPWR.t1095 646.071
R10292 VPWR.n529 VPWR.t1431 646.071
R10293 VPWR.n532 VPWR.t1175 646.071
R10294 VPWR.n533 VPWR.t1065 646.071
R10295 VPWR.n536 VPWR.t67 646.071
R10296 VPWR.n537 VPWR.t1489 646.071
R10297 VPWR.n540 VPWR.t1358 646.071
R10298 VPWR.n541 VPWR.t1659 646.071
R10299 VPWR.n544 VPWR.t1372 646.071
R10300 VPWR.n545 VPWR.t821 646.071
R10301 VPWR.n563 VPWR.t1591 646.071
R10302 VPWR.n547 VPWR.t1030 646.071
R10303 VPWR.n551 VPWR.t1535 646.071
R10304 VPWR.n555 VPWR.t41 646.071
R10305 VPWR.n559 VPWR.t1296 646.071
R10306 VPWR.n567 VPWR.t211 646.071
R10307 VPWR.n571 VPWR.t269 646.071
R10308 VPWR.n575 VPWR.t504 646.071
R10309 VPWR.n579 VPWR.t1900 646.071
R10310 VPWR.n583 VPWR.t192 646.071
R10311 VPWR.n587 VPWR.t89 646.071
R10312 VPWR.n591 VPWR.t1507 646.071
R10313 VPWR.n595 VPWR.t171 646.071
R10314 VPWR.n599 VPWR.t1473 646.071
R10315 VPWR.n603 VPWR.t440 646.071
R10316 VPWR.n546 VPWR.t939 646.071
R10317 VPWR.n633 VPWR.t1599 646.071
R10318 VPWR.n641 VPWR.t480 646.071
R10319 VPWR.n640 VPWR.t1545 646.071
R10320 VPWR.n637 VPWR.t1276 646.071
R10321 VPWR.n636 VPWR.t548 646.071
R10322 VPWR.n632 VPWR.t1813 646.071
R10323 VPWR.n629 VPWR.t1101 646.071
R10324 VPWR.n628 VPWR.t1392 646.071
R10325 VPWR.n625 VPWR.t371 646.071
R10326 VPWR.n624 VPWR.t356 646.071
R10327 VPWR.n621 VPWR.t113 646.071
R10328 VPWR.n620 VPWR.t249 646.071
R10329 VPWR.n617 VPWR.t1343 646.071
R10330 VPWR.n616 VPWR.t1143 646.071
R10331 VPWR.n613 VPWR.t460 646.071
R10332 VPWR.n612 VPWR.t674 646.071
R10333 VPWR.n686 VPWR.t1713 646.071
R10334 VPWR.n642 VPWR.t1239 646.071
R10335 VPWR.n698 VPWR.t1445 646.071
R10336 VPWR.n694 VPWR.t37 646.071
R10337 VPWR.n690 VPWR.t1923 646.071
R10338 VPWR.n682 VPWR.t1553 646.071
R10339 VPWR.n678 VPWR.t542 646.071
R10340 VPWR.n674 VPWR.t512 646.071
R10341 VPWR.n670 VPWR.t231 646.071
R10342 VPWR.n666 VPWR.t289 646.071
R10343 VPWR.n662 VPWR.t61 646.071
R10344 VPWR.n658 VPWR.t1497 646.071
R10345 VPWR.n654 VPWR.t1603 646.071
R10346 VPWR.n650 VPWR.t1081 646.071
R10347 VPWR.n646 VPWR.t1378 646.071
R10348 VPWR.n643 VPWR.t775 646.071
R10349 VPWR.n716 VPWR.t1698 646.071
R10350 VPWR.n708 VPWR.t1034 646.071
R10351 VPWR.n709 VPWR.t1692 646.071
R10352 VPWR.n712 VPWR.t1268 646.071
R10353 VPWR.n713 VPWR.t1057 646.071
R10354 VPWR.n717 VPWR.t1557 646.071
R10355 VPWR.n720 VPWR.t165 646.071
R10356 VPWR.n721 VPWR.t518 646.071
R10357 VPWR.n724 VPWR.t235 646.071
R10358 VPWR.n725 VPWR.t345 646.071
R10359 VPWR.n728 VPWR.t115 646.071
R10360 VPWR.n729 VPWR.t1617 646.071
R10361 VPWR.n732 VPWR.t1410 646.071
R10362 VPWR.n733 VPWR.t598 646.071
R10363 VPWR.n736 VPWR.t494 646.071
R10364 VPWR.n737 VPWR.t735 646.071
R10365 VPWR.n755 VPWR.t1701 646.071
R10366 VPWR.n739 VPWR.t333 646.071
R10367 VPWR.n743 VPWR.t1688 646.071
R10368 VPWR.n747 VPWR.t1880 646.071
R10369 VPWR.n751 VPWR.t1282 646.071
R10370 VPWR.n759 VPWR.t279 646.071
R10371 VPWR.n763 VPWR.t1093 646.071
R10372 VPWR.n767 VPWR.t1429 646.071
R10373 VPWR.n771 VPWR.t1173 646.071
R10374 VPWR.n775 VPWR.t1063 646.071
R10375 VPWR.n779 VPWR.t65 646.071
R10376 VPWR.n783 VPWR.t564 646.071
R10377 VPWR.n787 VPWR.t1356 646.071
R10378 VPWR.n791 VPWR.t1657 646.071
R10379 VPWR.n795 VPWR.t1370 646.071
R10380 VPWR.n738 VPWR.t837 646.071
R10381 VPWR.n825 VPWR.t1523 646.071
R10382 VPWR.n833 VPWR.t592 646.071
R10383 VPWR.n832 VPWR.t1547 646.071
R10384 VPWR.n829 VPWR.t27 646.071
R10385 VPWR.n828 VPWR.t550 646.071
R10386 VPWR.n824 VPWR.t1815 646.071
R10387 VPWR.n821 VPWR.t1103 646.071
R10388 VPWR.n820 VPWR.t1394 646.071
R10389 VPWR.n817 VPWR.t373 646.071
R10390 VPWR.n816 VPWR.t358 646.071
R10391 VPWR.n813 VPWR.t103 646.071
R10392 VPWR.n812 VPWR.t251 646.071
R10393 VPWR.n809 VPWR.t1345 646.071
R10394 VPWR.n808 VPWR.t1145 646.071
R10395 VPWR.n805 VPWR.t462 646.071
R10396 VPWR.n804 VPWR.t671 646.071
R10397 VPWR.n878 VPWR.t1257 646.071
R10398 VPWR.n834 VPWR.t331 646.071
R10399 VPWR.n890 VPWR.t1686 646.071
R10400 VPWR.n886 VPWR.t387 646.071
R10401 VPWR.n882 VPWR.t579 646.071
R10402 VPWR.n874 VPWR.t277 646.071
R10403 VPWR.n870 VPWR.t1089 646.071
R10404 VPWR.n866 VPWR.t1427 646.071
R10405 VPWR.n862 VPWR.t1171 646.071
R10406 VPWR.n858 VPWR.t1061 646.071
R10407 VPWR.n854 VPWR.t77 646.071
R10408 VPWR.n850 VPWR.t562 646.071
R10409 VPWR.n846 VPWR.t1354 646.071
R10410 VPWR.n842 VPWR.t1655 646.071
R10411 VPWR.n838 VPWR.t1366 646.071
R10412 VPWR.n835 VPWR.t846 646.071
R10413 VPWR.n908 VPWR.t1589 646.071
R10414 VPWR.n947 VPWR.t1707 646.071
R10415 VPWR.n1436 VPWR.t608 646.071
R10416 VPWR.n1149 VPWR.t786 646.071
R10417 VPWR.n367 VPWR.t552 646.071
R10418 VPWR.n329 VPWR.t137 646.071
R10419 VPWR.n306 VPWR.t1469 646.071
R10420 VPWR.n92 VPWR.t685 646.071
R10421 VPWR.n943 VPWR.t1290 646.071
R10422 VPWR.n1440 VPWR.t139 646.071
R10423 VPWR.n1153 VPWR.t950 646.071
R10424 VPWR.n909 VPWR.t209 646.071
R10425 VPWR.n951 VPWR.t283 646.071
R10426 VPWR.n1432 VPWR.t217 646.071
R10427 VPWR.n1145 VPWR.t816 646.071
R10428 VPWR.n383 VPWR.t1396 646.071
R10429 VPWR.n387 VPWR.t375 646.071
R10430 VPWR.n391 VPWR.t360 646.071
R10431 VPWR.n395 VPWR.t105 646.071
R10432 VPWR.n399 VPWR.t253 646.071
R10433 VPWR.n403 VPWR.t1347 646.071
R10434 VPWR.n407 VPWR.t1231 646.071
R10435 VPWR.n411 VPWR.t466 646.071
R10436 VPWR.n354 VPWR.t665 646.071
R10437 VPWR.n336 VPWR.t273 646.071
R10438 VPWR.n294 VPWR.t1457 646.071
R10439 VPWR.n81 VPWR.t695 646.071
R10440 VPWR.n955 VPWR.t538 646.071
R10441 VPWR.n1428 VPWR.t1625 646.071
R10442 VPWR.n1141 VPWR.t958 646.071
R10443 VPWR.n916 VPWR.t1898 646.071
R10444 VPWR.n917 VPWR.t190 646.071
R10445 VPWR.n920 VPWR.t87 646.071
R10446 VPWR.n921 VPWR.t1505 646.071
R10447 VPWR.n924 VPWR.t169 646.071
R10448 VPWR.n925 VPWR.t1471 646.071
R10449 VPWR.n928 VPWR.t436 646.071
R10450 VPWR.n929 VPWR.t947 646.071
R10451 VPWR.n959 VPWR.t1435 646.071
R10452 VPWR.n1424 VPWR.t508 646.071
R10453 VPWR.n1137 VPWR.t703 646.071
R10454 VPWR.n328 VPWR.t43 646.071
R10455 VPWR.n310 VPWR.t23 646.071
R10456 VPWR.n93 VPWR.t647 646.071
R10457 VPWR.n1444 VPWR.t45 646.071
R10458 VPWR.n1157 VPWR.t911 646.071
R10459 VPWR.n963 VPWR.t1177 646.071
R10460 VPWR.n1420 VPWR.t1906 646.071
R10461 VPWR.n1133 VPWR.t719 646.071
R10462 VPWR.n344 VPWR.t93 646.071
R10463 VPWR.n345 VPWR.t1509 646.071
R10464 VPWR.n348 VPWR.t173 646.071
R10465 VPWR.n349 VPWR.t1475 646.071
R10466 VPWR.n352 VPWR.t444 646.071
R10467 VPWR.n353 VPWR.t933 646.071
R10468 VPWR.n282 VPWR.t188 646.071
R10469 VPWR.n74 VPWR.t677 646.071
R10470 VPWR.n1412 VPWR.t299 646.071
R10471 VPWR.n1129 VPWR.t936 646.071
R10472 VPWR.n971 VPWR.t69 646.071
R10473 VPWR.n975 VPWR.t1493 646.071
R10474 VPWR.n979 VPWR.t1362 646.071
R10475 VPWR.n983 VPWR.t1487 646.071
R10476 VPWR.n987 VPWR.t1374 646.071
R10477 VPWR.n930 VPWR.t805 646.071
R10478 VPWR.n1455 VPWR.t1539 646.071
R10479 VPWR.n1161 VPWR.t895 646.071
R10480 VPWR.n278 VPWR.t99 646.071
R10481 VPWR.n69 VPWR.t711 646.071
R10482 VPWR.n1125 VPWR.t984 646.071
R10483 VPWR.n1017 VPWR.t1511 646.071
R10484 VPWR.n1121 VPWR.t727 646.071
R10485 VPWR.n270 VPWR.t1119 646.071
R10486 VPWR.n262 VPWR.t470 646.071
R10487 VPWR.n259 VPWR.t979 646.071
R10488 VPWR.n1026 VPWR.t874 646.071
R10489 VPWR.n1684 VPWR.t1073 646.071
R10490 VPWR.n1004 VPWR.t448 646.071
R10491 VPWR.n1000 VPWR.t916 646.071
R10492 VPWR.n1117 VPWR.t859 646.071
R10493 VPWR.n63 VPWR.t976 646.071
R10494 VPWR.n57 VPWR.t756 646.071
R10495 VPWR.n2245 VPWR.t1240 629.652
R10496 VPWR.n2246 VPWR.t176 629.652
R10497 VPWR.n2255 VPWR.t38 629.652
R10498 VPWR.n2256 VPWR.t1924 629.652
R10499 VPWR.n2265 VPWR.t1714 629.652
R10500 VPWR.n2266 VPWR.t1554 629.652
R10501 VPWR.n2275 VPWR.t1385 629.652
R10502 VPWR.n2276 VPWR.t513 629.652
R10503 VPWR.n2285 VPWR.t232 629.652
R10504 VPWR.n2286 VPWR.t290 629.652
R10505 VPWR.n2295 VPWR.t62 629.652
R10506 VPWR.n2296 VPWR.t1498 629.652
R10507 VPWR.n2305 VPWR.t1604 629.652
R10508 VPWR.n2306 VPWR.t1082 629.652
R10509 VPWR.n2315 VPWR.t1383 629.652
R10510 VPWR.n510 VPWR.t1021 629.652
R10511 VPWR.t1792 VPWR.n509 629.652
R10512 VPWR.t18 VPWR.n505 629.652
R10513 VPWR.t1466 VPWR.n501 629.652
R10514 VPWR.t1578 VPWR.n497 629.652
R10515 VPWR.t1512 VPWR.n493 629.652
R10516 VPWR.t1454 VPWR.n489 629.652
R10517 VPWR.t1865 VPWR.n485 629.652
R10518 VPWR.t1842 VPWR.n481 629.652
R10519 VPWR.t322 VPWR.n477 629.652
R10520 VPWR.t94 VPWR.n473 629.652
R10521 VPWR.t258 VPWR.n469 629.652
R10522 VPWR.t1116 VPWR.n465 629.652
R10523 VPWR.t1648 VPWR.n461 629.652
R10524 VPWR.t467 VPWR.n457 629.652
R10525 VPWR.n2217 VPWR.t334 629.652
R10526 VPWR.t1689 VPWR.n2216 629.652
R10527 VPWR.n2207 VPWR.t1881 629.652
R10528 VPWR.t1283 VPWR.n2206 629.652
R10529 VPWR.n2197 VPWR.t1702 629.652
R10530 VPWR.t280 VPWR.n2196 629.652
R10531 VPWR.n2187 VPWR.t1094 629.652
R10532 VPWR.t1430 VPWR.n2186 629.652
R10533 VPWR.n2177 VPWR.t1174 629.652
R10534 VPWR.t1064 VPWR.n2176 629.652
R10535 VPWR.n2167 VPWR.t66 629.652
R10536 VPWR.t1488 VPWR.n2166 629.652
R10537 VPWR.n2157 VPWR.t1357 629.652
R10538 VPWR.t1658 VPWR.n2156 629.652
R10539 VPWR.n2147 VPWR.t1371 629.652
R10540 VPWR.n550 VPWR.t1029 629.652
R10541 VPWR.n554 VPWR.t1534 629.652
R10542 VPWR.n558 VPWR.t40 629.652
R10543 VPWR.n562 VPWR.t1295 629.652
R10544 VPWR.n566 VPWR.t1590 629.652
R10545 VPWR.n570 VPWR.t210 629.652
R10546 VPWR.n574 VPWR.t268 629.652
R10547 VPWR.n578 VPWR.t503 629.652
R10548 VPWR.n582 VPWR.t1899 629.652
R10549 VPWR.n586 VPWR.t191 629.652
R10550 VPWR.n590 VPWR.t88 629.652
R10551 VPWR.n594 VPWR.t1506 629.652
R10552 VPWR.n598 VPWR.t170 629.652
R10553 VPWR.n602 VPWR.t1472 629.652
R10554 VPWR.n606 VPWR.t439 629.652
R10555 VPWR.n2049 VPWR.t479 629.652
R10556 VPWR.n2050 VPWR.t1544 629.652
R10557 VPWR.n2059 VPWR.t1275 629.652
R10558 VPWR.n2060 VPWR.t547 629.652
R10559 VPWR.n2069 VPWR.t1598 629.652
R10560 VPWR.n2070 VPWR.t1812 629.652
R10561 VPWR.n2079 VPWR.t1100 629.652
R10562 VPWR.n2080 VPWR.t1391 629.652
R10563 VPWR.n2089 VPWR.t370 629.652
R10564 VPWR.n2090 VPWR.t355 629.652
R10565 VPWR.n2099 VPWR.t112 629.652
R10566 VPWR.n2100 VPWR.t248 629.652
R10567 VPWR.n2109 VPWR.t1342 629.652
R10568 VPWR.n2110 VPWR.t1142 629.652
R10569 VPWR.n2119 VPWR.t459 629.652
R10570 VPWR.n702 VPWR.t1238 629.652
R10571 VPWR.t1444 VPWR.n701 629.652
R10572 VPWR.t36 VPWR.n697 629.652
R10573 VPWR.t1922 VPWR.n693 629.652
R10574 VPWR.t1712 VPWR.n689 629.652
R10575 VPWR.t1552 VPWR.n685 629.652
R10576 VPWR.t541 VPWR.n681 629.652
R10577 VPWR.t511 VPWR.n677 629.652
R10578 VPWR.t230 VPWR.n673 629.652
R10579 VPWR.t288 VPWR.n669 629.652
R10580 VPWR.t60 VPWR.n665 629.652
R10581 VPWR.t1496 VPWR.n661 629.652
R10582 VPWR.t1602 VPWR.n657 629.652
R10583 VPWR.t1080 VPWR.n653 629.652
R10584 VPWR.t1377 VPWR.n649 629.652
R10585 VPWR.n2021 VPWR.t1033 629.652
R10586 VPWR.t1691 VPWR.n2020 629.652
R10587 VPWR.n2011 VPWR.t1267 629.652
R10588 VPWR.t1056 VPWR.n2010 629.652
R10589 VPWR.n2001 VPWR.t1697 629.652
R10590 VPWR.t1556 VPWR.n2000 629.652
R10591 VPWR.n1991 VPWR.t164 629.652
R10592 VPWR.t517 VPWR.n1990 629.652
R10593 VPWR.n1981 VPWR.t234 629.652
R10594 VPWR.t344 VPWR.n1980 629.652
R10595 VPWR.n1971 VPWR.t114 629.652
R10596 VPWR.t1616 VPWR.n1970 629.652
R10597 VPWR.n1961 VPWR.t1409 629.652
R10598 VPWR.t597 VPWR.n1960 629.652
R10599 VPWR.n1951 VPWR.t493 629.652
R10600 VPWR.n742 VPWR.t332 629.652
R10601 VPWR.n746 VPWR.t1687 629.652
R10602 VPWR.n750 VPWR.t1879 629.652
R10603 VPWR.n754 VPWR.t1281 629.652
R10604 VPWR.n758 VPWR.t1700 629.652
R10605 VPWR.n762 VPWR.t278 629.652
R10606 VPWR.n766 VPWR.t1092 629.652
R10607 VPWR.n770 VPWR.t1428 629.652
R10608 VPWR.n774 VPWR.t1172 629.652
R10609 VPWR.n778 VPWR.t1062 629.652
R10610 VPWR.n782 VPWR.t64 629.652
R10611 VPWR.n786 VPWR.t563 629.652
R10612 VPWR.n790 VPWR.t1355 629.652
R10613 VPWR.n794 VPWR.t1656 629.652
R10614 VPWR.n798 VPWR.t1369 629.652
R10615 VPWR.n1853 VPWR.t591 629.652
R10616 VPWR.n1854 VPWR.t1546 629.652
R10617 VPWR.n1863 VPWR.t26 629.652
R10618 VPWR.n1864 VPWR.t549 629.652
R10619 VPWR.n1873 VPWR.t1522 629.652
R10620 VPWR.n1874 VPWR.t1814 629.652
R10621 VPWR.n1883 VPWR.t1102 629.652
R10622 VPWR.n1884 VPWR.t1393 629.652
R10623 VPWR.n1893 VPWR.t372 629.652
R10624 VPWR.n1894 VPWR.t357 629.652
R10625 VPWR.n1903 VPWR.t102 629.652
R10626 VPWR.n1904 VPWR.t250 629.652
R10627 VPWR.n1913 VPWR.t1344 629.652
R10628 VPWR.n1914 VPWR.t1144 629.652
R10629 VPWR.n1923 VPWR.t461 629.652
R10630 VPWR.n894 VPWR.t330 629.652
R10631 VPWR.t1685 VPWR.n893 629.652
R10632 VPWR.t386 VPWR.n889 629.652
R10633 VPWR.t578 VPWR.n885 629.652
R10634 VPWR.t1256 VPWR.n881 629.652
R10635 VPWR.t276 VPWR.n877 629.652
R10636 VPWR.t1088 VPWR.n873 629.652
R10637 VPWR.t1426 VPWR.n869 629.652
R10638 VPWR.t1170 VPWR.n865 629.652
R10639 VPWR.t1060 VPWR.n861 629.652
R10640 VPWR.t76 VPWR.n857 629.652
R10641 VPWR.t561 VPWR.n853 629.652
R10642 VPWR.t1353 VPWR.n849 629.652
R10643 VPWR.t1654 VPWR.n845 629.652
R10644 VPWR.t1365 VPWR.n841 629.652
R10645 VPWR.n358 VPWR.t593 629.652
R10646 VPWR.n362 VPWR.t1548 629.652
R10647 VPWR.n366 VPWR.t28 629.652
R10648 VPWR.n370 VPWR.t551 629.652
R10649 VPWR.n374 VPWR.t1524 629.652
R10650 VPWR.n378 VPWR.t1816 629.652
R10651 VPWR.n382 VPWR.t1106 629.652
R10652 VPWR.n386 VPWR.t1395 629.652
R10653 VPWR.n390 VPWR.t374 629.652
R10654 VPWR.n394 VPWR.t359 629.652
R10655 VPWR.n398 VPWR.t104 629.652
R10656 VPWR.n402 VPWR.t252 629.652
R10657 VPWR.n406 VPWR.t1346 629.652
R10658 VPWR.n410 VPWR.t1230 629.652
R10659 VPWR.n414 VPWR.t465 629.652
R10660 VPWR.n1825 VPWR.t1027 629.652
R10661 VPWR.t1802 VPWR.n1824 629.652
R10662 VPWR.n1815 VPWR.t24 629.652
R10663 VPWR.t1293 VPWR.n1814 629.652
R10664 VPWR.n1805 VPWR.t1588 629.652
R10665 VPWR.t208 VPWR.n1804 629.652
R10666 VPWR.n1795 VPWR.t264 629.652
R10667 VPWR.t501 VPWR.n1794 629.652
R10668 VPWR.n1785 VPWR.t1897 629.652
R10669 VPWR.t189 VPWR.n1784 629.652
R10670 VPWR.n1775 VPWR.t86 629.652
R10671 VPWR.t1504 VPWR.n1774 629.652
R10672 VPWR.n1765 VPWR.t168 629.652
R10673 VPWR.t1470 VPWR.n1764 629.652
R10674 VPWR.n1755 VPWR.t435 629.652
R10675 VPWR.n2413 VPWR.t1031 629.652
R10676 VPWR.t1536 VPWR.n2412 629.652
R10677 VPWR.n2403 VPWR.t42 629.652
R10678 VPWR.t136 VPWR.n2402 629.652
R10679 VPWR.n2393 VPWR.t1336 629.652
R10680 VPWR.t214 VPWR.n2392 629.652
R10681 VPWR.n2383 VPWR.t272 629.652
R10682 VPWR.t505 VPWR.n2382 629.652
R10683 VPWR.n2373 VPWR.t1903 629.652
R10684 VPWR.t193 VPWR.n2372 629.652
R10685 VPWR.n2363 VPWR.t92 629.652
R10686 VPWR.t1508 VPWR.n2362 629.652
R10687 VPWR.n2353 VPWR.t172 629.652
R10688 VPWR.t1474 VPWR.n2352 629.652
R10689 VPWR.n2343 VPWR.t443 629.652
R10690 VPWR.n934 VPWR.t1236 629.652
R10691 VPWR.n938 VPWR.t1438 629.652
R10692 VPWR.n942 VPWR.t1885 629.652
R10693 VPWR.n946 VPWR.t1289 629.652
R10694 VPWR.n950 VPWR.t1706 629.652
R10695 VPWR.n954 VPWR.t282 629.652
R10696 VPWR.n958 VPWR.t537 629.652
R10697 VPWR.n962 VPWR.t1434 629.652
R10698 VPWR.n966 VPWR.t1176 629.652
R10699 VPWR.n970 VPWR.t1068 629.652
R10700 VPWR.n974 VPWR.t68 629.652
R10701 VPWR.n978 VPWR.t1492 629.652
R10702 VPWR.n982 VPWR.t1361 629.652
R10703 VPWR.n986 VPWR.t1486 629.652
R10704 VPWR.n990 VPWR.t1373 629.652
R10705 VPWR.n318 VPWR.t1023 629.652
R10706 VPWR.t1794 VPWR.n317 629.652
R10707 VPWR.t22 VPWR.n313 629.652
R10708 VPWR.t1468 VPWR.n309 629.652
R10709 VPWR.t1580 VPWR.n305 629.652
R10710 VPWR.t1516 VPWR.n301 629.652
R10711 VPWR.t1456 VPWR.n297 629.652
R10712 VPWR.t1867 VPWR.n293 629.652
R10713 VPWR.t1891 VPWR.n289 629.652
R10714 VPWR.t187 VPWR.n285 629.652
R10715 VPWR.t98 VPWR.n281 629.652
R10716 VPWR.t262 VPWR.n277 629.652
R10717 VPWR.t1118 VPWR.n273 629.652
R10718 VPWR.t1650 VPWR.n269 629.652
R10719 VPWR.t469 VPWR.n265 629.652
R10720 VPWR.n1451 VPWR.t1848 629.652
R10721 VPWR.n1457 VPWR.t1538 629.652
R10722 VPWR.n1458 VPWR.t44 629.652
R10723 VPWR.n1470 VPWR.t138 629.652
R10724 VPWR.n1471 VPWR.t607 629.652
R10725 VPWR.n1484 VPWR.t216 629.652
R10726 VPWR.n1485 VPWR.t1624 629.652
R10727 VPWR.n1498 VPWR.t507 629.652
R10728 VPWR.n1499 VPWR.t1905 629.652
R10729 VPWR.n1514 VPWR.t298 629.652
R10730 VPWR.t78 VPWR.n1513 629.652
R10731 VPWR.n1697 VPWR.t1510 629.652
R10732 VPWR.t174 VPWR.n1696 629.652
R10733 VPWR.n1685 VPWR.t1072 629.652
R10734 VPWR.n1727 VPWR.t447 629.652
R10735 VPWR.n2442 VPWR.t777 629.652
R10736 VPWR.n2443 VPWR.t634 629.652
R10737 VPWR.n2454 VPWR.t646 629.652
R10738 VPWR.n2455 VPWR.t684 629.652
R10739 VPWR.n2466 VPWR.t902 629.652
R10740 VPWR.n2467 VPWR.t941 629.652
R10741 VPWR.n2478 VPWR.t694 629.652
R10742 VPWR.n2479 VPWR.t812 629.652
R10743 VPWR.n2490 VPWR.t828 629.652
R10744 VPWR.n2491 VPWR.t676 629.652
R10745 VPWR.n2502 VPWR.t710 629.652
R10746 VPWR.n2503 VPWR.t842 629.652
R10747 VPWR.n2514 VPWR.t975 629.652
R10748 VPWR.n2515 VPWR.t616 629.652
R10749 VPWR.n2526 VPWR.t755 629.652
R10750 VPWR.n1165 VPWR.t654 629.652
R10751 VPWR.t894 VPWR.n1164 629.652
R10752 VPWR.t910 VPWR.n1160 629.652
R10753 VPWR.t949 VPWR.n1156 629.652
R10754 VPWR.t785 VPWR.n1152 629.652
R10755 VPWR.t815 VPWR.n1148 629.652
R10756 VPWR.t957 VPWR.n1144 629.652
R10757 VPWR.t702 VPWR.n1140 629.652
R10758 VPWR.t718 VPWR.n1136 629.652
R10759 VPWR.t935 VPWR.n1132 629.652
R10760 VPWR.t983 VPWR.n1128 629.652
R10761 VPWR.t726 VPWR.n1124 629.652
R10762 VPWR.t858 VPWR.n1120 629.652
R10763 VPWR.n1676 VPWR.t873 629.652
R10764 VPWR.t626 VPWR.n1675 629.652
R10765 VPWR.n2772 VPWR.t1210 531.804
R10766 VPWR.n2791 VPWR.t1210 531.804
R10767 VPWR.n2787 VPWR.n2786 504.707
R10768 VPWR.t1818 VPWR.t1200 497.094
R10769 VPWR.t1240 VPWR.t1818 497.094
R10770 VPWR.t1878 VPWR.t1846 497.094
R10771 VPWR.t176 VPWR.t1878 497.094
R10772 VPWR.t1442 VPWR.t1877 497.094
R10773 VPWR.t1877 VPWR.t38 497.094
R10774 VPWR.t224 VPWR.t1887 497.094
R10775 VPWR.t1924 VPWR.t224 497.094
R10776 VPWR.t1464 VPWR.t382 497.094
R10777 VPWR.t382 VPWR.t1714 497.094
R10778 VPWR.t381 VPWR.t1710 497.094
R10779 VPWR.t1554 VPWR.t381 497.094
R10780 VPWR.t220 VPWR.t223 497.094
R10781 VPWR.t223 VPWR.t1385 497.094
R10782 VPWR.t1406 VPWR.t1628 497.094
R10783 VPWR.t513 VPWR.t1406 497.094
R10784 VPWR.t509 VPWR.t1405 497.094
R10785 VPWR.t1405 VPWR.t232 497.094
R10786 VPWR.t398 VPWR.t1909 497.094
R10787 VPWR.t290 VPWR.t398 497.094
R10788 VPWR.t1070 VPWR.t222 497.094
R10789 VPWR.t222 VPWR.t62 497.094
R10790 VPWR.t1404 VPWR.t82 497.094
R10791 VPWR.t1498 VPWR.t1404 497.094
R10792 VPWR.t1494 VPWR.t397 497.094
R10793 VPWR.t397 VPWR.t1604 497.094
R10794 VPWR.t396 VPWR.t1600 497.094
R10795 VPWR.t1082 VPWR.t396 497.094
R10796 VPWR.t1478 VPWR.t1819 497.094
R10797 VPWR.t1819 VPWR.t1383 497.094
R10798 VPWR.t383 VPWR.t451 497.094
R10799 VPWR.t766 VPWR.t383 497.094
R10800 VPWR.t328 VPWR.t1222 497.094
R10801 VPWR.t1021 VPWR.t328 497.094
R10802 VPWR.t1242 VPWR.t365 497.094
R10803 VPWR.t365 VPWR.t1792 497.094
R10804 VPWR.t1400 VPWR.t364 497.094
R10805 VPWR.t364 VPWR.t18 497.094
R10806 VPWR.t30 VPWR.t363 497.094
R10807 VPWR.t363 VPWR.t1466 497.094
R10808 VPWR.t1285 VPWR.t341 497.094
R10809 VPWR.t341 VPWR.t1578 497.094
R10810 VPWR.t1526 VPWR.t369 497.094
R10811 VPWR.t369 VPWR.t1512 497.094
R10812 VPWR.t1558 VPWR.t362 497.094
R10813 VPWR.t362 VPWR.t1454 497.094
R10814 VPWR.t425 VPWR.t327 497.094
R10815 VPWR.t327 VPWR.t1865 497.094
R10816 VPWR.t1861 VPWR.t326 497.094
R10817 VPWR.t326 VPWR.t1842 497.094
R10818 VPWR.t236 VPWR.t368 497.094
R10819 VPWR.t368 VPWR.t322 497.094
R10820 VPWR.t314 VPWR.t361 497.094
R10821 VPWR.t361 VPWR.t94 497.094
R10822 VPWR.t116 VPWR.t325 497.094
R10823 VPWR.t325 VPWR.t258 497.094
R10824 VPWR.t565 VPWR.t367 497.094
R10825 VPWR.t367 VPWR.t1116 497.094
R10826 VPWR.t1112 VPWR.t366 497.094
R10827 VPWR.t366 VPWR.t1648 497.094
R10828 VPWR.t1084 VPWR.t329 497.094
R10829 VPWR.t329 VPWR.t467 497.094
R10830 VPWR.t471 VPWR.t324 497.094
R10831 VPWR.t324 VPWR.t986 497.094
R10832 VPWR.t1334 VPWR.t1206 497.094
R10833 VPWR.t334 VPWR.t1334 497.094
R10834 VPWR.t1019 VPWR.t380 497.094
R10835 VPWR.t380 VPWR.t1689 497.094
R10836 VPWR.t379 VPWR.t1683 497.094
R10837 VPWR.t1881 VPWR.t379 497.094
R10838 VPWR.t997 VPWR.t378 497.094
R10839 VPWR.t378 VPWR.t1283 497.094
R10840 VPWR.t1329 VPWR.t584 497.094
R10841 VPWR.t1702 VPWR.t1329 497.094
R10842 VPWR.t1254 VPWR.t1325 497.094
R10843 VPWR.t1325 VPWR.t280 497.094
R10844 VPWR.t377 VPWR.t1520 497.094
R10845 VPWR.t1094 VPWR.t377 497.094
R10846 VPWR.t270 VPWR.t1333 497.094
R10847 VPWR.t1333 VPWR.t1430 497.094
R10848 VPWR.t1332 VPWR.t1424 497.094
R10849 VPWR.t1174 VPWR.t1332 497.094
R10850 VPWR.t1895 VPWR.t1324 497.094
R10851 VPWR.t1324 VPWR.t1064 497.094
R10852 VPWR.t376 VPWR.t304 497.094
R10853 VPWR.t66 VPWR.t376 497.094
R10854 VPWR.t84 VPWR.t1331 497.094
R10855 VPWR.t1331 VPWR.t1488 497.094
R10856 VPWR.t1323 VPWR.t423 497.094
R10857 VPWR.t1357 VPWR.t1323 497.094
R10858 VPWR.t1612 VPWR.t1322 497.094
R10859 VPWR.t1322 VPWR.t1658 497.094
R10860 VPWR.t1335 VPWR.t1646 497.094
R10861 VPWR.t1371 VPWR.t1335 497.094
R10862 VPWR.t441 VPWR.t1330 497.094
R10863 VPWR.t1330 VPWR.t820 497.094
R10864 VPWR.t296 VPWR.t1216 497.094
R10865 VPWR.t1029 VPWR.t296 497.094
R10866 VPWR.t1262 VPWR.t1037 497.094
R10867 VPWR.t1534 VPWR.t1262 497.094
R10868 VPWR.t1261 VPWR.t1798 497.094
R10869 VPWR.t40 VPWR.t1261 497.094
R10870 VPWR.t1260 VPWR.t16 497.094
R10871 VPWR.t1295 VPWR.t1260 497.094
R10872 VPWR.t340 VPWR.t1918 497.094
R10873 VPWR.t1590 VPWR.t340 497.094
R10874 VPWR.t1266 VPWR.t1584 497.094
R10875 VPWR.t210 VPWR.t1266 497.094
R10876 VPWR.t1259 VPWR.t1808 497.094
R10877 VPWR.t268 VPWR.t1259 497.094
R10878 VPWR.t295 VPWR.t431 497.094
R10879 VPWR.t503 VPWR.t295 497.094
R10880 VPWR.t294 VPWR.t497 497.094
R10881 VPWR.t1899 VPWR.t294 497.094
R10882 VPWR.t1265 VPWR.t242 497.094
R10883 VPWR.t191 VPWR.t1265 497.094
R10884 VPWR.t1258 VPWR.t320 497.094
R10885 VPWR.t88 VPWR.t1258 497.094
R10886 VPWR.t293 VPWR.t108 497.094
R10887 VPWR.t1506 VPWR.t293 497.094
R10888 VPWR.t1264 VPWR.t256 497.094
R10889 VPWR.t170 VPWR.t1264 497.094
R10890 VPWR.t1263 VPWR.t1122 497.094
R10891 VPWR.t1472 VPWR.t1263 497.094
R10892 VPWR.t297 VPWR.t601 497.094
R10893 VPWR.t439 VPWR.t297 497.094
R10894 VPWR.t292 VPWR.t457 497.094
R10895 VPWR.t938 VPWR.t292 497.094
R10896 VPWR.t183 VPWR.t1228 497.094
R10897 VPWR.t479 VPWR.t183 497.094
R10898 VPWR.t1076 VPWR.t336 497.094
R10899 VPWR.t1544 VPWR.t1076 497.094
R10900 VPWR.t1693 VPWR.t478 497.094
R10901 VPWR.t478 VPWR.t1275 497.094
R10902 VPWR.t477 VPWR.t1269 497.094
R10903 VPWR.t547 VPWR.t477 497.094
R10904 VPWR.t140 VPWR.t1138 497.094
R10905 VPWR.t1138 VPWR.t1598 497.094
R10906 VPWR.t1137 VPWR.t1592 497.094
R10907 VPWR.t1812 VPWR.t1137 497.094
R10908 VPWR.t284 VPWR.t476 497.094
R10909 VPWR.t476 VPWR.t1100 497.094
R10910 VPWR.t530 VPWR.t539 497.094
R10911 VPWR.t1391 VPWR.t530 497.094
R10912 VPWR.t519 VPWR.t529 497.094
R10913 VPWR.t529 VPWR.t370 497.094
R10914 VPWR.t1079 VPWR.t1178 497.094
R10915 VPWR.t355 VPWR.t1079 497.094
R10916 VPWR.t349 VPWR.t475 497.094
R10917 VPWR.t475 VPWR.t112 497.094
R10918 VPWR.t528 VPWR.t70 497.094
R10919 VPWR.t248 VPWR.t528 497.094
R10920 VPWR.t1108 VPWR.t1078 497.094
R10921 VPWR.t1078 VPWR.t1342 497.094
R10922 VPWR.t1077 VPWR.t1411 497.094
R10923 VPWR.t1142 VPWR.t1077 497.094
R10924 VPWR.t1480 VPWR.t184 497.094
R10925 VPWR.t184 VPWR.t459 497.094
R10926 VPWR.t1139 VPWR.t1375 497.094
R10927 VPWR.t673 VPWR.t1139 497.094
R10928 VPWR.t1661 VPWR.t1202 497.094
R10929 VPWR.t1238 VPWR.t1661 497.094
R10930 VPWR.t1844 VPWR.t522 497.094
R10931 VPWR.t522 VPWR.t1444 497.094
R10932 VPWR.t1440 VPWR.t521 497.094
R10933 VPWR.t521 VPWR.t36 497.094
R10934 VPWR.t1883 VPWR.t1328 497.094
R10935 VPWR.t1328 VPWR.t1922 497.094
R10936 VPWR.t1462 VPWR.t1838 497.094
R10937 VPWR.t1838 VPWR.t1712 497.094
R10938 VPWR.t1708 VPWR.t526 497.094
R10939 VPWR.t526 VPWR.t1552 497.094
R10940 VPWR.t218 VPWR.t1327 497.094
R10941 VPWR.t1327 VPWR.t541 497.094
R10942 VPWR.t1626 VPWR.t1660 497.094
R10943 VPWR.t1660 VPWR.t511 497.094
R10944 VPWR.t1436 VPWR.t1841 497.094
R10945 VPWR.t1841 VPWR.t230 497.094
R10946 VPWR.t1907 VPWR.t525 497.094
R10947 VPWR.t525 VPWR.t288 497.094
R10948 VPWR.t1066 VPWR.t1326 497.094
R10949 VPWR.t1326 VPWR.t60 497.094
R10950 VPWR.t80 VPWR.t1840 497.094
R10951 VPWR.t1840 VPWR.t1496 497.094
R10952 VPWR.t1490 VPWR.t524 497.094
R10953 VPWR.t524 VPWR.t1602 497.094
R10954 VPWR.t1363 VPWR.t523 497.094
R10955 VPWR.t523 VPWR.t1080 497.094
R10956 VPWR.t1476 VPWR.t1662 497.094
R10957 VPWR.t1662 VPWR.t1377 497.094
R10958 VPWR.t449 VPWR.t1839 497.094
R10959 VPWR.t1839 VPWR.t774 497.094
R10960 VPWR.t313 VPWR.t1198 497.094
R10961 VPWR.t1033 VPWR.t313 497.094
R10962 VPWR.t1850 VPWR.t1791 497.094
R10963 VPWR.t1791 VPWR.t1691 497.094
R10964 VPWR.t1790 VPWR.t178 497.094
R10965 VPWR.t1267 VPWR.t1790 497.094
R10966 VPWR.t56 VPWR.t1789 497.094
R10967 VPWR.t1789 VPWR.t1056 497.094
R10968 VPWR.t1397 VPWR.t1291 497.094
R10969 VPWR.t1697 VPWR.t1397 497.094
R10970 VPWR.t1695 VPWR.t309 497.094
R10971 VPWR.t309 VPWR.t1556 497.094
R10972 VPWR.t1788 VPWR.t46 497.094
R10973 VPWR.t164 VPWR.t1788 497.094
R10974 VPWR.t1090 VPWR.t312 497.094
R10975 VPWR.t312 VPWR.t517 497.094
R10976 VPWR.t311 VPWR.t515 497.094
R10977 VPWR.t234 VPWR.t311 497.094
R10978 VPWR.t1168 VPWR.t308 497.094
R10979 VPWR.t308 VPWR.t344 497.094
R10980 VPWR.t575 VPWR.t342 497.094
R10981 VPWR.t114 VPWR.t575 497.094
R10982 VPWR.t74 VPWR.t310 497.094
R10983 VPWR.t310 VPWR.t1616 497.094
R10984 VPWR.t307 VPWR.t1614 497.094
R10985 VPWR.t1409 VPWR.t307 497.094
R10986 VPWR.t1606 VPWR.t306 497.094
R10987 VPWR.t306 VPWR.t597 497.094
R10988 VPWR.t1399 VPWR.t1074 497.094
R10989 VPWR.t493 VPWR.t1399 497.094
R10990 VPWR.t1367 VPWR.t1398 497.094
R10991 VPWR.t1398 VPWR.t734 497.094
R10992 VPWR.t1306 VPWR.t1208 497.094
R10993 VPWR.t332 VPWR.t1306 497.094
R10994 VPWR.t150 VPWR.t1017 497.094
R10995 VPWR.t1687 VPWR.t150 497.094
R10996 VPWR.t149 VPWR.t1681 497.094
R10997 VPWR.t1879 VPWR.t149 497.094
R10998 VPWR.t1310 VPWR.t995 497.094
R10999 VPWR.t1281 VPWR.t1310 497.094
R11000 VPWR.t148 VPWR.t582 497.094
R11001 VPWR.t1700 VPWR.t148 497.094
R11002 VPWR.t147 VPWR.t1252 497.094
R11003 VPWR.t278 VPWR.t147 497.094
R11004 VPWR.t1309 VPWR.t1518 497.094
R11005 VPWR.t1092 VPWR.t1309 497.094
R11006 VPWR.t1305 VPWR.t266 497.094
R11007 VPWR.t1428 VPWR.t1305 497.094
R11008 VPWR.t1304 VPWR.t1422 497.094
R11009 VPWR.t1172 VPWR.t1304 497.094
R11010 VPWR.t146 VPWR.t1893 497.094
R11011 VPWR.t1062 VPWR.t146 497.094
R11012 VPWR.t1308 VPWR.t302 497.094
R11013 VPWR.t64 VPWR.t1308 497.094
R11014 VPWR.t1303 VPWR.t100 497.094
R11015 VPWR.t563 VPWR.t1303 497.094
R11016 VPWR.t145 VPWR.t421 497.094
R11017 VPWR.t1355 VPWR.t145 497.094
R11018 VPWR.t144 VPWR.t1610 497.094
R11019 VPWR.t1656 VPWR.t144 497.094
R11020 VPWR.t1307 VPWR.t1644 497.094
R11021 VPWR.t1369 VPWR.t1307 497.094
R11022 VPWR.t1302 VPWR.t437 497.094
R11023 VPWR.t836 VPWR.t1302 497.094
R11024 VPWR.t1098 VPWR.t1226 497.094
R11025 VPWR.t591 VPWR.t1098 497.094
R11026 VPWR.t1298 VPWR.t338 497.094
R11027 VPWR.t1546 VPWR.t1298 497.094
R11028 VPWR.t1540 VPWR.t1297 497.094
R11029 VPWR.t1297 VPWR.t26 497.094
R11030 VPWR.t1453 VPWR.t1271 497.094
R11031 VPWR.t549 VPWR.t1453 497.094
R11032 VPWR.t142 VPWR.t484 497.094
R11033 VPWR.t484 VPWR.t1522 497.094
R11034 VPWR.t483 VPWR.t1594 497.094
R11035 VPWR.t1814 VPWR.t483 497.094
R11036 VPWR.t286 VPWR.t1452 497.094
R11037 VPWR.t1452 VPWR.t1102 497.094
R11038 VPWR.t572 VPWR.t543 497.094
R11039 VPWR.t1393 VPWR.t572 497.094
R11040 VPWR.t1387 VPWR.t571 497.094
R11041 VPWR.t571 VPWR.t372 497.094
R11042 VPWR.t482 VPWR.t1180 497.094
R11043 VPWR.t357 VPWR.t482 497.094
R11044 VPWR.t351 VPWR.t1451 497.094
R11045 VPWR.t1451 VPWR.t102 497.094
R11046 VPWR.t570 VPWR.t72 497.094
R11047 VPWR.t250 VPWR.t570 497.094
R11048 VPWR.t1110 VPWR.t481 497.094
R11049 VPWR.t481 VPWR.t1344 497.094
R11050 VPWR.t1299 VPWR.t1413 497.094
R11051 VPWR.t1144 VPWR.t1299 497.094
R11052 VPWR.t1482 VPWR.t1099 497.094
R11053 VPWR.t1099 VPWR.t461 497.094
R11054 VPWR.t569 VPWR.t1379 497.094
R11055 VPWR.t670 VPWR.t569 497.094
R11056 VPWR.t1577 VPWR.t1212 497.094
R11057 VPWR.t330 VPWR.t1577 497.094
R11058 VPWR.t595 VPWR.t1680 497.094
R11059 VPWR.t1680 VPWR.t1685 497.094
R11060 VPWR.t1417 VPWR.t1679 497.094
R11061 VPWR.t1679 VPWR.t386 497.094
R11062 VPWR.t993 VPWR.t1678 497.094
R11063 VPWR.t1678 VPWR.t578 497.094
R11064 VPWR.t580 VPWR.t1572 497.094
R11065 VPWR.t1572 VPWR.t1256 497.094
R11066 VPWR.t1250 VPWR.t1280 497.094
R11067 VPWR.t1280 VPWR.t276 497.094
R11068 VPWR.t1514 VPWR.t1677 497.094
R11069 VPWR.t1677 VPWR.t1088 497.094
R11070 VPWR.t1458 VPWR.t1576 497.094
R11071 VPWR.t1576 VPWR.t1426 497.094
R11072 VPWR.t1420 VPWR.t1575 497.094
R11073 VPWR.t1575 VPWR.t1170 497.094
R11074 VPWR.t1889 VPWR.t1279 497.094
R11075 VPWR.t1279 VPWR.t1060 497.094
R11076 VPWR.t300 VPWR.t1676 497.094
R11077 VPWR.t1676 VPWR.t76 497.094
R11078 VPWR.t96 VPWR.t1574 497.094
R11079 VPWR.t1574 VPWR.t561 497.094
R11080 VPWR.t419 VPWR.t1278 497.094
R11081 VPWR.t1278 VPWR.t1353 497.094
R11082 VPWR.t1608 VPWR.t1277 497.094
R11083 VPWR.t1277 VPWR.t1654 497.094
R11084 VPWR.t1232 VPWR.t1675 497.094
R11085 VPWR.t1675 VPWR.t1365 497.094
R11086 VPWR.t433 VPWR.t1573 497.094
R11087 VPWR.t1573 VPWR.t845 497.094
R11088 VPWR.t151 VPWR.t1224 497.094
R11089 VPWR.t593 VPWR.t151 497.094
R11090 VPWR.t1047 VPWR.t1234 497.094
R11091 VPWR.t1548 VPWR.t1047 497.094
R11092 VPWR.t1046 VPWR.t1542 497.094
R11093 VPWR.t28 VPWR.t1046 497.094
R11094 VPWR.t1045 VPWR.t1273 497.094
R11095 VPWR.t551 VPWR.t1045 497.094
R11096 VPWR.t1160 VPWR.t576 497.094
R11097 VPWR.t1524 VPWR.t1160 497.094
R11098 VPWR.t1159 VPWR.t1596 497.094
R11099 VPWR.t1816 VPWR.t1159 497.094
R11100 VPWR.t1044 VPWR.t1550 497.094
R11101 VPWR.t1106 VPWR.t1044 497.094
R11102 VPWR.t999 VPWR.t545 497.094
R11103 VPWR.t1395 VPWR.t999 497.094
R11104 VPWR.t1163 VPWR.t1389 497.094
R11105 VPWR.t374 VPWR.t1163 497.094
R11106 VPWR.t1158 VPWR.t1182 497.094
R11107 VPWR.t359 VPWR.t1158 497.094
R11108 VPWR.t153 VPWR.t353 497.094
R11109 VPWR.t104 VPWR.t153 497.094
R11110 VPWR.t1162 VPWR.t58 497.094
R11111 VPWR.t252 VPWR.t1162 497.094
R11112 VPWR.t1049 VPWR.t246 497.094
R11113 VPWR.t1346 VPWR.t1049 497.094
R11114 VPWR.t1048 VPWR.t1415 497.094
R11115 VPWR.t1230 VPWR.t1048 497.094
R11116 VPWR.t152 VPWR.t1484 497.094
R11117 VPWR.t465 VPWR.t152 497.094
R11118 VPWR.t1161 VPWR.t1381 497.094
R11119 VPWR.t664 VPWR.t1161 497.094
R11120 VPWR.t1248 VPWR.t1218 497.094
R11121 VPWR.t1027 VPWR.t1248 497.094
R11122 VPWR.t1035 VPWR.t1566 497.094
R11123 VPWR.t1566 VPWR.t1802 497.094
R11124 VPWR.t1565 VPWR.t1796 497.094
R11125 VPWR.t24 VPWR.t1565 497.094
R11126 VPWR.t14 VPWR.t1564 497.094
R11127 VPWR.t1564 VPWR.t1293 497.094
R11128 VPWR.t1571 VPWR.t1916 497.094
R11129 VPWR.t1588 VPWR.t1571 497.094
R11130 VPWR.t1582 VPWR.t1570 497.094
R11131 VPWR.t1570 VPWR.t208 497.094
R11132 VPWR.t1563 VPWR.t1806 497.094
R11133 VPWR.t264 VPWR.t1563 497.094
R11134 VPWR.t429 VPWR.t1247 497.094
R11135 VPWR.t1247 VPWR.t501 497.094
R11136 VPWR.t1246 VPWR.t495 497.094
R11137 VPWR.t1897 VPWR.t1246 497.094
R11138 VPWR.t240 VPWR.t1569 497.094
R11139 VPWR.t1569 VPWR.t189 497.094
R11140 VPWR.t1562 VPWR.t318 497.094
R11141 VPWR.t86 VPWR.t1562 497.094
R11142 VPWR.t106 VPWR.t410 497.094
R11143 VPWR.t410 VPWR.t1504 497.094
R11144 VPWR.t1568 VPWR.t254 497.094
R11145 VPWR.t168 VPWR.t1568 497.094
R11146 VPWR.t1120 VPWR.t1567 497.094
R11147 VPWR.t1567 VPWR.t1470 497.094
R11148 VPWR.t1249 VPWR.t599 497.094
R11149 VPWR.t435 VPWR.t1249 497.094
R11150 VPWR.t455 VPWR.t409 497.094
R11151 VPWR.t409 VPWR.t946 497.094
R11152 VPWR.t590 VPWR.t1214 497.094
R11153 VPWR.t1031 VPWR.t590 497.094
R11154 VPWR.t1039 VPWR.t1824 497.094
R11155 VPWR.t1824 VPWR.t1536 497.094
R11156 VPWR.t492 VPWR.t1800 497.094
R11157 VPWR.t42 VPWR.t492 497.094
R11158 VPWR.t20 VPWR.t491 497.094
R11159 VPWR.t491 VPWR.t136 497.094
R11160 VPWR.t1829 VPWR.t1920 497.094
R11161 VPWR.t1336 VPWR.t1829 497.094
R11162 VPWR.t1586 VPWR.t1828 497.094
R11163 VPWR.t1828 VPWR.t214 497.094
R11164 VPWR.t490 VPWR.t1810 497.094
R11165 VPWR.t272 VPWR.t490 497.094
R11166 VPWR.t1104 VPWR.t589 497.094
R11167 VPWR.t589 VPWR.t505 497.094
R11168 VPWR.t588 VPWR.t499 497.094
R11169 VPWR.t1903 VPWR.t588 497.094
R11170 VPWR.t244 VPWR.t1827 497.094
R11171 VPWR.t1827 VPWR.t193 497.094
R11172 VPWR.t489 VPWR.t185 497.094
R11173 VPWR.t92 VPWR.t489 497.094
R11174 VPWR.t110 VPWR.t587 497.094
R11175 VPWR.t587 VPWR.t1508 497.094
R11176 VPWR.t1826 VPWR.t260 497.094
R11177 VPWR.t172 VPWR.t1826 497.094
R11178 VPWR.t1124 VPWR.t1825 497.094
R11179 VPWR.t1825 VPWR.t1474 497.094
R11180 VPWR.t488 VPWR.t1140 497.094
R11181 VPWR.t443 VPWR.t488 497.094
R11182 VPWR.t463 VPWR.t586 497.094
R11183 VPWR.t586 VPWR.t932 497.094
R11184 VPWR.t1531 VPWR.t1204 497.094
R11185 VPWR.t1236 VPWR.t1531 497.094
R11186 VPWR.t1533 VPWR.t1025 497.094
R11187 VPWR.t1438 VPWR.t1533 497.094
R11188 VPWR.t527 VPWR.t1407 497.094
R11189 VPWR.t1885 VPWR.t527 497.094
R11190 VPWR.t1674 VPWR.t384 497.094
R11191 VPWR.t1289 VPWR.t1674 497.094
R11192 VPWR.t1500 VPWR.t553 497.094
R11193 VPWR.t1706 VPWR.t1500 497.094
R11194 VPWR.t1341 VPWR.t1704 497.094
R11195 VPWR.t282 VPWR.t1341 497.094
R11196 VPWR.t1673 VPWR.t212 497.094
R11197 VPWR.t537 VPWR.t1673 497.094
R11198 VPWR.t1530 VPWR.t1622 497.094
R11199 VPWR.t1434 VPWR.t1530 497.094
R11200 VPWR.t1503 VPWR.t1432 497.094
R11201 VPWR.t1176 VPWR.t1503 497.094
R11202 VPWR.t1340 VPWR.t1901 497.094
R11203 VPWR.t1068 VPWR.t1340 497.094
R11204 VPWR.t1672 VPWR.t1058 497.094
R11205 VPWR.t68 VPWR.t1672 497.094
R11206 VPWR.t1502 VPWR.t90 497.094
R11207 VPWR.t1492 VPWR.t1502 497.094
R11208 VPWR.t1339 VPWR.t559 497.094
R11209 VPWR.t1361 VPWR.t1339 497.094
R11210 VPWR.t1338 VPWR.t1359 497.094
R11211 VPWR.t1486 VPWR.t1338 497.094
R11212 VPWR.t1532 VPWR.t1652 497.094
R11213 VPWR.t1373 VPWR.t1532 497.094
R11214 VPWR.t1501 VPWR.t445 497.094
R11215 VPWR.t804 VPWR.t1501 497.094
R11216 VPWR.t1664 VPWR.t1220 497.094
R11217 VPWR.t1023 VPWR.t1664 497.094
R11218 VPWR.t1244 VPWR.t1012 497.094
R11219 VPWR.t1012 VPWR.t1794 497.094
R11220 VPWR.t1402 VPWR.t1011 497.094
R11221 VPWR.t1011 VPWR.t22 497.094
R11222 VPWR.t12 VPWR.t1668 497.094
R11223 VPWR.t1668 VPWR.t1468 497.094
R11224 VPWR.t1287 VPWR.t1043 497.094
R11225 VPWR.t1043 VPWR.t1580 497.094
R11226 VPWR.t1528 VPWR.t1016 497.094
R11227 VPWR.t1016 VPWR.t1516 497.094
R11228 VPWR.t1560 VPWR.t1667 497.094
R11229 VPWR.t1667 VPWR.t1456 497.094
R11230 VPWR.t427 VPWR.t1663 497.094
R11231 VPWR.t1663 VPWR.t1867 497.094
R11232 VPWR.t1863 VPWR.t1313 497.094
R11233 VPWR.t1313 VPWR.t1891 497.094
R11234 VPWR.t238 VPWR.t1015 497.094
R11235 VPWR.t1015 VPWR.t187 497.094
R11236 VPWR.t316 VPWR.t1666 497.094
R11237 VPWR.t1666 VPWR.t98 497.094
R11238 VPWR.t118 VPWR.t1312 497.094
R11239 VPWR.t1312 VPWR.t262 497.094
R11240 VPWR.t567 VPWR.t1014 497.094
R11241 VPWR.t1014 VPWR.t1118 497.094
R11242 VPWR.t1114 VPWR.t1013 497.094
R11243 VPWR.t1013 VPWR.t1650 497.094
R11244 VPWR.t1086 VPWR.t1665 497.094
R11245 VPWR.t1665 VPWR.t469 497.094
R11246 VPWR.t473 VPWR.t1311 497.094
R11247 VPWR.t1311 VPWR.t978 497.094
R11248 VPWR.t823 VPWR.t825 497.094
R11249 VPWR.t1848 VPWR.t823 497.094
R11250 VPWR.t692 VPWR.t613 497.094
R11251 VPWR.t1538 VPWR.t692 497.094
R11252 VPWR.t705 VPWR.t707 497.094
R11253 VPWR.t44 VPWR.t705 497.094
R11254 VPWR.t747 VPWR.t745 497.094
R11255 VPWR.t745 VPWR.t138 497.094
R11256 VPWR.t965 VPWR.t967 497.094
R11257 VPWR.t607 VPWR.t965 497.094
R11258 VPWR.t610 VPWR.t624 497.094
R11259 VPWR.t624 VPWR.t216 497.094
R11260 VPWR.t750 VPWR.t752 497.094
R11261 VPWR.t1624 VPWR.t750 497.094
R11262 VPWR.t865 VPWR.t863 497.094
R11263 VPWR.t863 VPWR.t507 497.094
R11264 VPWR.t884 VPWR.t886 497.094
R11265 VPWR.t1905 VPWR.t884 497.094
R11266 VPWR.t641 VPWR.t639 497.094
R11267 VPWR.t639 VPWR.t298 497.094
R11268 VPWR.t771 VPWR.t769 497.094
R11269 VPWR.t769 VPWR.t78 497.094
R11270 VPWR.t897 VPWR.t892 497.094
R11271 VPWR.t892 VPWR.t1510 497.094
R11272 VPWR.t889 VPWR.t644 497.094
R11273 VPWR.t644 VPWR.t174 497.094
R11274 VPWR.t662 VPWR.t667 497.094
R11275 VPWR.t1072 VPWR.t662 497.094
R11276 VPWR.t809 VPWR.t807 497.094
R11277 VPWR.t807 VPWR.t447 497.094
R11278 VPWR.t921 VPWR.t923 497.094
R11279 VPWR.t915 VPWR.t921 497.094
R11280 VPWR.t780 VPWR.t782 497.094
R11281 VPWR.t777 VPWR.t780 497.094
R11282 VPWR.t637 VPWR.t929 497.094
R11283 VPWR.t634 VPWR.t637 497.094
R11284 VPWR.t651 VPWR.t649 497.094
R11285 VPWR.t649 VPWR.t646 497.094
R11286 VPWR.t687 VPWR.t689 497.094
R11287 VPWR.t684 VPWR.t687 497.094
R11288 VPWR.t907 VPWR.t905 497.094
R11289 VPWR.t905 VPWR.t902 497.094
R11290 VPWR.t944 VPWR.t926 497.094
R11291 VPWR.t941 VPWR.t944 497.094
R11292 VPWR.t699 VPWR.t697 497.094
R11293 VPWR.t697 VPWR.t694 497.094
R11294 VPWR.t793 VPWR.t795 497.094
R11295 VPWR.t812 VPWR.t793 497.094
R11296 VPWR.t831 VPWR.t834 497.094
R11297 VPWR.t834 VPWR.t828 497.094
R11298 VPWR.t970 VPWR.t972 497.094
R11299 VPWR.t676 VPWR.t970 497.094
R11300 VPWR.t715 VPWR.t713 497.094
R11301 VPWR.t713 VPWR.t710 497.094
R11302 VPWR.t848 VPWR.t850 497.094
R11303 VPWR.t842 VPWR.t848 497.094
R11304 VPWR.t881 VPWR.t981 497.094
R11305 VPWR.t981 VPWR.t975 497.094
R11306 VPWR.t619 VPWR.t621 497.094
R11307 VPWR.t616 VPWR.t619 497.094
R11308 VPWR.t760 VPWR.t758 497.094
R11309 VPWR.t758 VPWR.t755 497.094
R11310 VPWR.t868 VPWR.t870 497.094
R11311 VPWR.t839 VPWR.t868 497.094
R11312 VPWR.t657 VPWR.t659 497.094
R11313 VPWR.t654 VPWR.t657 497.094
R11314 VPWR.t801 VPWR.t900 497.094
R11315 VPWR.t900 VPWR.t894 497.094
R11316 VPWR.t918 VPWR.t913 497.094
R11317 VPWR.t913 VPWR.t910 497.094
R11318 VPWR.t954 VPWR.t952 497.094
R11319 VPWR.t952 VPWR.t949 497.094
R11320 VPWR.t790 VPWR.t788 497.094
R11321 VPWR.t788 VPWR.t785 497.094
R11322 VPWR.t798 VPWR.t818 497.094
R11323 VPWR.t818 VPWR.t815 497.094
R11324 VPWR.t962 VPWR.t960 497.094
R11325 VPWR.t960 VPWR.t957 497.094
R11326 VPWR.t681 VPWR.t679 497.094
R11327 VPWR.t679 VPWR.t702 497.094
R11328 VPWR.t723 VPWR.t721 497.094
R11329 VPWR.t721 VPWR.t718 497.094
R11330 VPWR.t855 VPWR.t853 497.094
R11331 VPWR.t853 VPWR.t935 497.094
R11332 VPWR.t991 VPWR.t989 497.094
R11333 VPWR.t989 VPWR.t983 497.094
R11334 VPWR.t731 VPWR.t729 497.094
R11335 VPWR.t729 VPWR.t726 497.094
R11336 VPWR.t763 VPWR.t861 497.094
R11337 VPWR.t861 VPWR.t858 497.094
R11338 VPWR.t878 VPWR.t876 497.094
R11339 VPWR.t876 VPWR.t873 497.094
R11340 VPWR.t631 VPWR.t629 497.094
R11341 VPWR.t629 VPWR.t626 497.094
R11342 VPWR.t740 VPWR.t742 497.094
R11343 VPWR.t737 VPWR.t740 497.094
R11344 VPWR.n2562 VPWR.t124 428.822
R11345 VPWR.n1166 VPWR.n1165 376.045
R11346 VPWR.n2442 VPWR.n2441 376.045
R11347 VPWR.n1451 VPWR.n1450 376.045
R11348 VPWR.n319 VPWR.n318 376.045
R11349 VPWR.n2504 VPWR.n2503 376.045
R11350 VPWR.n1513 VPWR.n1512 376.045
R11351 VPWR.n317 VPWR.n316 376.045
R11352 VPWR.n2444 VPWR.n2443 376.045
R11353 VPWR.n934 VPWR.n933 376.045
R11354 VPWR.n2414 VPWR.n2413 376.045
R11355 VPWR.n2412 VPWR.n2411 376.045
R11356 VPWR.n289 VPWR.n288 376.045
R11357 VPWR.n2490 VPWR.n2489 376.045
R11358 VPWR.n942 VPWR.n941 376.045
R11359 VPWR.n2382 VPWR.n2381 376.045
R11360 VPWR.n293 VPWR.n292 376.045
R11361 VPWR.n2480 VPWR.n2479 376.045
R11362 VPWR.n1826 VPWR.n1825 376.045
R11363 VPWR.n1824 VPWR.n1823 376.045
R11364 VPWR.n1816 VPWR.n1815 376.045
R11365 VPWR.n358 VPWR.n357 376.045
R11366 VPWR.n362 VPWR.n361 376.045
R11367 VPWR.n366 VPWR.n365 376.045
R11368 VPWR.n2392 VPWR.n2391 376.045
R11369 VPWR.n301 VPWR.n300 376.045
R11370 VPWR.n2468 VPWR.n2467 376.045
R11371 VPWR.n1814 VPWR.n1813 376.045
R11372 VPWR.n374 VPWR.n373 376.045
R11373 VPWR.n2394 VPWR.n2393 376.045
R11374 VPWR.n305 VPWR.n304 376.045
R11375 VPWR.n2466 VPWR.n2465 376.045
R11376 VPWR.n2245 VPWR.n2244 376.045
R11377 VPWR.n2247 VPWR.n2246 376.045
R11378 VPWR.n2255 VPWR.n2254 376.045
R11379 VPWR.n2257 VPWR.n2256 376.045
R11380 VPWR.n2267 VPWR.n2266 376.045
R11381 VPWR.n2275 VPWR.n2274 376.045
R11382 VPWR.n2277 VPWR.n2276 376.045
R11383 VPWR.n2285 VPWR.n2284 376.045
R11384 VPWR.n2287 VPWR.n2286 376.045
R11385 VPWR.n2295 VPWR.n2294 376.045
R11386 VPWR.n2297 VPWR.n2296 376.045
R11387 VPWR.n2305 VPWR.n2304 376.045
R11388 VPWR.n2307 VPWR.n2306 376.045
R11389 VPWR.n2315 VPWR.n2314 376.045
R11390 VPWR.n2265 VPWR.n2264 376.045
R11391 VPWR.n511 VPWR.n510 376.045
R11392 VPWR.n509 VPWR.n508 376.045
R11393 VPWR.n505 VPWR.n504 376.045
R11394 VPWR.n501 VPWR.n500 376.045
R11395 VPWR.n493 VPWR.n492 376.045
R11396 VPWR.n489 VPWR.n488 376.045
R11397 VPWR.n485 VPWR.n484 376.045
R11398 VPWR.n481 VPWR.n480 376.045
R11399 VPWR.n477 VPWR.n476 376.045
R11400 VPWR.n473 VPWR.n472 376.045
R11401 VPWR.n469 VPWR.n468 376.045
R11402 VPWR.n465 VPWR.n464 376.045
R11403 VPWR.n461 VPWR.n460 376.045
R11404 VPWR.n457 VPWR.n456 376.045
R11405 VPWR.n497 VPWR.n496 376.045
R11406 VPWR.n2218 VPWR.n2217 376.045
R11407 VPWR.n2216 VPWR.n2215 376.045
R11408 VPWR.n2208 VPWR.n2207 376.045
R11409 VPWR.n2206 VPWR.n2205 376.045
R11410 VPWR.n2196 VPWR.n2195 376.045
R11411 VPWR.n2188 VPWR.n2187 376.045
R11412 VPWR.n2186 VPWR.n2185 376.045
R11413 VPWR.n2178 VPWR.n2177 376.045
R11414 VPWR.n2176 VPWR.n2175 376.045
R11415 VPWR.n2168 VPWR.n2167 376.045
R11416 VPWR.n2166 VPWR.n2165 376.045
R11417 VPWR.n2158 VPWR.n2157 376.045
R11418 VPWR.n2156 VPWR.n2155 376.045
R11419 VPWR.n2148 VPWR.n2147 376.045
R11420 VPWR.n2198 VPWR.n2197 376.045
R11421 VPWR.n550 VPWR.n549 376.045
R11422 VPWR.n554 VPWR.n553 376.045
R11423 VPWR.n558 VPWR.n557 376.045
R11424 VPWR.n562 VPWR.n561 376.045
R11425 VPWR.n570 VPWR.n569 376.045
R11426 VPWR.n574 VPWR.n573 376.045
R11427 VPWR.n578 VPWR.n577 376.045
R11428 VPWR.n582 VPWR.n581 376.045
R11429 VPWR.n586 VPWR.n585 376.045
R11430 VPWR.n590 VPWR.n589 376.045
R11431 VPWR.n594 VPWR.n593 376.045
R11432 VPWR.n598 VPWR.n597 376.045
R11433 VPWR.n602 VPWR.n601 376.045
R11434 VPWR.n606 VPWR.n605 376.045
R11435 VPWR.n566 VPWR.n565 376.045
R11436 VPWR.n2049 VPWR.n2048 376.045
R11437 VPWR.n2051 VPWR.n2050 376.045
R11438 VPWR.n2059 VPWR.n2058 376.045
R11439 VPWR.n2061 VPWR.n2060 376.045
R11440 VPWR.n2071 VPWR.n2070 376.045
R11441 VPWR.n2079 VPWR.n2078 376.045
R11442 VPWR.n2081 VPWR.n2080 376.045
R11443 VPWR.n2089 VPWR.n2088 376.045
R11444 VPWR.n2091 VPWR.n2090 376.045
R11445 VPWR.n2099 VPWR.n2098 376.045
R11446 VPWR.n2101 VPWR.n2100 376.045
R11447 VPWR.n2109 VPWR.n2108 376.045
R11448 VPWR.n2111 VPWR.n2110 376.045
R11449 VPWR.n2119 VPWR.n2118 376.045
R11450 VPWR.n2069 VPWR.n2068 376.045
R11451 VPWR.n703 VPWR.n702 376.045
R11452 VPWR.n701 VPWR.n700 376.045
R11453 VPWR.n697 VPWR.n696 376.045
R11454 VPWR.n693 VPWR.n692 376.045
R11455 VPWR.n685 VPWR.n684 376.045
R11456 VPWR.n681 VPWR.n680 376.045
R11457 VPWR.n677 VPWR.n676 376.045
R11458 VPWR.n673 VPWR.n672 376.045
R11459 VPWR.n669 VPWR.n668 376.045
R11460 VPWR.n665 VPWR.n664 376.045
R11461 VPWR.n661 VPWR.n660 376.045
R11462 VPWR.n657 VPWR.n656 376.045
R11463 VPWR.n653 VPWR.n652 376.045
R11464 VPWR.n649 VPWR.n648 376.045
R11465 VPWR.n689 VPWR.n688 376.045
R11466 VPWR.n2022 VPWR.n2021 376.045
R11467 VPWR.n2020 VPWR.n2019 376.045
R11468 VPWR.n2012 VPWR.n2011 376.045
R11469 VPWR.n2010 VPWR.n2009 376.045
R11470 VPWR.n2000 VPWR.n1999 376.045
R11471 VPWR.n1992 VPWR.n1991 376.045
R11472 VPWR.n1990 VPWR.n1989 376.045
R11473 VPWR.n1982 VPWR.n1981 376.045
R11474 VPWR.n1980 VPWR.n1979 376.045
R11475 VPWR.n1972 VPWR.n1971 376.045
R11476 VPWR.n1970 VPWR.n1969 376.045
R11477 VPWR.n1962 VPWR.n1961 376.045
R11478 VPWR.n1960 VPWR.n1959 376.045
R11479 VPWR.n1952 VPWR.n1951 376.045
R11480 VPWR.n2002 VPWR.n2001 376.045
R11481 VPWR.n742 VPWR.n741 376.045
R11482 VPWR.n746 VPWR.n745 376.045
R11483 VPWR.n750 VPWR.n749 376.045
R11484 VPWR.n754 VPWR.n753 376.045
R11485 VPWR.n762 VPWR.n761 376.045
R11486 VPWR.n766 VPWR.n765 376.045
R11487 VPWR.n770 VPWR.n769 376.045
R11488 VPWR.n774 VPWR.n773 376.045
R11489 VPWR.n778 VPWR.n777 376.045
R11490 VPWR.n782 VPWR.n781 376.045
R11491 VPWR.n786 VPWR.n785 376.045
R11492 VPWR.n790 VPWR.n789 376.045
R11493 VPWR.n794 VPWR.n793 376.045
R11494 VPWR.n798 VPWR.n797 376.045
R11495 VPWR.n758 VPWR.n757 376.045
R11496 VPWR.n1853 VPWR.n1852 376.045
R11497 VPWR.n1855 VPWR.n1854 376.045
R11498 VPWR.n1863 VPWR.n1862 376.045
R11499 VPWR.n1865 VPWR.n1864 376.045
R11500 VPWR.n1875 VPWR.n1874 376.045
R11501 VPWR.n1883 VPWR.n1882 376.045
R11502 VPWR.n1885 VPWR.n1884 376.045
R11503 VPWR.n1893 VPWR.n1892 376.045
R11504 VPWR.n1895 VPWR.n1894 376.045
R11505 VPWR.n1903 VPWR.n1902 376.045
R11506 VPWR.n1905 VPWR.n1904 376.045
R11507 VPWR.n1913 VPWR.n1912 376.045
R11508 VPWR.n1915 VPWR.n1914 376.045
R11509 VPWR.n1923 VPWR.n1922 376.045
R11510 VPWR.n1873 VPWR.n1872 376.045
R11511 VPWR.n895 VPWR.n894 376.045
R11512 VPWR.n893 VPWR.n892 376.045
R11513 VPWR.n889 VPWR.n888 376.045
R11514 VPWR.n885 VPWR.n884 376.045
R11515 VPWR.n877 VPWR.n876 376.045
R11516 VPWR.n873 VPWR.n872 376.045
R11517 VPWR.n869 VPWR.n868 376.045
R11518 VPWR.n865 VPWR.n864 376.045
R11519 VPWR.n861 VPWR.n860 376.045
R11520 VPWR.n857 VPWR.n856 376.045
R11521 VPWR.n853 VPWR.n852 376.045
R11522 VPWR.n849 VPWR.n848 376.045
R11523 VPWR.n845 VPWR.n844 376.045
R11524 VPWR.n841 VPWR.n840 376.045
R11525 VPWR.n881 VPWR.n880 376.045
R11526 VPWR.n1806 VPWR.n1805 376.045
R11527 VPWR.n950 VPWR.n949 376.045
R11528 VPWR.n1472 VPWR.n1471 376.045
R11529 VPWR.n1152 VPWR.n1151 376.045
R11530 VPWR.n370 VPWR.n369 376.045
R11531 VPWR.n2402 VPWR.n2401 376.045
R11532 VPWR.n309 VPWR.n308 376.045
R11533 VPWR.n2456 VPWR.n2455 376.045
R11534 VPWR.n946 VPWR.n945 376.045
R11535 VPWR.n1470 VPWR.n1469 376.045
R11536 VPWR.n1156 VPWR.n1155 376.045
R11537 VPWR.n1804 VPWR.n1803 376.045
R11538 VPWR.n954 VPWR.n953 376.045
R11539 VPWR.n1484 VPWR.n1483 376.045
R11540 VPWR.n1148 VPWR.n1147 376.045
R11541 VPWR.n378 VPWR.n377 376.045
R11542 VPWR.n386 VPWR.n385 376.045
R11543 VPWR.n390 VPWR.n389 376.045
R11544 VPWR.n394 VPWR.n393 376.045
R11545 VPWR.n398 VPWR.n397 376.045
R11546 VPWR.n402 VPWR.n401 376.045
R11547 VPWR.n406 VPWR.n405 376.045
R11548 VPWR.n410 VPWR.n409 376.045
R11549 VPWR.n414 VPWR.n413 376.045
R11550 VPWR.n382 VPWR.n381 376.045
R11551 VPWR.n2384 VPWR.n2383 376.045
R11552 VPWR.n297 VPWR.n296 376.045
R11553 VPWR.n2478 VPWR.n2477 376.045
R11554 VPWR.n958 VPWR.n957 376.045
R11555 VPWR.n1486 VPWR.n1485 376.045
R11556 VPWR.n1144 VPWR.n1143 376.045
R11557 VPWR.n1796 VPWR.n1795 376.045
R11558 VPWR.n1786 VPWR.n1785 376.045
R11559 VPWR.n1784 VPWR.n1783 376.045
R11560 VPWR.n1776 VPWR.n1775 376.045
R11561 VPWR.n1774 VPWR.n1773 376.045
R11562 VPWR.n1766 VPWR.n1765 376.045
R11563 VPWR.n1764 VPWR.n1763 376.045
R11564 VPWR.n1756 VPWR.n1755 376.045
R11565 VPWR.n1794 VPWR.n1793 376.045
R11566 VPWR.n962 VPWR.n961 376.045
R11567 VPWR.n1498 VPWR.n1497 376.045
R11568 VPWR.n1140 VPWR.n1139 376.045
R11569 VPWR.n2404 VPWR.n2403 376.045
R11570 VPWR.n313 VPWR.n312 376.045
R11571 VPWR.n2454 VPWR.n2453 376.045
R11572 VPWR.n1459 VPWR.n1458 376.045
R11573 VPWR.n1160 VPWR.n1159 376.045
R11574 VPWR.n966 VPWR.n965 376.045
R11575 VPWR.n1500 VPWR.n1499 376.045
R11576 VPWR.n1136 VPWR.n1135 376.045
R11577 VPWR.n2374 VPWR.n2373 376.045
R11578 VPWR.n2364 VPWR.n2363 376.045
R11579 VPWR.n2362 VPWR.n2361 376.045
R11580 VPWR.n2354 VPWR.n2353 376.045
R11581 VPWR.n2352 VPWR.n2351 376.045
R11582 VPWR.n2344 VPWR.n2343 376.045
R11583 VPWR.n2372 VPWR.n2371 376.045
R11584 VPWR.n285 VPWR.n284 376.045
R11585 VPWR.n2492 VPWR.n2491 376.045
R11586 VPWR.n1515 VPWR.n1514 376.045
R11587 VPWR.n1132 VPWR.n1131 376.045
R11588 VPWR.n970 VPWR.n969 376.045
R11589 VPWR.n974 VPWR.n973 376.045
R11590 VPWR.n978 VPWR.n977 376.045
R11591 VPWR.n982 VPWR.n981 376.045
R11592 VPWR.n986 VPWR.n985 376.045
R11593 VPWR.n990 VPWR.n989 376.045
R11594 VPWR.n938 VPWR.n937 376.045
R11595 VPWR.n1457 VPWR.n1456 376.045
R11596 VPWR.n1164 VPWR.n1163 376.045
R11597 VPWR.n281 VPWR.n280 376.045
R11598 VPWR.n2502 VPWR.n2501 376.045
R11599 VPWR.n1128 VPWR.n1127 376.045
R11600 VPWR.n1698 VPWR.n1697 376.045
R11601 VPWR.n1124 VPWR.n1123 376.045
R11602 VPWR.n277 VPWR.n276 376.045
R11603 VPWR.n273 VPWR.n272 376.045
R11604 VPWR.n265 VPWR.n264 376.045
R11605 VPWR.n269 VPWR.n268 376.045
R11606 VPWR.n1677 VPWR.n1676 376.045
R11607 VPWR.n1686 VPWR.n1685 376.045
R11608 VPWR.n1727 VPWR.n1726 376.045
R11609 VPWR.n1696 VPWR.n1695 376.045
R11610 VPWR.n1120 VPWR.n1119 376.045
R11611 VPWR.n2514 VPWR.n2513 376.045
R11612 VPWR.n2516 VPWR.n2515 376.045
R11613 VPWR.n2526 VPWR.n2525 376.045
R11614 VPWR.n1675 VPWR.n1674 376.045
R11615 VPWR.n1278 VPWR.t606 342.841
R11616 VPWR.n1317 VPWR.t412 342.841
R11617 VPWR.n1354 VPWR.t54 342.841
R11618 VPWR.n2629 VPWR.t1914 342.841
R11619 VPWR.n2592 VPWR.t1190 342.841
R11620 VPWR.n2535 VPWR.t125 342.841
R11621 VPWR.n1278 VPWR.t206 342.839
R11622 VPWR.n1317 VPWR.t1822 342.839
R11623 VPWR.n1354 VPWR.t1316 342.839
R11624 VPWR.n2629 VPWR.t1637 342.839
R11625 VPWR.n2592 VPWR.t1618 342.839
R11626 VPWR.n2535 VPWR.t1870 342.839
R11627 VPWR.n2778 VPWR.n2760 339.212
R11628 VPWR.n1245 VPWR.t1448 338.488
R11629 VPWR.n2665 VPWR.t393 338.488
R11630 VPWR.n1254 VPWR.n1253 327.377
R11631 VPWR.n1247 VPWR.n1246 327.377
R11632 VPWR.n1261 VPWR.n1260 327.377
R11633 VPWR.n1291 VPWR.n1289 327.377
R11634 VPWR.n1284 VPWR.n1282 327.377
R11635 VPWR.n1299 VPWR.n1297 327.377
R11636 VPWR.n1330 VPWR.n1328 327.377
R11637 VPWR.n1323 VPWR.n1321 327.377
R11638 VPWR.n1338 VPWR.n1336 327.377
R11639 VPWR.n1367 VPWR.n1365 327.377
R11640 VPWR.n1360 VPWR.n1358 327.377
R11641 VPWR.n1375 VPWR.n1373 327.377
R11642 VPWR.n1263 VPWR.n1262 327.375
R11643 VPWR.n1291 VPWR.n1290 327.375
R11644 VPWR.n1284 VPWR.n1283 327.375
R11645 VPWR.n1299 VPWR.n1298 327.375
R11646 VPWR.n1330 VPWR.n1329 327.375
R11647 VPWR.n1323 VPWR.n1322 327.375
R11648 VPWR.n1338 VPWR.n1337 327.375
R11649 VPWR.n1367 VPWR.n1366 327.375
R11650 VPWR.n1360 VPWR.n1359 327.375
R11651 VPWR.n1375 VPWR.n1374 327.375
R11652 VPWR.n1 VPWR 325.546
R11653 VPWR.n2603 VPWR.t1636 322.262
R11654 VPWR.n2566 VPWR.t1189 322.262
R11655 VPWR.n2741 VPWR.n2740 321.642
R11656 VPWR.n2658 VPWR.n2648 320.976
R11657 VPWR.n2652 VPWR.n2651 320.976
R11658 VPWR.n2646 VPWR.n2645 320.976
R11659 VPWR.n2616 VPWR.n2615 320.976
R11660 VPWR.n2622 VPWR.n2611 320.976
R11661 VPWR.n2608 VPWR.n2607 320.976
R11662 VPWR.n2579 VPWR.n2578 320.976
R11663 VPWR.n2585 VPWR.n2574 320.976
R11664 VPWR.n2571 VPWR.n2570 320.976
R11665 VPWR.n2546 VPWR.n2542 320.976
R11666 VPWR.n2550 VPWR.n2549 320.976
R11667 VPWR.n2556 VPWR.n2538 320.976
R11668 VPWR.n2663 VPWR.n2644 320.976
R11669 VPWR.n2616 VPWR.n2614 320.976
R11670 VPWR.n2622 VPWR.n2610 320.976
R11671 VPWR.n2608 VPWR.n2606 320.976
R11672 VPWR.n2579 VPWR.n2577 320.976
R11673 VPWR.n2585 VPWR.n2573 320.976
R11674 VPWR.n2571 VPWR.n2569 320.976
R11675 VPWR.n2546 VPWR.n2541 320.976
R11676 VPWR.n2550 VPWR.n2548 320.976
R11677 VPWR.n2556 VPWR.n2537 320.976
R11678 VPWR.n2737 VPWR 319.627
R11679 VPWR.n6 VPWR.n5 316.245
R11680 VPWR.n1180 VPWR.n1178 316.245
R11681 VPWR.n1203 VPWR.n1201 316.245
R11682 VPWR.n1227 VPWR.n1225 316.245
R11683 VPWR.n2720 VPWR.n2719 316.245
R11684 VPWR.n2700 VPWR.n2699 316.245
R11685 VPWR.n2681 VPWR.n2680 316.245
R11686 VPWR.n1180 VPWR.n1179 316.245
R11687 VPWR.n1203 VPWR.n1202 316.245
R11688 VPWR.n1227 VPWR.n1226 316.245
R11689 VPWR.n2720 VPWR.n2718 316.245
R11690 VPWR.n2700 VPWR.n2698 316.245
R11691 VPWR.n2681 VPWR.n2679 316.245
R11692 VPWR.n2566 VPWR.t1096 313.87
R11693 VPWR.n10 VPWR.n4 310.502
R11694 VPWR.n1185 VPWR.n1177 310.502
R11695 VPWR.n1208 VPWR.n1200 310.502
R11696 VPWR.n1232 VPWR.n1224 310.502
R11697 VPWR.n2739 VPWR.n2738 310.502
R11698 VPWR.n2724 VPWR.n2723 310.502
R11699 VPWR.n2704 VPWR.n2703 310.502
R11700 VPWR.n2685 VPWR.n2684 310.502
R11701 VPWR.n1185 VPWR.n1184 310.5
R11702 VPWR.n1208 VPWR.n1207 310.5
R11703 VPWR.n1232 VPWR.n1231 310.5
R11704 VPWR.n2724 VPWR.n2722 310.5
R11705 VPWR.n2704 VPWR.n2702 310.5
R11706 VPWR.n2685 VPWR.n2683 310.5
R11707 VPWR.n2770 VPWR.n2769 279.341
R11708 VPWR.n2775 VPWR.n2774 279.341
R11709 VPWR.n1351 VPWR.t1630 255.905
R11710 VPWR.n2599 VPWR.t1097 255.905
R11711 VPWR.n1214 VPWR.t1352 255.904
R11712 VPWR.n1351 VPWR.t1858 255.904
R11713 VPWR.n2710 VPWR.t1133 255.904
R11714 VPWR.n2599 VPWR.t1631 255.904
R11715 VPWR.n1242 VPWR.t198 254.019
R11716 VPWR.n2671 VPWR.t534 254.019
R11717 VPWR.n1274 VPWR.t196 252.948
R11718 VPWR.n2673 VPWR.t532 252.948
R11719 VPWR.n1312 VPWR.t1055 250.722
R11720 VPWR.n2636 VPWR.t275 250.722
R11721 VPWR.n1249 VPWR.t10 249.901
R11722 VPWR.n1285 VPWR.t1002 249.901
R11723 VPWR.n1324 VPWR.t1784 249.901
R11724 VPWR.n1361 VPWR.t1004 249.901
R11725 VPWR.n2650 VPWR.t1767 249.901
R11726 VPWR.n2613 VPWR.t1764 249.901
R11727 VPWR.n2576 VPWR.t1778 249.901
R11728 VPWR.n2543 VPWR.t1732 249.901
R11729 VPWR.n1285 VPWR.t1836 249.901
R11730 VPWR.n1324 VPWR.t163 249.901
R11731 VPWR.n1361 VPWR.t1699 249.901
R11732 VPWR.n2613 VPWR.t1777 249.901
R11733 VPWR.n2576 VPWR.t1730 249.901
R11734 VPWR.n2543 VPWR.t1753 249.901
R11735 VPWR.n1192 VPWR.t1804 249.363
R11736 VPWR.n1277 VPWR.t485 249.363
R11737 VPWR.n2747 VPWR.t33 249.363
R11738 VPWR.n2731 VPWR.t1460 249.363
R11739 VPWR.n2634 VPWR.t1301 249.363
R11740 VPWR.n17 VPWR.t182 249.362
R11741 VPWR.n1192 VPWR.t453 249.362
R11742 VPWR.n2731 VPWR.t558 249.362
R11743 VPWR.t1348 VPWR.t181 248.599
R11744 VPWR.t407 VPWR.t1852 248.599
R11745 VPWR.t1852 VPWR.t1856 248.599
R11746 VPWR.t1856 VPWR.t403 248.599
R11747 VPWR.t403 VPWR.t346 248.599
R11748 VPWR.t346 VPWR.t0 248.599
R11749 VPWR.t0 VPWR.t1001 248.599
R11750 VPWR.t1001 VPWR.t1007 248.599
R11751 VPWR.t1832 VPWR.t1834 248.599
R11752 VPWR.t1834 VPWR.t9 248.599
R11753 VPWR.t1780 VPWR.t1756 248.599
R11754 VPWR.t1744 VPWR.t1780 248.599
R11755 VPWR.t1718 VPWR.t1744 248.599
R11756 VPWR.t390 VPWR.t1718 248.599
R11757 VPWR.t573 VPWR.t390 248.599
R11758 VPWR.t1154 VPWR.t573 248.599
R11759 VPWR.t1152 VPWR.t1154 248.599
R11760 VPWR.t1134 VPWR.t32 248.599
R11761 VPWR.t1724 VPWR.t1766 248.599
R11762 VPWR.t1772 VPWR.t1724 248.599
R11763 VPWR.n15 VPWR.t1349 247.394
R11764 VPWR.n1190 VPWR.t1351 247.394
R11765 VPWR.n2745 VPWR.t1135 247.394
R11766 VPWR.n2729 VPWR.t1129 247.394
R11767 VPWR.n1190 VPWR.t1350 247.394
R11768 VPWR.n2729 VPWR.t1131 247.394
R11769 VPWR.n1243 VPWR.t155 244.737
R11770 VPWR.n2666 VPWR.t1782 244.737
R11771 VPWR.n1313 VPWR.t1050 243.886
R11772 VPWR.n2637 VPWR.t1197 243.886
R11773 VPWR.n1216 VPWR.t180 243.512
R11774 VPWR.n1239 VPWR.t1805 243.512
R11775 VPWR.n1242 VPWR.t487 243.512
R11776 VPWR.n2712 VPWR.t35 243.512
R11777 VPWR.n2692 VPWR.t1461 243.512
R11778 VPWR.n2671 VPWR.t1127 243.512
R11779 VPWR.n1239 VPWR.t454 243.512
R11780 VPWR.n2692 VPWR.t556 243.512
R11781 VPWR.n1268 VPWR.t197 238.339
R11782 VPWR.n2641 VPWR.t533 238.339
R11783 VPWR.n2791 VPWR.t399 237.99
R11784 VPWR.n2603 VPWR.t1300 234.982
R11785 VPWR.t1830 VPWR.t1832 228.101
R11786 VPWR.t1750 VPWR.t1772 228.101
R11787 VPWR.n2737 VPWR 224.923
R11788 VPWR.n1 VPWR 219.004
R11789 VPWR.n1383 VPWR.n1382 214.613
R11790 VPWR.n1383 VPWR.n1381 214.613
R11791 VPWR.n1175 VPWR.n1174 214.326
R11792 VPWR.n1198 VPWR.n1197 214.326
R11793 VPWR.n1222 VPWR.n1221 214.326
R11794 VPWR.n1307 VPWR.n1306 214.326
R11795 VPWR.n1346 VPWR.n1345 214.326
R11796 VPWR.n1175 VPWR.n1173 214.326
R11797 VPWR.n1198 VPWR.n1196 214.326
R11798 VPWR.n1222 VPWR.n1220 214.326
R11799 VPWR.n1307 VPWR.n1305 214.326
R11800 VPWR.n1346 VPWR.n1344 214.326
R11801 VPWR.n2 VPWR.n1 213.119
R11802 VPWR.n2744 VPWR.n2737 213.119
R11803 VPWR VPWR.t1348 207.166
R11804 VPWR.n2776 VPWR.n2775 204.424
R11805 VPWR.n2766 VPWR.n2753 204.424
R11806 VPWR.n2769 VPWR.n2756 204.424
R11807 VPWR.n2780 VPWR.n2777 204.048
R11808 VPWR VPWR.t1152 201.246
R11809 VPWR.t9 VPWR 189.409
R11810 VPWR.n2677 VPWR 184.63
R11811 VPWR.n1268 VPWR 182.952
R11812 VPWR.n2696 VPWR 182.952
R11813 VPWR.n2716 VPWR 181.273
R11814 VPWR.t1096 VPWR 177.916
R11815 VPWR.n2784 VPWR.n2783 166.4
R11816 VPWR.n1706 VPWR.n1704 161.365
R11817 VPWR.n1009 VPWR.n1007 161.365
R11818 VPWR.n1523 VPWR.n1521 161.365
R11819 VPWR.n1528 VPWR.n1526 161.365
R11820 VPWR.n1533 VPWR.n1531 161.365
R11821 VPWR.n1538 VPWR.n1536 161.365
R11822 VPWR.n1543 VPWR.n1541 161.365
R11823 VPWR.n1548 VPWR.n1546 161.365
R11824 VPWR.n1553 VPWR.n1551 161.365
R11825 VPWR.n1558 VPWR.n1556 161.365
R11826 VPWR.n1563 VPWR.n1561 161.365
R11827 VPWR.n1398 VPWR.n1396 161.365
R11828 VPWR.n1393 VPWR.n1391 161.365
R11829 VPWR.n1711 VPWR.n1709 161.365
R11830 VPWR.n1719 VPWR.n1717 161.365
R11831 VPWR.n1715 VPWR.n1713 161.365
R11832 VPWR VPWR.n1075 161.363
R11833 VPWR VPWR.n103 161.363
R11834 VPWR VPWR.n53 161.363
R11835 VPWR VPWR.n51 161.363
R11836 VPWR VPWR.n49 161.363
R11837 VPWR VPWR.n47 161.363
R11838 VPWR VPWR.n45 161.363
R11839 VPWR VPWR.n43 161.363
R11840 VPWR VPWR.n41 161.363
R11841 VPWR VPWR.n39 161.363
R11842 VPWR VPWR.n37 161.363
R11843 VPWR VPWR.n35 161.363
R11844 VPWR VPWR.n33 161.363
R11845 VPWR VPWR.n31 161.363
R11846 VPWR VPWR.n29 161.363
R11847 VPWR VPWR.n27 161.363
R11848 VPWR VPWR.n25 161.363
R11849 VPWR VPWR.n23 161.363
R11850 VPWR.n1115 VPWR.n1114 161.3
R11851 VPWR.n1576 VPWR.n1575 161.3
R11852 VPWR.n1074 VPWR.n1073 161.3
R11853 VPWR.n1579 VPWR.n1578 161.3
R11854 VPWR.n1582 VPWR.n1581 161.3
R11855 VPWR.n1071 VPWR.n1070 161.3
R11856 VPWR.n1585 VPWR.n1584 161.3
R11857 VPWR.n1588 VPWR.n1587 161.3
R11858 VPWR.n1068 VPWR.n1067 161.3
R11859 VPWR.n1591 VPWR.n1590 161.3
R11860 VPWR.n1594 VPWR.n1593 161.3
R11861 VPWR.n1065 VPWR.n1064 161.3
R11862 VPWR.n1597 VPWR.n1596 161.3
R11863 VPWR.n1600 VPWR.n1599 161.3
R11864 VPWR.n1062 VPWR.n1061 161.3
R11865 VPWR.n1603 VPWR.n1602 161.3
R11866 VPWR.n1606 VPWR.n1605 161.3
R11867 VPWR.n1059 VPWR.n1058 161.3
R11868 VPWR.n1609 VPWR.n1608 161.3
R11869 VPWR.n1612 VPWR.n1611 161.3
R11870 VPWR.n1056 VPWR.n1055 161.3
R11871 VPWR.n1615 VPWR.n1614 161.3
R11872 VPWR.n1618 VPWR.n1617 161.3
R11873 VPWR.n1053 VPWR.n1052 161.3
R11874 VPWR.n1621 VPWR.n1620 161.3
R11875 VPWR.n1624 VPWR.n1623 161.3
R11876 VPWR.n1050 VPWR.n1049 161.3
R11877 VPWR.n1627 VPWR.n1626 161.3
R11878 VPWR.n1630 VPWR.n1629 161.3
R11879 VPWR.n1047 VPWR.n1046 161.3
R11880 VPWR.n1633 VPWR.n1632 161.3
R11881 VPWR.n1636 VPWR.n1635 161.3
R11882 VPWR.n1044 VPWR.n1043 161.3
R11883 VPWR.n1639 VPWR.n1638 161.3
R11884 VPWR.n1642 VPWR.n1641 161.3
R11885 VPWR.n1041 VPWR.n1040 161.3
R11886 VPWR.n1645 VPWR.n1644 161.3
R11887 VPWR.n1648 VPWR.n1647 161.3
R11888 VPWR.n1651 VPWR.n1650 161.3
R11889 VPWR.n1037 VPWR.n1036 161.3
R11890 VPWR.n1658 VPWR.n1657 161.3
R11891 VPWR.n1661 VPWR.n1660 161.3
R11892 VPWR.n1656 VPWR.n1655 161.3
R11893 VPWR.n1670 VPWR.n1669 161.3
R11894 VPWR.n1112 VPWR.n1111 161.3
R11895 VPWR.n1667 VPWR.n1666 161.3
R11896 VPWR.n1033 VPWR.n1032 161.3
R11897 VPWR.n121 VPWR.n120 161.3
R11898 VPWR.n114 VPWR.n113 161.3
R11899 VPWR.n117 VPWR.n116 161.3
R11900 VPWR.n112 VPWR.n111 161.3
R11901 VPWR.n131 VPWR.n130 161.3
R11902 VPWR.n123 VPWR.n122 161.3
R11903 VPWR.n108 VPWR.n107 161.3
R11904 VPWR.n105 VPWR.n104 161.3
R11905 VPWR.n256 VPWR.n255 161.3
R11906 VPWR.n253 VPWR.n252 161.3
R11907 VPWR.n101 VPWR.n100 161.3
R11908 VPWR.n243 VPWR.n242 161.3
R11909 VPWR.n246 VPWR.n245 161.3
R11910 VPWR.n241 VPWR.n240 161.3
R11911 VPWR.n233 VPWR.n232 161.3
R11912 VPWR.n236 VPWR.n235 161.3
R11913 VPWR.n231 VPWR.n230 161.3
R11914 VPWR.n223 VPWR.n222 161.3
R11915 VPWR.n226 VPWR.n225 161.3
R11916 VPWR.n221 VPWR.n220 161.3
R11917 VPWR.n213 VPWR.n212 161.3
R11918 VPWR.n216 VPWR.n215 161.3
R11919 VPWR.n211 VPWR.n210 161.3
R11920 VPWR.n203 VPWR.n202 161.3
R11921 VPWR.n206 VPWR.n205 161.3
R11922 VPWR.n201 VPWR.n200 161.3
R11923 VPWR.n193 VPWR.n192 161.3
R11924 VPWR.n196 VPWR.n195 161.3
R11925 VPWR.n191 VPWR.n190 161.3
R11926 VPWR.n183 VPWR.n182 161.3
R11927 VPWR.n186 VPWR.n185 161.3
R11928 VPWR.n181 VPWR.n180 161.3
R11929 VPWR.n173 VPWR.n172 161.3
R11930 VPWR.n176 VPWR.n175 161.3
R11931 VPWR.n171 VPWR.n170 161.3
R11932 VPWR.n163 VPWR.n162 161.3
R11933 VPWR.n166 VPWR.n165 161.3
R11934 VPWR.n161 VPWR.n160 161.3
R11935 VPWR.n153 VPWR.n152 161.3
R11936 VPWR.n156 VPWR.n155 161.3
R11937 VPWR.n151 VPWR.n150 161.3
R11938 VPWR.n143 VPWR.n142 161.3
R11939 VPWR.n146 VPWR.n145 161.3
R11940 VPWR.n141 VPWR.n140 161.3
R11941 VPWR.n133 VPWR.n132 161.3
R11942 VPWR.n136 VPWR.n135 161.3
R11943 VPWR.n126 VPWR.n125 161.3
R11944 VPWR.n1114 VPWR.t653 161.106
R11945 VPWR.n1575 VPWR.t800 161.106
R11946 VPWR.n1073 VPWR.t899 161.106
R11947 VPWR.n1578 VPWR.t893 161.106
R11948 VPWR.n1581 VPWR.t917 161.106
R11949 VPWR.n1070 VPWR.t912 161.106
R11950 VPWR.n1584 VPWR.t909 161.106
R11951 VPWR.n1587 VPWR.t953 161.106
R11952 VPWR.n1067 VPWR.t951 161.106
R11953 VPWR.n1590 VPWR.t948 161.106
R11954 VPWR.n1593 VPWR.t789 161.106
R11955 VPWR.n1064 VPWR.t787 161.106
R11956 VPWR.n1596 VPWR.t784 161.106
R11957 VPWR.n1599 VPWR.t797 161.106
R11958 VPWR.n1061 VPWR.t817 161.106
R11959 VPWR.n1602 VPWR.t814 161.106
R11960 VPWR.n1605 VPWR.t961 161.106
R11961 VPWR.n1058 VPWR.t959 161.106
R11962 VPWR.n1608 VPWR.t956 161.106
R11963 VPWR.n1611 VPWR.t680 161.106
R11964 VPWR.n1055 VPWR.t678 161.106
R11965 VPWR.n1614 VPWR.t701 161.106
R11966 VPWR.n1617 VPWR.t722 161.106
R11967 VPWR.n1052 VPWR.t720 161.106
R11968 VPWR.n1620 VPWR.t717 161.106
R11969 VPWR.n1623 VPWR.t854 161.106
R11970 VPWR.n1049 VPWR.t852 161.106
R11971 VPWR.n1626 VPWR.t934 161.106
R11972 VPWR.n1629 VPWR.t990 161.106
R11973 VPWR.n1046 VPWR.t988 161.106
R11974 VPWR.n1632 VPWR.t982 161.106
R11975 VPWR.n1635 VPWR.t730 161.106
R11976 VPWR.n1043 VPWR.t728 161.106
R11977 VPWR.n1638 VPWR.t725 161.106
R11978 VPWR.n1641 VPWR.t762 161.106
R11979 VPWR.n1040 VPWR.t860 161.106
R11980 VPWR.n1644 VPWR.t857 161.106
R11981 VPWR.n1647 VPWR.t877 161.106
R11982 VPWR.n1650 VPWR.t875 161.106
R11983 VPWR.n1036 VPWR.t872 161.106
R11984 VPWR.n1657 VPWR.t630 161.106
R11985 VPWR.n1660 VPWR.t628 161.106
R11986 VPWR.n1655 VPWR.t625 161.106
R11987 VPWR.n1669 VPWR.t741 161.106
R11988 VPWR.n1111 VPWR.t656 161.106
R11989 VPWR.n1075 VPWR.t658 161.106
R11990 VPWR.n1666 VPWR.t739 161.106
R11991 VPWR.n1032 VPWR.t736 161.106
R11992 VPWR.n120 VPWR.t754 161.106
R11993 VPWR.n113 VPWR.t869 161.106
R11994 VPWR.n116 VPWR.t867 161.106
R11995 VPWR.n111 VPWR.t838 161.106
R11996 VPWR.n130 VPWR.t615 161.106
R11997 VPWR.n122 VPWR.t759 161.106
R11998 VPWR.n107 VPWR.t779 161.106
R11999 VPWR.n103 VPWR.t781 161.106
R12000 VPWR.n104 VPWR.t776 161.106
R12001 VPWR.n255 VPWR.t928 161.106
R12002 VPWR.n252 VPWR.t636 161.106
R12003 VPWR.n100 VPWR.t633 161.106
R12004 VPWR.n242 VPWR.t650 161.106
R12005 VPWR.n245 VPWR.t648 161.106
R12006 VPWR.n240 VPWR.t645 161.106
R12007 VPWR.n232 VPWR.t688 161.106
R12008 VPWR.n235 VPWR.t686 161.106
R12009 VPWR.n230 VPWR.t683 161.106
R12010 VPWR.n222 VPWR.t906 161.106
R12011 VPWR.n225 VPWR.t904 161.106
R12012 VPWR.n220 VPWR.t901 161.106
R12013 VPWR.n212 VPWR.t925 161.106
R12014 VPWR.n215 VPWR.t943 161.106
R12015 VPWR.n210 VPWR.t940 161.106
R12016 VPWR.n202 VPWR.t698 161.106
R12017 VPWR.n205 VPWR.t696 161.106
R12018 VPWR.n200 VPWR.t693 161.106
R12019 VPWR.n192 VPWR.t794 161.106
R12020 VPWR.n195 VPWR.t792 161.106
R12021 VPWR.n190 VPWR.t811 161.106
R12022 VPWR.n182 VPWR.t830 161.106
R12023 VPWR.n185 VPWR.t833 161.106
R12024 VPWR.n180 VPWR.t827 161.106
R12025 VPWR.n172 VPWR.t971 161.106
R12026 VPWR.n175 VPWR.t969 161.106
R12027 VPWR.n170 VPWR.t675 161.106
R12028 VPWR.n162 VPWR.t714 161.106
R12029 VPWR.n165 VPWR.t712 161.106
R12030 VPWR.n160 VPWR.t709 161.106
R12031 VPWR.n152 VPWR.t849 161.106
R12032 VPWR.n155 VPWR.t847 161.106
R12033 VPWR.n150 VPWR.t841 161.106
R12034 VPWR.n142 VPWR.t880 161.106
R12035 VPWR.n145 VPWR.t980 161.106
R12036 VPWR.n140 VPWR.t974 161.106
R12037 VPWR.n1445 VPWR.t824 161.106
R12038 VPWR.n1704 VPWR.t643 161.106
R12039 VPWR.n1007 VPWR.t891 161.106
R12040 VPWR.n1521 VPWR.t768 161.106
R12041 VPWR.n1526 VPWR.t638 161.106
R12042 VPWR.n1531 VPWR.t883 161.106
R12043 VPWR.n1536 VPWR.t862 161.106
R12044 VPWR.n1541 VPWR.t749 161.106
R12045 VPWR.n1546 VPWR.t623 161.106
R12046 VPWR.n1551 VPWR.t964 161.106
R12047 VPWR.n1556 VPWR.t744 161.106
R12048 VPWR.n1561 VPWR.t704 161.106
R12049 VPWR.n1396 VPWR.t691 161.106
R12050 VPWR.n1391 VPWR.t822 161.106
R12051 VPWR.n1413 VPWR.t770 161.106
R12052 VPWR.n1433 VPWR.t966 161.106
R12053 VPWR.n1437 VPWR.t746 161.106
R12054 VPWR.n1429 VPWR.t609 161.106
R12055 VPWR.n1425 VPWR.t751 161.106
R12056 VPWR.n1421 VPWR.t864 161.106
R12057 VPWR.n1441 VPWR.t706 161.106
R12058 VPWR.n1417 VPWR.t885 161.106
R12059 VPWR.n1409 VPWR.t640 161.106
R12060 VPWR.n1452 VPWR.t612 161.106
R12061 VPWR.n1709 VPWR.t661 161.106
R12062 VPWR.n1717 VPWR.t806 161.106
R12063 VPWR.n1713 VPWR.t920 161.106
R12064 VPWR.n1014 VPWR.t896 161.106
R12065 VPWR.n1681 VPWR.t666 161.106
R12066 VPWR.n1001 VPWR.t808 161.106
R12067 VPWR.n997 VPWR.t922 161.106
R12068 VPWR.n1018 VPWR.t888 161.106
R12069 VPWR.n132 VPWR.t620 161.106
R12070 VPWR.n135 VPWR.t618 161.106
R12071 VPWR.n125 VPWR.t757 161.106
R12072 VPWR.n53 VPWR.t977 161.106
R12073 VPWR.n51 VPWR.t931 161.106
R12074 VPWR.n49 VPWR.t663 161.106
R12075 VPWR.n47 VPWR.t765 161.106
R12076 VPWR.n45 VPWR.t985 161.106
R12077 VPWR.n43 VPWR.t819 161.106
R12078 VPWR.n41 VPWR.t937 161.106
R12079 VPWR.n39 VPWR.t672 161.106
R12080 VPWR.n37 VPWR.t773 161.106
R12081 VPWR.n35 VPWR.t733 161.106
R12082 VPWR.n33 VPWR.t835 161.106
R12083 VPWR.n31 VPWR.t669 161.106
R12084 VPWR.n29 VPWR.t844 161.106
R12085 VPWR.n27 VPWR.t945 161.106
R12086 VPWR.n25 VPWR.t803 161.106
R12087 VPWR.n23 VPWR.t914 161.106
R12088 VPWR.n1114 VPWR.t2020 154.679
R12089 VPWR.n1575 VPWR.t1963 154.679
R12090 VPWR.n1073 VPWR.t1930 154.679
R12091 VPWR.n1578 VPWR.t1931 154.679
R12092 VPWR.n1581 VPWR.t2067 154.679
R12093 VPWR.n1070 VPWR.t2068 154.679
R12094 VPWR.n1584 VPWR.t2069 154.679
R12095 VPWR.n1587 VPWR.t2055 154.679
R12096 VPWR.n1067 VPWR.t2056 154.679
R12097 VPWR.n1590 VPWR.t2057 154.679
R12098 VPWR.n1593 VPWR.t1971 154.679
R12099 VPWR.n1064 VPWR.t1973 154.679
R12100 VPWR.n1596 VPWR.t1974 154.679
R12101 VPWR.n1599 VPWR.t1965 154.679
R12102 VPWR.n1061 VPWR.t1957 154.679
R12103 VPWR.n1602 VPWR.t1958 154.679
R12104 VPWR.n1605 VPWR.t2048 154.679
R12105 VPWR.n1058 VPWR.t2050 154.679
R12106 VPWR.n1608 VPWR.t2051 154.679
R12107 VPWR.n1611 VPWR.t2007 154.679
R12108 VPWR.n1055 VPWR.t2008 154.679
R12109 VPWR.n1614 VPWR.t2002 154.679
R12110 VPWR.n1617 VPWR.t1999 154.679
R12111 VPWR.n1052 VPWR.t2000 154.679
R12112 VPWR.n1620 VPWR.t2001 154.679
R12113 VPWR.n1623 VPWR.t1947 154.679
R12114 VPWR.n1049 VPWR.t1949 154.679
R12115 VPWR.n1626 VPWR.t2058 154.679
R12116 VPWR.n1629 VPWR.t2043 154.679
R12117 VPWR.n1046 VPWR.t2044 154.679
R12118 VPWR.n1632 VPWR.t2046 154.679
R12119 VPWR.n1635 VPWR.t1992 154.679
R12120 VPWR.n1043 VPWR.t1993 154.679
R12121 VPWR.n1638 VPWR.t1994 154.679
R12122 VPWR.n1641 VPWR.t1981 154.679
R12123 VPWR.n1040 VPWR.t1944 154.679
R12124 VPWR.n1644 VPWR.t1945 154.679
R12125 VPWR.n1647 VPWR.t1939 154.679
R12126 VPWR.n1650 VPWR.t1942 154.679
R12127 VPWR.n1036 VPWR.t1943 154.679
R12128 VPWR.n1657 VPWR.t2028 154.679
R12129 VPWR.n1660 VPWR.t2030 154.679
R12130 VPWR.n1655 VPWR.t2032 154.679
R12131 VPWR.n1669 VPWR.t1986 154.679
R12132 VPWR.n1111 VPWR.t2019 154.679
R12133 VPWR.n1075 VPWR.t2018 154.679
R12134 VPWR.n1666 VPWR.t1988 154.679
R12135 VPWR.n1032 VPWR.t1989 154.679
R12136 VPWR.n120 VPWR.t1997 154.679
R12137 VPWR.n113 VPWR.t1954 154.679
R12138 VPWR.n116 VPWR.t1955 154.679
R12139 VPWR.n111 VPWR.t1956 154.679
R12140 VPWR.n130 VPWR.t2054 154.679
R12141 VPWR.n122 VPWR.t1995 154.679
R12142 VPWR.n107 VPWR.t1984 154.679
R12143 VPWR.n103 VPWR.t1983 154.679
R12144 VPWR.n104 VPWR.t1985 154.679
R12145 VPWR.n255 VPWR.t1932 154.679
R12146 VPWR.n252 VPWR.t2040 154.679
R12147 VPWR.n100 VPWR.t2041 154.679
R12148 VPWR.n242 VPWR.t2033 154.679
R12149 VPWR.n245 VPWR.t2034 154.679
R12150 VPWR.n240 VPWR.t2035 154.679
R12151 VPWR.n232 VPWR.t2021 154.679
R12152 VPWR.n235 VPWR.t2022 154.679
R12153 VPWR.n230 VPWR.t2023 154.679
R12154 VPWR.n222 VPWR.t1934 154.679
R12155 VPWR.n225 VPWR.t1935 154.679
R12156 VPWR.n220 VPWR.t1936 154.679
R12157 VPWR.n212 VPWR.t1933 154.679
R12158 VPWR.n215 VPWR.t1926 154.679
R12159 VPWR.n210 VPWR.t1927 154.679
R12160 VPWR.n202 VPWR.t2014 154.679
R12161 VPWR.n205 VPWR.t2015 154.679
R12162 VPWR.n200 VPWR.t2016 154.679
R12163 VPWR.n192 VPWR.t1977 154.679
R12164 VPWR.n195 VPWR.t1978 154.679
R12165 VPWR.n190 VPWR.t1975 154.679
R12166 VPWR.n182 VPWR.t1966 154.679
R12167 VPWR.n185 VPWR.t1967 154.679
R12168 VPWR.n180 VPWR.t1968 154.679
R12169 VPWR.n172 VPWR.t2062 154.679
R12170 VPWR.n175 VPWR.t2063 154.679
R12171 VPWR.n170 VPWR.t2026 154.679
R12172 VPWR.n162 VPWR.t2009 154.679
R12173 VPWR.n165 VPWR.t2010 154.679
R12174 VPWR.n160 VPWR.t2011 154.679
R12175 VPWR.n152 VPWR.t1959 154.679
R12176 VPWR.n155 VPWR.t1960 154.679
R12177 VPWR.n150 VPWR.t1961 154.679
R12178 VPWR.n142 VPWR.t1950 154.679
R12179 VPWR.n145 VPWR.t2059 154.679
R12180 VPWR.n140 VPWR.t2061 154.679
R12181 VPWR.n1445 VPWR.t2065 154.679
R12182 VPWR.n1704 VPWR.t1987 154.679
R12183 VPWR.n1007 VPWR.t2037 154.679
R12184 VPWR.n1521 VPWR.t1940 154.679
R12185 VPWR.n1526 VPWR.t1991 154.679
R12186 VPWR.n1531 VPWR.t2039 154.679
R12187 VPWR.n1536 VPWR.t2049 154.679
R12188 VPWR.n1541 VPWR.t1948 154.679
R12189 VPWR.n1546 VPWR.t1998 154.679
R12190 VPWR.n1551 VPWR.t2006 154.679
R12191 VPWR.n1556 VPWR.t1952 154.679
R12192 VPWR.n1561 VPWR.t1964 154.679
R12193 VPWR.n1396 VPWR.t1972 154.679
R12194 VPWR.n1391 VPWR.t2066 154.679
R12195 VPWR.n1413 VPWR.t1938 154.679
R12196 VPWR.n1433 VPWR.t2005 154.679
R12197 VPWR.n1437 VPWR.t1951 154.679
R12198 VPWR.n1429 VPWR.t2004 154.679
R12199 VPWR.n1425 VPWR.t1946 154.679
R12200 VPWR.n1421 VPWR.t2047 154.679
R12201 VPWR.n1441 VPWR.t1962 154.679
R12202 VPWR.n1417 VPWR.t2038 154.679
R12203 VPWR.n1409 VPWR.t1990 154.679
R12204 VPWR.n1452 VPWR.t2003 154.679
R12205 VPWR.n1709 VPWR.t1982 154.679
R12206 VPWR.n1717 VPWR.t1929 154.679
R12207 VPWR.n1713 VPWR.t2029 154.679
R12208 VPWR.n1014 VPWR.t2036 154.679
R12209 VPWR.n1681 VPWR.t1980 154.679
R12210 VPWR.n1001 VPWR.t1928 154.679
R12211 VPWR.n997 VPWR.t2027 154.679
R12212 VPWR.n1018 VPWR.t2025 154.679
R12213 VPWR.n132 VPWR.t2052 154.679
R12214 VPWR.n135 VPWR.t2053 154.679
R12215 VPWR.n125 VPWR.t1996 154.679
R12216 VPWR.n53 VPWR.t1970 154.679
R12217 VPWR.n51 VPWR.t2064 154.679
R12218 VPWR.n49 VPWR.t2017 154.679
R12219 VPWR.n47 VPWR.t1941 154.679
R12220 VPWR.n45 VPWR.t2045 154.679
R12221 VPWR.n43 VPWR.t1969 154.679
R12222 VPWR.n41 VPWR.t2024 154.679
R12223 VPWR.n39 VPWR.t1979 154.679
R12224 VPWR.n37 VPWR.t1937 154.679
R12225 VPWR.n35 VPWR.t2042 154.679
R12226 VPWR.n33 VPWR.t2060 154.679
R12227 VPWR.n31 VPWR.t2013 154.679
R12228 VPWR.n29 VPWR.t1953 154.679
R12229 VPWR.n27 VPWR.t2012 154.679
R12230 VPWR.n25 VPWR.t1976 154.679
R12231 VPWR.n23 VPWR.t2031 154.679
R12232 VPWR.n1446 VPWR.n1445 152
R12233 VPWR.n1414 VPWR.n1413 152
R12234 VPWR.n1434 VPWR.n1433 152
R12235 VPWR.n1438 VPWR.n1437 152
R12236 VPWR.n1430 VPWR.n1429 152
R12237 VPWR.n1426 VPWR.n1425 152
R12238 VPWR.n1422 VPWR.n1421 152
R12239 VPWR.n1442 VPWR.n1441 152
R12240 VPWR.n1418 VPWR.n1417 152
R12241 VPWR.n1410 VPWR.n1409 152
R12242 VPWR.n1453 VPWR.n1452 152
R12243 VPWR.n1015 VPWR.n1014 152
R12244 VPWR.n1682 VPWR.n1681 152
R12245 VPWR.n1002 VPWR.n1001 152
R12246 VPWR.n998 VPWR.n997 152
R12247 VPWR.n1019 VPWR.n1018 152
R12248 VPWR.n2781 VPWR.n2780 150.213
R12249 VPWR.t401 VPWR.t1830 140.989
R12250 VPWR.t1735 VPWR.t1722 140.989
R12251 VPWR.t1762 VPWR.t1735 140.989
R12252 VPWR.t1737 VPWR.t1762 140.989
R12253 VPWR.t1051 VPWR.t1737 140.989
R12254 VPWR.t1638 VPWR.t1051 140.989
R12255 VPWR.t1166 VPWR.t1638 140.989
R12256 VPWR.t1164 VPWR.t1166 140.989
R12257 VPWR.t1128 VPWR.t557 140.989
R12258 VPWR.t1774 VPWR.t1741 140.989
R12259 VPWR.t1728 VPWR.t1774 140.989
R12260 VPWR.t1775 VPWR.t1728 140.989
R12261 VPWR.t535 VPWR.t1775 140.989
R12262 VPWR.t1150 VPWR.t535 140.989
R12263 VPWR.t1187 VPWR.t1150 140.989
R12264 VPWR.t1191 VPWR.t1187 140.989
R12265 VPWR.t1719 VPWR.t1760 140.989
R12266 VPWR.t1749 VPWR.t1719 140.989
R12267 VPWR.t1723 VPWR.t1749 140.989
R12268 VPWR.t128 VPWR.t1723 140.989
R12269 VPWR.t126 VPWR.t128 140.989
R12270 VPWR.t132 VPWR.t126 140.989
R12271 VPWR.t120 VPWR.t132 140.989
R12272 VPWR.t388 VPWR.t1750 140.989
R12273 VPWR.t1720 VPWR.t1763 140.989
R12274 VPWR.t1770 VPWR.t1720 140.989
R12275 VPWR.t1747 VPWR.t1770 140.989
R12276 VPWR.t1640 VPWR.t1747 140.989
R12277 VPWR.t1634 VPWR.t1640 140.989
R12278 VPWR.t1053 VPWR.t1634 140.989
R12279 VPWR.t1636 VPWR.t1053 140.989
R12280 VPWR.t1742 VPWR.t1729 140.989
R12281 VPWR.t1716 VPWR.t1742 140.989
R12282 VPWR.t1768 VPWR.t1716 140.989
R12283 VPWR.t1148 VPWR.t1768 140.989
R12284 VPWR.t1185 VPWR.t1148 140.989
R12285 VPWR.t1146 VPWR.t1185 140.989
R12286 VPWR.t1189 VPWR.t1146 140.989
R12287 VPWR.t1738 VPWR.t1731 140.989
R12288 VPWR.t1745 VPWR.t1738 140.989
R12289 VPWR.t1733 VPWR.t1745 140.989
R12290 VPWR.t130 VPWR.t1733 140.989
R12291 VPWR.t134 VPWR.t130 140.989
R12292 VPWR.t122 VPWR.t134 140.989
R12293 VPWR.t124 VPWR.t122 140.989
R12294 VPWR VPWR.n1381 133.312
R12295 VPWR.n2777 VPWR.n2776 129.13
R12296 VPWR.n2794 VPWR.n2755 129.13
R12297 VPWR.n2716 VPWR 127.562
R12298 VPWR.n2696 VPWR 127.562
R12299 VPWR.n2677 VPWR 127.562
R12300 VPWR VPWR.t1781 125.883
R12301 VPWR.n2641 VPWR 125.883
R12302 VPWR.t1130 VPWR.t555 120.849
R12303 VPWR.t486 VPWR.t195 117.492
R12304 VPWR.t1126 VPWR.t531 117.492
R12305 VPWR.t1196 VPWR 115.814
R12306 VPWR VPWR.t1164 114.135
R12307 VPWR VPWR.t1191 114.135
R12308 VPWR VPWR.t120 114.135
R12309 VPWR.n2795 VPWR.n2753 111.059
R12310 VPWR.t1446 VPWR 107.421
R12311 VPWR.n1269 VPWR.n1268 106.561
R12312 VPWR.n2717 VPWR.n2716 106.561
R12313 VPWR.n2697 VPWR.n2696 106.561
R12314 VPWR.n2678 VPWR.n2677 106.561
R12315 VPWR.n2642 VPWR.n2641 106.561
R12316 VPWR.n2604 VPWR.n2603 106.561
R12317 VPWR.n2567 VPWR.n2566 106.561
R12318 VPWR VPWR.t1134 106.543
R12319 VPWR VPWR.n1173 104.8
R12320 VPWR VPWR.n1196 104.8
R12321 VPWR VPWR.n1220 104.8
R12322 VPWR VPWR.n1305 104.8
R12323 VPWR VPWR.n1344 104.8
R12324 VPWR.n1382 VPWR 100.883
R12325 VPWR VPWR.t407 100.624
R12326 VPWR.t1859 VPWR.t399 97.9386
R12327 VPWR.n2795 VPWR.n2794 93.3652
R12328 VPWR.n1448 VPWR.n1447 91.7293
R12329 VPWR.n1416 VPWR.n1415 91.7293
R12330 VPWR.n1436 VPWR.n1435 91.7293
R12331 VPWR.n1440 VPWR.n1439 91.7293
R12332 VPWR.n1432 VPWR.n1431 91.7293
R12333 VPWR.n1428 VPWR.n1427 91.7293
R12334 VPWR.n1424 VPWR.n1423 91.7293
R12335 VPWR.n1444 VPWR.n1443 91.7293
R12336 VPWR.n1420 VPWR.n1419 91.7293
R12337 VPWR.n1412 VPWR.n1411 91.7293
R12338 VPWR.n1455 VPWR.n1454 91.7293
R12339 VPWR.n1017 VPWR.n1016 91.7293
R12340 VPWR.n1684 VPWR.n1683 91.7293
R12341 VPWR.n1004 VPWR.n1003 91.7293
R12342 VPWR.n1000 VPWR.n999 91.7293
R12343 VPWR.n1021 VPWR.n1020 91.7293
R12344 VPWR.n2783 VPWR.n2756 91.4829
R12345 VPWR.t1859 VPWR.n2778 90.0872
R12346 VPWR.t1766 VPWR 88.7855
R12347 VPWR.n1174 VPWR 79.407
R12348 VPWR.n1197 VPWR 79.407
R12349 VPWR.n1221 VPWR 79.407
R12350 VPWR.n1306 VPWR 79.407
R12351 VPWR.n1345 VPWR 79.407
R12352 VPWR.t1300 VPWR.t274 78.8874
R12353 VPWR.n2776 VPWR.n2754 74.9181
R12354 VPWR.n2794 VPWR.n2754 74.9181
R12355 VPWR.n2794 VPWR.n2793 74.9181
R12356 VPWR.n2793 VPWR.n2756 74.9181
R12357 VPWR.t154 VPWR.t1447 70.4952
R12358 VPWR.t1447 VPWR.t157 70.4952
R12359 VPWR.t157 VPWR.t1854 70.4952
R12360 VPWR.t1854 VPWR.t228 70.4952
R12361 VPWR.t228 VPWR.t405 70.4952
R12362 VPWR.t405 VPWR.t347 70.4952
R12363 VPWR.t347 VPWR.t401 70.4952
R12364 VPWR.t1754 VPWR.t388 70.4952
R12365 VPWR.t394 VPWR.t1754 70.4952
R12366 VPWR.t1726 VPWR.t394 70.4952
R12367 VPWR.t1156 VPWR.t1726 70.4952
R12368 VPWR.t1758 VPWR.t1156 70.4952
R12369 VPWR.t392 VPWR.t1758 70.4952
R12370 VPWR.t1781 VPWR.t392 70.4952
R12371 VPWR VPWR.t154 68.8168
R12372 VPWR.t1136 VPWR.t1132 68.8168
R12373 VPWR.t274 VPWR.t1196 62.103
R12374 VPWR VPWR.t1128 60.4245
R12375 VPWR.n2785 VPWR.n2778 59.762
R12376 VPWR.n2781 VPWR.n2755 53.8358
R12377 VPWR.t1132 VPWR.t34 52.0323
R12378 VPWR.t1419 VPWR 50.3539
R12379 VPWR VPWR.t1136 50.3539
R12380 VPWR VPWR.t1130 50.3539
R12381 VPWR.t1763 VPWR 50.3539
R12382 VPWR.t1729 VPWR 50.3539
R12383 VPWR.t1731 VPWR 50.3539
R12384 VPWR.n2790 VPWR.n2754 46.2505
R12385 VPWR.n2791 VPWR.n2790 46.2505
R12386 VPWR.n2771 VPWR.n2770 46.2505
R12387 VPWR.n2772 VPWR.n2771 46.2505
R12388 VPWR.n2774 VPWR.n2773 46.2505
R12389 VPWR.n2773 VPWR.n2772 46.2505
R12390 VPWR.n2780 VPWR.n2760 46.2505
R12391 VPWR.n2793 VPWR.n2792 46.2505
R12392 VPWR.n2792 VPWR.n2791 46.2505
R12393 VPWR.n2785 VPWR.n2784 46.2505
R12394 VPWR.n2782 VPWR.n2781 45.9299
R12395 VPWR.n2768 VPWR.n2766 44.8005
R12396 VPWR.n2766 VPWR.n2762 44.8005
R12397 VPWR.n2783 VPWR.n2779 37.0005
R12398 VPWR.n2779 VPWR.t399 37.0005
R12399 VPWR.n1238 VPWR.n1237 34.6358
R12400 VPWR.n1296 VPWR.n1280 34.6358
R12401 VPWR.n1301 VPWR.n1300 34.6358
R12402 VPWR.n1335 VPWR.n1319 34.6358
R12403 VPWR.n1340 VPWR.n1339 34.6358
R12404 VPWR.n1350 VPWR.n1316 34.6358
R12405 VPWR.n1372 VPWR.n1356 34.6358
R12406 VPWR.n1377 VPWR.n1376 34.6358
R12407 VPWR.n2691 VPWR.n2690 34.6358
R12408 VPWR.n2657 VPWR.n2649 34.6358
R12409 VPWR.n2664 VPWR.n2663 34.6358
R12410 VPWR.n2621 VPWR.n2612 34.6358
R12411 VPWR.n2624 VPWR.n2623 34.6358
R12412 VPWR.n2628 VPWR.n2627 34.6358
R12413 VPWR.n2584 VPWR.n2575 34.6358
R12414 VPWR.n2587 VPWR.n2586 34.6358
R12415 VPWR.n2591 VPWR.n2590 34.6358
R12416 VPWR.n2598 VPWR.n2597 34.6358
R12417 VPWR.n2551 VPWR.n2547 34.6358
R12418 VPWR.n2555 VPWR.n2539 34.6358
R12419 VPWR.n2558 VPWR.n2557 34.6358
R12420 VPWR.n1447 VPWR.n1446 33.9921
R12421 VPWR.n1415 VPWR.n1414 33.9921
R12422 VPWR.n1435 VPWR.n1434 33.9921
R12423 VPWR.n1439 VPWR.n1438 33.9921
R12424 VPWR.n1431 VPWR.n1430 33.9921
R12425 VPWR.n1427 VPWR.n1426 33.9921
R12426 VPWR.n1423 VPWR.n1422 33.9921
R12427 VPWR.n1443 VPWR.n1442 33.9921
R12428 VPWR.n1419 VPWR.n1418 33.9921
R12429 VPWR.n1411 VPWR.n1410 33.9921
R12430 VPWR.n1454 VPWR.n1453 33.9921
R12431 VPWR.n1016 VPWR.n1015 33.9921
R12432 VPWR.n1683 VPWR.n1682 33.9921
R12433 VPWR.n1003 VPWR.n1002 33.9921
R12434 VPWR.n999 VPWR.n998 33.9921
R12435 VPWR.n1020 VPWR.n1019 33.9921
R12436 VPWR.n1255 VPWR.n1254 32.0005
R12437 VPWR.n1292 VPWR.n1291 32.0005
R12438 VPWR.n1331 VPWR.n1330 32.0005
R12439 VPWR.n1368 VPWR.n1367 32.0005
R12440 VPWR.n2653 VPWR.n2652 30.8711
R12441 VPWR.n2617 VPWR.n2616 30.8711
R12442 VPWR.n2580 VPWR.n2579 30.8711
R12443 VPWR.n2546 VPWR.n2545 30.8711
R12444 VPWR.n2770 VPWR.n2768 30.1181
R12445 VPWR.n2774 VPWR.n2762 30.1181
R12446 VPWR.n2784 VPWR.n2782 28.9887
R12447 VPWR.n1264 VPWR.n1263 28.2358
R12448 VPWR.n5 VPWR.t1857 26.5955
R12449 VPWR.n5 VPWR.t404 26.5955
R12450 VPWR.n4 VPWR.t408 26.5955
R12451 VPWR.n4 VPWR.t1853 26.5955
R12452 VPWR.n1179 VPWR.t204 26.5955
R12453 VPWR.n1179 VPWR.t203 26.5955
R12454 VPWR.n1178 VPWR.t605 26.5955
R12455 VPWR.n1178 VPWR.t1041 26.5955
R12456 VPWR.n1184 VPWR.t199 26.5955
R12457 VPWR.n1184 VPWR.t205 26.5955
R12458 VPWR.n1177 VPWR.t166 26.5955
R12459 VPWR.n1177 VPWR.t604 26.5955
R12460 VPWR.n1202 VPWR.t1449 26.5955
R12461 VPWR.n1202 VPWR.t1450 26.5955
R12462 VPWR.n1201 VPWR.t413 26.5955
R12463 VPWR.n1201 VPWR.t411 26.5955
R12464 VPWR.n1207 VPWR.t1821 26.5955
R12465 VPWR.n1207 VPWR.t1823 26.5955
R12466 VPWR.n1200 VPWR.t416 26.5955
R12467 VPWR.n1200 VPWR.t414 26.5955
R12468 VPWR.n1226 VPWR.t1314 26.5955
R12469 VPWR.n1226 VPWR.t1321 26.5955
R12470 VPWR.n1225 VPWR.t52 26.5955
R12471 VPWR.n1225 VPWR.t51 26.5955
R12472 VPWR.n1231 VPWR.t1318 26.5955
R12473 VPWR.n1231 VPWR.t1315 26.5955
R12474 VPWR.n1224 VPWR.t55 26.5955
R12475 VPWR.n1224 VPWR.t53 26.5955
R12476 VPWR.n1253 VPWR.t1833 26.5955
R12477 VPWR.n1253 VPWR.t1835 26.5955
R12478 VPWR.n1246 VPWR.t402 26.5955
R12479 VPWR.n1246 VPWR.t1831 26.5955
R12480 VPWR.n1260 VPWR.t1855 26.5955
R12481 VPWR.n1260 VPWR.t406 26.5955
R12482 VPWR.n1262 VPWR.t158 26.5955
R12483 VPWR.n1262 VPWR.t229 26.5955
R12484 VPWR.n1290 VPWR.t1006 26.5955
R12485 VPWR.n1290 VPWR.t225 26.5955
R12486 VPWR.n1289 VPWR.t1669 26.5955
R12487 VPWR.n1289 VPWR.t3 26.5955
R12488 VPWR.n1283 VPWR.t207 26.5955
R12489 VPWR.n1283 VPWR.t1000 26.5955
R12490 VPWR.n1282 VPWR.t167 26.5955
R12491 VPWR.n1282 VPWR.t1786 26.5955
R12492 VPWR.n1298 VPWR.t202 26.5955
R12493 VPWR.n1298 VPWR.t201 26.5955
R12494 VPWR.n1297 VPWR.t1042 26.5955
R12495 VPWR.n1297 VPWR.t603 26.5955
R12496 VPWR.n1329 VPWR.t1785 26.5955
R12497 VPWR.n1329 VPWR.t1671 26.5955
R12498 VPWR.n1328 VPWR.t1008 26.5955
R12499 VPWR.n1328 VPWR.t227 26.5955
R12500 VPWR.n1322 VPWR.t1010 26.5955
R12501 VPWR.n1322 VPWR.t1837 26.5955
R12502 VPWR.n1321 VPWR.t417 26.5955
R12503 VPWR.n1321 VPWR.t1003 26.5955
R12504 VPWR.n1337 VPWR.t1009 26.5955
R12505 VPWR.n1337 VPWR.t1820 26.5955
R12506 VPWR.n1336 VPWR.t418 26.5955
R12507 VPWR.n1336 VPWR.t415 26.5955
R12508 VPWR.n1366 VPWR.t11 26.5955
R12509 VPWR.n1366 VPWR.t159 26.5955
R12510 VPWR.n1365 VPWR.t1670 26.5955
R12511 VPWR.n1365 VPWR.t5 26.5955
R12512 VPWR.n1359 VPWR.t1317 26.5955
R12513 VPWR.n1359 VPWR.t7 26.5955
R12514 VPWR.n1358 VPWR.t49 26.5955
R12515 VPWR.n1358 VPWR.t1787 26.5955
R12516 VPWR.n1374 VPWR.t1320 26.5955
R12517 VPWR.n1374 VPWR.t1319 26.5955
R12518 VPWR.n1373 VPWR.t50 26.5955
R12519 VPWR.n1373 VPWR.t48 26.5955
R12520 VPWR.n2738 VPWR.t1155 26.5955
R12521 VPWR.n2738 VPWR.t1153 26.5955
R12522 VPWR.n2740 VPWR.t391 26.5955
R12523 VPWR.n2740 VPWR.t574 26.5955
R12524 VPWR.n2718 VPWR.t1643 26.5955
R12525 VPWR.n2718 VPWR.t1639 26.5955
R12526 VPWR.n2719 VPWR.t1052 26.5955
R12527 VPWR.n2719 VPWR.t1913 26.5955
R12528 VPWR.n2722 VPWR.t1632 26.5955
R12529 VPWR.n2722 VPWR.t1633 26.5955
R12530 VPWR.n2723 VPWR.t1167 26.5955
R12531 VPWR.n2723 VPWR.t1165 26.5955
R12532 VPWR.n2698 VPWR.t536 26.5955
R12533 VPWR.n2698 VPWR.t1151 26.5955
R12534 VPWR.n2699 VPWR.t1184 26.5955
R12535 VPWR.n2699 VPWR.t1194 26.5955
R12536 VPWR.n2702 VPWR.t1621 26.5955
R12537 VPWR.n2702 VPWR.t1620 26.5955
R12538 VPWR.n2703 VPWR.t1188 26.5955
R12539 VPWR.n2703 VPWR.t1192 26.5955
R12540 VPWR.n2679 VPWR.t1874 26.5955
R12541 VPWR.n2679 VPWR.t1871 26.5955
R12542 VPWR.n2680 VPWR.t129 26.5955
R12543 VPWR.n2680 VPWR.t127 26.5955
R12544 VPWR.n2683 VPWR.t1875 26.5955
R12545 VPWR.n2683 VPWR.t1876 26.5955
R12546 VPWR.n2684 VPWR.t133 26.5955
R12547 VPWR.n2684 VPWR.t121 26.5955
R12548 VPWR.n2644 VPWR.t1727 26.5955
R12549 VPWR.n2644 VPWR.t1759 26.5955
R12550 VPWR.n2648 VPWR.t1751 26.5955
R12551 VPWR.n2648 VPWR.t389 26.5955
R12552 VPWR.n2651 VPWR.t1725 26.5955
R12553 VPWR.n2651 VPWR.t1773 26.5955
R12554 VPWR.n2645 VPWR.t395 26.5955
R12555 VPWR.n2645 VPWR.t1157 26.5955
R12556 VPWR.n2615 VPWR.t1721 26.5955
R12557 VPWR.n2615 VPWR.t1771 26.5955
R12558 VPWR.n2614 VPWR.t1740 26.5955
R12559 VPWR.n2614 VPWR.t1783 26.5955
R12560 VPWR.n2611 VPWR.t1748 26.5955
R12561 VPWR.n2611 VPWR.t1912 26.5955
R12562 VPWR.n2610 VPWR.t1765 26.5955
R12563 VPWR.n2610 VPWR.t1641 26.5955
R12564 VPWR.n2607 VPWR.t1915 26.5955
R12565 VPWR.n2607 VPWR.t1054 26.5955
R12566 VPWR.n2606 VPWR.t1635 26.5955
R12567 VPWR.n2606 VPWR.t1642 26.5955
R12568 VPWR.n2578 VPWR.t1743 26.5955
R12569 VPWR.n2578 VPWR.t1717 26.5955
R12570 VPWR.n2577 VPWR.t1761 26.5955
R12571 VPWR.n2577 VPWR.t1736 26.5955
R12572 VPWR.n2574 VPWR.t1769 26.5955
R12573 VPWR.n2574 VPWR.t1193 26.5955
R12574 VPWR.n2573 VPWR.t1779 26.5955
R12575 VPWR.n2573 VPWR.t1149 26.5955
R12576 VPWR.n2570 VPWR.t1186 26.5955
R12577 VPWR.n2570 VPWR.t1195 26.5955
R12578 VPWR.n2569 VPWR.t1619 26.5955
R12579 VPWR.n2569 VPWR.t1147 26.5955
R12580 VPWR.n2542 VPWR.t1739 26.5955
R12581 VPWR.n2542 VPWR.t1746 26.5955
R12582 VPWR.n2541 VPWR.t1776 26.5955
R12583 VPWR.n2541 VPWR.t1757 26.5955
R12584 VPWR.n2549 VPWR.t1752 26.5955
R12585 VPWR.n2549 VPWR.t131 26.5955
R12586 VPWR.n2548 VPWR.t1734 26.5955
R12587 VPWR.n2548 VPWR.t1872 26.5955
R12588 VPWR.n2538 VPWR.t135 26.5955
R12589 VPWR.n2538 VPWR.t123 26.5955
R12590 VPWR.n2537 VPWR.t1869 26.5955
R12591 VPWR.n2537 VPWR.t1873 26.5955
R12592 VPWR.n17 VPWR.n16 25.977
R12593 VPWR.n1192 VPWR.n1191 25.977
R12594 VPWR.n1252 VPWR.n1249 25.977
R12595 VPWR.n1288 VPWR.n1285 25.977
R12596 VPWR.n1311 VPWR.n1277 25.977
R12597 VPWR.n1327 VPWR.n1324 25.977
R12598 VPWR.n1364 VPWR.n1361 25.977
R12599 VPWR.n2747 VPWR.n2746 25.977
R12600 VPWR.n2731 VPWR.n2730 25.977
R12601 VPWR.n2653 VPWR.n2650 25.977
R12602 VPWR.n2617 VPWR.n2613 25.977
R12603 VPWR.n2635 VPWR.n2634 25.977
R12604 VPWR.n2580 VPWR.n2576 25.977
R12605 VPWR.n2545 VPWR.n2543 25.977
R12606 VPWR.n1274 VPWR.n1273 25.224
R12607 VPWR.n2673 VPWR.n2672 25.224
R12608 VPWR.n2658 VPWR.n2657 24.8476
R12609 VPWR.n2622 VPWR.n2621 24.8476
R12610 VPWR.n2585 VPWR.n2584 24.8476
R12611 VPWR.n2551 VPWR.n2550 24.8476
R12612 VPWR.n16 VPWR.n15 24.4711
R12613 VPWR.n1191 VPWR.n1190 24.4711
R12614 VPWR.n1254 VPWR.n1252 24.4711
R12615 VPWR.n1291 VPWR.n1288 24.4711
R12616 VPWR.n1330 VPWR.n1327 24.4711
R12617 VPWR.n1367 VPWR.n1364 24.4711
R12618 VPWR.n2746 VPWR.n2745 24.4711
R12619 VPWR.n2730 VPWR.n2729 24.4711
R12620 VPWR.n11 VPWR.n2 23.7181
R12621 VPWR.n1186 VPWR.n1175 23.7181
R12622 VPWR.n1209 VPWR.n1198 23.7181
R12623 VPWR.n1213 VPWR.n1198 23.7181
R12624 VPWR.n1233 VPWR.n1222 23.7181
R12625 VPWR.n1237 VPWR.n1222 23.7181
R12626 VPWR.n1269 VPWR.n1267 23.7181
R12627 VPWR.n1307 VPWR.n1304 23.7181
R12628 VPWR.n1346 VPWR.n1343 23.7181
R12629 VPWR.n1346 VPWR.n1316 23.7181
R12630 VPWR.n1383 VPWR.n1380 23.7181
R12631 VPWR.n2744 VPWR.n2743 23.7181
R12632 VPWR.n2725 VPWR.n2717 23.7181
R12633 VPWR.n2705 VPWR.n2697 23.7181
R12634 VPWR.n2709 VPWR.n2697 23.7181
R12635 VPWR.n2686 VPWR.n2678 23.7181
R12636 VPWR.n2690 VPWR.n2678 23.7181
R12637 VPWR.n2667 VPWR.n2642 23.7181
R12638 VPWR.n2630 VPWR.n2604 23.7181
R12639 VPWR.n2593 VPWR.n2567 23.7181
R12640 VPWR.n2597 VPWR.n2567 23.7181
R12641 VPWR.n2562 VPWR.n2561 23.7181
R12642 VPWR.t197 VPWR.t486 23.4987
R12643 VPWR.t533 VPWR.t1126 23.4987
R12644 VPWR.n2788 VPWR.n2777 23.1255
R12645 VPWR.n2788 VPWR.t1859 23.1255
R12646 VPWR.n2787 VPWR.n2755 23.1255
R12647 VPWR.t1859 VPWR.n2787 23.1255
R12648 VPWR.n11 VPWR.n10 22.9652
R12649 VPWR.n1186 VPWR.n1185 22.9652
R12650 VPWR.n1209 VPWR.n1208 22.9652
R12651 VPWR.n1233 VPWR.n1232 22.9652
R12652 VPWR.n2743 VPWR.n2739 22.9652
R12653 VPWR.n2725 VPWR.n2724 22.9652
R12654 VPWR.n2705 VPWR.n2704 22.9652
R12655 VPWR.n2686 VPWR.n2685 22.9652
R12656 VPWR.n1259 VPWR.n1247 22.2123
R12657 VPWR.n2660 VPWR.n2659 22.2123
R12658 VPWR.n10 VPWR.n3 21.4593
R12659 VPWR.n1185 VPWR.n1176 21.4593
R12660 VPWR.n1208 VPWR.n1199 21.4593
R12661 VPWR.n1232 VPWR.n1223 21.4593
R12662 VPWR.n1381 VPWR.t4 20.5957
R12663 VPWR.n1382 VPWR.t6 20.5957
R12664 VPWR.n1216 VPWR.n1215 19.9534
R12665 VPWR.n1239 VPWR.n1238 19.9534
R12666 VPWR.n1273 VPWR.n1242 19.9534
R12667 VPWR.n2712 VPWR.n2711 19.9534
R12668 VPWR.n2692 VPWR.n2691 19.9534
R12669 VPWR.n2672 VPWR.n2671 19.9534
R12670 VPWR.n2660 VPWR.n2646 18.824
R12671 VPWR.n2624 VPWR.n2608 18.824
R12672 VPWR.n2587 VPWR.n2571 18.824
R12673 VPWR.n2556 VPWR.n2555 18.824
R12674 VPWR.n1255 VPWR.n1247 18.4476
R12675 VPWR.n1292 VPWR.n1284 18.4476
R12676 VPWR.n1312 VPWR.n1311 18.4476
R12677 VPWR.n1331 VPWR.n1323 18.4476
R12678 VPWR.n1368 VPWR.n1360 18.4476
R12679 VPWR.n2636 VPWR.n2635 18.4476
R12680 VPWR.n1352 VPWR.n1351 17.5829
R12681 VPWR.n2600 VPWR.n2599 17.5829
R12682 VPWR.n6 VPWR.n3 16.9417
R12683 VPWR.n1180 VPWR.n1176 16.9417
R12684 VPWR.n1203 VPWR.n1199 16.9417
R12685 VPWR.n1227 VPWR.n1223 16.9417
R12686 VPWR.n2666 VPWR.n2665 16.5652
R12687 VPWR.n1245 VPWR.n1243 16.1887
R12688 VPWR.n1313 VPWR.n1312 16.1887
R12689 VPWR.n2637 VPWR.n2636 16.1887
R12690 VPWR.n1174 VPWR.t161 16.0935
R12691 VPWR.n1197 VPWR.t1005 16.0935
R12692 VPWR.n1221 VPWR.t1 16.0935
R12693 VPWR.n1306 VPWR.t200 16.0935
R12694 VPWR.n1345 VPWR.t162 16.0935
R12695 VPWR.n1173 VPWR.t156 16.0935
R12696 VPWR.n1196 VPWR.t160 16.0935
R12697 VPWR.n1220 VPWR.t8 16.0935
R12698 VPWR.n1305 VPWR.t2 16.0935
R12699 VPWR.n1344 VPWR.t226 16.0935
R12700 VPWR.n1264 VPWR.n1245 15.8123
R12701 VPWR.n2663 VPWR.n2646 15.8123
R12702 VPWR.n2665 VPWR.n2664 15.8123
R12703 VPWR.n2627 VPWR.n2608 15.8123
R12704 VPWR.n2590 VPWR.n2571 15.8123
R12705 VPWR.n2557 VPWR.n2556 15.8123
R12706 VPWR.n1269 VPWR.n1242 13.5534
R12707 VPWR.n2671 VPWR.n2642 13.5534
R12708 VPWR.n2775 VPWR.n2759 13.2148
R12709 VPWR.n2759 VPWR.t1210 13.2148
R12710 VPWR.n2763 VPWR.n2753 13.2148
R12711 VPWR.n2763 VPWR.t1210 13.2148
R12712 VPWR.n2769 VPWR.n2765 13.2148
R12713 VPWR.n2765 VPWR.t1210 13.2148
R12714 VPWR.n15 VPWR.n2 12.8005
R12715 VPWR.n1190 VPWR.n1175 12.8005
R12716 VPWR.n1307 VPWR.n1277 12.8005
R12717 VPWR.n2745 VPWR.n2744 12.8005
R12718 VPWR.n2729 VPWR.n2717 12.8005
R12719 VPWR.n2634 VPWR.n2604 12.8005
R12720 VPWR.n1261 VPWR.n1259 12.424
R12721 VPWR.n1299 VPWR.n1296 12.424
R12722 VPWR.n1338 VPWR.n1335 12.424
R12723 VPWR.n1375 VPWR.n1372 12.424
R12724 VPWR.n1215 VPWR.n1214 10.5417
R12725 VPWR.n1351 VPWR.n1350 10.5417
R12726 VPWR.n2711 VPWR.n2710 10.5417
R12727 VPWR.n2599 VPWR.n2598 10.5417
R12728 VPWR.n2623 VPWR.n2622 9.78874
R12729 VPWR.n2586 VPWR.n2585 9.78874
R12730 VPWR.n2550 VPWR.n2539 9.78874
R12731 VPWR.n1300 VPWR.n1299 9.41227
R12732 VPWR.n1304 VPWR.n1278 9.41227
R12733 VPWR.n1339 VPWR.n1338 9.41227
R12734 VPWR.n1343 VPWR.n1317 9.41227
R12735 VPWR.n1376 VPWR.n1375 9.41227
R12736 VPWR.n1380 VPWR.n1354 9.41227
R12737 VPWR.n2630 VPWR.n2629 9.41227
R12738 VPWR.n2593 VPWR.n2592 9.41227
R12739 VPWR.n2561 VPWR.n2535 9.41227
R12740 VPWR.n1446 VPWR 9.363
R12741 VPWR.n1414 VPWR 9.363
R12742 VPWR.n1434 VPWR 9.363
R12743 VPWR.n1438 VPWR 9.363
R12744 VPWR.n1430 VPWR 9.363
R12745 VPWR.n1426 VPWR 9.363
R12746 VPWR.n1422 VPWR 9.363
R12747 VPWR.n1442 VPWR 9.363
R12748 VPWR.n1418 VPWR 9.363
R12749 VPWR.n1410 VPWR 9.363
R12750 VPWR.n1453 VPWR 9.363
R12751 VPWR.n1015 VPWR 9.363
R12752 VPWR.n1682 VPWR 9.363
R12753 VPWR.n1002 VPWR 9.363
R12754 VPWR.n998 VPWR 9.363
R12755 VPWR.n1019 VPWR 9.363
R12756 VPWR.n1450 VPWR.n1449 9.33404
R12757 VPWR.n320 VPWR.n319 9.33404
R12758 VPWR.n1512 VPWR.n1511 9.33404
R12759 VPWR.n316 VPWR.n315 9.33404
R12760 VPWR.n933 VPWR.n932 9.33404
R12761 VPWR.n2415 VPWR.n2414 9.33404
R12762 VPWR.n2411 VPWR.n2410 9.33404
R12763 VPWR.n288 VPWR.n287 9.33404
R12764 VPWR.n941 VPWR.n940 9.33404
R12765 VPWR.n2381 VPWR.n2380 9.33404
R12766 VPWR.n292 VPWR.n291 9.33404
R12767 VPWR.n1827 VPWR.n1826 9.33404
R12768 VPWR.n1823 VPWR.n1822 9.33404
R12769 VPWR.n1817 VPWR.n1816 9.33404
R12770 VPWR.n357 VPWR.n356 9.33404
R12771 VPWR.n361 VPWR.n360 9.33404
R12772 VPWR.n365 VPWR.n364 9.33404
R12773 VPWR.n2391 VPWR.n2390 9.33404
R12774 VPWR.n300 VPWR.n299 9.33404
R12775 VPWR.n1813 VPWR.n1812 9.33404
R12776 VPWR.n373 VPWR.n372 9.33404
R12777 VPWR.n2395 VPWR.n2394 9.33404
R12778 VPWR.n304 VPWR.n303 9.33404
R12779 VPWR.n2244 VPWR.n2243 9.33404
R12780 VPWR.n2248 VPWR.n2247 9.33404
R12781 VPWR.n2254 VPWR.n2253 9.33404
R12782 VPWR.n2258 VPWR.n2257 9.33404
R12783 VPWR.n2268 VPWR.n2267 9.33404
R12784 VPWR.n2274 VPWR.n2273 9.33404
R12785 VPWR.n2278 VPWR.n2277 9.33404
R12786 VPWR.n2284 VPWR.n2283 9.33404
R12787 VPWR.n2288 VPWR.n2287 9.33404
R12788 VPWR.n2294 VPWR.n2293 9.33404
R12789 VPWR.n2298 VPWR.n2297 9.33404
R12790 VPWR.n2304 VPWR.n2303 9.33404
R12791 VPWR.n2308 VPWR.n2307 9.33404
R12792 VPWR.n2314 VPWR.n2313 9.33404
R12793 VPWR.n2317 VPWR.n2316 9.33404
R12794 VPWR.n2264 VPWR.n2263 9.33404
R12795 VPWR.n512 VPWR.n511 9.33404
R12796 VPWR.n508 VPWR.n507 9.33404
R12797 VPWR.n504 VPWR.n503 9.33404
R12798 VPWR.n500 VPWR.n499 9.33404
R12799 VPWR.n492 VPWR.n491 9.33404
R12800 VPWR.n488 VPWR.n487 9.33404
R12801 VPWR.n484 VPWR.n483 9.33404
R12802 VPWR.n480 VPWR.n479 9.33404
R12803 VPWR.n476 VPWR.n475 9.33404
R12804 VPWR.n472 VPWR.n471 9.33404
R12805 VPWR.n468 VPWR.n467 9.33404
R12806 VPWR.n464 VPWR.n463 9.33404
R12807 VPWR.n460 VPWR.n459 9.33404
R12808 VPWR.n456 VPWR.n455 9.33404
R12809 VPWR.n453 VPWR.n452 9.33404
R12810 VPWR.n496 VPWR.n495 9.33404
R12811 VPWR.n2219 VPWR.n2218 9.33404
R12812 VPWR.n2215 VPWR.n2214 9.33404
R12813 VPWR.n2209 VPWR.n2208 9.33404
R12814 VPWR.n2205 VPWR.n2204 9.33404
R12815 VPWR.n2195 VPWR.n2194 9.33404
R12816 VPWR.n2189 VPWR.n2188 9.33404
R12817 VPWR.n2185 VPWR.n2184 9.33404
R12818 VPWR.n2179 VPWR.n2178 9.33404
R12819 VPWR.n2175 VPWR.n2174 9.33404
R12820 VPWR.n2169 VPWR.n2168 9.33404
R12821 VPWR.n2165 VPWR.n2164 9.33404
R12822 VPWR.n2159 VPWR.n2158 9.33404
R12823 VPWR.n2155 VPWR.n2154 9.33404
R12824 VPWR.n2149 VPWR.n2148 9.33404
R12825 VPWR.n2146 VPWR.n2145 9.33404
R12826 VPWR.n2199 VPWR.n2198 9.33404
R12827 VPWR.n549 VPWR.n548 9.33404
R12828 VPWR.n553 VPWR.n552 9.33404
R12829 VPWR.n557 VPWR.n556 9.33404
R12830 VPWR.n561 VPWR.n560 9.33404
R12831 VPWR.n569 VPWR.n568 9.33404
R12832 VPWR.n573 VPWR.n572 9.33404
R12833 VPWR.n577 VPWR.n576 9.33404
R12834 VPWR.n581 VPWR.n580 9.33404
R12835 VPWR.n585 VPWR.n584 9.33404
R12836 VPWR.n589 VPWR.n588 9.33404
R12837 VPWR.n593 VPWR.n592 9.33404
R12838 VPWR.n597 VPWR.n596 9.33404
R12839 VPWR.n601 VPWR.n600 9.33404
R12840 VPWR.n605 VPWR.n604 9.33404
R12841 VPWR.n608 VPWR.n607 9.33404
R12842 VPWR.n565 VPWR.n564 9.33404
R12843 VPWR.n2048 VPWR.n2047 9.33404
R12844 VPWR.n2052 VPWR.n2051 9.33404
R12845 VPWR.n2058 VPWR.n2057 9.33404
R12846 VPWR.n2062 VPWR.n2061 9.33404
R12847 VPWR.n2072 VPWR.n2071 9.33404
R12848 VPWR.n2078 VPWR.n2077 9.33404
R12849 VPWR.n2082 VPWR.n2081 9.33404
R12850 VPWR.n2088 VPWR.n2087 9.33404
R12851 VPWR.n2092 VPWR.n2091 9.33404
R12852 VPWR.n2098 VPWR.n2097 9.33404
R12853 VPWR.n2102 VPWR.n2101 9.33404
R12854 VPWR.n2108 VPWR.n2107 9.33404
R12855 VPWR.n2112 VPWR.n2111 9.33404
R12856 VPWR.n2118 VPWR.n2117 9.33404
R12857 VPWR.n2121 VPWR.n2120 9.33404
R12858 VPWR.n2068 VPWR.n2067 9.33404
R12859 VPWR.n704 VPWR.n703 9.33404
R12860 VPWR.n700 VPWR.n699 9.33404
R12861 VPWR.n696 VPWR.n695 9.33404
R12862 VPWR.n692 VPWR.n691 9.33404
R12863 VPWR.n684 VPWR.n683 9.33404
R12864 VPWR.n680 VPWR.n679 9.33404
R12865 VPWR.n676 VPWR.n675 9.33404
R12866 VPWR.n672 VPWR.n671 9.33404
R12867 VPWR.n668 VPWR.n667 9.33404
R12868 VPWR.n664 VPWR.n663 9.33404
R12869 VPWR.n660 VPWR.n659 9.33404
R12870 VPWR.n656 VPWR.n655 9.33404
R12871 VPWR.n652 VPWR.n651 9.33404
R12872 VPWR.n648 VPWR.n647 9.33404
R12873 VPWR.n645 VPWR.n644 9.33404
R12874 VPWR.n688 VPWR.n687 9.33404
R12875 VPWR.n2023 VPWR.n2022 9.33404
R12876 VPWR.n2019 VPWR.n2018 9.33404
R12877 VPWR.n2013 VPWR.n2012 9.33404
R12878 VPWR.n2009 VPWR.n2008 9.33404
R12879 VPWR.n1999 VPWR.n1998 9.33404
R12880 VPWR.n1993 VPWR.n1992 9.33404
R12881 VPWR.n1989 VPWR.n1988 9.33404
R12882 VPWR.n1983 VPWR.n1982 9.33404
R12883 VPWR.n1979 VPWR.n1978 9.33404
R12884 VPWR.n1973 VPWR.n1972 9.33404
R12885 VPWR.n1969 VPWR.n1968 9.33404
R12886 VPWR.n1963 VPWR.n1962 9.33404
R12887 VPWR.n1959 VPWR.n1958 9.33404
R12888 VPWR.n1953 VPWR.n1952 9.33404
R12889 VPWR.n1950 VPWR.n1949 9.33404
R12890 VPWR.n2003 VPWR.n2002 9.33404
R12891 VPWR.n741 VPWR.n740 9.33404
R12892 VPWR.n745 VPWR.n744 9.33404
R12893 VPWR.n749 VPWR.n748 9.33404
R12894 VPWR.n753 VPWR.n752 9.33404
R12895 VPWR.n761 VPWR.n760 9.33404
R12896 VPWR.n765 VPWR.n764 9.33404
R12897 VPWR.n769 VPWR.n768 9.33404
R12898 VPWR.n773 VPWR.n772 9.33404
R12899 VPWR.n777 VPWR.n776 9.33404
R12900 VPWR.n781 VPWR.n780 9.33404
R12901 VPWR.n785 VPWR.n784 9.33404
R12902 VPWR.n789 VPWR.n788 9.33404
R12903 VPWR.n793 VPWR.n792 9.33404
R12904 VPWR.n797 VPWR.n796 9.33404
R12905 VPWR.n800 VPWR.n799 9.33404
R12906 VPWR.n757 VPWR.n756 9.33404
R12907 VPWR.n1852 VPWR.n1851 9.33404
R12908 VPWR.n1856 VPWR.n1855 9.33404
R12909 VPWR.n1862 VPWR.n1861 9.33404
R12910 VPWR.n1866 VPWR.n1865 9.33404
R12911 VPWR.n1876 VPWR.n1875 9.33404
R12912 VPWR.n1882 VPWR.n1881 9.33404
R12913 VPWR.n1886 VPWR.n1885 9.33404
R12914 VPWR.n1892 VPWR.n1891 9.33404
R12915 VPWR.n1896 VPWR.n1895 9.33404
R12916 VPWR.n1902 VPWR.n1901 9.33404
R12917 VPWR.n1906 VPWR.n1905 9.33404
R12918 VPWR.n1912 VPWR.n1911 9.33404
R12919 VPWR.n1916 VPWR.n1915 9.33404
R12920 VPWR.n1922 VPWR.n1921 9.33404
R12921 VPWR.n1925 VPWR.n1924 9.33404
R12922 VPWR.n1872 VPWR.n1871 9.33404
R12923 VPWR.n896 VPWR.n895 9.33404
R12924 VPWR.n892 VPWR.n891 9.33404
R12925 VPWR.n888 VPWR.n887 9.33404
R12926 VPWR.n884 VPWR.n883 9.33404
R12927 VPWR.n876 VPWR.n875 9.33404
R12928 VPWR.n872 VPWR.n871 9.33404
R12929 VPWR.n868 VPWR.n867 9.33404
R12930 VPWR.n864 VPWR.n863 9.33404
R12931 VPWR.n860 VPWR.n859 9.33404
R12932 VPWR.n856 VPWR.n855 9.33404
R12933 VPWR.n852 VPWR.n851 9.33404
R12934 VPWR.n848 VPWR.n847 9.33404
R12935 VPWR.n844 VPWR.n843 9.33404
R12936 VPWR.n840 VPWR.n839 9.33404
R12937 VPWR.n837 VPWR.n836 9.33404
R12938 VPWR.n880 VPWR.n879 9.33404
R12939 VPWR.n1807 VPWR.n1806 9.33404
R12940 VPWR.n949 VPWR.n948 9.33404
R12941 VPWR.n1473 VPWR.n1472 9.33404
R12942 VPWR.n369 VPWR.n368 9.33404
R12943 VPWR.n2401 VPWR.n2400 9.33404
R12944 VPWR.n308 VPWR.n307 9.33404
R12945 VPWR.n945 VPWR.n944 9.33404
R12946 VPWR.n1469 VPWR.n1468 9.33404
R12947 VPWR.n1803 VPWR.n1802 9.33404
R12948 VPWR.n953 VPWR.n952 9.33404
R12949 VPWR.n1483 VPWR.n1482 9.33404
R12950 VPWR.n377 VPWR.n376 9.33404
R12951 VPWR.n385 VPWR.n384 9.33404
R12952 VPWR.n389 VPWR.n388 9.33404
R12953 VPWR.n393 VPWR.n392 9.33404
R12954 VPWR.n397 VPWR.n396 9.33404
R12955 VPWR.n401 VPWR.n400 9.33404
R12956 VPWR.n405 VPWR.n404 9.33404
R12957 VPWR.n409 VPWR.n408 9.33404
R12958 VPWR.n413 VPWR.n412 9.33404
R12959 VPWR.n416 VPWR.n415 9.33404
R12960 VPWR.n381 VPWR.n380 9.33404
R12961 VPWR.n2385 VPWR.n2384 9.33404
R12962 VPWR.n296 VPWR.n295 9.33404
R12963 VPWR.n957 VPWR.n956 9.33404
R12964 VPWR.n1487 VPWR.n1486 9.33404
R12965 VPWR.n1797 VPWR.n1796 9.33404
R12966 VPWR.n1787 VPWR.n1786 9.33404
R12967 VPWR.n1783 VPWR.n1782 9.33404
R12968 VPWR.n1777 VPWR.n1776 9.33404
R12969 VPWR.n1773 VPWR.n1772 9.33404
R12970 VPWR.n1767 VPWR.n1766 9.33404
R12971 VPWR.n1763 VPWR.n1762 9.33404
R12972 VPWR.n1757 VPWR.n1756 9.33404
R12973 VPWR.n1754 VPWR.n1753 9.33404
R12974 VPWR.n1793 VPWR.n1792 9.33404
R12975 VPWR.n961 VPWR.n960 9.33404
R12976 VPWR.n1497 VPWR.n1496 9.33404
R12977 VPWR.n2405 VPWR.n2404 9.33404
R12978 VPWR.n312 VPWR.n311 9.33404
R12979 VPWR.n1460 VPWR.n1459 9.33404
R12980 VPWR.n965 VPWR.n964 9.33404
R12981 VPWR.n1501 VPWR.n1500 9.33404
R12982 VPWR.n2375 VPWR.n2374 9.33404
R12983 VPWR.n2365 VPWR.n2364 9.33404
R12984 VPWR.n2361 VPWR.n2360 9.33404
R12985 VPWR.n2355 VPWR.n2354 9.33404
R12986 VPWR.n2351 VPWR.n2350 9.33404
R12987 VPWR.n2345 VPWR.n2344 9.33404
R12988 VPWR.n2342 VPWR.n2341 9.33404
R12989 VPWR.n2371 VPWR.n2370 9.33404
R12990 VPWR.n284 VPWR.n283 9.33404
R12991 VPWR.n1516 VPWR.n1515 9.33404
R12992 VPWR.n969 VPWR.n968 9.33404
R12993 VPWR.n973 VPWR.n972 9.33404
R12994 VPWR.n977 VPWR.n976 9.33404
R12995 VPWR.n981 VPWR.n980 9.33404
R12996 VPWR.n985 VPWR.n984 9.33404
R12997 VPWR.n989 VPWR.n988 9.33404
R12998 VPWR.n992 VPWR.n991 9.33404
R12999 VPWR.n937 VPWR.n936 9.33404
R13000 VPWR.n1456 VPWR.n1169 9.33404
R13001 VPWR.n280 VPWR.n279 9.33404
R13002 VPWR.n1699 VPWR.n1698 9.33404
R13003 VPWR.n276 VPWR.n275 9.33404
R13004 VPWR.n272 VPWR.n271 9.33404
R13005 VPWR.n264 VPWR.n263 9.33404
R13006 VPWR.n261 VPWR.n260 9.33404
R13007 VPWR.n268 VPWR.n267 9.33404
R13008 VPWR.n1687 VPWR.n1686 9.33404
R13009 VPWR.n1726 VPWR.n1725 9.33404
R13010 VPWR.n1729 VPWR.n1728 9.33404
R13011 VPWR.n1695 VPWR.n1694 9.33404
R13012 VPWR.n2650 VPWR 9.32394
R13013 VPWR.n2613 VPWR 9.32394
R13014 VPWR.n2576 VPWR 9.32394
R13015 VPWR VPWR.n2543 9.32394
R13016 VPWR.n18 VPWR.n17 9.3005
R13017 VPWR.n15 VPWR.n14 9.3005
R13018 VPWR.n13 VPWR.n2 9.3005
R13019 VPWR.n10 VPWR.n9 9.3005
R13020 VPWR.n8 VPWR.n3 9.3005
R13021 VPWR.n12 VPWR.n11 9.3005
R13022 VPWR.n16 VPWR.n0 9.3005
R13023 VPWR.n1193 VPWR.n1192 9.3005
R13024 VPWR.n1190 VPWR.n1189 9.3005
R13025 VPWR.n1188 VPWR.n1175 9.3005
R13026 VPWR.n1185 VPWR.n1183 9.3005
R13027 VPWR.n1182 VPWR.n1176 9.3005
R13028 VPWR.n1187 VPWR.n1186 9.3005
R13029 VPWR.n1191 VPWR.n1172 9.3005
R13030 VPWR.n1217 VPWR.n1216 9.3005
R13031 VPWR.n1211 VPWR.n1198 9.3005
R13032 VPWR.n1208 VPWR.n1206 9.3005
R13033 VPWR.n1205 VPWR.n1199 9.3005
R13034 VPWR.n1210 VPWR.n1209 9.3005
R13035 VPWR.n1213 VPWR.n1212 9.3005
R13036 VPWR.n1215 VPWR.n1195 9.3005
R13037 VPWR.n1240 VPWR.n1239 9.3005
R13038 VPWR.n1235 VPWR.n1222 9.3005
R13039 VPWR.n1232 VPWR.n1230 9.3005
R13040 VPWR.n1229 VPWR.n1223 9.3005
R13041 VPWR.n1234 VPWR.n1233 9.3005
R13042 VPWR.n1237 VPWR.n1236 9.3005
R13043 VPWR.n1238 VPWR.n1219 9.3005
R13044 VPWR.n1271 VPWR.n1242 9.3005
R13045 VPWR.n1270 VPWR.n1269 9.3005
R13046 VPWR.n1250 VPWR.n1249 9.3005
R13047 VPWR.n1252 VPWR.n1251 9.3005
R13048 VPWR.n1254 VPWR.n1248 9.3005
R13049 VPWR.n1256 VPWR.n1255 9.3005
R13050 VPWR.n1257 VPWR.n1247 9.3005
R13051 VPWR.n1259 VPWR.n1258 9.3005
R13052 VPWR.n1263 VPWR.n1244 9.3005
R13053 VPWR.n1265 VPWR.n1264 9.3005
R13054 VPWR.n1267 VPWR.n1266 9.3005
R13055 VPWR.n1273 VPWR.n1272 9.3005
R13056 VPWR.n1275 VPWR.n1274 9.3005
R13057 VPWR.n1314 VPWR.n1313 9.3005
R13058 VPWR.n1309 VPWR.n1277 9.3005
R13059 VPWR.n1308 VPWR.n1307 9.3005
R13060 VPWR.n1286 VPWR.n1285 9.3005
R13061 VPWR.n1288 VPWR.n1287 9.3005
R13062 VPWR.n1291 VPWR.n1281 9.3005
R13063 VPWR.n1293 VPWR.n1292 9.3005
R13064 VPWR.n1294 VPWR.n1280 9.3005
R13065 VPWR.n1296 VPWR.n1295 9.3005
R13066 VPWR.n1300 VPWR.n1279 9.3005
R13067 VPWR.n1302 VPWR.n1301 9.3005
R13068 VPWR.n1304 VPWR.n1303 9.3005
R13069 VPWR.n1311 VPWR.n1310 9.3005
R13070 VPWR.n1347 VPWR.n1346 9.3005
R13071 VPWR.n1325 VPWR.n1324 9.3005
R13072 VPWR.n1327 VPWR.n1326 9.3005
R13073 VPWR.n1330 VPWR.n1320 9.3005
R13074 VPWR.n1332 VPWR.n1331 9.3005
R13075 VPWR.n1333 VPWR.n1319 9.3005
R13076 VPWR.n1335 VPWR.n1334 9.3005
R13077 VPWR.n1339 VPWR.n1318 9.3005
R13078 VPWR.n1341 VPWR.n1340 9.3005
R13079 VPWR.n1343 VPWR.n1342 9.3005
R13080 VPWR.n1348 VPWR.n1316 9.3005
R13081 VPWR.n1350 VPWR.n1349 9.3005
R13082 VPWR.n1384 VPWR.n1383 9.3005
R13083 VPWR.n1362 VPWR.n1361 9.3005
R13084 VPWR.n1364 VPWR.n1363 9.3005
R13085 VPWR.n1367 VPWR.n1357 9.3005
R13086 VPWR.n1369 VPWR.n1368 9.3005
R13087 VPWR.n1370 VPWR.n1356 9.3005
R13088 VPWR.n1372 VPWR.n1371 9.3005
R13089 VPWR.n1376 VPWR.n1355 9.3005
R13090 VPWR.n1378 VPWR.n1377 9.3005
R13091 VPWR.n1380 VPWR.n1379 9.3005
R13092 VPWR.n2743 VPWR.n2742 9.3005
R13093 VPWR.n2744 VPWR.n2736 9.3005
R13094 VPWR.n2745 VPWR.n2735 9.3005
R13095 VPWR.n2746 VPWR.n2734 9.3005
R13096 VPWR.n2748 VPWR.n2747 9.3005
R13097 VPWR.n2732 VPWR.n2731 9.3005
R13098 VPWR.n2726 VPWR.n2725 9.3005
R13099 VPWR.n2727 VPWR.n2717 9.3005
R13100 VPWR.n2729 VPWR.n2728 9.3005
R13101 VPWR.n2730 VPWR.n2715 9.3005
R13102 VPWR.n2713 VPWR.n2712 9.3005
R13103 VPWR.n2711 VPWR.n2695 9.3005
R13104 VPWR.n2706 VPWR.n2705 9.3005
R13105 VPWR.n2707 VPWR.n2697 9.3005
R13106 VPWR.n2709 VPWR.n2708 9.3005
R13107 VPWR.n2693 VPWR.n2692 9.3005
R13108 VPWR.n2687 VPWR.n2686 9.3005
R13109 VPWR.n2688 VPWR.n2678 9.3005
R13110 VPWR.n2690 VPWR.n2689 9.3005
R13111 VPWR.n2691 VPWR.n2676 9.3005
R13112 VPWR.n2674 VPWR.n2673 9.3005
R13113 VPWR.n2654 VPWR.n2653 9.3005
R13114 VPWR.n2655 VPWR.n2649 9.3005
R13115 VPWR.n2657 VPWR.n2656 9.3005
R13116 VPWR.n2659 VPWR.n2647 9.3005
R13117 VPWR.n2661 VPWR.n2660 9.3005
R13118 VPWR.n2663 VPWR.n2662 9.3005
R13119 VPWR.n2664 VPWR.n2643 9.3005
R13120 VPWR.n2668 VPWR.n2667 9.3005
R13121 VPWR.n2669 VPWR.n2642 9.3005
R13122 VPWR.n2671 VPWR.n2670 9.3005
R13123 VPWR.n2672 VPWR.n2640 9.3005
R13124 VPWR.n2638 VPWR.n2637 9.3005
R13125 VPWR.n2618 VPWR.n2617 9.3005
R13126 VPWR.n2619 VPWR.n2612 9.3005
R13127 VPWR.n2621 VPWR.n2620 9.3005
R13128 VPWR.n2623 VPWR.n2609 9.3005
R13129 VPWR.n2625 VPWR.n2624 9.3005
R13130 VPWR.n2627 VPWR.n2626 9.3005
R13131 VPWR.n2628 VPWR.n2605 9.3005
R13132 VPWR.n2631 VPWR.n2630 9.3005
R13133 VPWR.n2632 VPWR.n2604 9.3005
R13134 VPWR.n2634 VPWR.n2633 9.3005
R13135 VPWR.n2635 VPWR.n2602 9.3005
R13136 VPWR.n2581 VPWR.n2580 9.3005
R13137 VPWR.n2582 VPWR.n2575 9.3005
R13138 VPWR.n2584 VPWR.n2583 9.3005
R13139 VPWR.n2586 VPWR.n2572 9.3005
R13140 VPWR.n2588 VPWR.n2587 9.3005
R13141 VPWR.n2590 VPWR.n2589 9.3005
R13142 VPWR.n2591 VPWR.n2568 9.3005
R13143 VPWR.n2594 VPWR.n2593 9.3005
R13144 VPWR.n2595 VPWR.n2567 9.3005
R13145 VPWR.n2597 VPWR.n2596 9.3005
R13146 VPWR.n2598 VPWR.n2565 9.3005
R13147 VPWR.n2563 VPWR.n2562 9.3005
R13148 VPWR.n2545 VPWR.n2544 9.3005
R13149 VPWR.n2547 VPWR.n2540 9.3005
R13150 VPWR.n2552 VPWR.n2551 9.3005
R13151 VPWR.n2553 VPWR.n2539 9.3005
R13152 VPWR.n2555 VPWR.n2554 9.3005
R13153 VPWR.n2557 VPWR.n2536 9.3005
R13154 VPWR.n2559 VPWR.n2558 9.3005
R13155 VPWR.n2561 VPWR.n2560 9.3005
R13156 VPWR.n2441 VPWR.n2440 9.3005
R13157 VPWR.n2505 VPWR.n2504 9.3005
R13158 VPWR.n2445 VPWR.n2444 9.3005
R13159 VPWR.n2489 VPWR.n2488 9.3005
R13160 VPWR.n2481 VPWR.n2480 9.3005
R13161 VPWR.n2469 VPWR.n2468 9.3005
R13162 VPWR.n2465 VPWR.n2464 9.3005
R13163 VPWR.n1151 VPWR.n1150 9.3005
R13164 VPWR.n2457 VPWR.n2456 9.3005
R13165 VPWR.n1155 VPWR.n1154 9.3005
R13166 VPWR.n1147 VPWR.n1146 9.3005
R13167 VPWR.n2477 VPWR.n2476 9.3005
R13168 VPWR.n1143 VPWR.n1142 9.3005
R13169 VPWR.n1139 VPWR.n1138 9.3005
R13170 VPWR.n2453 VPWR.n2452 9.3005
R13171 VPWR.n1159 VPWR.n1158 9.3005
R13172 VPWR.n1135 VPWR.n1134 9.3005
R13173 VPWR.n2493 VPWR.n2492 9.3005
R13174 VPWR.n1131 VPWR.n1130 9.3005
R13175 VPWR.n1163 VPWR.n1162 9.3005
R13176 VPWR.n2501 VPWR.n2500 9.3005
R13177 VPWR.n1127 VPWR.n1126 9.3005
R13178 VPWR.n1123 VPWR.n1122 9.3005
R13179 VPWR.n1678 VPWR.n1677 9.3005
R13180 VPWR.n1119 VPWR.n1118 9.3005
R13181 VPWR.n2513 VPWR.n2512 9.3005
R13182 VPWR.n2517 VPWR.n2516 9.3005
R13183 VPWR.n2528 VPWR.n2527 9.3005
R13184 VPWR.n2525 VPWR.n2524 9.3005
R13185 VPWR.n1674 VPWR.n1673 9.3005
R13186 VPWR.n1030 VPWR.n1029 9.3005
R13187 VPWR.n1167 VPWR.n1166 9.3005
R13188 VPWR.n1214 VPWR.n1213 8.28285
R13189 VPWR.n2710 VPWR.n2709 8.28285
R13190 VPWR.n1110 VPWR.n1109 8.25914
R13191 VPWR.n1665 VPWR.n1664 8.25914
R13192 VPWR.n250 VPWR.n110 8.25914
R13193 VPWR.n129 VPWR.n119 8.25914
R13194 VPWR.n1716 VPWR.n1715 7.91351
R13195 VPWR.n1707 VPWR.n1706 7.9105
R13196 VPWR.n1010 VPWR.n1009 7.9105
R13197 VPWR.n1524 VPWR.n1523 7.9105
R13198 VPWR.n1529 VPWR.n1528 7.9105
R13199 VPWR.n1534 VPWR.n1533 7.9105
R13200 VPWR.n1539 VPWR.n1538 7.9105
R13201 VPWR.n1544 VPWR.n1543 7.9105
R13202 VPWR.n1549 VPWR.n1548 7.9105
R13203 VPWR.n1554 VPWR.n1553 7.9105
R13204 VPWR.n1559 VPWR.n1558 7.9105
R13205 VPWR.n1564 VPWR.n1563 7.9105
R13206 VPWR.n1399 VPWR.n1398 7.9105
R13207 VPWR.n1394 VPWR.n1393 7.9105
R13208 VPWR.n1712 VPWR.n1711 7.9105
R13209 VPWR.n1720 VPWR.n1719 7.9105
R13210 VPWR.n251 VPWR.n250 7.9105
R13211 VPWR.n249 VPWR.n248 7.9105
R13212 VPWR.n239 VPWR.n238 7.9105
R13213 VPWR.n229 VPWR.n228 7.9105
R13214 VPWR.n219 VPWR.n218 7.9105
R13215 VPWR.n209 VPWR.n208 7.9105
R13216 VPWR.n199 VPWR.n198 7.9105
R13217 VPWR.n189 VPWR.n188 7.9105
R13218 VPWR.n179 VPWR.n178 7.9105
R13219 VPWR.n169 VPWR.n168 7.9105
R13220 VPWR.n159 VPWR.n158 7.9105
R13221 VPWR.n149 VPWR.n148 7.9105
R13222 VPWR.n139 VPWR.n138 7.9105
R13223 VPWR.n129 VPWR.n128 7.9105
R13224 VPWR.n1664 VPWR.n1663 7.9105
R13225 VPWR.n1654 VPWR.n1653 7.9105
R13226 VPWR.n1039 VPWR.n1035 7.9105
R13227 VPWR.n1079 VPWR.n1078 7.9105
R13228 VPWR.n1082 VPWR.n1081 7.9105
R13229 VPWR.n1085 VPWR.n1084 7.9105
R13230 VPWR.n1088 VPWR.n1087 7.9105
R13231 VPWR.n1091 VPWR.n1090 7.9105
R13232 VPWR.n1094 VPWR.n1093 7.9105
R13233 VPWR.n1097 VPWR.n1096 7.9105
R13234 VPWR.n1100 VPWR.n1099 7.9105
R13235 VPWR.n1103 VPWR.n1102 7.9105
R13236 VPWR.n1106 VPWR.n1105 7.9105
R13237 VPWR.n1109 VPWR.n1108 7.9105
R13238 VPWR.n26 VPWR.n24 7.86657
R13239 VPWR.n7 VPWR.n6 7.56315
R13240 VPWR.n1181 VPWR.n1180 7.56315
R13241 VPWR.n1204 VPWR.n1203 7.56315
R13242 VPWR.n1228 VPWR.n1227 7.56315
R13243 VPWR.n2741 VPWR.n2739 6.4511
R13244 VPWR.n2724 VPWR.n2721 6.4511
R13245 VPWR.n2704 VPWR.n2701 6.4511
R13246 VPWR.n2685 VPWR.n2682 6.4511
R13247 VPWR.n1301 VPWR.n1278 6.4005
R13248 VPWR.n1340 VPWR.n1317 6.4005
R13249 VPWR.n1377 VPWR.n1354 6.4005
R13250 VPWR.n2659 VPWR.n2658 6.4005
R13251 VPWR.n2629 VPWR.n2628 6.4005
R13252 VPWR.n2592 VPWR.n2591 6.4005
R13253 VPWR.n2558 VPWR.n2535 6.4005
R13254 VPWR.n1166 VPWR.n1116 6.04494
R13255 VPWR.n2441 VPWR.n99 6.04494
R13256 VPWR.n1450 VPWR.n1448 6.04494
R13257 VPWR.n319 VPWR.n258 6.04494
R13258 VPWR.n2504 VPWR.n68 6.04494
R13259 VPWR.n1512 VPWR.n1416 6.04494
R13260 VPWR.n316 VPWR.n314 6.04494
R13261 VPWR.n2444 VPWR.n98 6.04494
R13262 VPWR.n933 VPWR.n931 6.04494
R13263 VPWR.n2414 VPWR.n324 6.04494
R13264 VPWR.n2411 VPWR.n325 6.04494
R13265 VPWR.n288 VPWR.n286 6.04494
R13266 VPWR.n2489 VPWR.n75 6.04494
R13267 VPWR.n941 VPWR.n939 6.04494
R13268 VPWR.n2381 VPWR.n337 6.04494
R13269 VPWR.n292 VPWR.n290 6.04494
R13270 VPWR.n2480 VPWR.n80 6.04494
R13271 VPWR.n1826 VPWR.n900 6.04494
R13272 VPWR.n1823 VPWR.n901 6.04494
R13273 VPWR.n1816 VPWR.n904 6.04494
R13274 VPWR.n357 VPWR.n355 6.04494
R13275 VPWR.n361 VPWR.n359 6.04494
R13276 VPWR.n365 VPWR.n363 6.04494
R13277 VPWR.n2391 VPWR.n333 6.04494
R13278 VPWR.n300 VPWR.n298 6.04494
R13279 VPWR.n2468 VPWR.n86 6.04494
R13280 VPWR.n1813 VPWR.n905 6.04494
R13281 VPWR.n373 VPWR.n371 6.04494
R13282 VPWR.n2394 VPWR.n332 6.04494
R13283 VPWR.n304 VPWR.n302 6.04494
R13284 VPWR.n2465 VPWR.n87 6.04494
R13285 VPWR.n2244 VPWR.n449 6.04494
R13286 VPWR.n2247 VPWR.n448 6.04494
R13287 VPWR.n2254 VPWR.n445 6.04494
R13288 VPWR.n2257 VPWR.n444 6.04494
R13289 VPWR.n2267 VPWR.n440 6.04494
R13290 VPWR.n2274 VPWR.n437 6.04494
R13291 VPWR.n2277 VPWR.n436 6.04494
R13292 VPWR.n2284 VPWR.n433 6.04494
R13293 VPWR.n2287 VPWR.n432 6.04494
R13294 VPWR.n2294 VPWR.n429 6.04494
R13295 VPWR.n2297 VPWR.n428 6.04494
R13296 VPWR.n2304 VPWR.n425 6.04494
R13297 VPWR.n2307 VPWR.n424 6.04494
R13298 VPWR.n2314 VPWR.n421 6.04494
R13299 VPWR.n2316 VPWR.n420 6.04494
R13300 VPWR.n2264 VPWR.n441 6.04494
R13301 VPWR.n511 VPWR.n450 6.04494
R13302 VPWR.n508 VPWR.n506 6.04494
R13303 VPWR.n504 VPWR.n502 6.04494
R13304 VPWR.n500 VPWR.n498 6.04494
R13305 VPWR.n492 VPWR.n490 6.04494
R13306 VPWR.n488 VPWR.n486 6.04494
R13307 VPWR.n484 VPWR.n482 6.04494
R13308 VPWR.n480 VPWR.n478 6.04494
R13309 VPWR.n476 VPWR.n474 6.04494
R13310 VPWR.n472 VPWR.n470 6.04494
R13311 VPWR.n468 VPWR.n466 6.04494
R13312 VPWR.n464 VPWR.n462 6.04494
R13313 VPWR.n460 VPWR.n458 6.04494
R13314 VPWR.n456 VPWR.n454 6.04494
R13315 VPWR.n453 VPWR.n451 6.04494
R13316 VPWR.n496 VPWR.n494 6.04494
R13317 VPWR.n2218 VPWR.n516 6.04494
R13318 VPWR.n2215 VPWR.n517 6.04494
R13319 VPWR.n2208 VPWR.n520 6.04494
R13320 VPWR.n2205 VPWR.n521 6.04494
R13321 VPWR.n2195 VPWR.n525 6.04494
R13322 VPWR.n2188 VPWR.n528 6.04494
R13323 VPWR.n2185 VPWR.n529 6.04494
R13324 VPWR.n2178 VPWR.n532 6.04494
R13325 VPWR.n2175 VPWR.n533 6.04494
R13326 VPWR.n2168 VPWR.n536 6.04494
R13327 VPWR.n2165 VPWR.n537 6.04494
R13328 VPWR.n2158 VPWR.n540 6.04494
R13329 VPWR.n2155 VPWR.n541 6.04494
R13330 VPWR.n2148 VPWR.n544 6.04494
R13331 VPWR.n2146 VPWR.n545 6.04494
R13332 VPWR.n2198 VPWR.n524 6.04494
R13333 VPWR.n549 VPWR.n547 6.04494
R13334 VPWR.n553 VPWR.n551 6.04494
R13335 VPWR.n557 VPWR.n555 6.04494
R13336 VPWR.n561 VPWR.n559 6.04494
R13337 VPWR.n569 VPWR.n567 6.04494
R13338 VPWR.n573 VPWR.n571 6.04494
R13339 VPWR.n577 VPWR.n575 6.04494
R13340 VPWR.n581 VPWR.n579 6.04494
R13341 VPWR.n585 VPWR.n583 6.04494
R13342 VPWR.n589 VPWR.n587 6.04494
R13343 VPWR.n593 VPWR.n591 6.04494
R13344 VPWR.n597 VPWR.n595 6.04494
R13345 VPWR.n601 VPWR.n599 6.04494
R13346 VPWR.n605 VPWR.n603 6.04494
R13347 VPWR.n607 VPWR.n546 6.04494
R13348 VPWR.n565 VPWR.n563 6.04494
R13349 VPWR.n2048 VPWR.n641 6.04494
R13350 VPWR.n2051 VPWR.n640 6.04494
R13351 VPWR.n2058 VPWR.n637 6.04494
R13352 VPWR.n2061 VPWR.n636 6.04494
R13353 VPWR.n2071 VPWR.n632 6.04494
R13354 VPWR.n2078 VPWR.n629 6.04494
R13355 VPWR.n2081 VPWR.n628 6.04494
R13356 VPWR.n2088 VPWR.n625 6.04494
R13357 VPWR.n2091 VPWR.n624 6.04494
R13358 VPWR.n2098 VPWR.n621 6.04494
R13359 VPWR.n2101 VPWR.n620 6.04494
R13360 VPWR.n2108 VPWR.n617 6.04494
R13361 VPWR.n2111 VPWR.n616 6.04494
R13362 VPWR.n2118 VPWR.n613 6.04494
R13363 VPWR.n2120 VPWR.n612 6.04494
R13364 VPWR.n2068 VPWR.n633 6.04494
R13365 VPWR.n703 VPWR.n642 6.04494
R13366 VPWR.n700 VPWR.n698 6.04494
R13367 VPWR.n696 VPWR.n694 6.04494
R13368 VPWR.n692 VPWR.n690 6.04494
R13369 VPWR.n684 VPWR.n682 6.04494
R13370 VPWR.n680 VPWR.n678 6.04494
R13371 VPWR.n676 VPWR.n674 6.04494
R13372 VPWR.n672 VPWR.n670 6.04494
R13373 VPWR.n668 VPWR.n666 6.04494
R13374 VPWR.n664 VPWR.n662 6.04494
R13375 VPWR.n660 VPWR.n658 6.04494
R13376 VPWR.n656 VPWR.n654 6.04494
R13377 VPWR.n652 VPWR.n650 6.04494
R13378 VPWR.n648 VPWR.n646 6.04494
R13379 VPWR.n645 VPWR.n643 6.04494
R13380 VPWR.n688 VPWR.n686 6.04494
R13381 VPWR.n2022 VPWR.n708 6.04494
R13382 VPWR.n2019 VPWR.n709 6.04494
R13383 VPWR.n2012 VPWR.n712 6.04494
R13384 VPWR.n2009 VPWR.n713 6.04494
R13385 VPWR.n1999 VPWR.n717 6.04494
R13386 VPWR.n1992 VPWR.n720 6.04494
R13387 VPWR.n1989 VPWR.n721 6.04494
R13388 VPWR.n1982 VPWR.n724 6.04494
R13389 VPWR.n1979 VPWR.n725 6.04494
R13390 VPWR.n1972 VPWR.n728 6.04494
R13391 VPWR.n1969 VPWR.n729 6.04494
R13392 VPWR.n1962 VPWR.n732 6.04494
R13393 VPWR.n1959 VPWR.n733 6.04494
R13394 VPWR.n1952 VPWR.n736 6.04494
R13395 VPWR.n1950 VPWR.n737 6.04494
R13396 VPWR.n2002 VPWR.n716 6.04494
R13397 VPWR.n741 VPWR.n739 6.04494
R13398 VPWR.n745 VPWR.n743 6.04494
R13399 VPWR.n749 VPWR.n747 6.04494
R13400 VPWR.n753 VPWR.n751 6.04494
R13401 VPWR.n761 VPWR.n759 6.04494
R13402 VPWR.n765 VPWR.n763 6.04494
R13403 VPWR.n769 VPWR.n767 6.04494
R13404 VPWR.n773 VPWR.n771 6.04494
R13405 VPWR.n777 VPWR.n775 6.04494
R13406 VPWR.n781 VPWR.n779 6.04494
R13407 VPWR.n785 VPWR.n783 6.04494
R13408 VPWR.n789 VPWR.n787 6.04494
R13409 VPWR.n793 VPWR.n791 6.04494
R13410 VPWR.n797 VPWR.n795 6.04494
R13411 VPWR.n799 VPWR.n738 6.04494
R13412 VPWR.n757 VPWR.n755 6.04494
R13413 VPWR.n1852 VPWR.n833 6.04494
R13414 VPWR.n1855 VPWR.n832 6.04494
R13415 VPWR.n1862 VPWR.n829 6.04494
R13416 VPWR.n1865 VPWR.n828 6.04494
R13417 VPWR.n1875 VPWR.n824 6.04494
R13418 VPWR.n1882 VPWR.n821 6.04494
R13419 VPWR.n1885 VPWR.n820 6.04494
R13420 VPWR.n1892 VPWR.n817 6.04494
R13421 VPWR.n1895 VPWR.n816 6.04494
R13422 VPWR.n1902 VPWR.n813 6.04494
R13423 VPWR.n1905 VPWR.n812 6.04494
R13424 VPWR.n1912 VPWR.n809 6.04494
R13425 VPWR.n1915 VPWR.n808 6.04494
R13426 VPWR.n1922 VPWR.n805 6.04494
R13427 VPWR.n1924 VPWR.n804 6.04494
R13428 VPWR.n1872 VPWR.n825 6.04494
R13429 VPWR.n895 VPWR.n834 6.04494
R13430 VPWR.n892 VPWR.n890 6.04494
R13431 VPWR.n888 VPWR.n886 6.04494
R13432 VPWR.n884 VPWR.n882 6.04494
R13433 VPWR.n876 VPWR.n874 6.04494
R13434 VPWR.n872 VPWR.n870 6.04494
R13435 VPWR.n868 VPWR.n866 6.04494
R13436 VPWR.n864 VPWR.n862 6.04494
R13437 VPWR.n860 VPWR.n858 6.04494
R13438 VPWR.n856 VPWR.n854 6.04494
R13439 VPWR.n852 VPWR.n850 6.04494
R13440 VPWR.n848 VPWR.n846 6.04494
R13441 VPWR.n844 VPWR.n842 6.04494
R13442 VPWR.n840 VPWR.n838 6.04494
R13443 VPWR.n837 VPWR.n835 6.04494
R13444 VPWR.n880 VPWR.n878 6.04494
R13445 VPWR.n1806 VPWR.n908 6.04494
R13446 VPWR.n949 VPWR.n947 6.04494
R13447 VPWR.n1472 VPWR.n1436 6.04494
R13448 VPWR.n1151 VPWR.n1149 6.04494
R13449 VPWR.n369 VPWR.n367 6.04494
R13450 VPWR.n2401 VPWR.n329 6.04494
R13451 VPWR.n308 VPWR.n306 6.04494
R13452 VPWR.n2456 VPWR.n92 6.04494
R13453 VPWR.n945 VPWR.n943 6.04494
R13454 VPWR.n1469 VPWR.n1440 6.04494
R13455 VPWR.n1155 VPWR.n1153 6.04494
R13456 VPWR.n1803 VPWR.n909 6.04494
R13457 VPWR.n953 VPWR.n951 6.04494
R13458 VPWR.n1483 VPWR.n1432 6.04494
R13459 VPWR.n1147 VPWR.n1145 6.04494
R13460 VPWR.n377 VPWR.n375 6.04494
R13461 VPWR.n385 VPWR.n383 6.04494
R13462 VPWR.n389 VPWR.n387 6.04494
R13463 VPWR.n393 VPWR.n391 6.04494
R13464 VPWR.n397 VPWR.n395 6.04494
R13465 VPWR.n401 VPWR.n399 6.04494
R13466 VPWR.n405 VPWR.n403 6.04494
R13467 VPWR.n409 VPWR.n407 6.04494
R13468 VPWR.n413 VPWR.n411 6.04494
R13469 VPWR.n415 VPWR.n354 6.04494
R13470 VPWR.n381 VPWR.n379 6.04494
R13471 VPWR.n2384 VPWR.n336 6.04494
R13472 VPWR.n296 VPWR.n294 6.04494
R13473 VPWR.n2477 VPWR.n81 6.04494
R13474 VPWR.n957 VPWR.n955 6.04494
R13475 VPWR.n1486 VPWR.n1428 6.04494
R13476 VPWR.n1143 VPWR.n1141 6.04494
R13477 VPWR.n1796 VPWR.n912 6.04494
R13478 VPWR.n1786 VPWR.n916 6.04494
R13479 VPWR.n1783 VPWR.n917 6.04494
R13480 VPWR.n1776 VPWR.n920 6.04494
R13481 VPWR.n1773 VPWR.n921 6.04494
R13482 VPWR.n1766 VPWR.n924 6.04494
R13483 VPWR.n1763 VPWR.n925 6.04494
R13484 VPWR.n1756 VPWR.n928 6.04494
R13485 VPWR.n1754 VPWR.n929 6.04494
R13486 VPWR.n1793 VPWR.n913 6.04494
R13487 VPWR.n961 VPWR.n959 6.04494
R13488 VPWR.n1497 VPWR.n1424 6.04494
R13489 VPWR.n1139 VPWR.n1137 6.04494
R13490 VPWR.n2404 VPWR.n328 6.04494
R13491 VPWR.n312 VPWR.n310 6.04494
R13492 VPWR.n2453 VPWR.n93 6.04494
R13493 VPWR.n1459 VPWR.n1444 6.04494
R13494 VPWR.n1159 VPWR.n1157 6.04494
R13495 VPWR.n965 VPWR.n963 6.04494
R13496 VPWR.n1500 VPWR.n1420 6.04494
R13497 VPWR.n1135 VPWR.n1133 6.04494
R13498 VPWR.n2374 VPWR.n340 6.04494
R13499 VPWR.n2364 VPWR.n344 6.04494
R13500 VPWR.n2361 VPWR.n345 6.04494
R13501 VPWR.n2354 VPWR.n348 6.04494
R13502 VPWR.n2351 VPWR.n349 6.04494
R13503 VPWR.n2344 VPWR.n352 6.04494
R13504 VPWR.n2342 VPWR.n353 6.04494
R13505 VPWR.n2371 VPWR.n341 6.04494
R13506 VPWR.n284 VPWR.n282 6.04494
R13507 VPWR.n2492 VPWR.n74 6.04494
R13508 VPWR.n1515 VPWR.n1412 6.04494
R13509 VPWR.n1131 VPWR.n1129 6.04494
R13510 VPWR.n969 VPWR.n967 6.04494
R13511 VPWR.n973 VPWR.n971 6.04494
R13512 VPWR.n977 VPWR.n975 6.04494
R13513 VPWR.n981 VPWR.n979 6.04494
R13514 VPWR.n985 VPWR.n983 6.04494
R13515 VPWR.n989 VPWR.n987 6.04494
R13516 VPWR.n991 VPWR.n930 6.04494
R13517 VPWR.n937 VPWR.n935 6.04494
R13518 VPWR.n1456 VPWR.n1455 6.04494
R13519 VPWR.n1163 VPWR.n1161 6.04494
R13520 VPWR.n280 VPWR.n278 6.04494
R13521 VPWR.n2501 VPWR.n69 6.04494
R13522 VPWR.n1127 VPWR.n1125 6.04494
R13523 VPWR.n1698 VPWR.n1017 6.04494
R13524 VPWR.n1123 VPWR.n1121 6.04494
R13525 VPWR.n276 VPWR.n274 6.04494
R13526 VPWR.n272 VPWR.n270 6.04494
R13527 VPWR.n264 VPWR.n262 6.04494
R13528 VPWR.n261 VPWR.n259 6.04494
R13529 VPWR.n268 VPWR.n266 6.04494
R13530 VPWR.n1677 VPWR.n1026 6.04494
R13531 VPWR.n1686 VPWR.n1684 6.04494
R13532 VPWR.n1726 VPWR.n1004 6.04494
R13533 VPWR.n1728 VPWR.n1000 6.04494
R13534 VPWR.n1695 VPWR.n1021 6.04494
R13535 VPWR.n1119 VPWR.n1117 6.04494
R13536 VPWR.n2513 VPWR.n63 6.04494
R13537 VPWR.n2516 VPWR.n62 6.04494
R13538 VPWR.n2525 VPWR.n57 6.04494
R13539 VPWR.n2527 VPWR.n56 6.04494
R13540 VPWR.n1674 VPWR.n1027 6.04494
R13541 VPWR.n1029 VPWR.n1028 6.04494
R13542 VPWR.n2721 VPWR.n2720 5.39628
R13543 VPWR.n2701 VPWR.n2700 5.39628
R13544 VPWR.n2682 VPWR.n2681 5.39628
R13545 VPWR.n54 VPWR 4.71698
R13546 VPWR.n52 VPWR 4.71698
R13547 VPWR.n50 VPWR 4.71698
R13548 VPWR.n48 VPWR 4.71698
R13549 VPWR.n46 VPWR 4.71698
R13550 VPWR.n44 VPWR 4.71698
R13551 VPWR.n42 VPWR 4.71698
R13552 VPWR.n40 VPWR 4.71698
R13553 VPWR.n38 VPWR 4.71698
R13554 VPWR.n36 VPWR 4.71698
R13555 VPWR.n34 VPWR 4.71698
R13556 VPWR.n32 VPWR 4.71698
R13557 VPWR.n30 VPWR 4.71698
R13558 VPWR.n28 VPWR 4.71698
R13559 VPWR.n26 VPWR 4.71698
R13560 VPWR.n1385 VPWR.n1384 4.55954
R13561 VPWR.n2507 VPWR.n2506 4.5005
R13562 VPWR.n2447 VPWR.n2446 4.5005
R13563 VPWR.n2487 VPWR.n2486 4.5005
R13564 VPWR.n287 VPWR.n77 4.5005
R13565 VPWR.n2483 VPWR.n2482 4.5005
R13566 VPWR.n291 VPWR.n78 4.5005
R13567 VPWR.n2471 VPWR.n2470 4.5005
R13568 VPWR.n299 VPWR.n84 4.5005
R13569 VPWR.n2390 VPWR.n2389 4.5005
R13570 VPWR.n2463 VPWR.n2462 4.5005
R13571 VPWR.n303 VPWR.n89 4.5005
R13572 VPWR.n2396 VPWR.n2395 4.5005
R13573 VPWR.n1476 VPWR.n1063 4.5005
R13574 VPWR.n1475 VPWR.n1473 4.5005
R13575 VPWR.n948 VPWR.n907 4.5005
R13576 VPWR.n1808 VPWR.n1807 4.5005
R13577 VPWR.n879 VPWR.n826 4.5005
R13578 VPWR.n1871 VPWR.n1870 4.5005
R13579 VPWR.n756 VPWR.n715 4.5005
R13580 VPWR.n2004 VPWR.n2003 4.5005
R13581 VPWR.n687 VPWR.n634 4.5005
R13582 VPWR.n2067 VPWR.n2066 4.5005
R13583 VPWR.n564 VPWR.n523 4.5005
R13584 VPWR.n2200 VPWR.n2199 4.5005
R13585 VPWR.n495 VPWR.n442 4.5005
R13586 VPWR.n2263 VPWR.n2262 4.5005
R13587 VPWR.n372 VPWR.n331 4.5005
R13588 VPWR.n2459 VPWR.n2458 4.5005
R13589 VPWR.n307 VPWR.n90 4.5005
R13590 VPWR.n2400 VPWR.n2399 4.5005
R13591 VPWR.n368 VPWR.n330 4.5005
R13592 VPWR.n2259 VPWR.n2258 4.5005
R13593 VPWR.n499 VPWR.n443 4.5005
R13594 VPWR.n2204 VPWR.n2203 4.5005
R13595 VPWR.n560 VPWR.n522 4.5005
R13596 VPWR.n2063 VPWR.n2062 4.5005
R13597 VPWR.n691 VPWR.n635 4.5005
R13598 VPWR.n2008 VPWR.n2007 4.5005
R13599 VPWR.n752 VPWR.n714 4.5005
R13600 VPWR.n1867 VPWR.n1866 4.5005
R13601 VPWR.n883 VPWR.n827 4.5005
R13602 VPWR.n1465 VPWR.n1066 4.5005
R13603 VPWR.n1468 VPWR.n1467 4.5005
R13604 VPWR.n944 VPWR.n906 4.5005
R13605 VPWR.n1812 VPWR.n1811 4.5005
R13606 VPWR.n1479 VPWR.n1060 4.5005
R13607 VPWR.n1482 VPWR.n1481 4.5005
R13608 VPWR.n952 VPWR.n910 4.5005
R13609 VPWR.n1802 VPWR.n1801 4.5005
R13610 VPWR.n875 VPWR.n823 4.5005
R13611 VPWR.n1877 VPWR.n1876 4.5005
R13612 VPWR.n760 VPWR.n718 4.5005
R13613 VPWR.n1998 VPWR.n1997 4.5005
R13614 VPWR.n683 VPWR.n631 4.5005
R13615 VPWR.n2073 VPWR.n2072 4.5005
R13616 VPWR.n568 VPWR.n526 4.5005
R13617 VPWR.n2194 VPWR.n2193 4.5005
R13618 VPWR.n491 VPWR.n439 4.5005
R13619 VPWR.n2269 VPWR.n2268 4.5005
R13620 VPWR.n376 VPWR.n334 4.5005
R13621 VPWR.n2475 VPWR.n2474 4.5005
R13622 VPWR.n295 VPWR.n83 4.5005
R13623 VPWR.n2386 VPWR.n2385 4.5005
R13624 VPWR.n380 VPWR.n335 4.5005
R13625 VPWR.n2273 VPWR.n2272 4.5005
R13626 VPWR.n487 VPWR.n438 4.5005
R13627 VPWR.n2190 VPWR.n2189 4.5005
R13628 VPWR.n572 VPWR.n527 4.5005
R13629 VPWR.n2077 VPWR.n2076 4.5005
R13630 VPWR.n679 VPWR.n630 4.5005
R13631 VPWR.n1994 VPWR.n1993 4.5005
R13632 VPWR.n764 VPWR.n719 4.5005
R13633 VPWR.n1881 VPWR.n1880 4.5005
R13634 VPWR.n871 VPWR.n822 4.5005
R13635 VPWR.n1490 VPWR.n1057 4.5005
R13636 VPWR.n1489 VPWR.n1487 4.5005
R13637 VPWR.n956 VPWR.n911 4.5005
R13638 VPWR.n1798 VPWR.n1797 4.5005
R13639 VPWR.n1493 VPWR.n1054 4.5005
R13640 VPWR.n1496 VPWR.n1495 4.5005
R13641 VPWR.n960 VPWR.n914 4.5005
R13642 VPWR.n1792 VPWR.n1791 4.5005
R13643 VPWR.n867 VPWR.n819 4.5005
R13644 VPWR.n1887 VPWR.n1886 4.5005
R13645 VPWR.n768 VPWR.n722 4.5005
R13646 VPWR.n1988 VPWR.n1987 4.5005
R13647 VPWR.n675 VPWR.n627 4.5005
R13648 VPWR.n2083 VPWR.n2082 4.5005
R13649 VPWR.n576 VPWR.n530 4.5005
R13650 VPWR.n2184 VPWR.n2183 4.5005
R13651 VPWR.n483 VPWR.n435 4.5005
R13652 VPWR.n2279 VPWR.n2278 4.5005
R13653 VPWR.n384 VPWR.n338 4.5005
R13654 VPWR.n2380 VPWR.n2379 4.5005
R13655 VPWR.n2451 VPWR.n2450 4.5005
R13656 VPWR.n311 VPWR.n95 4.5005
R13657 VPWR.n2406 VPWR.n2405 4.5005
R13658 VPWR.n364 VPWR.n327 4.5005
R13659 VPWR.n2253 VPWR.n2252 4.5005
R13660 VPWR.n503 VPWR.n446 4.5005
R13661 VPWR.n2210 VPWR.n2209 4.5005
R13662 VPWR.n556 VPWR.n519 4.5005
R13663 VPWR.n2057 VPWR.n2056 4.5005
R13664 VPWR.n695 VPWR.n638 4.5005
R13665 VPWR.n2014 VPWR.n2013 4.5005
R13666 VPWR.n748 VPWR.n711 4.5005
R13667 VPWR.n1861 VPWR.n1860 4.5005
R13668 VPWR.n887 VPWR.n830 4.5005
R13669 VPWR.n1818 VPWR.n1817 4.5005
R13670 VPWR.n1462 VPWR.n1069 4.5005
R13671 VPWR.n1461 VPWR.n1460 4.5005
R13672 VPWR.n940 VPWR.n903 4.5005
R13673 VPWR.n1504 VPWR.n1051 4.5005
R13674 VPWR.n1503 VPWR.n1501 4.5005
R13675 VPWR.n964 VPWR.n915 4.5005
R13676 VPWR.n1788 VPWR.n1787 4.5005
R13677 VPWR.n863 VPWR.n818 4.5005
R13678 VPWR.n1891 VPWR.n1890 4.5005
R13679 VPWR.n772 VPWR.n723 4.5005
R13680 VPWR.n1984 VPWR.n1983 4.5005
R13681 VPWR.n671 VPWR.n626 4.5005
R13682 VPWR.n2087 VPWR.n2086 4.5005
R13683 VPWR.n580 VPWR.n531 4.5005
R13684 VPWR.n2180 VPWR.n2179 4.5005
R13685 VPWR.n479 VPWR.n434 4.5005
R13686 VPWR.n2283 VPWR.n2282 4.5005
R13687 VPWR.n388 VPWR.n339 4.5005
R13688 VPWR.n2376 VPWR.n2375 4.5005
R13689 VPWR.n2495 VPWR.n2494 4.5005
R13690 VPWR.n283 VPWR.n72 4.5005
R13691 VPWR.n2370 VPWR.n2369 4.5005
R13692 VPWR.n392 VPWR.n342 4.5005
R13693 VPWR.n2289 VPWR.n2288 4.5005
R13694 VPWR.n475 VPWR.n431 4.5005
R13695 VPWR.n2174 VPWR.n2173 4.5005
R13696 VPWR.n584 VPWR.n534 4.5005
R13697 VPWR.n2093 VPWR.n2092 4.5005
R13698 VPWR.n667 VPWR.n623 4.5005
R13699 VPWR.n1978 VPWR.n1977 4.5005
R13700 VPWR.n776 VPWR.n726 4.5005
R13701 VPWR.n1897 VPWR.n1896 4.5005
R13702 VPWR.n859 VPWR.n815 4.5005
R13703 VPWR.n1782 VPWR.n1781 4.5005
R13704 VPWR.n1408 VPWR.n1048 4.5005
R13705 VPWR.n1517 VPWR.n1516 4.5005
R13706 VPWR.n968 VPWR.n918 4.5005
R13707 VPWR.n1569 VPWR.n1072 4.5005
R13708 VPWR.n1568 VPWR.n1169 4.5005
R13709 VPWR.n936 VPWR.n902 4.5005
R13710 VPWR.n1822 VPWR.n1821 4.5005
R13711 VPWR.n891 VPWR.n831 4.5005
R13712 VPWR.n1857 VPWR.n1856 4.5005
R13713 VPWR.n744 VPWR.n710 4.5005
R13714 VPWR.n2018 VPWR.n2017 4.5005
R13715 VPWR.n699 VPWR.n639 4.5005
R13716 VPWR.n2053 VPWR.n2052 4.5005
R13717 VPWR.n552 VPWR.n518 4.5005
R13718 VPWR.n2214 VPWR.n2213 4.5005
R13719 VPWR.n507 VPWR.n447 4.5005
R13720 VPWR.n2249 VPWR.n2248 4.5005
R13721 VPWR.n360 VPWR.n326 4.5005
R13722 VPWR.n2410 VPWR.n2409 4.5005
R13723 VPWR.n315 VPWR.n96 4.5005
R13724 VPWR.n2499 VPWR.n2498 4.5005
R13725 VPWR.n279 VPWR.n71 4.5005
R13726 VPWR.n2366 VPWR.n2365 4.5005
R13727 VPWR.n396 VPWR.n343 4.5005
R13728 VPWR.n2293 VPWR.n2292 4.5005
R13729 VPWR.n471 VPWR.n430 4.5005
R13730 VPWR.n2170 VPWR.n2169 4.5005
R13731 VPWR.n588 VPWR.n535 4.5005
R13732 VPWR.n2097 VPWR.n2096 4.5005
R13733 VPWR.n663 VPWR.n622 4.5005
R13734 VPWR.n1974 VPWR.n1973 4.5005
R13735 VPWR.n780 VPWR.n727 4.5005
R13736 VPWR.n1901 VPWR.n1900 4.5005
R13737 VPWR.n855 VPWR.n814 4.5005
R13738 VPWR.n1778 VPWR.n1777 4.5005
R13739 VPWR.n972 VPWR.n919 4.5005
R13740 VPWR.n1509 VPWR.n1045 4.5005
R13741 VPWR.n1511 VPWR.n1510 4.5005
R13742 VPWR.n1042 VPWR.n1013 4.5005
R13743 VPWR.n1700 VPWR.n1699 4.5005
R13744 VPWR.n976 VPWR.n922 4.5005
R13745 VPWR.n1772 VPWR.n1771 4.5005
R13746 VPWR.n851 VPWR.n811 4.5005
R13747 VPWR.n1907 VPWR.n1906 4.5005
R13748 VPWR.n784 VPWR.n730 4.5005
R13749 VPWR.n1968 VPWR.n1967 4.5005
R13750 VPWR.n659 VPWR.n619 4.5005
R13751 VPWR.n2103 VPWR.n2102 4.5005
R13752 VPWR.n592 VPWR.n538 4.5005
R13753 VPWR.n2164 VPWR.n2163 4.5005
R13754 VPWR.n467 VPWR.n427 4.5005
R13755 VPWR.n2299 VPWR.n2298 4.5005
R13756 VPWR.n400 VPWR.n346 4.5005
R13757 VPWR.n2360 VPWR.n2359 4.5005
R13758 VPWR.n275 VPWR.n66 4.5005
R13759 VPWR.n267 VPWR.n60 4.5005
R13760 VPWR.n2350 VPWR.n2349 4.5005
R13761 VPWR.n408 VPWR.n350 4.5005
R13762 VPWR.n2309 VPWR.n2308 4.5005
R13763 VPWR.n459 VPWR.n423 4.5005
R13764 VPWR.n2154 VPWR.n2153 4.5005
R13765 VPWR.n600 VPWR.n542 4.5005
R13766 VPWR.n2113 VPWR.n2112 4.5005
R13767 VPWR.n651 VPWR.n615 4.5005
R13768 VPWR.n1958 VPWR.n1957 4.5005
R13769 VPWR.n792 VPWR.n734 4.5005
R13770 VPWR.n1917 VPWR.n1916 4.5005
R13771 VPWR.n843 VPWR.n807 4.5005
R13772 VPWR.n1762 VPWR.n1761 4.5005
R13773 VPWR.n984 VPWR.n926 4.5005
R13774 VPWR.n1689 VPWR.n1679 4.5005
R13775 VPWR.n1688 VPWR.n1687 4.5005
R13776 VPWR.n1692 VPWR.n1022 4.5005
R13777 VPWR.n1694 VPWR.n1693 4.5005
R13778 VPWR.n980 VPWR.n923 4.5005
R13779 VPWR.n1768 VPWR.n1767 4.5005
R13780 VPWR.n847 VPWR.n810 4.5005
R13781 VPWR.n1911 VPWR.n1910 4.5005
R13782 VPWR.n788 VPWR.n731 4.5005
R13783 VPWR.n1964 VPWR.n1963 4.5005
R13784 VPWR.n655 VPWR.n618 4.5005
R13785 VPWR.n2107 VPWR.n2106 4.5005
R13786 VPWR.n596 VPWR.n539 4.5005
R13787 VPWR.n2160 VPWR.n2159 4.5005
R13788 VPWR.n463 VPWR.n426 4.5005
R13789 VPWR.n2303 VPWR.n2302 4.5005
R13790 VPWR.n404 VPWR.n347 4.5005
R13791 VPWR.n2356 VPWR.n2355 4.5005
R13792 VPWR.n271 VPWR.n65 4.5005
R13793 VPWR.n2511 VPWR.n2510 4.5005
R13794 VPWR.n2519 VPWR.n2518 4.5005
R13795 VPWR.n2523 VPWR.n2522 4.5005
R13796 VPWR.n263 VPWR.n59 4.5005
R13797 VPWR.n2346 VPWR.n2345 4.5005
R13798 VPWR.n412 VPWR.n351 4.5005
R13799 VPWR.n2313 VPWR.n2312 4.5005
R13800 VPWR.n455 VPWR.n422 4.5005
R13801 VPWR.n2150 VPWR.n2149 4.5005
R13802 VPWR.n604 VPWR.n543 4.5005
R13803 VPWR.n2117 VPWR.n2116 4.5005
R13804 VPWR.n647 VPWR.n614 4.5005
R13805 VPWR.n1954 VPWR.n1953 4.5005
R13806 VPWR.n796 VPWR.n735 4.5005
R13807 VPWR.n1921 VPWR.n1920 4.5005
R13808 VPWR.n839 VPWR.n806 4.5005
R13809 VPWR.n1758 VPWR.n1757 4.5005
R13810 VPWR.n988 VPWR.n927 4.5005
R13811 VPWR.n1725 VPWR.n1724 4.5005
R13812 VPWR.n1672 VPWR.n1005 4.5005
R13813 VPWR.n1573 VPWR.n1572 4.5005
R13814 VPWR.n1449 VPWR.n1168 4.5005
R13815 VPWR.n932 VPWR.n899 4.5005
R13816 VPWR.n1828 VPWR.n1827 4.5005
R13817 VPWR.n897 VPWR.n896 4.5005
R13818 VPWR.n1851 VPWR.n1850 4.5005
R13819 VPWR.n740 VPWR.n707 4.5005
R13820 VPWR.n2024 VPWR.n2023 4.5005
R13821 VPWR.n705 VPWR.n704 4.5005
R13822 VPWR.n2047 VPWR.n2046 4.5005
R13823 VPWR.n548 VPWR.n515 4.5005
R13824 VPWR.n2220 VPWR.n2219 4.5005
R13825 VPWR.n513 VPWR.n512 4.5005
R13826 VPWR.n2243 VPWR.n2242 4.5005
R13827 VPWR.n356 VPWR.n323 4.5005
R13828 VPWR.n2416 VPWR.n2415 4.5005
R13829 VPWR.n321 VPWR.n320 4.5005
R13830 VPWR.n2439 VPWR.n2438 4.5005
R13831 VPWR.n2530 VPWR.n2529 4.5005
R13832 VPWR.n260 VPWR.n22 4.5005
R13833 VPWR.n2341 VPWR.n2340 4.5005
R13834 VPWR.n417 VPWR.n416 4.5005
R13835 VPWR.n2318 VPWR.n2317 4.5005
R13836 VPWR.n452 VPWR.n419 4.5005
R13837 VPWR.n2145 VPWR.n2144 4.5005
R13838 VPWR.n609 VPWR.n608 4.5005
R13839 VPWR.n2122 VPWR.n2121 4.5005
R13840 VPWR.n644 VPWR.n611 4.5005
R13841 VPWR.n1949 VPWR.n1948 4.5005
R13842 VPWR.n801 VPWR.n800 4.5005
R13843 VPWR.n1926 VPWR.n1925 4.5005
R13844 VPWR.n836 VPWR.n803 4.5005
R13845 VPWR.n1753 VPWR.n1752 4.5005
R13846 VPWR.n993 VPWR.n992 4.5005
R13847 VPWR.n1730 VPWR.n1729 4.5005
R13848 VPWR.n1031 VPWR.n996 4.5005
R13849 VPWR.n2564 VPWR 4.49965
R13850 VPWR.n19 VPWR.n18 4.20017
R13851 VPWR.n1194 VPWR.n1193 4.20017
R13852 VPWR.n1218 VPWR.n1217 4.20017
R13853 VPWR.n1241 VPWR.n1240 4.20017
R13854 VPWR.n1276 VPWR.n1275 4.20017
R13855 VPWR.n1315 VPWR.n1314 4.20017
R13856 VPWR.n1353 VPWR.n1352 4.20017
R13857 VPWR.n2749 VPWR 4.14027
R13858 VPWR.n2733 VPWR 4.14027
R13859 VPWR.n2714 VPWR 4.14027
R13860 VPWR.n2694 VPWR 4.14027
R13861 VPWR.n2675 VPWR 4.14027
R13862 VPWR.n2639 VPWR 4.14027
R13863 VPWR.n2601 VPWR 4.14027
R13864 VPWR.n55 VPWR.n54 4.00943
R13865 VPWR.n2652 VPWR.n2649 3.76521
R13866 VPWR.n2616 VPWR.n2612 3.76521
R13867 VPWR.n2579 VPWR.n2575 3.76521
R13868 VPWR.n2547 VPWR.n2546 3.76521
R13869 VPWR.n1842 VPWR.n826 3.4105
R13870 VPWR.n1870 VPWR.n1869 3.4105
R13871 VPWR.n1933 VPWR.n715 3.4105
R13872 VPWR.n2005 VPWR.n2004 3.4105
R13873 VPWR.n2038 VPWR.n634 3.4105
R13874 VPWR.n2066 VPWR.n2065 3.4105
R13875 VPWR.n2129 VPWR.n523 3.4105
R13876 VPWR.n2201 VPWR.n2200 3.4105
R13877 VPWR.n2234 VPWR.n442 3.4105
R13878 VPWR.n2262 VPWR.n2261 3.4105
R13879 VPWR.n2325 VPWR.n331 3.4105
R13880 VPWR.n2324 VPWR.n330 3.4105
R13881 VPWR.n2260 VPWR.n2259 3.4105
R13882 VPWR.n2235 VPWR.n443 3.4105
R13883 VPWR.n2203 VPWR.n2202 3.4105
R13884 VPWR.n2128 VPWR.n522 3.4105
R13885 VPWR.n2064 VPWR.n2063 3.4105
R13886 VPWR.n2039 VPWR.n635 3.4105
R13887 VPWR.n2007 VPWR.n2006 3.4105
R13888 VPWR.n1932 VPWR.n714 3.4105
R13889 VPWR.n1868 VPWR.n1867 3.4105
R13890 VPWR.n1843 VPWR.n827 3.4105
R13891 VPWR.n1811 VPWR.n1810 3.4105
R13892 VPWR.n1809 VPWR.n1808 3.4105
R13893 VPWR.n1801 VPWR.n1800 3.4105
R13894 VPWR.n1841 VPWR.n823 3.4105
R13895 VPWR.n1878 VPWR.n1877 3.4105
R13896 VPWR.n1934 VPWR.n718 3.4105
R13897 VPWR.n1997 VPWR.n1996 3.4105
R13898 VPWR.n2037 VPWR.n631 3.4105
R13899 VPWR.n2074 VPWR.n2073 3.4105
R13900 VPWR.n2130 VPWR.n526 3.4105
R13901 VPWR.n2193 VPWR.n2192 3.4105
R13902 VPWR.n2233 VPWR.n439 3.4105
R13903 VPWR.n2270 VPWR.n2269 3.4105
R13904 VPWR.n2326 VPWR.n334 3.4105
R13905 VPWR.n2327 VPWR.n335 3.4105
R13906 VPWR.n2272 VPWR.n2271 3.4105
R13907 VPWR.n2232 VPWR.n438 3.4105
R13908 VPWR.n2191 VPWR.n2190 3.4105
R13909 VPWR.n2131 VPWR.n527 3.4105
R13910 VPWR.n2076 VPWR.n2075 3.4105
R13911 VPWR.n2036 VPWR.n630 3.4105
R13912 VPWR.n1995 VPWR.n1994 3.4105
R13913 VPWR.n1935 VPWR.n719 3.4105
R13914 VPWR.n1880 VPWR.n1879 3.4105
R13915 VPWR.n1840 VPWR.n822 3.4105
R13916 VPWR.n1799 VPWR.n1798 3.4105
R13917 VPWR.n1791 VPWR.n1790 3.4105
R13918 VPWR.n1839 VPWR.n819 3.4105
R13919 VPWR.n1888 VPWR.n1887 3.4105
R13920 VPWR.n1936 VPWR.n722 3.4105
R13921 VPWR.n1987 VPWR.n1986 3.4105
R13922 VPWR.n2035 VPWR.n627 3.4105
R13923 VPWR.n2084 VPWR.n2083 3.4105
R13924 VPWR.n2132 VPWR.n530 3.4105
R13925 VPWR.n2183 VPWR.n2182 3.4105
R13926 VPWR.n2231 VPWR.n435 3.4105
R13927 VPWR.n2280 VPWR.n2279 3.4105
R13928 VPWR.n2328 VPWR.n338 3.4105
R13929 VPWR.n2379 VPWR.n2378 3.4105
R13930 VPWR.n2387 VPWR.n2386 3.4105
R13931 VPWR.n2389 VPWR.n2388 3.4105
R13932 VPWR.n2397 VPWR.n2396 3.4105
R13933 VPWR.n2399 VPWR.n2398 3.4105
R13934 VPWR.n2407 VPWR.n2406 3.4105
R13935 VPWR.n2323 VPWR.n327 3.4105
R13936 VPWR.n2252 VPWR.n2251 3.4105
R13937 VPWR.n2236 VPWR.n446 3.4105
R13938 VPWR.n2211 VPWR.n2210 3.4105
R13939 VPWR.n2127 VPWR.n519 3.4105
R13940 VPWR.n2056 VPWR.n2055 3.4105
R13941 VPWR.n2040 VPWR.n638 3.4105
R13942 VPWR.n2015 VPWR.n2014 3.4105
R13943 VPWR.n1931 VPWR.n711 3.4105
R13944 VPWR.n1860 VPWR.n1859 3.4105
R13945 VPWR.n1844 VPWR.n830 3.4105
R13946 VPWR.n1819 VPWR.n1818 3.4105
R13947 VPWR.n1735 VPWR.n903 3.4105
R13948 VPWR.n1736 VPWR.n906 3.4105
R13949 VPWR.n1737 VPWR.n907 3.4105
R13950 VPWR.n1738 VPWR.n910 3.4105
R13951 VPWR.n1739 VPWR.n911 3.4105
R13952 VPWR.n1740 VPWR.n914 3.4105
R13953 VPWR.n1741 VPWR.n915 3.4105
R13954 VPWR.n1789 VPWR.n1788 3.4105
R13955 VPWR.n1838 VPWR.n818 3.4105
R13956 VPWR.n1890 VPWR.n1889 3.4105
R13957 VPWR.n1937 VPWR.n723 3.4105
R13958 VPWR.n1985 VPWR.n1984 3.4105
R13959 VPWR.n2034 VPWR.n626 3.4105
R13960 VPWR.n2086 VPWR.n2085 3.4105
R13961 VPWR.n2133 VPWR.n531 3.4105
R13962 VPWR.n2181 VPWR.n2180 3.4105
R13963 VPWR.n2230 VPWR.n434 3.4105
R13964 VPWR.n2282 VPWR.n2281 3.4105
R13965 VPWR.n2329 VPWR.n339 3.4105
R13966 VPWR.n2377 VPWR.n2376 3.4105
R13967 VPWR.n2369 VPWR.n2368 3.4105
R13968 VPWR.n2330 VPWR.n342 3.4105
R13969 VPWR.n2290 VPWR.n2289 3.4105
R13970 VPWR.n2229 VPWR.n431 3.4105
R13971 VPWR.n2173 VPWR.n2172 3.4105
R13972 VPWR.n2134 VPWR.n534 3.4105
R13973 VPWR.n2094 VPWR.n2093 3.4105
R13974 VPWR.n2033 VPWR.n623 3.4105
R13975 VPWR.n1977 VPWR.n1976 3.4105
R13976 VPWR.n1938 VPWR.n726 3.4105
R13977 VPWR.n1898 VPWR.n1897 3.4105
R13978 VPWR.n1837 VPWR.n815 3.4105
R13979 VPWR.n1781 VPWR.n1780 3.4105
R13980 VPWR.n1742 VPWR.n918 3.4105
R13981 VPWR.n1734 VPWR.n902 3.4105
R13982 VPWR.n1821 VPWR.n1820 3.4105
R13983 VPWR.n1845 VPWR.n831 3.4105
R13984 VPWR.n1858 VPWR.n1857 3.4105
R13985 VPWR.n1930 VPWR.n710 3.4105
R13986 VPWR.n2017 VPWR.n2016 3.4105
R13987 VPWR.n2041 VPWR.n639 3.4105
R13988 VPWR.n2054 VPWR.n2053 3.4105
R13989 VPWR.n2126 VPWR.n518 3.4105
R13990 VPWR.n2213 VPWR.n2212 3.4105
R13991 VPWR.n2237 VPWR.n447 3.4105
R13992 VPWR.n2250 VPWR.n2249 3.4105
R13993 VPWR.n2322 VPWR.n326 3.4105
R13994 VPWR.n2409 VPWR.n2408 3.4105
R13995 VPWR.n2433 VPWR.n96 3.4105
R13996 VPWR.n2432 VPWR.n95 3.4105
R13997 VPWR.n2431 VPWR.n90 3.4105
R13998 VPWR.n2430 VPWR.n89 3.4105
R13999 VPWR.n2429 VPWR.n84 3.4105
R14000 VPWR.n2428 VPWR.n83 3.4105
R14001 VPWR.n2427 VPWR.n78 3.4105
R14002 VPWR.n2426 VPWR.n77 3.4105
R14003 VPWR.n2425 VPWR.n72 3.4105
R14004 VPWR.n2424 VPWR.n71 3.4105
R14005 VPWR.n2367 VPWR.n2366 3.4105
R14006 VPWR.n2331 VPWR.n343 3.4105
R14007 VPWR.n2292 VPWR.n2291 3.4105
R14008 VPWR.n2228 VPWR.n430 3.4105
R14009 VPWR.n2171 VPWR.n2170 3.4105
R14010 VPWR.n2135 VPWR.n535 3.4105
R14011 VPWR.n2096 VPWR.n2095 3.4105
R14012 VPWR.n2032 VPWR.n622 3.4105
R14013 VPWR.n1975 VPWR.n1974 3.4105
R14014 VPWR.n1939 VPWR.n727 3.4105
R14015 VPWR.n1900 VPWR.n1899 3.4105
R14016 VPWR.n1836 VPWR.n814 3.4105
R14017 VPWR.n1779 VPWR.n1778 3.4105
R14018 VPWR.n1743 VPWR.n919 3.4105
R14019 VPWR.n1510 VPWR.n1407 3.4105
R14020 VPWR.n1518 VPWR.n1517 3.4105
R14021 VPWR.n1503 VPWR.n1502 3.4105
R14022 VPWR.n1495 VPWR.n1494 3.4105
R14023 VPWR.n1489 VPWR.n1488 3.4105
R14024 VPWR.n1481 VPWR.n1480 3.4105
R14025 VPWR.n1475 VPWR.n1474 3.4105
R14026 VPWR.n1467 VPWR.n1466 3.4105
R14027 VPWR.n1461 VPWR.n1171 3.4105
R14028 VPWR.n1568 VPWR.n1567 3.4105
R14029 VPWR.n1701 VPWR.n1700 3.4105
R14030 VPWR.n1744 VPWR.n922 3.4105
R14031 VPWR.n1771 VPWR.n1770 3.4105
R14032 VPWR.n1835 VPWR.n811 3.4105
R14033 VPWR.n1908 VPWR.n1907 3.4105
R14034 VPWR.n1940 VPWR.n730 3.4105
R14035 VPWR.n1967 VPWR.n1966 3.4105
R14036 VPWR.n2031 VPWR.n619 3.4105
R14037 VPWR.n2104 VPWR.n2103 3.4105
R14038 VPWR.n2136 VPWR.n538 3.4105
R14039 VPWR.n2163 VPWR.n2162 3.4105
R14040 VPWR.n2227 VPWR.n427 3.4105
R14041 VPWR.n2300 VPWR.n2299 3.4105
R14042 VPWR.n2332 VPWR.n346 3.4105
R14043 VPWR.n2359 VPWR.n2358 3.4105
R14044 VPWR.n2423 VPWR.n66 3.4105
R14045 VPWR.n2421 VPWR.n60 3.4105
R14046 VPWR.n2349 VPWR.n2348 3.4105
R14047 VPWR.n2334 VPWR.n350 3.4105
R14048 VPWR.n2310 VPWR.n2309 3.4105
R14049 VPWR.n2225 VPWR.n423 3.4105
R14050 VPWR.n2153 VPWR.n2152 3.4105
R14051 VPWR.n2138 VPWR.n542 3.4105
R14052 VPWR.n2114 VPWR.n2113 3.4105
R14053 VPWR.n2029 VPWR.n615 3.4105
R14054 VPWR.n1957 VPWR.n1956 3.4105
R14055 VPWR.n1942 VPWR.n734 3.4105
R14056 VPWR.n1918 VPWR.n1917 3.4105
R14057 VPWR.n1833 VPWR.n807 3.4105
R14058 VPWR.n1761 VPWR.n1760 3.4105
R14059 VPWR.n1746 VPWR.n926 3.4105
R14060 VPWR.n1688 VPWR.n1680 3.4105
R14061 VPWR.n1693 VPWR.n1011 3.4105
R14062 VPWR.n1745 VPWR.n923 3.4105
R14063 VPWR.n1769 VPWR.n1768 3.4105
R14064 VPWR.n1834 VPWR.n810 3.4105
R14065 VPWR.n1910 VPWR.n1909 3.4105
R14066 VPWR.n1941 VPWR.n731 3.4105
R14067 VPWR.n1965 VPWR.n1964 3.4105
R14068 VPWR.n2030 VPWR.n618 3.4105
R14069 VPWR.n2106 VPWR.n2105 3.4105
R14070 VPWR.n2137 VPWR.n539 3.4105
R14071 VPWR.n2161 VPWR.n2160 3.4105
R14072 VPWR.n2226 VPWR.n426 3.4105
R14073 VPWR.n2302 VPWR.n2301 3.4105
R14074 VPWR.n2333 VPWR.n347 3.4105
R14075 VPWR.n2357 VPWR.n2356 3.4105
R14076 VPWR.n2422 VPWR.n65 3.4105
R14077 VPWR.n2420 VPWR.n59 3.4105
R14078 VPWR.n2347 VPWR.n2346 3.4105
R14079 VPWR.n2335 VPWR.n351 3.4105
R14080 VPWR.n2312 VPWR.n2311 3.4105
R14081 VPWR.n2224 VPWR.n422 3.4105
R14082 VPWR.n2151 VPWR.n2150 3.4105
R14083 VPWR.n2139 VPWR.n543 3.4105
R14084 VPWR.n2116 VPWR.n2115 3.4105
R14085 VPWR.n2028 VPWR.n614 3.4105
R14086 VPWR.n1955 VPWR.n1954 3.4105
R14087 VPWR.n1943 VPWR.n735 3.4105
R14088 VPWR.n1920 VPWR.n1919 3.4105
R14089 VPWR.n1832 VPWR.n806 3.4105
R14090 VPWR.n1759 VPWR.n1758 3.4105
R14091 VPWR.n1747 VPWR.n927 3.4105
R14092 VPWR.n1724 VPWR.n1723 3.4105
R14093 VPWR.n1389 VPWR.n1168 3.4105
R14094 VPWR.n1733 VPWR.n899 3.4105
R14095 VPWR.n1829 VPWR.n1828 3.4105
R14096 VPWR.n1846 VPWR.n897 3.4105
R14097 VPWR.n1850 VPWR.n1849 3.4105
R14098 VPWR.n1929 VPWR.n707 3.4105
R14099 VPWR.n2025 VPWR.n2024 3.4105
R14100 VPWR.n2042 VPWR.n705 3.4105
R14101 VPWR.n2046 VPWR.n2045 3.4105
R14102 VPWR.n2125 VPWR.n515 3.4105
R14103 VPWR.n2221 VPWR.n2220 3.4105
R14104 VPWR.n2238 VPWR.n513 3.4105
R14105 VPWR.n2242 VPWR.n2241 3.4105
R14106 VPWR.n2321 VPWR.n323 3.4105
R14107 VPWR.n2417 VPWR.n2416 3.4105
R14108 VPWR.n2434 VPWR.n321 3.4105
R14109 VPWR.n2438 VPWR.n2437 3.4105
R14110 VPWR.n2448 VPWR.n2447 3.4105
R14111 VPWR.n2450 VPWR.n2449 3.4105
R14112 VPWR.n2460 VPWR.n2459 3.4105
R14113 VPWR.n2462 VPWR.n2461 3.4105
R14114 VPWR.n2472 VPWR.n2471 3.4105
R14115 VPWR.n2474 VPWR.n2473 3.4105
R14116 VPWR.n2484 VPWR.n2483 3.4105
R14117 VPWR.n2486 VPWR.n2485 3.4105
R14118 VPWR.n2496 VPWR.n2495 3.4105
R14119 VPWR.n2498 VPWR.n2497 3.4105
R14120 VPWR.n2508 VPWR.n2507 3.4105
R14121 VPWR.n2510 VPWR.n2509 3.4105
R14122 VPWR.n2520 VPWR.n2519 3.4105
R14123 VPWR.n2522 VPWR.n2521 3.4105
R14124 VPWR.n2531 VPWR.n2530 3.4105
R14125 VPWR.n2419 VPWR.n22 3.4105
R14126 VPWR.n2340 VPWR.n2339 3.4105
R14127 VPWR.n2336 VPWR.n417 3.4105
R14128 VPWR.n2319 VPWR.n2318 3.4105
R14129 VPWR.n2223 VPWR.n419 3.4105
R14130 VPWR.n2144 VPWR.n2143 3.4105
R14131 VPWR.n2140 VPWR.n609 3.4105
R14132 VPWR.n2123 VPWR.n2122 3.4105
R14133 VPWR.n2027 VPWR.n611 3.4105
R14134 VPWR.n1948 VPWR.n1947 3.4105
R14135 VPWR.n1944 VPWR.n801 3.4105
R14136 VPWR.n1927 VPWR.n1926 3.4105
R14137 VPWR.n1831 VPWR.n803 3.4105
R14138 VPWR.n1752 VPWR.n1751 3.4105
R14139 VPWR.n1748 VPWR.n993 3.4105
R14140 VPWR.n1731 VPWR.n1730 3.4105
R14141 VPWR.n1023 VPWR.n996 3.4105
R14142 VPWR.n1024 VPWR.n1005 3.4105
R14143 VPWR.n1690 VPWR.n1689 3.4105
R14144 VPWR.n1692 VPWR.n1691 3.4105
R14145 VPWR.n1507 VPWR.n1013 3.4105
R14146 VPWR.n1509 VPWR.n1508 3.4105
R14147 VPWR.n1506 VPWR.n1408 3.4105
R14148 VPWR.n1505 VPWR.n1504 3.4105
R14149 VPWR.n1493 VPWR.n1492 3.4105
R14150 VPWR.n1491 VPWR.n1490 3.4105
R14151 VPWR.n1479 VPWR.n1478 3.4105
R14152 VPWR.n1477 VPWR.n1476 3.4105
R14153 VPWR.n1465 VPWR.n1464 3.4105
R14154 VPWR.n1463 VPWR.n1462 3.4105
R14155 VPWR.n1570 VPWR.n1569 3.4105
R14156 VPWR.n1572 VPWR.n1571 3.4105
R14157 VPWR.n1284 VPWR.n1280 3.38874
R14158 VPWR.n1323 VPWR.n1319 3.38874
R14159 VPWR.n1360 VPWR.n1356 3.38874
R14160 VPWR.n28 VPWR.n26 3.36657
R14161 VPWR.n30 VPWR.n28 3.36657
R14162 VPWR.n32 VPWR.n30 3.36657
R14163 VPWR.n34 VPWR.n32 3.36657
R14164 VPWR.n36 VPWR.n34 3.36657
R14165 VPWR.n38 VPWR.n36 3.36657
R14166 VPWR.n40 VPWR.n38 3.36657
R14167 VPWR.n42 VPWR.n40 3.36657
R14168 VPWR.n44 VPWR.n42 3.36657
R14169 VPWR.n46 VPWR.n44 3.36657
R14170 VPWR.n48 VPWR.n46 3.36657
R14171 VPWR.n50 VPWR.n48 3.36657
R14172 VPWR.n52 VPWR.n50 3.36657
R14173 VPWR.n54 VPWR.n52 3.36657
R14174 VPWR.t195 VPWR.t1419 3.35739
R14175 VPWR.t531 VPWR.t1446 3.35739
R14176 VPWR.n2507 VPWR.n66 3.28012
R14177 VPWR.n2447 VPWR.n96 3.28012
R14178 VPWR.n2486 VPWR.n77 3.28012
R14179 VPWR.n2376 VPWR.n77 3.28012
R14180 VPWR.n2483 VPWR.n78 3.28012
R14181 VPWR.n2379 VPWR.n78 3.28012
R14182 VPWR.n2471 VPWR.n84 3.28012
R14183 VPWR.n2389 VPWR.n84 3.28012
R14184 VPWR.n2389 VPWR.n334 3.28012
R14185 VPWR.n2462 VPWR.n89 3.28012
R14186 VPWR.n2396 VPWR.n89 3.28012
R14187 VPWR.n2396 VPWR.n331 3.28012
R14188 VPWR.n1476 VPWR.n1475 3.28012
R14189 VPWR.n1475 VPWR.n907 3.28012
R14190 VPWR.n1808 VPWR.n907 3.28012
R14191 VPWR.n1808 VPWR.n826 3.28012
R14192 VPWR.n1870 VPWR.n826 3.28012
R14193 VPWR.n1870 VPWR.n715 3.28012
R14194 VPWR.n2004 VPWR.n715 3.28012
R14195 VPWR.n2004 VPWR.n634 3.28012
R14196 VPWR.n2066 VPWR.n634 3.28012
R14197 VPWR.n2066 VPWR.n523 3.28012
R14198 VPWR.n2200 VPWR.n523 3.28012
R14199 VPWR.n2200 VPWR.n442 3.28012
R14200 VPWR.n2262 VPWR.n442 3.28012
R14201 VPWR.n2262 VPWR.n331 3.28012
R14202 VPWR.n2459 VPWR.n90 3.28012
R14203 VPWR.n2399 VPWR.n90 3.28012
R14204 VPWR.n2399 VPWR.n330 3.28012
R14205 VPWR.n2259 VPWR.n330 3.28012
R14206 VPWR.n2259 VPWR.n443 3.28012
R14207 VPWR.n2203 VPWR.n443 3.28012
R14208 VPWR.n2203 VPWR.n522 3.28012
R14209 VPWR.n2063 VPWR.n522 3.28012
R14210 VPWR.n2063 VPWR.n635 3.28012
R14211 VPWR.n2007 VPWR.n635 3.28012
R14212 VPWR.n2007 VPWR.n714 3.28012
R14213 VPWR.n1867 VPWR.n714 3.28012
R14214 VPWR.n1867 VPWR.n827 3.28012
R14215 VPWR.n1811 VPWR.n827 3.28012
R14216 VPWR.n1467 VPWR.n1465 3.28012
R14217 VPWR.n1467 VPWR.n906 3.28012
R14218 VPWR.n1811 VPWR.n906 3.28012
R14219 VPWR.n1481 VPWR.n1479 3.28012
R14220 VPWR.n1481 VPWR.n910 3.28012
R14221 VPWR.n1801 VPWR.n910 3.28012
R14222 VPWR.n1801 VPWR.n823 3.28012
R14223 VPWR.n1877 VPWR.n823 3.28012
R14224 VPWR.n1877 VPWR.n718 3.28012
R14225 VPWR.n1997 VPWR.n718 3.28012
R14226 VPWR.n1997 VPWR.n631 3.28012
R14227 VPWR.n2073 VPWR.n631 3.28012
R14228 VPWR.n2073 VPWR.n526 3.28012
R14229 VPWR.n2193 VPWR.n526 3.28012
R14230 VPWR.n2193 VPWR.n439 3.28012
R14231 VPWR.n2269 VPWR.n439 3.28012
R14232 VPWR.n2269 VPWR.n334 3.28012
R14233 VPWR.n2474 VPWR.n83 3.28012
R14234 VPWR.n2386 VPWR.n83 3.28012
R14235 VPWR.n2386 VPWR.n335 3.28012
R14236 VPWR.n2272 VPWR.n335 3.28012
R14237 VPWR.n2272 VPWR.n438 3.28012
R14238 VPWR.n2190 VPWR.n438 3.28012
R14239 VPWR.n2190 VPWR.n527 3.28012
R14240 VPWR.n2076 VPWR.n527 3.28012
R14241 VPWR.n2076 VPWR.n630 3.28012
R14242 VPWR.n1994 VPWR.n630 3.28012
R14243 VPWR.n1994 VPWR.n719 3.28012
R14244 VPWR.n1880 VPWR.n719 3.28012
R14245 VPWR.n1880 VPWR.n822 3.28012
R14246 VPWR.n1798 VPWR.n822 3.28012
R14247 VPWR.n1490 VPWR.n1489 3.28012
R14248 VPWR.n1489 VPWR.n911 3.28012
R14249 VPWR.n1798 VPWR.n911 3.28012
R14250 VPWR.n1495 VPWR.n1493 3.28012
R14251 VPWR.n1495 VPWR.n914 3.28012
R14252 VPWR.n1791 VPWR.n914 3.28012
R14253 VPWR.n1791 VPWR.n819 3.28012
R14254 VPWR.n1887 VPWR.n819 3.28012
R14255 VPWR.n1887 VPWR.n722 3.28012
R14256 VPWR.n1987 VPWR.n722 3.28012
R14257 VPWR.n1987 VPWR.n627 3.28012
R14258 VPWR.n2083 VPWR.n627 3.28012
R14259 VPWR.n2083 VPWR.n530 3.28012
R14260 VPWR.n2183 VPWR.n530 3.28012
R14261 VPWR.n2183 VPWR.n435 3.28012
R14262 VPWR.n2279 VPWR.n435 3.28012
R14263 VPWR.n2279 VPWR.n338 3.28012
R14264 VPWR.n2379 VPWR.n338 3.28012
R14265 VPWR.n2450 VPWR.n95 3.28012
R14266 VPWR.n2406 VPWR.n95 3.28012
R14267 VPWR.n2406 VPWR.n327 3.28012
R14268 VPWR.n2252 VPWR.n327 3.28012
R14269 VPWR.n2252 VPWR.n446 3.28012
R14270 VPWR.n2210 VPWR.n446 3.28012
R14271 VPWR.n2210 VPWR.n519 3.28012
R14272 VPWR.n2056 VPWR.n519 3.28012
R14273 VPWR.n2056 VPWR.n638 3.28012
R14274 VPWR.n2014 VPWR.n638 3.28012
R14275 VPWR.n2014 VPWR.n711 3.28012
R14276 VPWR.n1860 VPWR.n711 3.28012
R14277 VPWR.n1860 VPWR.n830 3.28012
R14278 VPWR.n1818 VPWR.n830 3.28012
R14279 VPWR.n1818 VPWR.n903 3.28012
R14280 VPWR.n1462 VPWR.n1461 3.28012
R14281 VPWR.n1461 VPWR.n903 3.28012
R14282 VPWR.n1504 VPWR.n1503 3.28012
R14283 VPWR.n1503 VPWR.n915 3.28012
R14284 VPWR.n1788 VPWR.n915 3.28012
R14285 VPWR.n1788 VPWR.n818 3.28012
R14286 VPWR.n1890 VPWR.n818 3.28012
R14287 VPWR.n1890 VPWR.n723 3.28012
R14288 VPWR.n1984 VPWR.n723 3.28012
R14289 VPWR.n1984 VPWR.n626 3.28012
R14290 VPWR.n2086 VPWR.n626 3.28012
R14291 VPWR.n2086 VPWR.n531 3.28012
R14292 VPWR.n2180 VPWR.n531 3.28012
R14293 VPWR.n2180 VPWR.n434 3.28012
R14294 VPWR.n2282 VPWR.n434 3.28012
R14295 VPWR.n2282 VPWR.n339 3.28012
R14296 VPWR.n2376 VPWR.n339 3.28012
R14297 VPWR.n2495 VPWR.n72 3.28012
R14298 VPWR.n2369 VPWR.n72 3.28012
R14299 VPWR.n2369 VPWR.n342 3.28012
R14300 VPWR.n2289 VPWR.n342 3.28012
R14301 VPWR.n2289 VPWR.n431 3.28012
R14302 VPWR.n2173 VPWR.n431 3.28012
R14303 VPWR.n2173 VPWR.n534 3.28012
R14304 VPWR.n2093 VPWR.n534 3.28012
R14305 VPWR.n2093 VPWR.n623 3.28012
R14306 VPWR.n1977 VPWR.n623 3.28012
R14307 VPWR.n1977 VPWR.n726 3.28012
R14308 VPWR.n1897 VPWR.n726 3.28012
R14309 VPWR.n1897 VPWR.n815 3.28012
R14310 VPWR.n1781 VPWR.n815 3.28012
R14311 VPWR.n1781 VPWR.n918 3.28012
R14312 VPWR.n1517 VPWR.n1408 3.28012
R14313 VPWR.n1517 VPWR.n918 3.28012
R14314 VPWR.n1569 VPWR.n1568 3.28012
R14315 VPWR.n1568 VPWR.n902 3.28012
R14316 VPWR.n1821 VPWR.n902 3.28012
R14317 VPWR.n1821 VPWR.n831 3.28012
R14318 VPWR.n1857 VPWR.n831 3.28012
R14319 VPWR.n1857 VPWR.n710 3.28012
R14320 VPWR.n2017 VPWR.n710 3.28012
R14321 VPWR.n2017 VPWR.n639 3.28012
R14322 VPWR.n2053 VPWR.n639 3.28012
R14323 VPWR.n2053 VPWR.n518 3.28012
R14324 VPWR.n2213 VPWR.n518 3.28012
R14325 VPWR.n2213 VPWR.n447 3.28012
R14326 VPWR.n2249 VPWR.n447 3.28012
R14327 VPWR.n2249 VPWR.n326 3.28012
R14328 VPWR.n2409 VPWR.n326 3.28012
R14329 VPWR.n2409 VPWR.n96 3.28012
R14330 VPWR.n2498 VPWR.n71 3.28012
R14331 VPWR.n2366 VPWR.n71 3.28012
R14332 VPWR.n2366 VPWR.n343 3.28012
R14333 VPWR.n2292 VPWR.n343 3.28012
R14334 VPWR.n2292 VPWR.n430 3.28012
R14335 VPWR.n2170 VPWR.n430 3.28012
R14336 VPWR.n2170 VPWR.n535 3.28012
R14337 VPWR.n2096 VPWR.n535 3.28012
R14338 VPWR.n2096 VPWR.n622 3.28012
R14339 VPWR.n1974 VPWR.n622 3.28012
R14340 VPWR.n1974 VPWR.n727 3.28012
R14341 VPWR.n1900 VPWR.n727 3.28012
R14342 VPWR.n1900 VPWR.n814 3.28012
R14343 VPWR.n1778 VPWR.n814 3.28012
R14344 VPWR.n1778 VPWR.n919 3.28012
R14345 VPWR.n1510 VPWR.n919 3.28012
R14346 VPWR.n1510 VPWR.n1509 3.28012
R14347 VPWR.n1700 VPWR.n1013 3.28012
R14348 VPWR.n1700 VPWR.n922 3.28012
R14349 VPWR.n1771 VPWR.n922 3.28012
R14350 VPWR.n1771 VPWR.n811 3.28012
R14351 VPWR.n1907 VPWR.n811 3.28012
R14352 VPWR.n1907 VPWR.n730 3.28012
R14353 VPWR.n1967 VPWR.n730 3.28012
R14354 VPWR.n1967 VPWR.n619 3.28012
R14355 VPWR.n2103 VPWR.n619 3.28012
R14356 VPWR.n2103 VPWR.n538 3.28012
R14357 VPWR.n2163 VPWR.n538 3.28012
R14358 VPWR.n2163 VPWR.n427 3.28012
R14359 VPWR.n2299 VPWR.n427 3.28012
R14360 VPWR.n2299 VPWR.n346 3.28012
R14361 VPWR.n2359 VPWR.n346 3.28012
R14362 VPWR.n2359 VPWR.n66 3.28012
R14363 VPWR.n2519 VPWR.n60 3.28012
R14364 VPWR.n2349 VPWR.n60 3.28012
R14365 VPWR.n2349 VPWR.n350 3.28012
R14366 VPWR.n2309 VPWR.n350 3.28012
R14367 VPWR.n2309 VPWR.n423 3.28012
R14368 VPWR.n2153 VPWR.n423 3.28012
R14369 VPWR.n2153 VPWR.n542 3.28012
R14370 VPWR.n2113 VPWR.n542 3.28012
R14371 VPWR.n2113 VPWR.n615 3.28012
R14372 VPWR.n1957 VPWR.n615 3.28012
R14373 VPWR.n1957 VPWR.n734 3.28012
R14374 VPWR.n1917 VPWR.n734 3.28012
R14375 VPWR.n1917 VPWR.n807 3.28012
R14376 VPWR.n1761 VPWR.n807 3.28012
R14377 VPWR.n1761 VPWR.n926 3.28012
R14378 VPWR.n1688 VPWR.n926 3.28012
R14379 VPWR.n1689 VPWR.n1688 3.28012
R14380 VPWR.n1693 VPWR.n1692 3.28012
R14381 VPWR.n1693 VPWR.n923 3.28012
R14382 VPWR.n1768 VPWR.n923 3.28012
R14383 VPWR.n1768 VPWR.n810 3.28012
R14384 VPWR.n1910 VPWR.n810 3.28012
R14385 VPWR.n1910 VPWR.n731 3.28012
R14386 VPWR.n1964 VPWR.n731 3.28012
R14387 VPWR.n1964 VPWR.n618 3.28012
R14388 VPWR.n2106 VPWR.n618 3.28012
R14389 VPWR.n2106 VPWR.n539 3.28012
R14390 VPWR.n2160 VPWR.n539 3.28012
R14391 VPWR.n2160 VPWR.n426 3.28012
R14392 VPWR.n2302 VPWR.n426 3.28012
R14393 VPWR.n2302 VPWR.n347 3.28012
R14394 VPWR.n2356 VPWR.n347 3.28012
R14395 VPWR.n2356 VPWR.n65 3.28012
R14396 VPWR.n2510 VPWR.n65 3.28012
R14397 VPWR.n2522 VPWR.n59 3.28012
R14398 VPWR.n2346 VPWR.n59 3.28012
R14399 VPWR.n2346 VPWR.n351 3.28012
R14400 VPWR.n2312 VPWR.n351 3.28012
R14401 VPWR.n2312 VPWR.n422 3.28012
R14402 VPWR.n2150 VPWR.n422 3.28012
R14403 VPWR.n2150 VPWR.n543 3.28012
R14404 VPWR.n2116 VPWR.n543 3.28012
R14405 VPWR.n2116 VPWR.n614 3.28012
R14406 VPWR.n1954 VPWR.n614 3.28012
R14407 VPWR.n1954 VPWR.n735 3.28012
R14408 VPWR.n1920 VPWR.n735 3.28012
R14409 VPWR.n1920 VPWR.n806 3.28012
R14410 VPWR.n1758 VPWR.n806 3.28012
R14411 VPWR.n1758 VPWR.n927 3.28012
R14412 VPWR.n1724 VPWR.n927 3.28012
R14413 VPWR.n1724 VPWR.n1005 3.28012
R14414 VPWR.n1572 VPWR.n1168 3.28012
R14415 VPWR.n1168 VPWR.n899 3.28012
R14416 VPWR.n1828 VPWR.n899 3.28012
R14417 VPWR.n1828 VPWR.n897 3.28012
R14418 VPWR.n1850 VPWR.n897 3.28012
R14419 VPWR.n1850 VPWR.n707 3.28012
R14420 VPWR.n2024 VPWR.n707 3.28012
R14421 VPWR.n2024 VPWR.n705 3.28012
R14422 VPWR.n2046 VPWR.n705 3.28012
R14423 VPWR.n2046 VPWR.n515 3.28012
R14424 VPWR.n2220 VPWR.n515 3.28012
R14425 VPWR.n2220 VPWR.n513 3.28012
R14426 VPWR.n2242 VPWR.n513 3.28012
R14427 VPWR.n2242 VPWR.n323 3.28012
R14428 VPWR.n2416 VPWR.n323 3.28012
R14429 VPWR.n2416 VPWR.n321 3.28012
R14430 VPWR.n2438 VPWR.n321 3.28012
R14431 VPWR.n2340 VPWR.n22 3.28012
R14432 VPWR.n2340 VPWR.n417 3.28012
R14433 VPWR.n2318 VPWR.n417 3.28012
R14434 VPWR.n2318 VPWR.n419 3.28012
R14435 VPWR.n2144 VPWR.n419 3.28012
R14436 VPWR.n2144 VPWR.n609 3.28012
R14437 VPWR.n2122 VPWR.n609 3.28012
R14438 VPWR.n2122 VPWR.n611 3.28012
R14439 VPWR.n1948 VPWR.n611 3.28012
R14440 VPWR.n1948 VPWR.n801 3.28012
R14441 VPWR.n1926 VPWR.n801 3.28012
R14442 VPWR.n1926 VPWR.n803 3.28012
R14443 VPWR.n1752 VPWR.n803 3.28012
R14444 VPWR.n1752 VPWR.n993 3.28012
R14445 VPWR.n1730 VPWR.n993 3.28012
R14446 VPWR.n1730 VPWR.n996 3.28012
R14447 VPWR.n2530 VPWR.n22 3.26393
R14448 VPWR.n2768 VPWR.n2767 3.1005
R14449 VPWR.n2762 VPWR.n2761 3.1005
R14450 VPWR.n2782 VPWR.n2751 3.1005
R14451 VPWR.n1263 VPWR.n1261 3.01226
R14452 VPWR.n2799 VPWR 2.83761
R14453 VPWR.n1267 VPWR.n1243 2.63579
R14454 VPWR.n2667 VPWR.n2666 2.25932
R14455 VPWR.n1386 VPWR.n1385 2.01514
R14456 VPWR.n1386 VPWR.n994 1.65255
R14457 VPWR.n2320 VPWR.n2319 1.32852
R14458 VPWR.n2223 VPWR.n418 1.32852
R14459 VPWR.n2143 VPWR.n2142 1.32852
R14460 VPWR.n2141 VPWR.n2140 1.32852
R14461 VPWR.n2124 VPWR.n2123 1.32852
R14462 VPWR.n2027 VPWR.n610 1.32852
R14463 VPWR.n1947 VPWR.n1946 1.32852
R14464 VPWR.n1945 VPWR.n1944 1.32852
R14465 VPWR.n1928 VPWR.n1927 1.32852
R14466 VPWR.n1831 VPWR.n802 1.32852
R14467 VPWR.n2337 VPWR.n2336 1.32852
R14468 VPWR.n1751 VPWR.n1750 1.32852
R14469 VPWR.n2339 VPWR.n2338 1.32852
R14470 VPWR.n1749 VPWR.n1748 1.32852
R14471 VPWR.n2419 VPWR.n21 1.32852
R14472 VPWR.n1732 VPWR.n1731 1.32852
R14473 VPWR.n2532 VPWR.n2531 1.32852
R14474 VPWR.n1023 VPWR.n994 1.32852
R14475 VPWR.n2418 VPWR 1.25994
R14476 VPWR VPWR.n322 1.25994
R14477 VPWR VPWR.n2240 1.25994
R14478 VPWR.n2239 VPWR 1.25994
R14479 VPWR.n2222 VPWR 1.25994
R14480 VPWR VPWR.n514 1.25994
R14481 VPWR VPWR.n2044 1.25994
R14482 VPWR.n2043 VPWR 1.25994
R14483 VPWR.n2026 VPWR 1.25994
R14484 VPWR VPWR.n706 1.25994
R14485 VPWR VPWR.n1848 1.25994
R14486 VPWR.n1847 VPWR 1.25994
R14487 VPWR.n1830 VPWR 1.25994
R14488 VPWR VPWR.n898 1.25994
R14489 VPWR.n2435 VPWR 1.25994
R14490 VPWR VPWR.n1388 1.25994
R14491 VPWR VPWR.n2436 1.25994
R14492 VPWR.n1387 VPWR 1.25994
R14493 VPWR.n2533 VPWR.n2532 1.144
R14494 VPWR.n2797 VPWR.n2796 0.936724
R14495 VPWR.n2796 VPWR.n2752 0.925245
R14496 VPWR VPWR.n2799 0.812229
R14497 VPWR.n133 VPWR.n64 0.682492
R14498 VPWR.n143 VPWR.n67 0.682492
R14499 VPWR.n153 VPWR.n70 0.682492
R14500 VPWR.n163 VPWR.n73 0.682492
R14501 VPWR.n173 VPWR.n76 0.682492
R14502 VPWR.n183 VPWR.n79 0.682492
R14503 VPWR.n193 VPWR.n82 0.682492
R14504 VPWR.n203 VPWR.n85 0.682492
R14505 VPWR.n213 VPWR.n88 0.682492
R14506 VPWR.n223 VPWR.n91 0.682492
R14507 VPWR.n233 VPWR.n94 0.682492
R14508 VPWR.n243 VPWR.n97 0.682492
R14509 VPWR.n257 VPWR.n256 0.682492
R14510 VPWR.n123 VPWR.n61 0.682492
R14511 VPWR.n114 VPWR.n58 0.682492
R14512 VPWR.n1671 VPWR.n1670 0.682492
R14513 VPWR.n1658 VPWR.n1025 0.682492
R14514 VPWR.n1648 VPWR.n1646 0.682492
R14515 VPWR.n1642 VPWR.n1640 0.682492
R14516 VPWR.n1636 VPWR.n1634 0.682492
R14517 VPWR.n1630 VPWR.n1628 0.682492
R14518 VPWR.n1624 VPWR.n1622 0.682492
R14519 VPWR.n1618 VPWR.n1616 0.682492
R14520 VPWR.n1612 VPWR.n1610 0.682492
R14521 VPWR.n1606 VPWR.n1604 0.682492
R14522 VPWR.n1600 VPWR.n1598 0.682492
R14523 VPWR.n1594 VPWR.n1592 0.682492
R14524 VPWR.n1588 VPWR.n1586 0.682492
R14525 VPWR.n1582 VPWR.n1580 0.682492
R14526 VPWR.n1576 VPWR.n1574 0.682492
R14527 VPWR.n2742 VPWR.n2741 0.672385
R14528 VPWR.n2726 VPWR.n2721 0.672385
R14529 VPWR.n2706 VPWR.n2701 0.672385
R14530 VPWR.n2687 VPWR.n2682 0.672385
R14531 VPWR.n7 VPWR 0.63497
R14532 VPWR.n1181 VPWR 0.63497
R14533 VPWR.n1204 VPWR 0.63497
R14534 VPWR.n1228 VPWR 0.63497
R14535 VPWR.n24 VPWR 0.485653
R14536 VPWR.n2529 VPWR 0.468942
R14537 VPWR VPWR.n1031 0.468942
R14538 VPWR.n2439 VPWR.n257 0.460321
R14539 VPWR.n2506 VPWR.n67 0.460321
R14540 VPWR.n2446 VPWR.n97 0.460321
R14541 VPWR.n2487 VPWR.n76 0.460321
R14542 VPWR.n2482 VPWR.n79 0.460321
R14543 VPWR.n2470 VPWR.n85 0.460321
R14544 VPWR.n2463 VPWR.n88 0.460321
R14545 VPWR.n1598 VPWR.n1063 0.460321
R14546 VPWR.n2458 VPWR.n91 0.460321
R14547 VPWR.n1592 VPWR.n1066 0.460321
R14548 VPWR.n1604 VPWR.n1060 0.460321
R14549 VPWR.n2475 VPWR.n82 0.460321
R14550 VPWR.n1610 VPWR.n1057 0.460321
R14551 VPWR.n1616 VPWR.n1054 0.460321
R14552 VPWR.n2451 VPWR.n94 0.460321
R14553 VPWR.n1586 VPWR.n1069 0.460321
R14554 VPWR.n1622 VPWR.n1051 0.460321
R14555 VPWR.n2494 VPWR.n73 0.460321
R14556 VPWR.n1628 VPWR.n1048 0.460321
R14557 VPWR.n1580 VPWR.n1072 0.460321
R14558 VPWR.n2499 VPWR.n70 0.460321
R14559 VPWR.n1634 VPWR.n1045 0.460321
R14560 VPWR.n1640 VPWR.n1042 0.460321
R14561 VPWR.n1679 VPWR.n1025 0.460321
R14562 VPWR.n1646 VPWR.n1022 0.460321
R14563 VPWR.n2511 VPWR.n64 0.460321
R14564 VPWR.n2518 VPWR.n61 0.460321
R14565 VPWR.n2523 VPWR.n58 0.460321
R14566 VPWR.n1672 VPWR.n1671 0.460321
R14567 VPWR.n1574 VPWR.n1573 0.460321
R14568 VPWR.n2750 VPWR.n2749 0.442692
R14569 VPWR.n2796 VPWR.n2795 0.388
R14570 VPWR.n1109 VPWR.n1106 0.349144
R14571 VPWR.n1106 VPWR.n1103 0.349144
R14572 VPWR.n1103 VPWR.n1100 0.349144
R14573 VPWR.n1100 VPWR.n1097 0.349144
R14574 VPWR.n1097 VPWR.n1094 0.349144
R14575 VPWR.n1094 VPWR.n1091 0.349144
R14576 VPWR.n1091 VPWR.n1088 0.349144
R14577 VPWR.n1088 VPWR.n1085 0.349144
R14578 VPWR.n1085 VPWR.n1082 0.349144
R14579 VPWR.n1082 VPWR.n1079 0.349144
R14580 VPWR.n1079 VPWR.n1035 0.349144
R14581 VPWR.n1654 VPWR.n1035 0.349144
R14582 VPWR.n1664 VPWR.n1654 0.349144
R14583 VPWR.n250 VPWR.n249 0.349144
R14584 VPWR.n249 VPWR.n239 0.349144
R14585 VPWR.n239 VPWR.n229 0.349144
R14586 VPWR.n229 VPWR.n219 0.349144
R14587 VPWR.n219 VPWR.n209 0.349144
R14588 VPWR.n209 VPWR.n199 0.349144
R14589 VPWR.n199 VPWR.n189 0.349144
R14590 VPWR.n189 VPWR.n179 0.349144
R14591 VPWR.n179 VPWR.n169 0.349144
R14592 VPWR.n169 VPWR.n159 0.349144
R14593 VPWR.n159 VPWR.n149 0.349144
R14594 VPWR.n149 VPWR.n139 0.349144
R14595 VPWR.n139 VPWR.n129 0.349144
R14596 VPWR.n1395 VPWR.n1394 0.346131
R14597 VPWR.n1565 VPWR.n1399 0.346131
R14598 VPWR.n1564 VPWR.n1560 0.346131
R14599 VPWR.n1559 VPWR.n1555 0.346131
R14600 VPWR.n1554 VPWR.n1550 0.346131
R14601 VPWR.n1549 VPWR.n1545 0.346131
R14602 VPWR.n1544 VPWR.n1540 0.346131
R14603 VPWR.n1539 VPWR.n1535 0.346131
R14604 VPWR.n1534 VPWR.n1530 0.346131
R14605 VPWR.n1529 VPWR.n1525 0.346131
R14606 VPWR.n1524 VPWR.n1520 0.346131
R14607 VPWR.n1703 VPWR.n1010 0.346131
R14608 VPWR.n1720 VPWR.n1716 0.346131
R14609 VPWR.n1721 VPWR.n1712 0.346131
R14610 VPWR.n1708 VPWR.n1707 0.346131
R14611 VPWR.n2798 VPWR.n2797 0.304571
R14612 VPWR.n2530 VPWR.n55 0.300179
R14613 VPWR.n55 VPWR 0.2505
R14614 VPWR VPWR.n2417 0.249238
R14615 VPWR.n2408 VPWR 0.249238
R14616 VPWR VPWR.n2407 0.249238
R14617 VPWR.n2321 VPWR 0.249238
R14618 VPWR.n2322 VPWR 0.249238
R14619 VPWR.n2323 VPWR 0.249238
R14620 VPWR.n2324 VPWR 0.249238
R14621 VPWR.n2241 VPWR 0.249238
R14622 VPWR.n2250 VPWR 0.249238
R14623 VPWR.n2251 VPWR 0.249238
R14624 VPWR.n2260 VPWR 0.249238
R14625 VPWR.n2261 VPWR 0.249238
R14626 VPWR.n2319 VPWR 0.249238
R14627 VPWR.n2311 VPWR 0.249238
R14628 VPWR.n2310 VPWR 0.249238
R14629 VPWR.n2301 VPWR 0.249238
R14630 VPWR.n2300 VPWR 0.249238
R14631 VPWR.n2291 VPWR 0.249238
R14632 VPWR.n2290 VPWR 0.249238
R14633 VPWR.n2281 VPWR 0.249238
R14634 VPWR.n2280 VPWR 0.249238
R14635 VPWR.n2271 VPWR 0.249238
R14636 VPWR.n2270 VPWR 0.249238
R14637 VPWR VPWR.n2238 0.249238
R14638 VPWR VPWR.n2237 0.249238
R14639 VPWR VPWR.n2236 0.249238
R14640 VPWR VPWR.n2235 0.249238
R14641 VPWR VPWR.n2234 0.249238
R14642 VPWR VPWR.n2223 0.249238
R14643 VPWR VPWR.n2224 0.249238
R14644 VPWR VPWR.n2225 0.249238
R14645 VPWR VPWR.n2226 0.249238
R14646 VPWR VPWR.n2227 0.249238
R14647 VPWR VPWR.n2228 0.249238
R14648 VPWR VPWR.n2229 0.249238
R14649 VPWR VPWR.n2230 0.249238
R14650 VPWR VPWR.n2231 0.249238
R14651 VPWR VPWR.n2232 0.249238
R14652 VPWR VPWR.n2233 0.249238
R14653 VPWR VPWR.n2221 0.249238
R14654 VPWR.n2212 VPWR 0.249238
R14655 VPWR VPWR.n2211 0.249238
R14656 VPWR.n2202 VPWR 0.249238
R14657 VPWR VPWR.n2201 0.249238
R14658 VPWR.n2143 VPWR 0.249238
R14659 VPWR VPWR.n2151 0.249238
R14660 VPWR.n2152 VPWR 0.249238
R14661 VPWR VPWR.n2161 0.249238
R14662 VPWR.n2162 VPWR 0.249238
R14663 VPWR VPWR.n2171 0.249238
R14664 VPWR.n2172 VPWR 0.249238
R14665 VPWR VPWR.n2181 0.249238
R14666 VPWR.n2182 VPWR 0.249238
R14667 VPWR VPWR.n2191 0.249238
R14668 VPWR.n2192 VPWR 0.249238
R14669 VPWR.n2125 VPWR 0.249238
R14670 VPWR.n2126 VPWR 0.249238
R14671 VPWR.n2127 VPWR 0.249238
R14672 VPWR.n2128 VPWR 0.249238
R14673 VPWR.n2129 VPWR 0.249238
R14674 VPWR.n2140 VPWR 0.249238
R14675 VPWR.n2139 VPWR 0.249238
R14676 VPWR.n2138 VPWR 0.249238
R14677 VPWR.n2137 VPWR 0.249238
R14678 VPWR.n2136 VPWR 0.249238
R14679 VPWR.n2135 VPWR 0.249238
R14680 VPWR.n2134 VPWR 0.249238
R14681 VPWR.n2133 VPWR 0.249238
R14682 VPWR.n2132 VPWR 0.249238
R14683 VPWR.n2131 VPWR 0.249238
R14684 VPWR.n2130 VPWR 0.249238
R14685 VPWR.n2045 VPWR 0.249238
R14686 VPWR.n2054 VPWR 0.249238
R14687 VPWR.n2055 VPWR 0.249238
R14688 VPWR.n2064 VPWR 0.249238
R14689 VPWR.n2065 VPWR 0.249238
R14690 VPWR.n2123 VPWR 0.249238
R14691 VPWR.n2115 VPWR 0.249238
R14692 VPWR.n2114 VPWR 0.249238
R14693 VPWR.n2105 VPWR 0.249238
R14694 VPWR.n2104 VPWR 0.249238
R14695 VPWR.n2095 VPWR 0.249238
R14696 VPWR.n2094 VPWR 0.249238
R14697 VPWR.n2085 VPWR 0.249238
R14698 VPWR.n2084 VPWR 0.249238
R14699 VPWR.n2075 VPWR 0.249238
R14700 VPWR.n2074 VPWR 0.249238
R14701 VPWR VPWR.n2042 0.249238
R14702 VPWR VPWR.n2041 0.249238
R14703 VPWR VPWR.n2040 0.249238
R14704 VPWR VPWR.n2039 0.249238
R14705 VPWR VPWR.n2038 0.249238
R14706 VPWR VPWR.n2027 0.249238
R14707 VPWR VPWR.n2028 0.249238
R14708 VPWR VPWR.n2029 0.249238
R14709 VPWR VPWR.n2030 0.249238
R14710 VPWR VPWR.n2031 0.249238
R14711 VPWR VPWR.n2032 0.249238
R14712 VPWR VPWR.n2033 0.249238
R14713 VPWR VPWR.n2034 0.249238
R14714 VPWR VPWR.n2035 0.249238
R14715 VPWR VPWR.n2036 0.249238
R14716 VPWR VPWR.n2037 0.249238
R14717 VPWR VPWR.n2025 0.249238
R14718 VPWR.n2016 VPWR 0.249238
R14719 VPWR VPWR.n2015 0.249238
R14720 VPWR.n2006 VPWR 0.249238
R14721 VPWR VPWR.n2005 0.249238
R14722 VPWR.n1947 VPWR 0.249238
R14723 VPWR VPWR.n1955 0.249238
R14724 VPWR.n1956 VPWR 0.249238
R14725 VPWR VPWR.n1965 0.249238
R14726 VPWR.n1966 VPWR 0.249238
R14727 VPWR VPWR.n1975 0.249238
R14728 VPWR.n1976 VPWR 0.249238
R14729 VPWR VPWR.n1985 0.249238
R14730 VPWR.n1986 VPWR 0.249238
R14731 VPWR VPWR.n1995 0.249238
R14732 VPWR.n1996 VPWR 0.249238
R14733 VPWR.n1929 VPWR 0.249238
R14734 VPWR.n1930 VPWR 0.249238
R14735 VPWR.n1931 VPWR 0.249238
R14736 VPWR.n1932 VPWR 0.249238
R14737 VPWR.n1933 VPWR 0.249238
R14738 VPWR.n1944 VPWR 0.249238
R14739 VPWR.n1943 VPWR 0.249238
R14740 VPWR.n1942 VPWR 0.249238
R14741 VPWR.n1941 VPWR 0.249238
R14742 VPWR.n1940 VPWR 0.249238
R14743 VPWR.n1939 VPWR 0.249238
R14744 VPWR.n1938 VPWR 0.249238
R14745 VPWR.n1937 VPWR 0.249238
R14746 VPWR.n1936 VPWR 0.249238
R14747 VPWR.n1935 VPWR 0.249238
R14748 VPWR.n1934 VPWR 0.249238
R14749 VPWR.n1849 VPWR 0.249238
R14750 VPWR.n1858 VPWR 0.249238
R14751 VPWR.n1859 VPWR 0.249238
R14752 VPWR.n1868 VPWR 0.249238
R14753 VPWR.n1869 VPWR 0.249238
R14754 VPWR.n1927 VPWR 0.249238
R14755 VPWR.n1919 VPWR 0.249238
R14756 VPWR.n1918 VPWR 0.249238
R14757 VPWR.n1909 VPWR 0.249238
R14758 VPWR.n1908 VPWR 0.249238
R14759 VPWR.n1899 VPWR 0.249238
R14760 VPWR.n1898 VPWR 0.249238
R14761 VPWR.n1889 VPWR 0.249238
R14762 VPWR.n1888 VPWR 0.249238
R14763 VPWR.n1879 VPWR 0.249238
R14764 VPWR.n1878 VPWR 0.249238
R14765 VPWR VPWR.n1846 0.249238
R14766 VPWR VPWR.n1845 0.249238
R14767 VPWR VPWR.n1844 0.249238
R14768 VPWR VPWR.n1843 0.249238
R14769 VPWR VPWR.n1842 0.249238
R14770 VPWR VPWR.n1831 0.249238
R14771 VPWR VPWR.n1832 0.249238
R14772 VPWR VPWR.n1833 0.249238
R14773 VPWR VPWR.n1834 0.249238
R14774 VPWR VPWR.n1835 0.249238
R14775 VPWR VPWR.n1836 0.249238
R14776 VPWR VPWR.n1837 0.249238
R14777 VPWR VPWR.n1838 0.249238
R14778 VPWR VPWR.n1839 0.249238
R14779 VPWR VPWR.n1840 0.249238
R14780 VPWR VPWR.n1841 0.249238
R14781 VPWR.n2336 VPWR 0.249238
R14782 VPWR.n2335 VPWR 0.249238
R14783 VPWR.n2334 VPWR 0.249238
R14784 VPWR.n2333 VPWR 0.249238
R14785 VPWR.n2332 VPWR 0.249238
R14786 VPWR.n2331 VPWR 0.249238
R14787 VPWR.n2330 VPWR 0.249238
R14788 VPWR.n2329 VPWR 0.249238
R14789 VPWR.n2328 VPWR 0.249238
R14790 VPWR.n2327 VPWR 0.249238
R14791 VPWR.n2326 VPWR 0.249238
R14792 VPWR.n2325 VPWR 0.249238
R14793 VPWR VPWR.n1829 0.249238
R14794 VPWR.n1820 VPWR 0.249238
R14795 VPWR VPWR.n1819 0.249238
R14796 VPWR.n1810 VPWR 0.249238
R14797 VPWR VPWR.n1809 0.249238
R14798 VPWR.n1800 VPWR 0.249238
R14799 VPWR.n1751 VPWR 0.249238
R14800 VPWR VPWR.n1759 0.249238
R14801 VPWR.n1760 VPWR 0.249238
R14802 VPWR VPWR.n1769 0.249238
R14803 VPWR.n1770 VPWR 0.249238
R14804 VPWR VPWR.n1779 0.249238
R14805 VPWR.n1780 VPWR 0.249238
R14806 VPWR VPWR.n1789 0.249238
R14807 VPWR.n1790 VPWR 0.249238
R14808 VPWR VPWR.n1799 0.249238
R14809 VPWR.n2339 VPWR 0.249238
R14810 VPWR VPWR.n2347 0.249238
R14811 VPWR.n2348 VPWR 0.249238
R14812 VPWR VPWR.n2357 0.249238
R14813 VPWR.n2358 VPWR 0.249238
R14814 VPWR VPWR.n2367 0.249238
R14815 VPWR.n2368 VPWR 0.249238
R14816 VPWR VPWR.n2377 0.249238
R14817 VPWR.n2378 VPWR 0.249238
R14818 VPWR VPWR.n2387 0.249238
R14819 VPWR.n2388 VPWR 0.249238
R14820 VPWR VPWR.n2397 0.249238
R14821 VPWR.n2398 VPWR 0.249238
R14822 VPWR.n1733 VPWR 0.249238
R14823 VPWR.n1734 VPWR 0.249238
R14824 VPWR.n1735 VPWR 0.249238
R14825 VPWR.n1736 VPWR 0.249238
R14826 VPWR.n1737 VPWR 0.249238
R14827 VPWR.n1738 VPWR 0.249238
R14828 VPWR.n1739 VPWR 0.249238
R14829 VPWR.n1740 VPWR 0.249238
R14830 VPWR.n1741 VPWR 0.249238
R14831 VPWR.n1748 VPWR 0.249238
R14832 VPWR.n1747 VPWR 0.249238
R14833 VPWR.n1746 VPWR 0.249238
R14834 VPWR.n1745 VPWR 0.249238
R14835 VPWR.n1744 VPWR 0.249238
R14836 VPWR.n1743 VPWR 0.249238
R14837 VPWR.n1742 VPWR 0.249238
R14838 VPWR VPWR.n2434 0.249238
R14839 VPWR VPWR.n2433 0.249238
R14840 VPWR VPWR.n2432 0.249238
R14841 VPWR VPWR.n2431 0.249238
R14842 VPWR VPWR.n2430 0.249238
R14843 VPWR VPWR.n2429 0.249238
R14844 VPWR VPWR.n2428 0.249238
R14845 VPWR VPWR.n2427 0.249238
R14846 VPWR VPWR.n2426 0.249238
R14847 VPWR VPWR.n2425 0.249238
R14848 VPWR VPWR.n2424 0.249238
R14849 VPWR VPWR.n2419 0.249238
R14850 VPWR VPWR.n2420 0.249238
R14851 VPWR VPWR.n2421 0.249238
R14852 VPWR VPWR.n2422 0.249238
R14853 VPWR VPWR.n2423 0.249238
R14854 VPWR.n2437 VPWR 0.249238
R14855 VPWR.n2448 VPWR 0.249238
R14856 VPWR.n2449 VPWR 0.249238
R14857 VPWR.n2460 VPWR 0.249238
R14858 VPWR.n2461 VPWR 0.249238
R14859 VPWR.n2472 VPWR 0.249238
R14860 VPWR.n2473 VPWR 0.249238
R14861 VPWR.n2484 VPWR 0.249238
R14862 VPWR.n2485 VPWR 0.249238
R14863 VPWR.n2496 VPWR 0.249238
R14864 VPWR.n2497 VPWR 0.249238
R14865 VPWR.n2508 VPWR 0.249238
R14866 VPWR.n2509 VPWR 0.249238
R14867 VPWR.n2520 VPWR 0.249238
R14868 VPWR.n2521 VPWR 0.249238
R14869 VPWR.n2531 VPWR 0.249238
R14870 VPWR VPWR.n1023 0.249238
R14871 VPWR VPWR.n1024 0.249238
R14872 VPWR VPWR.n1690 0.249238
R14873 VPWR.n1691 VPWR 0.249238
R14874 VPWR VPWR.n1507 0.249238
R14875 VPWR.n1508 VPWR 0.249238
R14876 VPWR.n1506 VPWR 0.249238
R14877 VPWR.n1505 VPWR 0.249238
R14878 VPWR.n1492 VPWR 0.249238
R14879 VPWR.n1491 VPWR 0.249238
R14880 VPWR.n1478 VPWR 0.249238
R14881 VPWR.n1477 VPWR 0.249238
R14882 VPWR.n1464 VPWR 0.249238
R14883 VPWR.n1463 VPWR 0.249238
R14884 VPWR VPWR.n1570 0.249238
R14885 VPWR.n1571 VPWR 0.249238
R14886 VPWR.n2797 VPWR.n2751 0.245065
R14887 VPWR.n1115 VPWR.n1113 0.217699
R14888 VPWR.n134 VPWR.n131 0.217699
R14889 VPWR.n144 VPWR.n141 0.217699
R14890 VPWR.n154 VPWR.n151 0.217699
R14891 VPWR.n164 VPWR.n161 0.217699
R14892 VPWR.n174 VPWR.n171 0.217699
R14893 VPWR.n184 VPWR.n181 0.217699
R14894 VPWR.n194 VPWR.n191 0.217699
R14895 VPWR.n204 VPWR.n201 0.217699
R14896 VPWR.n214 VPWR.n211 0.217699
R14897 VPWR.n224 VPWR.n221 0.217699
R14898 VPWR.n234 VPWR.n231 0.217699
R14899 VPWR.n244 VPWR.n241 0.217699
R14900 VPWR.n254 VPWR.n101 0.217699
R14901 VPWR.n106 VPWR.n105 0.217699
R14902 VPWR.n124 VPWR.n121 0.217699
R14903 VPWR.n115 VPWR.n112 0.217699
R14904 VPWR.n1668 VPWR.n1033 0.217699
R14905 VPWR.n1659 VPWR.n1656 0.217699
R14906 VPWR.n1649 VPWR.n1037 0.217699
R14907 VPWR.n1645 VPWR.n1643 0.217699
R14908 VPWR.n1639 VPWR.n1637 0.217699
R14909 VPWR.n1633 VPWR.n1631 0.217699
R14910 VPWR.n1627 VPWR.n1625 0.217699
R14911 VPWR.n1621 VPWR.n1619 0.217699
R14912 VPWR.n1615 VPWR.n1613 0.217699
R14913 VPWR.n1609 VPWR.n1607 0.217699
R14914 VPWR.n1603 VPWR.n1601 0.217699
R14915 VPWR.n1597 VPWR.n1595 0.217699
R14916 VPWR.n1591 VPWR.n1589 0.217699
R14917 VPWR.n1585 VPWR.n1583 0.217699
R14918 VPWR.n1579 VPWR.n1577 0.217699
R14919 VPWR.n2749 VPWR.n2733 0.213567
R14920 VPWR.n2733 VPWR.n2714 0.213567
R14921 VPWR.n2714 VPWR.n2694 0.213567
R14922 VPWR.n2694 VPWR.n2675 0.213567
R14923 VPWR.n2675 VPWR.n2639 0.213567
R14924 VPWR.n2639 VPWR.n2601 0.213567
R14925 VPWR.n2601 VPWR.n2564 0.213567
R14926 VPWR.n1385 VPWR.n1353 0.213567
R14927 VPWR.n1353 VPWR.n1315 0.213567
R14928 VPWR.n1315 VPWR.n1276 0.213567
R14929 VPWR.n1276 VPWR.n1241 0.213567
R14930 VPWR.n1241 VPWR.n1218 0.213567
R14931 VPWR.n1218 VPWR.n1194 0.213567
R14932 VPWR.n1194 VPWR.n19 0.213567
R14933 VPWR VPWR.n2798 0.204304
R14934 VPWR.n1387 VPWR.n1386 0.182233
R14935 VPWR.n1388 VPWR.n1387 0.154425
R14936 VPWR.n1388 VPWR.n898 0.154425
R14937 VPWR.n1830 VPWR.n898 0.154425
R14938 VPWR.n1847 VPWR.n1830 0.154425
R14939 VPWR.n1848 VPWR.n1847 0.154425
R14940 VPWR.n1848 VPWR.n706 0.154425
R14941 VPWR.n2026 VPWR.n706 0.154425
R14942 VPWR.n2043 VPWR.n2026 0.154425
R14943 VPWR.n2044 VPWR.n2043 0.154425
R14944 VPWR.n2044 VPWR.n514 0.154425
R14945 VPWR.n2222 VPWR.n514 0.154425
R14946 VPWR.n2239 VPWR.n2222 0.154425
R14947 VPWR.n2240 VPWR.n2239 0.154425
R14948 VPWR.n2240 VPWR.n322 0.154425
R14949 VPWR.n2418 VPWR.n322 0.154425
R14950 VPWR.n2435 VPWR.n2418 0.154425
R14951 VPWR.n2436 VPWR.n2435 0.154425
R14952 VPWR.n1732 VPWR.n994 0.154425
R14953 VPWR.n1749 VPWR.n1732 0.154425
R14954 VPWR.n1750 VPWR.n1749 0.154425
R14955 VPWR.n1750 VPWR.n802 0.154425
R14956 VPWR.n1928 VPWR.n802 0.154425
R14957 VPWR.n1945 VPWR.n1928 0.154425
R14958 VPWR.n1946 VPWR.n1945 0.154425
R14959 VPWR.n1946 VPWR.n610 0.154425
R14960 VPWR.n2124 VPWR.n610 0.154425
R14961 VPWR.n2141 VPWR.n2124 0.154425
R14962 VPWR.n2142 VPWR.n2141 0.154425
R14963 VPWR.n2142 VPWR.n418 0.154425
R14964 VPWR.n2320 VPWR.n418 0.154425
R14965 VPWR.n2337 VPWR.n2320 0.154425
R14966 VPWR.n2338 VPWR.n2337 0.154425
R14967 VPWR.n2338 VPWR.n21 0.154425
R14968 VPWR.n2532 VPWR.n21 0.154425
R14969 VPWR.n8 VPWR.n7 0.147771
R14970 VPWR.n1182 VPWR.n1181 0.147771
R14971 VPWR.n1205 VPWR.n1204 0.147771
R14972 VPWR.n1229 VPWR.n1228 0.147771
R14973 VPWR.n2799 VPWR.n2750 0.127988
R14974 VPWR.n2761 VPWR.n2752 0.1255
R14975 VPWR.n2767 VPWR.n2752 0.1255
R14976 VPWR.n18 VPWR.n0 0.120292
R14977 VPWR.n14 VPWR.n0 0.120292
R14978 VPWR.n9 VPWR.n8 0.120292
R14979 VPWR.n1193 VPWR.n1172 0.120292
R14980 VPWR.n1189 VPWR.n1172 0.120292
R14981 VPWR.n1183 VPWR.n1182 0.120292
R14982 VPWR.n1217 VPWR.n1195 0.120292
R14983 VPWR.n1212 VPWR.n1195 0.120292
R14984 VPWR.n1206 VPWR.n1205 0.120292
R14985 VPWR.n1240 VPWR.n1219 0.120292
R14986 VPWR.n1236 VPWR.n1219 0.120292
R14987 VPWR.n1230 VPWR.n1229 0.120292
R14988 VPWR.n1272 VPWR.n1271 0.120292
R14989 VPWR.n1265 VPWR.n1244 0.120292
R14990 VPWR.n1258 VPWR.n1244 0.120292
R14991 VPWR.n1258 VPWR.n1257 0.120292
R14992 VPWR.n1256 VPWR.n1248 0.120292
R14993 VPWR.n1251 VPWR.n1248 0.120292
R14994 VPWR.n1251 VPWR.n1250 0.120292
R14995 VPWR.n1310 VPWR.n1309 0.120292
R14996 VPWR.n1303 VPWR.n1302 0.120292
R14997 VPWR.n1302 VPWR.n1279 0.120292
R14998 VPWR.n1295 VPWR.n1279 0.120292
R14999 VPWR.n1295 VPWR.n1294 0.120292
R15000 VPWR.n1294 VPWR.n1293 0.120292
R15001 VPWR.n1293 VPWR.n1281 0.120292
R15002 VPWR.n1287 VPWR.n1281 0.120292
R15003 VPWR.n1287 VPWR.n1286 0.120292
R15004 VPWR.n1349 VPWR.n1348 0.120292
R15005 VPWR.n1342 VPWR.n1341 0.120292
R15006 VPWR.n1341 VPWR.n1318 0.120292
R15007 VPWR.n1334 VPWR.n1318 0.120292
R15008 VPWR.n1334 VPWR.n1333 0.120292
R15009 VPWR.n1333 VPWR.n1332 0.120292
R15010 VPWR.n1332 VPWR.n1320 0.120292
R15011 VPWR.n1326 VPWR.n1320 0.120292
R15012 VPWR.n1326 VPWR.n1325 0.120292
R15013 VPWR.n1379 VPWR.n1378 0.120292
R15014 VPWR.n1378 VPWR.n1355 0.120292
R15015 VPWR.n1371 VPWR.n1355 0.120292
R15016 VPWR.n1371 VPWR.n1370 0.120292
R15017 VPWR.n1370 VPWR.n1369 0.120292
R15018 VPWR.n1369 VPWR.n1357 0.120292
R15019 VPWR.n1363 VPWR.n1357 0.120292
R15020 VPWR.n1363 VPWR.n1362 0.120292
R15021 VPWR.n2748 VPWR.n2734 0.120292
R15022 VPWR.n2732 VPWR.n2715 0.120292
R15023 VPWR.n2713 VPWR.n2695 0.120292
R15024 VPWR.n2693 VPWR.n2676 0.120292
R15025 VPWR.n2655 VPWR.n2654 0.120292
R15026 VPWR.n2656 VPWR.n2655 0.120292
R15027 VPWR.n2656 VPWR.n2647 0.120292
R15028 VPWR.n2661 VPWR.n2647 0.120292
R15029 VPWR.n2662 VPWR.n2661 0.120292
R15030 VPWR.n2662 VPWR.n2643 0.120292
R15031 VPWR.n2668 VPWR.n2643 0.120292
R15032 VPWR.n2670 VPWR.n2640 0.120292
R15033 VPWR.n2674 VPWR.n2640 0.120292
R15034 VPWR.n2619 VPWR.n2618 0.120292
R15035 VPWR.n2620 VPWR.n2619 0.120292
R15036 VPWR.n2620 VPWR.n2609 0.120292
R15037 VPWR.n2625 VPWR.n2609 0.120292
R15038 VPWR.n2626 VPWR.n2625 0.120292
R15039 VPWR.n2626 VPWR.n2605 0.120292
R15040 VPWR.n2631 VPWR.n2605 0.120292
R15041 VPWR.n2633 VPWR.n2602 0.120292
R15042 VPWR.n2638 VPWR.n2602 0.120292
R15043 VPWR.n2582 VPWR.n2581 0.120292
R15044 VPWR.n2583 VPWR.n2582 0.120292
R15045 VPWR.n2583 VPWR.n2572 0.120292
R15046 VPWR.n2588 VPWR.n2572 0.120292
R15047 VPWR.n2589 VPWR.n2588 0.120292
R15048 VPWR.n2589 VPWR.n2568 0.120292
R15049 VPWR.n2594 VPWR.n2568 0.120292
R15050 VPWR.n2596 VPWR.n2565 0.120292
R15051 VPWR.n2600 VPWR.n2565 0.120292
R15052 VPWR.n2544 VPWR.n2540 0.120292
R15053 VPWR.n2552 VPWR.n2540 0.120292
R15054 VPWR.n2553 VPWR.n2552 0.120292
R15055 VPWR.n2554 VPWR.n2553 0.120292
R15056 VPWR.n2554 VPWR.n2536 0.120292
R15057 VPWR.n2559 VPWR.n2536 0.120292
R15058 VPWR.n2560 VPWR.n2559 0.120292
R15059 VPWR.n1701 VPWR.n1012 0.108238
R15060 VPWR.n1519 VPWR.n1407 0.108238
R15061 VPWR.n1518 VPWR.n1406 0.108238
R15062 VPWR.n1502 VPWR.n1405 0.108238
R15063 VPWR.n1494 VPWR.n1404 0.108238
R15064 VPWR.n1488 VPWR.n1403 0.108238
R15065 VPWR.n1480 VPWR.n1402 0.108238
R15066 VPWR.n1474 VPWR.n1401 0.108238
R15067 VPWR.n1466 VPWR.n1400 0.108238
R15068 VPWR.n1566 VPWR.n1171 0.108238
R15069 VPWR.n1567 VPWR.n1170 0.108238
R15070 VPWR.n1390 VPWR.n1389 0.108238
R15071 VPWR.n1731 VPWR.n995 0.108238
R15072 VPWR.n1702 VPWR.n1011 0.108238
R15073 VPWR.n1680 VPWR.n1006 0.108238
R15074 VPWR.n1723 VPWR.n1722 0.108238
R15075 VPWR.n2417 VPWR 0.100405
R15076 VPWR.n2408 VPWR 0.100405
R15077 VPWR VPWR.n2321 0.100405
R15078 VPWR VPWR.n2322 0.100405
R15079 VPWR VPWR.n2323 0.100405
R15080 VPWR.n2241 VPWR 0.100405
R15081 VPWR VPWR.n2250 0.100405
R15082 VPWR.n2251 VPWR 0.100405
R15083 VPWR VPWR.n2260 0.100405
R15084 VPWR.n2311 VPWR 0.100405
R15085 VPWR VPWR.n2310 0.100405
R15086 VPWR.n2301 VPWR 0.100405
R15087 VPWR VPWR.n2300 0.100405
R15088 VPWR.n2291 VPWR 0.100405
R15089 VPWR VPWR.n2290 0.100405
R15090 VPWR.n2281 VPWR 0.100405
R15091 VPWR VPWR.n2280 0.100405
R15092 VPWR.n2271 VPWR 0.100405
R15093 VPWR VPWR.n2270 0.100405
R15094 VPWR.n2261 VPWR 0.100405
R15095 VPWR.n2238 VPWR 0.100405
R15096 VPWR.n2237 VPWR 0.100405
R15097 VPWR.n2236 VPWR 0.100405
R15098 VPWR.n2235 VPWR 0.100405
R15099 VPWR.n2224 VPWR 0.100405
R15100 VPWR.n2225 VPWR 0.100405
R15101 VPWR.n2226 VPWR 0.100405
R15102 VPWR.n2227 VPWR 0.100405
R15103 VPWR.n2228 VPWR 0.100405
R15104 VPWR.n2229 VPWR 0.100405
R15105 VPWR.n2230 VPWR 0.100405
R15106 VPWR.n2231 VPWR 0.100405
R15107 VPWR.n2232 VPWR 0.100405
R15108 VPWR.n2233 VPWR 0.100405
R15109 VPWR.n2234 VPWR 0.100405
R15110 VPWR.n2221 VPWR 0.100405
R15111 VPWR.n2212 VPWR 0.100405
R15112 VPWR.n2211 VPWR 0.100405
R15113 VPWR.n2202 VPWR 0.100405
R15114 VPWR.n2151 VPWR 0.100405
R15115 VPWR.n2152 VPWR 0.100405
R15116 VPWR.n2161 VPWR 0.100405
R15117 VPWR.n2162 VPWR 0.100405
R15118 VPWR.n2171 VPWR 0.100405
R15119 VPWR.n2172 VPWR 0.100405
R15120 VPWR.n2181 VPWR 0.100405
R15121 VPWR.n2182 VPWR 0.100405
R15122 VPWR.n2191 VPWR 0.100405
R15123 VPWR.n2192 VPWR 0.100405
R15124 VPWR.n2201 VPWR 0.100405
R15125 VPWR VPWR.n2125 0.100405
R15126 VPWR VPWR.n2126 0.100405
R15127 VPWR VPWR.n2127 0.100405
R15128 VPWR VPWR.n2128 0.100405
R15129 VPWR VPWR.n2139 0.100405
R15130 VPWR VPWR.n2138 0.100405
R15131 VPWR VPWR.n2137 0.100405
R15132 VPWR VPWR.n2136 0.100405
R15133 VPWR VPWR.n2135 0.100405
R15134 VPWR VPWR.n2134 0.100405
R15135 VPWR VPWR.n2133 0.100405
R15136 VPWR VPWR.n2132 0.100405
R15137 VPWR VPWR.n2131 0.100405
R15138 VPWR VPWR.n2130 0.100405
R15139 VPWR VPWR.n2129 0.100405
R15140 VPWR.n2045 VPWR 0.100405
R15141 VPWR VPWR.n2054 0.100405
R15142 VPWR.n2055 VPWR 0.100405
R15143 VPWR VPWR.n2064 0.100405
R15144 VPWR.n2115 VPWR 0.100405
R15145 VPWR VPWR.n2114 0.100405
R15146 VPWR.n2105 VPWR 0.100405
R15147 VPWR VPWR.n2104 0.100405
R15148 VPWR.n2095 VPWR 0.100405
R15149 VPWR VPWR.n2094 0.100405
R15150 VPWR.n2085 VPWR 0.100405
R15151 VPWR VPWR.n2084 0.100405
R15152 VPWR.n2075 VPWR 0.100405
R15153 VPWR VPWR.n2074 0.100405
R15154 VPWR.n2065 VPWR 0.100405
R15155 VPWR.n2042 VPWR 0.100405
R15156 VPWR.n2041 VPWR 0.100405
R15157 VPWR.n2040 VPWR 0.100405
R15158 VPWR.n2039 VPWR 0.100405
R15159 VPWR.n2028 VPWR 0.100405
R15160 VPWR.n2029 VPWR 0.100405
R15161 VPWR.n2030 VPWR 0.100405
R15162 VPWR.n2031 VPWR 0.100405
R15163 VPWR.n2032 VPWR 0.100405
R15164 VPWR.n2033 VPWR 0.100405
R15165 VPWR.n2034 VPWR 0.100405
R15166 VPWR.n2035 VPWR 0.100405
R15167 VPWR.n2036 VPWR 0.100405
R15168 VPWR.n2037 VPWR 0.100405
R15169 VPWR.n2038 VPWR 0.100405
R15170 VPWR.n2025 VPWR 0.100405
R15171 VPWR.n2016 VPWR 0.100405
R15172 VPWR.n2015 VPWR 0.100405
R15173 VPWR.n2006 VPWR 0.100405
R15174 VPWR.n1955 VPWR 0.100405
R15175 VPWR.n1956 VPWR 0.100405
R15176 VPWR.n1965 VPWR 0.100405
R15177 VPWR.n1966 VPWR 0.100405
R15178 VPWR.n1975 VPWR 0.100405
R15179 VPWR.n1976 VPWR 0.100405
R15180 VPWR.n1985 VPWR 0.100405
R15181 VPWR.n1986 VPWR 0.100405
R15182 VPWR.n1995 VPWR 0.100405
R15183 VPWR.n1996 VPWR 0.100405
R15184 VPWR.n2005 VPWR 0.100405
R15185 VPWR VPWR.n1929 0.100405
R15186 VPWR VPWR.n1930 0.100405
R15187 VPWR VPWR.n1931 0.100405
R15188 VPWR VPWR.n1932 0.100405
R15189 VPWR VPWR.n1943 0.100405
R15190 VPWR VPWR.n1942 0.100405
R15191 VPWR VPWR.n1941 0.100405
R15192 VPWR VPWR.n1940 0.100405
R15193 VPWR VPWR.n1939 0.100405
R15194 VPWR VPWR.n1938 0.100405
R15195 VPWR VPWR.n1937 0.100405
R15196 VPWR VPWR.n1936 0.100405
R15197 VPWR VPWR.n1935 0.100405
R15198 VPWR VPWR.n1934 0.100405
R15199 VPWR VPWR.n1933 0.100405
R15200 VPWR.n1849 VPWR 0.100405
R15201 VPWR VPWR.n1858 0.100405
R15202 VPWR.n1859 VPWR 0.100405
R15203 VPWR VPWR.n1868 0.100405
R15204 VPWR.n1919 VPWR 0.100405
R15205 VPWR VPWR.n1918 0.100405
R15206 VPWR.n1909 VPWR 0.100405
R15207 VPWR VPWR.n1908 0.100405
R15208 VPWR.n1899 VPWR 0.100405
R15209 VPWR VPWR.n1898 0.100405
R15210 VPWR.n1889 VPWR 0.100405
R15211 VPWR VPWR.n1888 0.100405
R15212 VPWR.n1879 VPWR 0.100405
R15213 VPWR VPWR.n1878 0.100405
R15214 VPWR.n1869 VPWR 0.100405
R15215 VPWR.n1846 VPWR 0.100405
R15216 VPWR.n1845 VPWR 0.100405
R15217 VPWR.n1844 VPWR 0.100405
R15218 VPWR.n1843 VPWR 0.100405
R15219 VPWR.n1832 VPWR 0.100405
R15220 VPWR.n1833 VPWR 0.100405
R15221 VPWR.n1834 VPWR 0.100405
R15222 VPWR.n1835 VPWR 0.100405
R15223 VPWR.n1836 VPWR 0.100405
R15224 VPWR.n1837 VPWR 0.100405
R15225 VPWR.n1838 VPWR 0.100405
R15226 VPWR.n1839 VPWR 0.100405
R15227 VPWR.n1840 VPWR 0.100405
R15228 VPWR.n1841 VPWR 0.100405
R15229 VPWR.n1842 VPWR 0.100405
R15230 VPWR VPWR.n2335 0.100405
R15231 VPWR VPWR.n2334 0.100405
R15232 VPWR VPWR.n2333 0.100405
R15233 VPWR VPWR.n2332 0.100405
R15234 VPWR VPWR.n2331 0.100405
R15235 VPWR VPWR.n2330 0.100405
R15236 VPWR VPWR.n2329 0.100405
R15237 VPWR VPWR.n2328 0.100405
R15238 VPWR VPWR.n2327 0.100405
R15239 VPWR VPWR.n2326 0.100405
R15240 VPWR VPWR.n2325 0.100405
R15241 VPWR VPWR.n2324 0.100405
R15242 VPWR.n1829 VPWR 0.100405
R15243 VPWR.n1820 VPWR 0.100405
R15244 VPWR.n1819 VPWR 0.100405
R15245 VPWR.n1810 VPWR 0.100405
R15246 VPWR.n1809 VPWR 0.100405
R15247 VPWR.n1759 VPWR 0.100405
R15248 VPWR.n1760 VPWR 0.100405
R15249 VPWR.n1769 VPWR 0.100405
R15250 VPWR.n1770 VPWR 0.100405
R15251 VPWR.n1779 VPWR 0.100405
R15252 VPWR.n1780 VPWR 0.100405
R15253 VPWR.n1789 VPWR 0.100405
R15254 VPWR.n1790 VPWR 0.100405
R15255 VPWR.n1799 VPWR 0.100405
R15256 VPWR.n1800 VPWR 0.100405
R15257 VPWR.n2347 VPWR 0.100405
R15258 VPWR.n2348 VPWR 0.100405
R15259 VPWR.n2357 VPWR 0.100405
R15260 VPWR.n2358 VPWR 0.100405
R15261 VPWR.n2367 VPWR 0.100405
R15262 VPWR.n2368 VPWR 0.100405
R15263 VPWR.n2377 VPWR 0.100405
R15264 VPWR.n2378 VPWR 0.100405
R15265 VPWR.n2387 VPWR 0.100405
R15266 VPWR.n2388 VPWR 0.100405
R15267 VPWR.n2397 VPWR 0.100405
R15268 VPWR.n2398 VPWR 0.100405
R15269 VPWR.n2407 VPWR 0.100405
R15270 VPWR VPWR.n1733 0.100405
R15271 VPWR VPWR.n1734 0.100405
R15272 VPWR VPWR.n1735 0.100405
R15273 VPWR VPWR.n1736 0.100405
R15274 VPWR VPWR.n1737 0.100405
R15275 VPWR VPWR.n1738 0.100405
R15276 VPWR VPWR.n1739 0.100405
R15277 VPWR VPWR.n1740 0.100405
R15278 VPWR VPWR.n1747 0.100405
R15279 VPWR VPWR.n1746 0.100405
R15280 VPWR VPWR.n1745 0.100405
R15281 VPWR VPWR.n1744 0.100405
R15282 VPWR VPWR.n1743 0.100405
R15283 VPWR VPWR.n1742 0.100405
R15284 VPWR VPWR.n1741 0.100405
R15285 VPWR.n2434 VPWR 0.100405
R15286 VPWR.n2433 VPWR 0.100405
R15287 VPWR.n2432 VPWR 0.100405
R15288 VPWR.n2431 VPWR 0.100405
R15289 VPWR.n2430 VPWR 0.100405
R15290 VPWR.n2429 VPWR 0.100405
R15291 VPWR.n2428 VPWR 0.100405
R15292 VPWR.n2427 VPWR 0.100405
R15293 VPWR.n2426 VPWR 0.100405
R15294 VPWR.n2425 VPWR 0.100405
R15295 VPWR.n2420 VPWR 0.100405
R15296 VPWR.n2421 VPWR 0.100405
R15297 VPWR.n2422 VPWR 0.100405
R15298 VPWR.n2423 VPWR 0.100405
R15299 VPWR.n2424 VPWR 0.100405
R15300 VPWR.n1407 VPWR 0.100405
R15301 VPWR VPWR.n1518 0.100405
R15302 VPWR.n1502 VPWR 0.100405
R15303 VPWR.n1494 VPWR 0.100405
R15304 VPWR.n1488 VPWR 0.100405
R15305 VPWR.n1480 VPWR 0.100405
R15306 VPWR.n1474 VPWR 0.100405
R15307 VPWR.n1466 VPWR 0.100405
R15308 VPWR VPWR.n1171 0.100405
R15309 VPWR.n1567 VPWR 0.100405
R15310 VPWR.n1389 VPWR 0.100405
R15311 VPWR.n1011 VPWR 0.100405
R15312 VPWR.n1680 VPWR 0.100405
R15313 VPWR.n1723 VPWR 0.100405
R15314 VPWR VPWR.n1701 0.100405
R15315 VPWR.n2437 VPWR 0.100405
R15316 VPWR VPWR.n2448 0.100405
R15317 VPWR.n2449 VPWR 0.100405
R15318 VPWR VPWR.n2460 0.100405
R15319 VPWR.n2461 VPWR 0.100405
R15320 VPWR VPWR.n2472 0.100405
R15321 VPWR.n2473 VPWR 0.100405
R15322 VPWR VPWR.n2484 0.100405
R15323 VPWR.n2485 VPWR 0.100405
R15324 VPWR VPWR.n2496 0.100405
R15325 VPWR.n2497 VPWR 0.100405
R15326 VPWR VPWR.n2508 0.100405
R15327 VPWR.n2509 VPWR 0.100405
R15328 VPWR VPWR.n2520 0.100405
R15329 VPWR.n2521 VPWR 0.100405
R15330 VPWR.n1024 VPWR 0.100405
R15331 VPWR.n1690 VPWR 0.100405
R15332 VPWR.n1691 VPWR 0.100405
R15333 VPWR.n1507 VPWR 0.100405
R15334 VPWR.n1508 VPWR 0.100405
R15335 VPWR VPWR.n1506 0.100405
R15336 VPWR VPWR.n1505 0.100405
R15337 VPWR.n1492 VPWR 0.100405
R15338 VPWR VPWR.n1491 0.100405
R15339 VPWR.n1478 VPWR 0.100405
R15340 VPWR VPWR.n1477 0.100405
R15341 VPWR.n1464 VPWR 0.100405
R15342 VPWR VPWR.n1463 0.100405
R15343 VPWR.n1570 VPWR 0.100405
R15344 VPWR.n1571 VPWR 0.100405
R15345 VPWR VPWR.n2734 0.0994583
R15346 VPWR VPWR.n2715 0.0994583
R15347 VPWR VPWR.n1265 0.0981562
R15348 VPWR.n1310 VPWR 0.0981562
R15349 VPWR.n1349 VPWR 0.0981562
R15350 VPWR.n9 VPWR 0.0968542
R15351 VPWR.n1183 VPWR 0.0968542
R15352 VPWR.n1206 VPWR 0.0968542
R15353 VPWR.n1230 VPWR 0.0968542
R15354 VPWR.n1272 VPWR 0.0968542
R15355 VPWR VPWR.n2695 0.0968542
R15356 VPWR VPWR.n2676 0.0968542
R15357 VPWR.n2654 VPWR 0.0968542
R15358 VPWR.n2618 VPWR 0.0968542
R15359 VPWR.n2581 VPWR 0.0968542
R15360 VPWR.n2544 VPWR 0.0968542
R15361 VPWR VPWR.n1012 0.0945
R15362 VPWR.n1519 VPWR 0.0945
R15363 VPWR VPWR.n1406 0.0945
R15364 VPWR VPWR.n1405 0.0945
R15365 VPWR VPWR.n1404 0.0945
R15366 VPWR VPWR.n1403 0.0945
R15367 VPWR VPWR.n1402 0.0945
R15368 VPWR VPWR.n1401 0.0945
R15369 VPWR.n1400 VPWR 0.0945
R15370 VPWR VPWR.n1566 0.0945
R15371 VPWR VPWR.n1170 0.0945
R15372 VPWR.n1390 VPWR 0.0945
R15373 VPWR VPWR.n1006 0.0945
R15374 VPWR.n1722 VPWR 0.0945
R15375 VPWR VPWR.n995 0.0945
R15376 VPWR.n1702 VPWR 0.0945
R15377 VPWR.n2534 VPWR 0.0849042
R15378 VPWR.n1394 VPWR.n1390 0.0740128
R15379 VPWR.n1113 VPWR 0.0737759
R15380 VPWR.n106 VPWR 0.0737759
R15381 VPWR.n134 VPWR 0.0737759
R15382 VPWR.n144 VPWR 0.0737759
R15383 VPWR.n154 VPWR 0.0737759
R15384 VPWR.n164 VPWR 0.0737759
R15385 VPWR.n174 VPWR 0.0737759
R15386 VPWR.n184 VPWR 0.0737759
R15387 VPWR.n194 VPWR 0.0737759
R15388 VPWR.n204 VPWR 0.0737759
R15389 VPWR.n214 VPWR 0.0737759
R15390 VPWR.n224 VPWR 0.0737759
R15391 VPWR.n234 VPWR 0.0737759
R15392 VPWR.n244 VPWR 0.0737759
R15393 VPWR VPWR.n254 0.0737759
R15394 VPWR.n124 VPWR 0.0737759
R15395 VPWR.n115 VPWR 0.0737759
R15396 VPWR VPWR.n1668 0.0737759
R15397 VPWR.n1659 VPWR 0.0737759
R15398 VPWR.n1649 VPWR 0.0737759
R15399 VPWR.n1643 VPWR 0.0737759
R15400 VPWR.n1637 VPWR 0.0737759
R15401 VPWR.n1631 VPWR 0.0737759
R15402 VPWR.n1625 VPWR 0.0737759
R15403 VPWR.n1619 VPWR 0.0737759
R15404 VPWR.n1613 VPWR 0.0737759
R15405 VPWR.n1607 VPWR 0.0737759
R15406 VPWR.n1601 VPWR 0.0737759
R15407 VPWR.n1595 VPWR 0.0737759
R15408 VPWR.n1589 VPWR 0.0737759
R15409 VPWR.n1583 VPWR 0.0737759
R15410 VPWR.n1577 VPWR 0.0737759
R15411 VPWR.n1520 VPWR.n1012 0.071
R15412 VPWR.n1525 VPWR.n1519 0.071
R15413 VPWR.n1530 VPWR.n1406 0.071
R15414 VPWR.n1535 VPWR.n1405 0.071
R15415 VPWR.n1540 VPWR.n1404 0.071
R15416 VPWR.n1545 VPWR.n1403 0.071
R15417 VPWR.n1550 VPWR.n1402 0.071
R15418 VPWR.n1555 VPWR.n1401 0.071
R15419 VPWR.n1560 VPWR.n1400 0.071
R15420 VPWR.n1566 VPWR.n1565 0.071
R15421 VPWR.n1395 VPWR.n1170 0.071
R15422 VPWR.n1708 VPWR.n1006 0.071
R15423 VPWR.n1722 VPWR.n1721 0.071
R15424 VPWR.n1716 VPWR.n995 0.071
R15425 VPWR.n1703 VPWR.n1702 0.071
R15426 VPWR.n1112 VPWR.n1110 0.0645244
R15427 VPWR.n138 VPWR.n136 0.0645244
R15428 VPWR.n148 VPWR.n146 0.0645244
R15429 VPWR.n158 VPWR.n156 0.0645244
R15430 VPWR.n168 VPWR.n166 0.0645244
R15431 VPWR.n178 VPWR.n176 0.0645244
R15432 VPWR.n188 VPWR.n186 0.0645244
R15433 VPWR.n198 VPWR.n196 0.0645244
R15434 VPWR.n208 VPWR.n206 0.0645244
R15435 VPWR.n218 VPWR.n216 0.0645244
R15436 VPWR.n228 VPWR.n226 0.0645244
R15437 VPWR.n238 VPWR.n236 0.0645244
R15438 VPWR.n248 VPWR.n246 0.0645244
R15439 VPWR.n253 VPWR.n251 0.0645244
R15440 VPWR.n110 VPWR.n108 0.0645244
R15441 VPWR.n128 VPWR.n126 0.0645244
R15442 VPWR.n119 VPWR.n117 0.0645244
R15443 VPWR.n1667 VPWR.n1665 0.0645244
R15444 VPWR.n1663 VPWR.n1661 0.0645244
R15445 VPWR.n1653 VPWR.n1651 0.0645244
R15446 VPWR.n1041 VPWR.n1039 0.0645244
R15447 VPWR.n1078 VPWR.n1044 0.0645244
R15448 VPWR.n1081 VPWR.n1047 0.0645244
R15449 VPWR.n1084 VPWR.n1050 0.0645244
R15450 VPWR.n1087 VPWR.n1053 0.0645244
R15451 VPWR.n1090 VPWR.n1056 0.0645244
R15452 VPWR.n1093 VPWR.n1059 0.0645244
R15453 VPWR.n1096 VPWR.n1062 0.0645244
R15454 VPWR.n1099 VPWR.n1065 0.0645244
R15455 VPWR.n1102 VPWR.n1068 0.0645244
R15456 VPWR.n1105 VPWR.n1071 0.0645244
R15457 VPWR.n1108 VPWR.n1074 0.0645244
R15458 VPWR VPWR.n133 0.063
R15459 VPWR.n141 VPWR 0.063
R15460 VPWR VPWR.n143 0.063
R15461 VPWR.n151 VPWR 0.063
R15462 VPWR VPWR.n153 0.063
R15463 VPWR.n161 VPWR 0.063
R15464 VPWR VPWR.n163 0.063
R15465 VPWR.n171 VPWR 0.063
R15466 VPWR VPWR.n173 0.063
R15467 VPWR.n181 VPWR 0.063
R15468 VPWR VPWR.n183 0.063
R15469 VPWR.n191 VPWR 0.063
R15470 VPWR VPWR.n193 0.063
R15471 VPWR.n201 VPWR 0.063
R15472 VPWR VPWR.n203 0.063
R15473 VPWR.n211 VPWR 0.063
R15474 VPWR VPWR.n213 0.063
R15475 VPWR.n221 VPWR 0.063
R15476 VPWR VPWR.n223 0.063
R15477 VPWR.n231 VPWR 0.063
R15478 VPWR VPWR.n233 0.063
R15479 VPWR.n241 VPWR 0.063
R15480 VPWR VPWR.n243 0.063
R15481 VPWR.n101 VPWR 0.063
R15482 VPWR.n256 VPWR 0.063
R15483 VPWR.n105 VPWR 0.063
R15484 VPWR VPWR.n123 0.063
R15485 VPWR.n131 VPWR 0.063
R15486 VPWR.n112 VPWR 0.063
R15487 VPWR VPWR.n114 0.063
R15488 VPWR.n121 VPWR 0.063
R15489 VPWR.n1033 VPWR 0.063
R15490 VPWR.n1670 VPWR 0.063
R15491 VPWR.n1656 VPWR 0.063
R15492 VPWR VPWR.n1658 0.063
R15493 VPWR.n1037 VPWR 0.063
R15494 VPWR VPWR.n1648 0.063
R15495 VPWR VPWR.n1645 0.063
R15496 VPWR VPWR.n1642 0.063
R15497 VPWR VPWR.n1639 0.063
R15498 VPWR VPWR.n1636 0.063
R15499 VPWR VPWR.n1633 0.063
R15500 VPWR VPWR.n1630 0.063
R15501 VPWR VPWR.n1627 0.063
R15502 VPWR VPWR.n1624 0.063
R15503 VPWR VPWR.n1621 0.063
R15504 VPWR VPWR.n1618 0.063
R15505 VPWR VPWR.n1615 0.063
R15506 VPWR VPWR.n1612 0.063
R15507 VPWR VPWR.n1609 0.063
R15508 VPWR VPWR.n1606 0.063
R15509 VPWR VPWR.n1603 0.063
R15510 VPWR VPWR.n1600 0.063
R15511 VPWR VPWR.n1597 0.063
R15512 VPWR VPWR.n1594 0.063
R15513 VPWR VPWR.n1591 0.063
R15514 VPWR VPWR.n1588 0.063
R15515 VPWR VPWR.n1585 0.063
R15516 VPWR VPWR.n1582 0.063
R15517 VPWR VPWR.n1579 0.063
R15518 VPWR VPWR.n1576 0.063
R15519 VPWR VPWR.n1115 0.063
R15520 VPWR VPWR.n13 0.0603958
R15521 VPWR VPWR.n12 0.0603958
R15522 VPWR VPWR.n1188 0.0603958
R15523 VPWR VPWR.n1187 0.0603958
R15524 VPWR VPWR.n1211 0.0603958
R15525 VPWR VPWR.n1210 0.0603958
R15526 VPWR VPWR.n1235 0.0603958
R15527 VPWR VPWR.n1234 0.0603958
R15528 VPWR.n1271 VPWR 0.0603958
R15529 VPWR VPWR.n1270 0.0603958
R15530 VPWR.n1266 VPWR 0.0603958
R15531 VPWR.n1257 VPWR 0.0603958
R15532 VPWR VPWR.n1256 0.0603958
R15533 VPWR.n1309 VPWR 0.0603958
R15534 VPWR VPWR.n1308 0.0603958
R15535 VPWR.n1303 VPWR 0.0603958
R15536 VPWR.n1348 VPWR 0.0603958
R15537 VPWR VPWR.n1347 0.0603958
R15538 VPWR.n1342 VPWR 0.0603958
R15539 VPWR.n1379 VPWR 0.0603958
R15540 VPWR VPWR.n2736 0.0603958
R15541 VPWR VPWR.n2735 0.0603958
R15542 VPWR VPWR.n2748 0.0603958
R15543 VPWR.n2727 VPWR 0.0603958
R15544 VPWR.n2728 VPWR 0.0603958
R15545 VPWR VPWR.n2732 0.0603958
R15546 VPWR.n2707 VPWR 0.0603958
R15547 VPWR.n2708 VPWR 0.0603958
R15548 VPWR VPWR.n2713 0.0603958
R15549 VPWR.n2688 VPWR 0.0603958
R15550 VPWR.n2689 VPWR 0.0603958
R15551 VPWR VPWR.n2693 0.0603958
R15552 VPWR.n2669 VPWR 0.0603958
R15553 VPWR.n2670 VPWR 0.0603958
R15554 VPWR VPWR.n2631 0.0603958
R15555 VPWR.n2632 VPWR 0.0603958
R15556 VPWR.n2633 VPWR 0.0603958
R15557 VPWR VPWR.n2594 0.0603958
R15558 VPWR.n2595 VPWR 0.0603958
R15559 VPWR.n2596 VPWR 0.0603958
R15560 VPWR.n2560 VPWR 0.0603958
R15561 VPWR.n2563 VPWR 0.0603958
R15562 VPWR.n1110 VPWR.n1076 0.0599512
R15563 VPWR.n1706 VPWR.n1705 0.0599512
R15564 VPWR.n1009 VPWR.n1008 0.0599512
R15565 VPWR.n1523 VPWR.n1522 0.0599512
R15566 VPWR.n1528 VPWR.n1527 0.0599512
R15567 VPWR.n1533 VPWR.n1532 0.0599512
R15568 VPWR.n1538 VPWR.n1537 0.0599512
R15569 VPWR.n1543 VPWR.n1542 0.0599512
R15570 VPWR.n1548 VPWR.n1547 0.0599512
R15571 VPWR.n1553 VPWR.n1552 0.0599512
R15572 VPWR.n1558 VPWR.n1557 0.0599512
R15573 VPWR.n1563 VPWR.n1562 0.0599512
R15574 VPWR.n1398 VPWR.n1397 0.0599512
R15575 VPWR.n1393 VPWR.n1392 0.0599512
R15576 VPWR.n1711 VPWR.n1710 0.0599512
R15577 VPWR.n1719 VPWR.n1718 0.0599512
R15578 VPWR.n1715 VPWR.n1714 0.0599512
R15579 VPWR.n138 VPWR.n137 0.0599512
R15580 VPWR.n148 VPWR.n147 0.0599512
R15581 VPWR.n158 VPWR.n157 0.0599512
R15582 VPWR.n168 VPWR.n167 0.0599512
R15583 VPWR.n178 VPWR.n177 0.0599512
R15584 VPWR.n188 VPWR.n187 0.0599512
R15585 VPWR.n198 VPWR.n197 0.0599512
R15586 VPWR.n208 VPWR.n207 0.0599512
R15587 VPWR.n218 VPWR.n217 0.0599512
R15588 VPWR.n228 VPWR.n227 0.0599512
R15589 VPWR.n238 VPWR.n237 0.0599512
R15590 VPWR.n248 VPWR.n247 0.0599512
R15591 VPWR.n251 VPWR.n102 0.0599512
R15592 VPWR.n110 VPWR.n109 0.0599512
R15593 VPWR.n128 VPWR.n127 0.0599512
R15594 VPWR.n119 VPWR.n118 0.0599512
R15595 VPWR.n1665 VPWR.n1034 0.0599512
R15596 VPWR.n1663 VPWR.n1662 0.0599512
R15597 VPWR.n1653 VPWR.n1652 0.0599512
R15598 VPWR.n1039 VPWR.n1038 0.0599512
R15599 VPWR.n1078 VPWR.n1077 0.0599512
R15600 VPWR.n1081 VPWR.n1080 0.0599512
R15601 VPWR.n1084 VPWR.n1083 0.0599512
R15602 VPWR.n1087 VPWR.n1086 0.0599512
R15603 VPWR.n1090 VPWR.n1089 0.0599512
R15604 VPWR.n1093 VPWR.n1092 0.0599512
R15605 VPWR.n1096 VPWR.n1095 0.0599512
R15606 VPWR.n1099 VPWR.n1098 0.0599512
R15607 VPWR.n1102 VPWR.n1101 0.0599512
R15608 VPWR.n1105 VPWR.n1104 0.0599512
R15609 VPWR.n1108 VPWR.n1107 0.0599512
R15610 VPWR.n1107 VPWR 0.0469286
R15611 VPWR.n1104 VPWR 0.0469286
R15612 VPWR.n1101 VPWR 0.0469286
R15613 VPWR.n1098 VPWR 0.0469286
R15614 VPWR.n1095 VPWR 0.0469286
R15615 VPWR.n1092 VPWR 0.0469286
R15616 VPWR.n1089 VPWR 0.0469286
R15617 VPWR.n1086 VPWR 0.0469286
R15618 VPWR.n1083 VPWR 0.0469286
R15619 VPWR.n1080 VPWR 0.0469286
R15620 VPWR.n1077 VPWR 0.0469286
R15621 VPWR.n1038 VPWR 0.0469286
R15622 VPWR.n1652 VPWR 0.0469286
R15623 VPWR.n1662 VPWR 0.0469286
R15624 VPWR.n1076 VPWR 0.0469286
R15625 VPWR.n1034 VPWR 0.0469286
R15626 VPWR.n118 VPWR 0.0469286
R15627 VPWR.n109 VPWR 0.0469286
R15628 VPWR.n102 VPWR 0.0469286
R15629 VPWR.n247 VPWR 0.0469286
R15630 VPWR.n237 VPWR 0.0469286
R15631 VPWR.n227 VPWR 0.0469286
R15632 VPWR.n217 VPWR 0.0469286
R15633 VPWR.n207 VPWR 0.0469286
R15634 VPWR.n197 VPWR 0.0469286
R15635 VPWR.n187 VPWR 0.0469286
R15636 VPWR.n177 VPWR 0.0469286
R15637 VPWR.n167 VPWR 0.0469286
R15638 VPWR.n157 VPWR 0.0469286
R15639 VPWR.n147 VPWR 0.0469286
R15640 VPWR.n1705 VPWR 0.0469286
R15641 VPWR.n1008 VPWR 0.0469286
R15642 VPWR.n1522 VPWR 0.0469286
R15643 VPWR.n1527 VPWR 0.0469286
R15644 VPWR.n1532 VPWR 0.0469286
R15645 VPWR.n1537 VPWR 0.0469286
R15646 VPWR.n1542 VPWR 0.0469286
R15647 VPWR.n1547 VPWR 0.0469286
R15648 VPWR.n1552 VPWR 0.0469286
R15649 VPWR.n1557 VPWR 0.0469286
R15650 VPWR.n1562 VPWR 0.0469286
R15651 VPWR.n1397 VPWR 0.0469286
R15652 VPWR.n1392 VPWR 0.0469286
R15653 VPWR.n1710 VPWR 0.0469286
R15654 VPWR.n1718 VPWR 0.0469286
R15655 VPWR.n1714 VPWR 0.0469286
R15656 VPWR.n137 VPWR 0.0469286
R15657 VPWR.n127 VPWR 0.0469286
R15658 VPWR.n1076 VPWR 0.0401341
R15659 VPWR.n1705 VPWR 0.0401341
R15660 VPWR.n1008 VPWR 0.0401341
R15661 VPWR.n1522 VPWR 0.0401341
R15662 VPWR.n1527 VPWR 0.0401341
R15663 VPWR.n1532 VPWR 0.0401341
R15664 VPWR.n1537 VPWR 0.0401341
R15665 VPWR.n1542 VPWR 0.0401341
R15666 VPWR.n1547 VPWR 0.0401341
R15667 VPWR.n1552 VPWR 0.0401341
R15668 VPWR.n1557 VPWR 0.0401341
R15669 VPWR.n1562 VPWR 0.0401341
R15670 VPWR.n1397 VPWR 0.0401341
R15671 VPWR.n1392 VPWR 0.0401341
R15672 VPWR.n1710 VPWR 0.0401341
R15673 VPWR.n1718 VPWR 0.0401341
R15674 VPWR.n1714 VPWR 0.0401341
R15675 VPWR.n137 VPWR 0.0401341
R15676 VPWR.n147 VPWR 0.0401341
R15677 VPWR.n157 VPWR 0.0401341
R15678 VPWR.n167 VPWR 0.0401341
R15679 VPWR.n177 VPWR 0.0401341
R15680 VPWR.n187 VPWR 0.0401341
R15681 VPWR.n197 VPWR 0.0401341
R15682 VPWR.n207 VPWR 0.0401341
R15683 VPWR.n217 VPWR 0.0401341
R15684 VPWR.n227 VPWR 0.0401341
R15685 VPWR.n237 VPWR 0.0401341
R15686 VPWR.n247 VPWR 0.0401341
R15687 VPWR.n102 VPWR 0.0401341
R15688 VPWR.n109 VPWR 0.0401341
R15689 VPWR.n127 VPWR 0.0401341
R15690 VPWR.n118 VPWR 0.0401341
R15691 VPWR.n1034 VPWR 0.0401341
R15692 VPWR.n1662 VPWR 0.0401341
R15693 VPWR.n1652 VPWR 0.0401341
R15694 VPWR.n1038 VPWR 0.0401341
R15695 VPWR.n1077 VPWR 0.0401341
R15696 VPWR.n1080 VPWR 0.0401341
R15697 VPWR.n1083 VPWR 0.0401341
R15698 VPWR.n1086 VPWR 0.0401341
R15699 VPWR.n1089 VPWR 0.0401341
R15700 VPWR.n1092 VPWR 0.0401341
R15701 VPWR.n1095 VPWR 0.0401341
R15702 VPWR.n1098 VPWR 0.0401341
R15703 VPWR.n1101 VPWR 0.0401341
R15704 VPWR.n1104 VPWR 0.0401341
R15705 VPWR.n1107 VPWR 0.0401341
R15706 VPWR.n13 VPWR 0.0382604
R15707 VPWR.n1188 VPWR 0.0382604
R15708 VPWR.n1211 VPWR 0.0382604
R15709 VPWR.n1235 VPWR 0.0382604
R15710 VPWR.n1270 VPWR 0.0382604
R15711 VPWR.n1308 VPWR 0.0382604
R15712 VPWR.n1347 VPWR 0.0382604
R15713 VPWR.n1384 VPWR 0.0382604
R15714 VPWR.n2440 VPWR 0.0377024
R15715 VPWR.n2505 VPWR 0.0377024
R15716 VPWR.n2445 VPWR 0.0377024
R15717 VPWR.n2488 VPWR 0.0377024
R15718 VPWR.n2481 VPWR 0.0377024
R15719 VPWR.n2469 VPWR 0.0377024
R15720 VPWR.n2464 VPWR 0.0377024
R15721 VPWR.n1150 VPWR 0.0377024
R15722 VPWR.n2457 VPWR 0.0377024
R15723 VPWR.n1154 VPWR 0.0377024
R15724 VPWR.n1146 VPWR 0.0377024
R15725 VPWR.n2476 VPWR 0.0377024
R15726 VPWR.n1142 VPWR 0.0377024
R15727 VPWR.n1138 VPWR 0.0377024
R15728 VPWR.n2452 VPWR 0.0377024
R15729 VPWR.n1158 VPWR 0.0377024
R15730 VPWR.n1134 VPWR 0.0377024
R15731 VPWR.n2493 VPWR 0.0377024
R15732 VPWR.n1130 VPWR 0.0377024
R15733 VPWR.n1162 VPWR 0.0377024
R15734 VPWR.n2500 VPWR 0.0377024
R15735 VPWR.n1126 VPWR 0.0377024
R15736 VPWR.n1122 VPWR 0.0377024
R15737 VPWR.n1678 VPWR 0.0377024
R15738 VPWR.n1118 VPWR 0.0377024
R15739 VPWR.n2512 VPWR 0.0377024
R15740 VPWR.n2517 VPWR 0.0377024
R15741 VPWR.n2528 VPWR 0.0377024
R15742 VPWR.n2524 VPWR 0.0377024
R15743 VPWR.n1673 VPWR 0.0377024
R15744 VPWR.n1030 VPWR 0.0377024
R15745 VPWR.n1167 VPWR 0.0377024
R15746 VPWR.n20 VPWR 0.0375125
R15747 VPWR.n20 VPWR 0.0373589
R15748 VPWR.n2564 VPWR.n2534 0.0320292
R15749 VPWR.n2736 VPWR 0.03175
R15750 VPWR VPWR.n2727 0.03175
R15751 VPWR VPWR.n2707 0.03175
R15752 VPWR VPWR.n2688 0.03175
R15753 VPWR VPWR.n2669 0.03175
R15754 VPWR VPWR.n2632 0.03175
R15755 VPWR VPWR.n2595 0.03175
R15756 VPWR VPWR.n2563 0.03175
R15757 VPWR.n2534 VPWR.n2533 0.0240975
R15758 VPWR.n2533 VPWR.n20 0.0240975
R15759 VPWR.n2750 VPWR 0.024
R15760 VPWR.n14 VPWR 0.0239375
R15761 VPWR.n12 VPWR 0.0239375
R15762 VPWR.n1189 VPWR 0.0239375
R15763 VPWR.n1187 VPWR 0.0239375
R15764 VPWR.n1210 VPWR 0.0239375
R15765 VPWR.n1234 VPWR 0.0239375
R15766 VPWR.n2689 VPWR 0.0239375
R15767 VPWR.n1449 VPWR 0.0233659
R15768 VPWR.n320 VPWR 0.0233659
R15769 VPWR.n1511 VPWR 0.0233659
R15770 VPWR.n315 VPWR 0.0233659
R15771 VPWR.n932 VPWR 0.0233659
R15772 VPWR.n2415 VPWR 0.0233659
R15773 VPWR.n2410 VPWR 0.0233659
R15774 VPWR.n287 VPWR 0.0233659
R15775 VPWR.n940 VPWR 0.0233659
R15776 VPWR.n2380 VPWR 0.0233659
R15777 VPWR.n291 VPWR 0.0233659
R15778 VPWR.n1827 VPWR 0.0233659
R15779 VPWR.n1822 VPWR 0.0233659
R15780 VPWR.n1817 VPWR 0.0233659
R15781 VPWR.n356 VPWR 0.0233659
R15782 VPWR.n360 VPWR 0.0233659
R15783 VPWR.n364 VPWR 0.0233659
R15784 VPWR.n2390 VPWR 0.0233659
R15785 VPWR.n299 VPWR 0.0233659
R15786 VPWR.n1812 VPWR 0.0233659
R15787 VPWR.n372 VPWR 0.0233659
R15788 VPWR.n2395 VPWR 0.0233659
R15789 VPWR.n303 VPWR 0.0233659
R15790 VPWR.n2243 VPWR 0.0233659
R15791 VPWR.n2248 VPWR 0.0233659
R15792 VPWR.n2253 VPWR 0.0233659
R15793 VPWR.n2258 VPWR 0.0233659
R15794 VPWR.n2268 VPWR 0.0233659
R15795 VPWR.n2273 VPWR 0.0233659
R15796 VPWR.n2278 VPWR 0.0233659
R15797 VPWR.n2283 VPWR 0.0233659
R15798 VPWR.n2288 VPWR 0.0233659
R15799 VPWR.n2293 VPWR 0.0233659
R15800 VPWR.n2298 VPWR 0.0233659
R15801 VPWR.n2303 VPWR 0.0233659
R15802 VPWR.n2308 VPWR 0.0233659
R15803 VPWR.n2313 VPWR 0.0233659
R15804 VPWR.n2317 VPWR 0.0233659
R15805 VPWR.n2263 VPWR 0.0233659
R15806 VPWR.n512 VPWR 0.0233659
R15807 VPWR.n507 VPWR 0.0233659
R15808 VPWR.n503 VPWR 0.0233659
R15809 VPWR.n499 VPWR 0.0233659
R15810 VPWR.n491 VPWR 0.0233659
R15811 VPWR.n487 VPWR 0.0233659
R15812 VPWR.n483 VPWR 0.0233659
R15813 VPWR.n479 VPWR 0.0233659
R15814 VPWR.n475 VPWR 0.0233659
R15815 VPWR.n471 VPWR 0.0233659
R15816 VPWR.n467 VPWR 0.0233659
R15817 VPWR.n463 VPWR 0.0233659
R15818 VPWR.n459 VPWR 0.0233659
R15819 VPWR.n455 VPWR 0.0233659
R15820 VPWR.n452 VPWR 0.0233659
R15821 VPWR.n495 VPWR 0.0233659
R15822 VPWR.n2219 VPWR 0.0233659
R15823 VPWR.n2214 VPWR 0.0233659
R15824 VPWR.n2209 VPWR 0.0233659
R15825 VPWR.n2204 VPWR 0.0233659
R15826 VPWR.n2194 VPWR 0.0233659
R15827 VPWR.n2189 VPWR 0.0233659
R15828 VPWR.n2184 VPWR 0.0233659
R15829 VPWR.n2179 VPWR 0.0233659
R15830 VPWR.n2174 VPWR 0.0233659
R15831 VPWR.n2169 VPWR 0.0233659
R15832 VPWR.n2164 VPWR 0.0233659
R15833 VPWR.n2159 VPWR 0.0233659
R15834 VPWR.n2154 VPWR 0.0233659
R15835 VPWR.n2149 VPWR 0.0233659
R15836 VPWR.n2145 VPWR 0.0233659
R15837 VPWR.n2199 VPWR 0.0233659
R15838 VPWR.n548 VPWR 0.0233659
R15839 VPWR.n552 VPWR 0.0233659
R15840 VPWR.n556 VPWR 0.0233659
R15841 VPWR.n560 VPWR 0.0233659
R15842 VPWR.n568 VPWR 0.0233659
R15843 VPWR.n572 VPWR 0.0233659
R15844 VPWR.n576 VPWR 0.0233659
R15845 VPWR.n580 VPWR 0.0233659
R15846 VPWR.n584 VPWR 0.0233659
R15847 VPWR.n588 VPWR 0.0233659
R15848 VPWR.n592 VPWR 0.0233659
R15849 VPWR.n596 VPWR 0.0233659
R15850 VPWR.n600 VPWR 0.0233659
R15851 VPWR.n604 VPWR 0.0233659
R15852 VPWR.n608 VPWR 0.0233659
R15853 VPWR.n564 VPWR 0.0233659
R15854 VPWR.n2047 VPWR 0.0233659
R15855 VPWR.n2052 VPWR 0.0233659
R15856 VPWR.n2057 VPWR 0.0233659
R15857 VPWR.n2062 VPWR 0.0233659
R15858 VPWR.n2072 VPWR 0.0233659
R15859 VPWR.n2077 VPWR 0.0233659
R15860 VPWR.n2082 VPWR 0.0233659
R15861 VPWR.n2087 VPWR 0.0233659
R15862 VPWR.n2092 VPWR 0.0233659
R15863 VPWR.n2097 VPWR 0.0233659
R15864 VPWR.n2102 VPWR 0.0233659
R15865 VPWR.n2107 VPWR 0.0233659
R15866 VPWR.n2112 VPWR 0.0233659
R15867 VPWR.n2117 VPWR 0.0233659
R15868 VPWR.n2121 VPWR 0.0233659
R15869 VPWR.n2067 VPWR 0.0233659
R15870 VPWR.n704 VPWR 0.0233659
R15871 VPWR.n699 VPWR 0.0233659
R15872 VPWR.n695 VPWR 0.0233659
R15873 VPWR.n691 VPWR 0.0233659
R15874 VPWR.n683 VPWR 0.0233659
R15875 VPWR.n679 VPWR 0.0233659
R15876 VPWR.n675 VPWR 0.0233659
R15877 VPWR.n671 VPWR 0.0233659
R15878 VPWR.n667 VPWR 0.0233659
R15879 VPWR.n663 VPWR 0.0233659
R15880 VPWR.n659 VPWR 0.0233659
R15881 VPWR.n655 VPWR 0.0233659
R15882 VPWR.n651 VPWR 0.0233659
R15883 VPWR.n647 VPWR 0.0233659
R15884 VPWR.n644 VPWR 0.0233659
R15885 VPWR.n687 VPWR 0.0233659
R15886 VPWR.n2023 VPWR 0.0233659
R15887 VPWR.n2018 VPWR 0.0233659
R15888 VPWR.n2013 VPWR 0.0233659
R15889 VPWR.n2008 VPWR 0.0233659
R15890 VPWR.n1998 VPWR 0.0233659
R15891 VPWR.n1993 VPWR 0.0233659
R15892 VPWR.n1988 VPWR 0.0233659
R15893 VPWR.n1983 VPWR 0.0233659
R15894 VPWR.n1978 VPWR 0.0233659
R15895 VPWR.n1973 VPWR 0.0233659
R15896 VPWR.n1968 VPWR 0.0233659
R15897 VPWR.n1963 VPWR 0.0233659
R15898 VPWR.n1958 VPWR 0.0233659
R15899 VPWR.n1953 VPWR 0.0233659
R15900 VPWR.n1949 VPWR 0.0233659
R15901 VPWR.n2003 VPWR 0.0233659
R15902 VPWR.n740 VPWR 0.0233659
R15903 VPWR.n744 VPWR 0.0233659
R15904 VPWR.n748 VPWR 0.0233659
R15905 VPWR.n752 VPWR 0.0233659
R15906 VPWR.n760 VPWR 0.0233659
R15907 VPWR.n764 VPWR 0.0233659
R15908 VPWR.n768 VPWR 0.0233659
R15909 VPWR.n772 VPWR 0.0233659
R15910 VPWR.n776 VPWR 0.0233659
R15911 VPWR.n780 VPWR 0.0233659
R15912 VPWR.n784 VPWR 0.0233659
R15913 VPWR.n788 VPWR 0.0233659
R15914 VPWR.n792 VPWR 0.0233659
R15915 VPWR.n796 VPWR 0.0233659
R15916 VPWR.n800 VPWR 0.0233659
R15917 VPWR.n756 VPWR 0.0233659
R15918 VPWR.n1851 VPWR 0.0233659
R15919 VPWR.n1856 VPWR 0.0233659
R15920 VPWR.n1861 VPWR 0.0233659
R15921 VPWR.n1866 VPWR 0.0233659
R15922 VPWR.n1876 VPWR 0.0233659
R15923 VPWR.n1881 VPWR 0.0233659
R15924 VPWR.n1886 VPWR 0.0233659
R15925 VPWR.n1891 VPWR 0.0233659
R15926 VPWR.n1896 VPWR 0.0233659
R15927 VPWR.n1901 VPWR 0.0233659
R15928 VPWR.n1906 VPWR 0.0233659
R15929 VPWR.n1911 VPWR 0.0233659
R15930 VPWR.n1916 VPWR 0.0233659
R15931 VPWR.n1921 VPWR 0.0233659
R15932 VPWR.n1925 VPWR 0.0233659
R15933 VPWR.n1871 VPWR 0.0233659
R15934 VPWR.n896 VPWR 0.0233659
R15935 VPWR.n891 VPWR 0.0233659
R15936 VPWR.n887 VPWR 0.0233659
R15937 VPWR.n883 VPWR 0.0233659
R15938 VPWR.n875 VPWR 0.0233659
R15939 VPWR.n871 VPWR 0.0233659
R15940 VPWR.n867 VPWR 0.0233659
R15941 VPWR.n863 VPWR 0.0233659
R15942 VPWR.n859 VPWR 0.0233659
R15943 VPWR.n855 VPWR 0.0233659
R15944 VPWR.n851 VPWR 0.0233659
R15945 VPWR.n847 VPWR 0.0233659
R15946 VPWR.n843 VPWR 0.0233659
R15947 VPWR.n839 VPWR 0.0233659
R15948 VPWR.n836 VPWR 0.0233659
R15949 VPWR.n879 VPWR 0.0233659
R15950 VPWR.n1807 VPWR 0.0233659
R15951 VPWR.n948 VPWR 0.0233659
R15952 VPWR.n1473 VPWR 0.0233659
R15953 VPWR.n368 VPWR 0.0233659
R15954 VPWR.n2400 VPWR 0.0233659
R15955 VPWR.n307 VPWR 0.0233659
R15956 VPWR.n944 VPWR 0.0233659
R15957 VPWR.n1468 VPWR 0.0233659
R15958 VPWR.n1802 VPWR 0.0233659
R15959 VPWR.n952 VPWR 0.0233659
R15960 VPWR.n1482 VPWR 0.0233659
R15961 VPWR.n376 VPWR 0.0233659
R15962 VPWR.n384 VPWR 0.0233659
R15963 VPWR.n388 VPWR 0.0233659
R15964 VPWR.n392 VPWR 0.0233659
R15965 VPWR.n396 VPWR 0.0233659
R15966 VPWR.n400 VPWR 0.0233659
R15967 VPWR.n404 VPWR 0.0233659
R15968 VPWR.n408 VPWR 0.0233659
R15969 VPWR.n412 VPWR 0.0233659
R15970 VPWR.n416 VPWR 0.0233659
R15971 VPWR.n380 VPWR 0.0233659
R15972 VPWR.n2385 VPWR 0.0233659
R15973 VPWR.n295 VPWR 0.0233659
R15974 VPWR.n956 VPWR 0.0233659
R15975 VPWR.n1487 VPWR 0.0233659
R15976 VPWR.n1797 VPWR 0.0233659
R15977 VPWR.n1787 VPWR 0.0233659
R15978 VPWR.n1782 VPWR 0.0233659
R15979 VPWR.n1777 VPWR 0.0233659
R15980 VPWR.n1772 VPWR 0.0233659
R15981 VPWR.n1767 VPWR 0.0233659
R15982 VPWR.n1762 VPWR 0.0233659
R15983 VPWR.n1757 VPWR 0.0233659
R15984 VPWR.n1753 VPWR 0.0233659
R15985 VPWR.n1792 VPWR 0.0233659
R15986 VPWR.n960 VPWR 0.0233659
R15987 VPWR.n1496 VPWR 0.0233659
R15988 VPWR.n2405 VPWR 0.0233659
R15989 VPWR.n311 VPWR 0.0233659
R15990 VPWR.n1460 VPWR 0.0233659
R15991 VPWR.n964 VPWR 0.0233659
R15992 VPWR.n1501 VPWR 0.0233659
R15993 VPWR.n2375 VPWR 0.0233659
R15994 VPWR.n2365 VPWR 0.0233659
R15995 VPWR.n2360 VPWR 0.0233659
R15996 VPWR.n2355 VPWR 0.0233659
R15997 VPWR.n2350 VPWR 0.0233659
R15998 VPWR.n2345 VPWR 0.0233659
R15999 VPWR.n2341 VPWR 0.0233659
R16000 VPWR.n2370 VPWR 0.0233659
R16001 VPWR.n283 VPWR 0.0233659
R16002 VPWR.n1516 VPWR 0.0233659
R16003 VPWR.n968 VPWR 0.0233659
R16004 VPWR.n972 VPWR 0.0233659
R16005 VPWR.n976 VPWR 0.0233659
R16006 VPWR.n980 VPWR 0.0233659
R16007 VPWR.n984 VPWR 0.0233659
R16008 VPWR.n988 VPWR 0.0233659
R16009 VPWR.n992 VPWR 0.0233659
R16010 VPWR.n936 VPWR 0.0233659
R16011 VPWR.n1169 VPWR 0.0233659
R16012 VPWR.n279 VPWR 0.0233659
R16013 VPWR.n1699 VPWR 0.0233659
R16014 VPWR.n275 VPWR 0.0233659
R16015 VPWR.n271 VPWR 0.0233659
R16016 VPWR.n263 VPWR 0.0233659
R16017 VPWR.n260 VPWR 0.0233659
R16018 VPWR.n267 VPWR 0.0233659
R16019 VPWR.n1687 VPWR 0.0233659
R16020 VPWR.n1725 VPWR 0.0233659
R16021 VPWR.n1729 VPWR 0.0233659
R16022 VPWR.n1694 VPWR 0.0233659
R16023 VPWR.n1275 VPWR 0.0226354
R16024 VPWR.n1266 VPWR 0.0226354
R16025 VPWR.n1352 VPWR 0.0226354
R16026 VPWR.n2708 VPWR 0.0226354
R16027 VPWR VPWR.n2668 0.0226354
R16028 VPWR VPWR.n2638 0.0226354
R16029 VPWR VPWR.n2600 0.0226354
R16030 VPWR.n1212 VPWR 0.0213333
R16031 VPWR.n1236 VPWR 0.0213333
R16032 VPWR.n1250 VPWR 0.0213333
R16033 VPWR.n1314 VPWR 0.0213333
R16034 VPWR.n1286 VPWR 0.0213333
R16035 VPWR.n1325 VPWR 0.0213333
R16036 VPWR.n1362 VPWR 0.0213333
R16037 VPWR.n2742 VPWR 0.0213333
R16038 VPWR.n2735 VPWR 0.0213333
R16039 VPWR VPWR.n2726 0.0213333
R16040 VPWR.n2728 VPWR 0.0213333
R16041 VPWR VPWR.n2706 0.0213333
R16042 VPWR VPWR.n2687 0.0213333
R16043 VPWR VPWR.n2674 0.0213333
R16044 VPWR.n2436 VPWR 0.0196917
R16045 VPWR VPWR.n19 0.0099
R16046 VPWR.n1113 VPWR.n1112 0.00964634
R16047 VPWR.n136 VPWR.n134 0.00964634
R16048 VPWR.n146 VPWR.n144 0.00964634
R16049 VPWR.n156 VPWR.n154 0.00964634
R16050 VPWR.n166 VPWR.n164 0.00964634
R16051 VPWR.n176 VPWR.n174 0.00964634
R16052 VPWR.n186 VPWR.n184 0.00964634
R16053 VPWR.n196 VPWR.n194 0.00964634
R16054 VPWR.n206 VPWR.n204 0.00964634
R16055 VPWR.n216 VPWR.n214 0.00964634
R16056 VPWR.n226 VPWR.n224 0.00964634
R16057 VPWR.n236 VPWR.n234 0.00964634
R16058 VPWR.n246 VPWR.n244 0.00964634
R16059 VPWR.n254 VPWR.n253 0.00964634
R16060 VPWR.n108 VPWR.n106 0.00964634
R16061 VPWR.n126 VPWR.n124 0.00964634
R16062 VPWR.n117 VPWR.n115 0.00964634
R16063 VPWR.n1668 VPWR.n1667 0.00964634
R16064 VPWR.n1661 VPWR.n1659 0.00964634
R16065 VPWR.n1651 VPWR.n1649 0.00964634
R16066 VPWR.n1643 VPWR.n1041 0.00964634
R16067 VPWR.n1637 VPWR.n1044 0.00964634
R16068 VPWR.n1631 VPWR.n1047 0.00964634
R16069 VPWR.n1625 VPWR.n1050 0.00964634
R16070 VPWR.n1619 VPWR.n1053 0.00964634
R16071 VPWR.n1613 VPWR.n1056 0.00964634
R16072 VPWR.n1607 VPWR.n1059 0.00964634
R16073 VPWR.n1601 VPWR.n1062 0.00964634
R16074 VPWR.n1595 VPWR.n1065 0.00964634
R16075 VPWR.n1589 VPWR.n1068 0.00964634
R16076 VPWR.n1583 VPWR.n1071 0.00964634
R16077 VPWR.n1577 VPWR.n1074 0.00964634
R16078 VPWR VPWR.n64 0.00912069
R16079 VPWR VPWR.n67 0.00912069
R16080 VPWR VPWR.n70 0.00912069
R16081 VPWR VPWR.n73 0.00912069
R16082 VPWR VPWR.n76 0.00912069
R16083 VPWR VPWR.n79 0.00912069
R16084 VPWR VPWR.n82 0.00912069
R16085 VPWR VPWR.n85 0.00912069
R16086 VPWR VPWR.n88 0.00912069
R16087 VPWR VPWR.n91 0.00912069
R16088 VPWR VPWR.n94 0.00912069
R16089 VPWR VPWR.n97 0.00912069
R16090 VPWR.n257 VPWR 0.00912069
R16091 VPWR VPWR.n61 0.00912069
R16092 VPWR VPWR.n58 0.00912069
R16093 VPWR.n1671 VPWR 0.00912069
R16094 VPWR VPWR.n1025 0.00912069
R16095 VPWR.n1646 VPWR 0.00912069
R16096 VPWR.n1640 VPWR 0.00912069
R16097 VPWR.n1634 VPWR 0.00912069
R16098 VPWR.n1628 VPWR 0.00912069
R16099 VPWR.n1622 VPWR 0.00912069
R16100 VPWR.n1616 VPWR 0.00912069
R16101 VPWR.n1610 VPWR 0.00912069
R16102 VPWR.n1604 VPWR 0.00912069
R16103 VPWR.n1598 VPWR 0.00912069
R16104 VPWR.n1592 VPWR 0.00912069
R16105 VPWR.n1586 VPWR 0.00912069
R16106 VPWR.n1580 VPWR 0.00912069
R16107 VPWR.n1574 VPWR 0.00912069
R16108 VPWR.n24 VPWR 0.00744444
R16109 VPWR.n1399 VPWR.n1395 0.00351282
R16110 VPWR.n1565 VPWR.n1564 0.00351282
R16111 VPWR.n1560 VPWR.n1559 0.00351282
R16112 VPWR.n1555 VPWR.n1554 0.00351282
R16113 VPWR.n1550 VPWR.n1549 0.00351282
R16114 VPWR.n1545 VPWR.n1544 0.00351282
R16115 VPWR.n1540 VPWR.n1539 0.00351282
R16116 VPWR.n1535 VPWR.n1534 0.00351282
R16117 VPWR.n1530 VPWR.n1529 0.00351282
R16118 VPWR.n1525 VPWR.n1524 0.00351282
R16119 VPWR.n1520 VPWR.n1010 0.00351282
R16120 VPWR.n1721 VPWR.n1720 0.00351282
R16121 VPWR.n1712 VPWR.n1708 0.00351282
R16122 VPWR.n1707 VPWR.n1703 0.00351282
R16123 VPWR.n2440 VPWR.n2439 0.00347619
R16124 VPWR.n2506 VPWR.n2505 0.00347619
R16125 VPWR.n2446 VPWR.n2445 0.00347619
R16126 VPWR.n2488 VPWR.n2487 0.00347619
R16127 VPWR.n2482 VPWR.n2481 0.00347619
R16128 VPWR.n2470 VPWR.n2469 0.00347619
R16129 VPWR.n2464 VPWR.n2463 0.00347619
R16130 VPWR.n1150 VPWR.n1063 0.00347619
R16131 VPWR.n2458 VPWR.n2457 0.00347619
R16132 VPWR.n1154 VPWR.n1066 0.00347619
R16133 VPWR.n1146 VPWR.n1060 0.00347619
R16134 VPWR.n2476 VPWR.n2475 0.00347619
R16135 VPWR.n1142 VPWR.n1057 0.00347619
R16136 VPWR.n1138 VPWR.n1054 0.00347619
R16137 VPWR.n2452 VPWR.n2451 0.00347619
R16138 VPWR.n1158 VPWR.n1069 0.00347619
R16139 VPWR.n1134 VPWR.n1051 0.00347619
R16140 VPWR.n2494 VPWR.n2493 0.00347619
R16141 VPWR.n1130 VPWR.n1048 0.00347619
R16142 VPWR.n1162 VPWR.n1072 0.00347619
R16143 VPWR.n2500 VPWR.n2499 0.00347619
R16144 VPWR.n1126 VPWR.n1045 0.00347619
R16145 VPWR.n1122 VPWR.n1042 0.00347619
R16146 VPWR.n1679 VPWR.n1678 0.00347619
R16147 VPWR.n1118 VPWR.n1022 0.00347619
R16148 VPWR.n2512 VPWR.n2511 0.00347619
R16149 VPWR.n2518 VPWR.n2517 0.00347619
R16150 VPWR.n2529 VPWR.n2528 0.00347619
R16151 VPWR.n2524 VPWR.n2523 0.00347619
R16152 VPWR.n1673 VPWR.n1672 0.00347619
R16153 VPWR.n1031 VPWR.n1030 0.00347619
R16154 VPWR.n1573 VPWR.n1167 0.00347619
R16155 XThC.Tn[10].n71 XThC.Tn[10].n70 256.104
R16156 XThC.Tn[10].n75 XThC.Tn[10].n74 243.679
R16157 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16158 XThC.Tn[10].n75 XThC.Tn[10].n73 205.28
R16159 XThC.Tn[10].n71 XThC.Tn[10].n69 202.095
R16160 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16161 XThC.Tn[10].n65 XThC.Tn[10].n63 161.365
R16162 XThC.Tn[10].n61 XThC.Tn[10].n59 161.365
R16163 XThC.Tn[10].n57 XThC.Tn[10].n55 161.365
R16164 XThC.Tn[10].n53 XThC.Tn[10].n51 161.365
R16165 XThC.Tn[10].n49 XThC.Tn[10].n47 161.365
R16166 XThC.Tn[10].n45 XThC.Tn[10].n43 161.365
R16167 XThC.Tn[10].n41 XThC.Tn[10].n39 161.365
R16168 XThC.Tn[10].n37 XThC.Tn[10].n35 161.365
R16169 XThC.Tn[10].n33 XThC.Tn[10].n31 161.365
R16170 XThC.Tn[10].n29 XThC.Tn[10].n27 161.365
R16171 XThC.Tn[10].n25 XThC.Tn[10].n23 161.365
R16172 XThC.Tn[10].n21 XThC.Tn[10].n19 161.365
R16173 XThC.Tn[10].n17 XThC.Tn[10].n15 161.365
R16174 XThC.Tn[10].n13 XThC.Tn[10].n11 161.365
R16175 XThC.Tn[10].n9 XThC.Tn[10].n7 161.365
R16176 XThC.Tn[10].n6 XThC.Tn[10].n4 161.365
R16177 XThC.Tn[10].n63 XThC.Tn[10].t30 161.106
R16178 XThC.Tn[10].n59 XThC.Tn[10].t42 161.106
R16179 XThC.Tn[10].n55 XThC.Tn[10].t40 161.106
R16180 XThC.Tn[10].n51 XThC.Tn[10].t39 161.106
R16181 XThC.Tn[10].n47 XThC.Tn[10].t20 161.106
R16182 XThC.Tn[10].n43 XThC.Tn[10].t17 161.106
R16183 XThC.Tn[10].n39 XThC.Tn[10].t37 161.106
R16184 XThC.Tn[10].n35 XThC.Tn[10].t28 161.106
R16185 XThC.Tn[10].n31 XThC.Tn[10].t26 161.106
R16186 XThC.Tn[10].n27 XThC.Tn[10].t15 161.106
R16187 XThC.Tn[10].n23 XThC.Tn[10].t36 161.106
R16188 XThC.Tn[10].n19 XThC.Tn[10].t25 161.106
R16189 XThC.Tn[10].n15 XThC.Tn[10].t14 161.106
R16190 XThC.Tn[10].n11 XThC.Tn[10].t13 161.106
R16191 XThC.Tn[10].n7 XThC.Tn[10].t32 161.106
R16192 XThC.Tn[10].n4 XThC.Tn[10].t22 161.106
R16193 XThC.Tn[10].n63 XThC.Tn[10].t18 154.679
R16194 XThC.Tn[10].n59 XThC.Tn[10].t29 154.679
R16195 XThC.Tn[10].n55 XThC.Tn[10].t27 154.679
R16196 XThC.Tn[10].n51 XThC.Tn[10].t24 154.679
R16197 XThC.Tn[10].n47 XThC.Tn[10].t38 154.679
R16198 XThC.Tn[10].n43 XThC.Tn[10].t35 154.679
R16199 XThC.Tn[10].n39 XThC.Tn[10].t23 154.679
R16200 XThC.Tn[10].n35 XThC.Tn[10].t16 154.679
R16201 XThC.Tn[10].n31 XThC.Tn[10].t12 154.679
R16202 XThC.Tn[10].n27 XThC.Tn[10].t34 154.679
R16203 XThC.Tn[10].n23 XThC.Tn[10].t21 154.679
R16204 XThC.Tn[10].n19 XThC.Tn[10].t43 154.679
R16205 XThC.Tn[10].n15 XThC.Tn[10].t33 154.679
R16206 XThC.Tn[10].n11 XThC.Tn[10].t31 154.679
R16207 XThC.Tn[10].n7 XThC.Tn[10].t19 154.679
R16208 XThC.Tn[10].n4 XThC.Tn[10].t41 154.679
R16209 XThC.Tn[10].n69 XThC.Tn[10].t4 26.5955
R16210 XThC.Tn[10].n69 XThC.Tn[10].t3 26.5955
R16211 XThC.Tn[10].n70 XThC.Tn[10].t6 26.5955
R16212 XThC.Tn[10].n70 XThC.Tn[10].t9 26.5955
R16213 XThC.Tn[10].n73 XThC.Tn[10].t11 26.5955
R16214 XThC.Tn[10].n73 XThC.Tn[10].t10 26.5955
R16215 XThC.Tn[10].n74 XThC.Tn[10].t0 26.5955
R16216 XThC.Tn[10].n74 XThC.Tn[10].t8 26.5955
R16217 XThC.Tn[10].n1 XThC.Tn[10].t7 24.9236
R16218 XThC.Tn[10].n1 XThC.Tn[10].t2 24.9236
R16219 XThC.Tn[10].n0 XThC.Tn[10].t1 24.9236
R16220 XThC.Tn[10].n0 XThC.Tn[10].t5 24.9236
R16221 XThC.Tn[10] XThC.Tn[10].n75 22.9652
R16222 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16223 XThC.Tn[10].n72 XThC.Tn[10].n71 13.9299
R16224 XThC.Tn[10] XThC.Tn[10].n72 13.9299
R16225 XThC.Tn[10] XThC.Tn[10].n6 8.0245
R16226 XThC.Tn[10].n66 XThC.Tn[10].n65 7.9105
R16227 XThC.Tn[10].n62 XThC.Tn[10].n61 7.9105
R16228 XThC.Tn[10].n58 XThC.Tn[10].n57 7.9105
R16229 XThC.Tn[10].n54 XThC.Tn[10].n53 7.9105
R16230 XThC.Tn[10].n50 XThC.Tn[10].n49 7.9105
R16231 XThC.Tn[10].n46 XThC.Tn[10].n45 7.9105
R16232 XThC.Tn[10].n42 XThC.Tn[10].n41 7.9105
R16233 XThC.Tn[10].n38 XThC.Tn[10].n37 7.9105
R16234 XThC.Tn[10].n34 XThC.Tn[10].n33 7.9105
R16235 XThC.Tn[10].n30 XThC.Tn[10].n29 7.9105
R16236 XThC.Tn[10].n26 XThC.Tn[10].n25 7.9105
R16237 XThC.Tn[10].n22 XThC.Tn[10].n21 7.9105
R16238 XThC.Tn[10].n18 XThC.Tn[10].n17 7.9105
R16239 XThC.Tn[10].n14 XThC.Tn[10].n13 7.9105
R16240 XThC.Tn[10].n10 XThC.Tn[10].n9 7.9105
R16241 XThC.Tn[10].n68 XThC.Tn[10].n67 7.40985
R16242 XThC.Tn[10].n67 XThC.Tn[10] 4.38575
R16243 XThC.Tn[10].n72 XThC.Tn[10].n68 2.99115
R16244 XThC.Tn[10].n72 XThC.Tn[10] 2.87153
R16245 XThC.Tn[10].n3 XThC.Tn[10] 2.688
R16246 XThC.Tn[10].n68 XThC.Tn[10] 2.2734
R16247 XThC.Tn[10].n67 XThC.Tn[10].n3 0.244922
R16248 XThC.Tn[10].n10 XThC.Tn[10] 0.235138
R16249 XThC.Tn[10].n14 XThC.Tn[10] 0.235138
R16250 XThC.Tn[10].n18 XThC.Tn[10] 0.235138
R16251 XThC.Tn[10].n22 XThC.Tn[10] 0.235138
R16252 XThC.Tn[10].n26 XThC.Tn[10] 0.235138
R16253 XThC.Tn[10].n30 XThC.Tn[10] 0.235138
R16254 XThC.Tn[10].n34 XThC.Tn[10] 0.235138
R16255 XThC.Tn[10].n38 XThC.Tn[10] 0.235138
R16256 XThC.Tn[10].n42 XThC.Tn[10] 0.235138
R16257 XThC.Tn[10].n46 XThC.Tn[10] 0.235138
R16258 XThC.Tn[10].n50 XThC.Tn[10] 0.235138
R16259 XThC.Tn[10].n54 XThC.Tn[10] 0.235138
R16260 XThC.Tn[10].n58 XThC.Tn[10] 0.235138
R16261 XThC.Tn[10].n62 XThC.Tn[10] 0.235138
R16262 XThC.Tn[10].n66 XThC.Tn[10] 0.235138
R16263 XThC.Tn[10].n3 XThC.Tn[10] 0.141947
R16264 XThC.Tn[10] XThC.Tn[10].n10 0.114505
R16265 XThC.Tn[10] XThC.Tn[10].n14 0.114505
R16266 XThC.Tn[10] XThC.Tn[10].n18 0.114505
R16267 XThC.Tn[10] XThC.Tn[10].n22 0.114505
R16268 XThC.Tn[10] XThC.Tn[10].n26 0.114505
R16269 XThC.Tn[10] XThC.Tn[10].n30 0.114505
R16270 XThC.Tn[10] XThC.Tn[10].n34 0.114505
R16271 XThC.Tn[10] XThC.Tn[10].n38 0.114505
R16272 XThC.Tn[10] XThC.Tn[10].n42 0.114505
R16273 XThC.Tn[10] XThC.Tn[10].n46 0.114505
R16274 XThC.Tn[10] XThC.Tn[10].n50 0.114505
R16275 XThC.Tn[10] XThC.Tn[10].n54 0.114505
R16276 XThC.Tn[10] XThC.Tn[10].n58 0.114505
R16277 XThC.Tn[10] XThC.Tn[10].n62 0.114505
R16278 XThC.Tn[10] XThC.Tn[10].n66 0.114505
R16279 XThC.Tn[10].n65 XThC.Tn[10].n64 0.0599512
R16280 XThC.Tn[10].n61 XThC.Tn[10].n60 0.0599512
R16281 XThC.Tn[10].n57 XThC.Tn[10].n56 0.0599512
R16282 XThC.Tn[10].n53 XThC.Tn[10].n52 0.0599512
R16283 XThC.Tn[10].n49 XThC.Tn[10].n48 0.0599512
R16284 XThC.Tn[10].n45 XThC.Tn[10].n44 0.0599512
R16285 XThC.Tn[10].n41 XThC.Tn[10].n40 0.0599512
R16286 XThC.Tn[10].n37 XThC.Tn[10].n36 0.0599512
R16287 XThC.Tn[10].n33 XThC.Tn[10].n32 0.0599512
R16288 XThC.Tn[10].n29 XThC.Tn[10].n28 0.0599512
R16289 XThC.Tn[10].n25 XThC.Tn[10].n24 0.0599512
R16290 XThC.Tn[10].n21 XThC.Tn[10].n20 0.0599512
R16291 XThC.Tn[10].n17 XThC.Tn[10].n16 0.0599512
R16292 XThC.Tn[10].n13 XThC.Tn[10].n12 0.0599512
R16293 XThC.Tn[10].n9 XThC.Tn[10].n8 0.0599512
R16294 XThC.Tn[10].n6 XThC.Tn[10].n5 0.0599512
R16295 XThC.Tn[10].n64 XThC.Tn[10] 0.0469286
R16296 XThC.Tn[10].n60 XThC.Tn[10] 0.0469286
R16297 XThC.Tn[10].n56 XThC.Tn[10] 0.0469286
R16298 XThC.Tn[10].n52 XThC.Tn[10] 0.0469286
R16299 XThC.Tn[10].n48 XThC.Tn[10] 0.0469286
R16300 XThC.Tn[10].n44 XThC.Tn[10] 0.0469286
R16301 XThC.Tn[10].n40 XThC.Tn[10] 0.0469286
R16302 XThC.Tn[10].n36 XThC.Tn[10] 0.0469286
R16303 XThC.Tn[10].n32 XThC.Tn[10] 0.0469286
R16304 XThC.Tn[10].n28 XThC.Tn[10] 0.0469286
R16305 XThC.Tn[10].n24 XThC.Tn[10] 0.0469286
R16306 XThC.Tn[10].n20 XThC.Tn[10] 0.0469286
R16307 XThC.Tn[10].n16 XThC.Tn[10] 0.0469286
R16308 XThC.Tn[10].n12 XThC.Tn[10] 0.0469286
R16309 XThC.Tn[10].n8 XThC.Tn[10] 0.0469286
R16310 XThC.Tn[10].n5 XThC.Tn[10] 0.0469286
R16311 XThC.Tn[10].n64 XThC.Tn[10] 0.0401341
R16312 XThC.Tn[10].n60 XThC.Tn[10] 0.0401341
R16313 XThC.Tn[10].n56 XThC.Tn[10] 0.0401341
R16314 XThC.Tn[10].n52 XThC.Tn[10] 0.0401341
R16315 XThC.Tn[10].n48 XThC.Tn[10] 0.0401341
R16316 XThC.Tn[10].n44 XThC.Tn[10] 0.0401341
R16317 XThC.Tn[10].n40 XThC.Tn[10] 0.0401341
R16318 XThC.Tn[10].n36 XThC.Tn[10] 0.0401341
R16319 XThC.Tn[10].n32 XThC.Tn[10] 0.0401341
R16320 XThC.Tn[10].n28 XThC.Tn[10] 0.0401341
R16321 XThC.Tn[10].n24 XThC.Tn[10] 0.0401341
R16322 XThC.Tn[10].n20 XThC.Tn[10] 0.0401341
R16323 XThC.Tn[10].n16 XThC.Tn[10] 0.0401341
R16324 XThC.Tn[10].n12 XThC.Tn[10] 0.0401341
R16325 XThC.Tn[10].n8 XThC.Tn[10] 0.0401341
R16326 XThC.Tn[10].n5 XThC.Tn[10] 0.0401341
R16327 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R16328 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R16329 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R16330 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R16331 XThR.Tn[14].n87 XThR.Tn[14].n85 202.094
R16332 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R16333 XThR.Tn[14] XThR.Tn[14].n78 161.363
R16334 XThR.Tn[14] XThR.Tn[14].n73 161.363
R16335 XThR.Tn[14] XThR.Tn[14].n68 161.363
R16336 XThR.Tn[14] XThR.Tn[14].n63 161.363
R16337 XThR.Tn[14] XThR.Tn[14].n58 161.363
R16338 XThR.Tn[14] XThR.Tn[14].n53 161.363
R16339 XThR.Tn[14] XThR.Tn[14].n48 161.363
R16340 XThR.Tn[14] XThR.Tn[14].n43 161.363
R16341 XThR.Tn[14] XThR.Tn[14].n38 161.363
R16342 XThR.Tn[14] XThR.Tn[14].n33 161.363
R16343 XThR.Tn[14] XThR.Tn[14].n28 161.363
R16344 XThR.Tn[14] XThR.Tn[14].n23 161.363
R16345 XThR.Tn[14] XThR.Tn[14].n18 161.363
R16346 XThR.Tn[14] XThR.Tn[14].n13 161.363
R16347 XThR.Tn[14] XThR.Tn[14].n8 161.363
R16348 XThR.Tn[14] XThR.Tn[14].n6 161.363
R16349 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R16350 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R16351 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R16352 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R16353 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R16354 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R16355 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R16356 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R16357 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R16358 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R16359 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R16360 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R16361 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R16362 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R16363 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R16364 XThR.Tn[14].n79 XThR.Tn[14].t14 161.106
R16365 XThR.Tn[14].n78 XThR.Tn[14].t30 161.106
R16366 XThR.Tn[14].n74 XThR.Tn[14].t21 161.106
R16367 XThR.Tn[14].n73 XThR.Tn[14].t40 161.106
R16368 XThR.Tn[14].n69 XThR.Tn[14].t64 161.106
R16369 XThR.Tn[14].n68 XThR.Tn[14].t22 161.106
R16370 XThR.Tn[14].n64 XThR.Tn[14].t46 161.106
R16371 XThR.Tn[14].n63 XThR.Tn[14].t65 161.106
R16372 XThR.Tn[14].n59 XThR.Tn[14].t12 161.106
R16373 XThR.Tn[14].n58 XThR.Tn[14].t28 161.106
R16374 XThR.Tn[14].n54 XThR.Tn[14].t37 161.106
R16375 XThR.Tn[14].n53 XThR.Tn[14].t56 161.106
R16376 XThR.Tn[14].n49 XThR.Tn[14].t16 161.106
R16377 XThR.Tn[14].n48 XThR.Tn[14].t36 161.106
R16378 XThR.Tn[14].n44 XThR.Tn[14].t60 161.106
R16379 XThR.Tn[14].n43 XThR.Tn[14].t17 161.106
R16380 XThR.Tn[14].n39 XThR.Tn[14].t45 161.106
R16381 XThR.Tn[14].n38 XThR.Tn[14].t61 161.106
R16382 XThR.Tn[14].n34 XThR.Tn[14].t51 161.106
R16383 XThR.Tn[14].n33 XThR.Tn[14].t68 161.106
R16384 XThR.Tn[14].n29 XThR.Tn[14].t35 161.106
R16385 XThR.Tn[14].n28 XThR.Tn[14].t53 161.106
R16386 XThR.Tn[14].n24 XThR.Tn[14].t63 161.106
R16387 XThR.Tn[14].n23 XThR.Tn[14].t20 161.106
R16388 XThR.Tn[14].n19 XThR.Tn[14].t32 161.106
R16389 XThR.Tn[14].n18 XThR.Tn[14].t49 161.106
R16390 XThR.Tn[14].n14 XThR.Tn[14].t15 161.106
R16391 XThR.Tn[14].n13 XThR.Tn[14].t33 161.106
R16392 XThR.Tn[14].n9 XThR.Tn[14].t42 161.106
R16393 XThR.Tn[14].n8 XThR.Tn[14].t59 161.106
R16394 XThR.Tn[14].n6 XThR.Tn[14].t43 161.106
R16395 XThR.Tn[14].n79 XThR.Tn[14].t31 154.679
R16396 XThR.Tn[14].n78 XThR.Tn[14].t48 154.679
R16397 XThR.Tn[14].n74 XThR.Tn[14].t71 154.679
R16398 XThR.Tn[14].n73 XThR.Tn[14].t27 154.679
R16399 XThR.Tn[14].n69 XThR.Tn[14].t55 154.679
R16400 XThR.Tn[14].n68 XThR.Tn[14].t72 154.679
R16401 XThR.Tn[14].n64 XThR.Tn[14].t23 154.679
R16402 XThR.Tn[14].n63 XThR.Tn[14].t41 154.679
R16403 XThR.Tn[14].n59 XThR.Tn[14].t66 154.679
R16404 XThR.Tn[14].n58 XThR.Tn[14].t24 154.679
R16405 XThR.Tn[14].n54 XThR.Tn[14].t29 154.679
R16406 XThR.Tn[14].n53 XThR.Tn[14].t47 154.679
R16407 XThR.Tn[14].n49 XThR.Tn[14].t57 154.679
R16408 XThR.Tn[14].n48 XThR.Tn[14].t73 154.679
R16409 XThR.Tn[14].n44 XThR.Tn[14].t39 154.679
R16410 XThR.Tn[14].n43 XThR.Tn[14].t58 154.679
R16411 XThR.Tn[14].n39 XThR.Tn[14].t18 154.679
R16412 XThR.Tn[14].n38 XThR.Tn[14].t38 154.679
R16413 XThR.Tn[14].n34 XThR.Tn[14].t62 154.679
R16414 XThR.Tn[14].n33 XThR.Tn[14].t19 154.679
R16415 XThR.Tn[14].n29 XThR.Tn[14].t69 154.679
R16416 XThR.Tn[14].n28 XThR.Tn[14].t26 154.679
R16417 XThR.Tn[14].n24 XThR.Tn[14].t54 154.679
R16418 XThR.Tn[14].n23 XThR.Tn[14].t70 154.679
R16419 XThR.Tn[14].n19 XThR.Tn[14].t25 154.679
R16420 XThR.Tn[14].n18 XThR.Tn[14].t44 154.679
R16421 XThR.Tn[14].n14 XThR.Tn[14].t50 154.679
R16422 XThR.Tn[14].n13 XThR.Tn[14].t67 154.679
R16423 XThR.Tn[14].n9 XThR.Tn[14].t34 154.679
R16424 XThR.Tn[14].n8 XThR.Tn[14].t52 154.679
R16425 XThR.Tn[14].n6 XThR.Tn[14].t13 154.679
R16426 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R16427 XThR.Tn[14].n86 XThR.Tn[14].t0 26.5955
R16428 XThR.Tn[14].n86 XThR.Tn[14].t1 26.5955
R16429 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R16430 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R16431 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R16432 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R16433 XThR.Tn[14].n85 XThR.Tn[14].t2 26.5955
R16434 XThR.Tn[14].n85 XThR.Tn[14].t3 26.5955
R16435 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R16436 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R16437 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R16438 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R16439 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R16440 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R16441 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R16442 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R16443 XThR.Tn[14] XThR.Tn[14].n7 5.34871
R16444 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R16445 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R16446 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R16447 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R16448 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R16449 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R16450 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R16451 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R16452 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R16453 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R16454 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R16455 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R16456 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R16457 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R16458 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R16459 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R16460 XThR.Tn[14].n12 XThR.Tn[14] 2.51836
R16461 XThR.Tn[14].n17 XThR.Tn[14] 2.51836
R16462 XThR.Tn[14].n22 XThR.Tn[14] 2.51836
R16463 XThR.Tn[14].n27 XThR.Tn[14] 2.51836
R16464 XThR.Tn[14].n32 XThR.Tn[14] 2.51836
R16465 XThR.Tn[14].n37 XThR.Tn[14] 2.51836
R16466 XThR.Tn[14].n42 XThR.Tn[14] 2.51836
R16467 XThR.Tn[14].n47 XThR.Tn[14] 2.51836
R16468 XThR.Tn[14].n52 XThR.Tn[14] 2.51836
R16469 XThR.Tn[14].n57 XThR.Tn[14] 2.51836
R16470 XThR.Tn[14].n62 XThR.Tn[14] 2.51836
R16471 XThR.Tn[14].n67 XThR.Tn[14] 2.51836
R16472 XThR.Tn[14].n72 XThR.Tn[14] 2.51836
R16473 XThR.Tn[14].n77 XThR.Tn[14] 2.51836
R16474 XThR.Tn[14].n82 XThR.Tn[14] 2.51836
R16475 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R16476 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R16477 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R16478 XThR.Tn[14] XThR.Tn[14].n12 0.848714
R16479 XThR.Tn[14] XThR.Tn[14].n17 0.848714
R16480 XThR.Tn[14] XThR.Tn[14].n22 0.848714
R16481 XThR.Tn[14] XThR.Tn[14].n27 0.848714
R16482 XThR.Tn[14] XThR.Tn[14].n32 0.848714
R16483 XThR.Tn[14] XThR.Tn[14].n37 0.848714
R16484 XThR.Tn[14] XThR.Tn[14].n42 0.848714
R16485 XThR.Tn[14] XThR.Tn[14].n47 0.848714
R16486 XThR.Tn[14] XThR.Tn[14].n52 0.848714
R16487 XThR.Tn[14] XThR.Tn[14].n57 0.848714
R16488 XThR.Tn[14] XThR.Tn[14].n62 0.848714
R16489 XThR.Tn[14] XThR.Tn[14].n67 0.848714
R16490 XThR.Tn[14] XThR.Tn[14].n72 0.848714
R16491 XThR.Tn[14] XThR.Tn[14].n77 0.848714
R16492 XThR.Tn[14] XThR.Tn[14].n82 0.848714
R16493 XThR.Tn[14].n7 XThR.Tn[14] 0.485653
R16494 XThR.Tn[14].n80 XThR.Tn[14] 0.21482
R16495 XThR.Tn[14].n75 XThR.Tn[14] 0.21482
R16496 XThR.Tn[14].n70 XThR.Tn[14] 0.21482
R16497 XThR.Tn[14].n65 XThR.Tn[14] 0.21482
R16498 XThR.Tn[14].n60 XThR.Tn[14] 0.21482
R16499 XThR.Tn[14].n55 XThR.Tn[14] 0.21482
R16500 XThR.Tn[14].n50 XThR.Tn[14] 0.21482
R16501 XThR.Tn[14].n45 XThR.Tn[14] 0.21482
R16502 XThR.Tn[14].n40 XThR.Tn[14] 0.21482
R16503 XThR.Tn[14].n35 XThR.Tn[14] 0.21482
R16504 XThR.Tn[14].n30 XThR.Tn[14] 0.21482
R16505 XThR.Tn[14].n25 XThR.Tn[14] 0.21482
R16506 XThR.Tn[14].n20 XThR.Tn[14] 0.21482
R16507 XThR.Tn[14].n15 XThR.Tn[14] 0.21482
R16508 XThR.Tn[14].n10 XThR.Tn[14] 0.21482
R16509 XThR.Tn[14].n81 XThR.Tn[14] 0.0608448
R16510 XThR.Tn[14].n76 XThR.Tn[14] 0.0608448
R16511 XThR.Tn[14].n71 XThR.Tn[14] 0.0608448
R16512 XThR.Tn[14].n66 XThR.Tn[14] 0.0608448
R16513 XThR.Tn[14].n61 XThR.Tn[14] 0.0608448
R16514 XThR.Tn[14].n56 XThR.Tn[14] 0.0608448
R16515 XThR.Tn[14].n51 XThR.Tn[14] 0.0608448
R16516 XThR.Tn[14].n46 XThR.Tn[14] 0.0608448
R16517 XThR.Tn[14].n41 XThR.Tn[14] 0.0608448
R16518 XThR.Tn[14].n36 XThR.Tn[14] 0.0608448
R16519 XThR.Tn[14].n31 XThR.Tn[14] 0.0608448
R16520 XThR.Tn[14].n26 XThR.Tn[14] 0.0608448
R16521 XThR.Tn[14].n21 XThR.Tn[14] 0.0608448
R16522 XThR.Tn[14].n16 XThR.Tn[14] 0.0608448
R16523 XThR.Tn[14].n11 XThR.Tn[14] 0.0608448
R16524 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R16525 XThR.Tn[14] XThR.Tn[14].n83 0.038
R16526 XThR.Tn[14].n7 XThR.Tn[14] 0.00744444
R16527 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00265517
R16528 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00265517
R16529 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00265517
R16530 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00265517
R16531 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00265517
R16532 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00265517
R16533 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00265517
R16534 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00265517
R16535 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00265517
R16536 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00265517
R16537 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00265517
R16538 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00265517
R16539 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00265517
R16540 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00265517
R16541 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00265517
R16542 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R16543 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R16544 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R16545 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R16546 XThR.Tn[8].n87 XThR.Tn[8].n85 202.094
R16547 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R16548 XThR.Tn[8] XThR.Tn[8].n78 161.363
R16549 XThR.Tn[8] XThR.Tn[8].n73 161.363
R16550 XThR.Tn[8] XThR.Tn[8].n68 161.363
R16551 XThR.Tn[8] XThR.Tn[8].n63 161.363
R16552 XThR.Tn[8] XThR.Tn[8].n58 161.363
R16553 XThR.Tn[8] XThR.Tn[8].n53 161.363
R16554 XThR.Tn[8] XThR.Tn[8].n48 161.363
R16555 XThR.Tn[8] XThR.Tn[8].n43 161.363
R16556 XThR.Tn[8] XThR.Tn[8].n38 161.363
R16557 XThR.Tn[8] XThR.Tn[8].n33 161.363
R16558 XThR.Tn[8] XThR.Tn[8].n28 161.363
R16559 XThR.Tn[8] XThR.Tn[8].n23 161.363
R16560 XThR.Tn[8] XThR.Tn[8].n18 161.363
R16561 XThR.Tn[8] XThR.Tn[8].n13 161.363
R16562 XThR.Tn[8] XThR.Tn[8].n8 161.363
R16563 XThR.Tn[8] XThR.Tn[8].n6 161.363
R16564 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R16565 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R16566 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R16567 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R16568 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R16569 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R16570 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R16571 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R16572 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R16573 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R16574 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R16575 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R16576 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R16577 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R16578 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R16579 XThR.Tn[8].n79 XThR.Tn[8].t60 161.106
R16580 XThR.Tn[8].n78 XThR.Tn[8].t19 161.106
R16581 XThR.Tn[8].n74 XThR.Tn[8].t66 161.106
R16582 XThR.Tn[8].n73 XThR.Tn[8].t27 161.106
R16583 XThR.Tn[8].n69 XThR.Tn[8].t49 161.106
R16584 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R16585 XThR.Tn[8].n64 XThR.Tn[8].t32 161.106
R16586 XThR.Tn[8].n63 XThR.Tn[8].t52 161.106
R16587 XThR.Tn[8].n59 XThR.Tn[8].t58 161.106
R16588 XThR.Tn[8].n58 XThR.Tn[8].t16 161.106
R16589 XThR.Tn[8].n54 XThR.Tn[8].t21 161.106
R16590 XThR.Tn[8].n53 XThR.Tn[8].t43 161.106
R16591 XThR.Tn[8].n49 XThR.Tn[8].t64 161.106
R16592 XThR.Tn[8].n48 XThR.Tn[8].t24 161.106
R16593 XThR.Tn[8].n44 XThR.Tn[8].t46 161.106
R16594 XThR.Tn[8].n43 XThR.Tn[8].t68 161.106
R16595 XThR.Tn[8].n39 XThR.Tn[8].t30 161.106
R16596 XThR.Tn[8].n38 XThR.Tn[8].t51 161.106
R16597 XThR.Tn[8].n34 XThR.Tn[8].t35 161.106
R16598 XThR.Tn[8].n33 XThR.Tn[8].t56 161.106
R16599 XThR.Tn[8].n29 XThR.Tn[8].t20 161.106
R16600 XThR.Tn[8].n28 XThR.Tn[8].t42 161.106
R16601 XThR.Tn[8].n24 XThR.Tn[8].t48 161.106
R16602 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R16603 XThR.Tn[8].n19 XThR.Tn[8].t17 161.106
R16604 XThR.Tn[8].n18 XThR.Tn[8].t40 161.106
R16605 XThR.Tn[8].n14 XThR.Tn[8].t62 161.106
R16606 XThR.Tn[8].n13 XThR.Tn[8].t23 161.106
R16607 XThR.Tn[8].n9 XThR.Tn[8].t25 161.106
R16608 XThR.Tn[8].n8 XThR.Tn[8].t45 161.106
R16609 XThR.Tn[8].n6 XThR.Tn[8].t29 161.106
R16610 XThR.Tn[8].n79 XThR.Tn[8].t15 154.679
R16611 XThR.Tn[8].n78 XThR.Tn[8].t37 154.679
R16612 XThR.Tn[8].n74 XThR.Tn[8].t54 154.679
R16613 XThR.Tn[8].n73 XThR.Tn[8].t13 154.679
R16614 XThR.Tn[8].n69 XThR.Tn[8].t38 154.679
R16615 XThR.Tn[8].n68 XThR.Tn[8].t59 154.679
R16616 XThR.Tn[8].n64 XThR.Tn[8].t67 154.679
R16617 XThR.Tn[8].n63 XThR.Tn[8].t28 154.679
R16618 XThR.Tn[8].n59 XThR.Tn[8].t50 154.679
R16619 XThR.Tn[8].n58 XThR.Tn[8].t72 154.679
R16620 XThR.Tn[8].n54 XThR.Tn[8].t14 154.679
R16621 XThR.Tn[8].n53 XThR.Tn[8].t33 154.679
R16622 XThR.Tn[8].n49 XThR.Tn[8].t39 154.679
R16623 XThR.Tn[8].n48 XThR.Tn[8].t61 154.679
R16624 XThR.Tn[8].n44 XThR.Tn[8].t22 154.679
R16625 XThR.Tn[8].n43 XThR.Tn[8].t44 154.679
R16626 XThR.Tn[8].n39 XThR.Tn[8].t65 154.679
R16627 XThR.Tn[8].n38 XThR.Tn[8].t26 154.679
R16628 XThR.Tn[8].n34 XThR.Tn[8].t47 154.679
R16629 XThR.Tn[8].n33 XThR.Tn[8].t69 154.679
R16630 XThR.Tn[8].n29 XThR.Tn[8].t53 154.679
R16631 XThR.Tn[8].n28 XThR.Tn[8].t12 154.679
R16632 XThR.Tn[8].n24 XThR.Tn[8].t36 154.679
R16633 XThR.Tn[8].n23 XThR.Tn[8].t57 154.679
R16634 XThR.Tn[8].n19 XThR.Tn[8].t73 154.679
R16635 XThR.Tn[8].n18 XThR.Tn[8].t31 154.679
R16636 XThR.Tn[8].n14 XThR.Tn[8].t34 154.679
R16637 XThR.Tn[8].n13 XThR.Tn[8].t55 154.679
R16638 XThR.Tn[8].n9 XThR.Tn[8].t18 154.679
R16639 XThR.Tn[8].n8 XThR.Tn[8].t41 154.679
R16640 XThR.Tn[8].n6 XThR.Tn[8].t63 154.679
R16641 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R16642 XThR.Tn[8].n86 XThR.Tn[8].t7 26.5955
R16643 XThR.Tn[8].n86 XThR.Tn[8].t1 26.5955
R16644 XThR.Tn[8].n0 XThR.Tn[8].t10 26.5955
R16645 XThR.Tn[8].n0 XThR.Tn[8].t8 26.5955
R16646 XThR.Tn[8].n1 XThR.Tn[8].t11 26.5955
R16647 XThR.Tn[8].n1 XThR.Tn[8].t9 26.5955
R16648 XThR.Tn[8].n85 XThR.Tn[8].t0 26.5955
R16649 XThR.Tn[8].n85 XThR.Tn[8].t2 26.5955
R16650 XThR.Tn[8].n4 XThR.Tn[8].t4 24.9236
R16651 XThR.Tn[8].n4 XThR.Tn[8].t6 24.9236
R16652 XThR.Tn[8].n3 XThR.Tn[8].t3 24.9236
R16653 XThR.Tn[8].n3 XThR.Tn[8].t5 24.9236
R16654 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R16655 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R16656 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R16657 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R16658 XThR.Tn[8] XThR.Tn[8].n7 5.34871
R16659 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R16660 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R16661 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R16662 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R16663 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R16664 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R16665 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R16666 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R16667 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R16668 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R16669 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R16670 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R16671 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R16672 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R16673 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R16674 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R16675 XThR.Tn[8].n12 XThR.Tn[8] 2.51836
R16676 XThR.Tn[8].n17 XThR.Tn[8] 2.51836
R16677 XThR.Tn[8].n22 XThR.Tn[8] 2.51836
R16678 XThR.Tn[8].n27 XThR.Tn[8] 2.51836
R16679 XThR.Tn[8].n32 XThR.Tn[8] 2.51836
R16680 XThR.Tn[8].n37 XThR.Tn[8] 2.51836
R16681 XThR.Tn[8].n42 XThR.Tn[8] 2.51836
R16682 XThR.Tn[8].n47 XThR.Tn[8] 2.51836
R16683 XThR.Tn[8].n52 XThR.Tn[8] 2.51836
R16684 XThR.Tn[8].n57 XThR.Tn[8] 2.51836
R16685 XThR.Tn[8].n62 XThR.Tn[8] 2.51836
R16686 XThR.Tn[8].n67 XThR.Tn[8] 2.51836
R16687 XThR.Tn[8].n72 XThR.Tn[8] 2.51836
R16688 XThR.Tn[8].n77 XThR.Tn[8] 2.51836
R16689 XThR.Tn[8].n82 XThR.Tn[8] 2.51836
R16690 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R16691 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R16692 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R16693 XThR.Tn[8] XThR.Tn[8].n12 0.848714
R16694 XThR.Tn[8] XThR.Tn[8].n17 0.848714
R16695 XThR.Tn[8] XThR.Tn[8].n22 0.848714
R16696 XThR.Tn[8] XThR.Tn[8].n27 0.848714
R16697 XThR.Tn[8] XThR.Tn[8].n32 0.848714
R16698 XThR.Tn[8] XThR.Tn[8].n37 0.848714
R16699 XThR.Tn[8] XThR.Tn[8].n42 0.848714
R16700 XThR.Tn[8] XThR.Tn[8].n47 0.848714
R16701 XThR.Tn[8] XThR.Tn[8].n52 0.848714
R16702 XThR.Tn[8] XThR.Tn[8].n57 0.848714
R16703 XThR.Tn[8] XThR.Tn[8].n62 0.848714
R16704 XThR.Tn[8] XThR.Tn[8].n67 0.848714
R16705 XThR.Tn[8] XThR.Tn[8].n72 0.848714
R16706 XThR.Tn[8] XThR.Tn[8].n77 0.848714
R16707 XThR.Tn[8] XThR.Tn[8].n82 0.848714
R16708 XThR.Tn[8].n7 XThR.Tn[8] 0.485653
R16709 XThR.Tn[8].n80 XThR.Tn[8] 0.21482
R16710 XThR.Tn[8].n75 XThR.Tn[8] 0.21482
R16711 XThR.Tn[8].n70 XThR.Tn[8] 0.21482
R16712 XThR.Tn[8].n65 XThR.Tn[8] 0.21482
R16713 XThR.Tn[8].n60 XThR.Tn[8] 0.21482
R16714 XThR.Tn[8].n55 XThR.Tn[8] 0.21482
R16715 XThR.Tn[8].n50 XThR.Tn[8] 0.21482
R16716 XThR.Tn[8].n45 XThR.Tn[8] 0.21482
R16717 XThR.Tn[8].n40 XThR.Tn[8] 0.21482
R16718 XThR.Tn[8].n35 XThR.Tn[8] 0.21482
R16719 XThR.Tn[8].n30 XThR.Tn[8] 0.21482
R16720 XThR.Tn[8].n25 XThR.Tn[8] 0.21482
R16721 XThR.Tn[8].n20 XThR.Tn[8] 0.21482
R16722 XThR.Tn[8].n15 XThR.Tn[8] 0.21482
R16723 XThR.Tn[8].n10 XThR.Tn[8] 0.21482
R16724 XThR.Tn[8].n81 XThR.Tn[8] 0.0608448
R16725 XThR.Tn[8].n76 XThR.Tn[8] 0.0608448
R16726 XThR.Tn[8].n71 XThR.Tn[8] 0.0608448
R16727 XThR.Tn[8].n66 XThR.Tn[8] 0.0608448
R16728 XThR.Tn[8].n61 XThR.Tn[8] 0.0608448
R16729 XThR.Tn[8].n56 XThR.Tn[8] 0.0608448
R16730 XThR.Tn[8].n51 XThR.Tn[8] 0.0608448
R16731 XThR.Tn[8].n46 XThR.Tn[8] 0.0608448
R16732 XThR.Tn[8].n41 XThR.Tn[8] 0.0608448
R16733 XThR.Tn[8].n36 XThR.Tn[8] 0.0608448
R16734 XThR.Tn[8].n31 XThR.Tn[8] 0.0608448
R16735 XThR.Tn[8].n26 XThR.Tn[8] 0.0608448
R16736 XThR.Tn[8].n21 XThR.Tn[8] 0.0608448
R16737 XThR.Tn[8].n16 XThR.Tn[8] 0.0608448
R16738 XThR.Tn[8].n11 XThR.Tn[8] 0.0608448
R16739 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R16740 XThR.Tn[8] XThR.Tn[8].n83 0.038
R16741 XThR.Tn[8].n7 XThR.Tn[8] 0.00744444
R16742 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00265517
R16743 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00265517
R16744 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00265517
R16745 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00265517
R16746 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00265517
R16747 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00265517
R16748 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00265517
R16749 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00265517
R16750 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00265517
R16751 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00265517
R16752 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00265517
R16753 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00265517
R16754 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00265517
R16755 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00265517
R16756 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00265517
R16757 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R16758 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R16759 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R16760 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R16761 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R16762 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R16763 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R16764 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R16765 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R16766 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R16767 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R16768 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R16769 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R16770 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R16771 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R16772 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R16773 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R16774 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R16775 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R16776 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R16777 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R16778 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R16779 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R16780 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R16781 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R16782 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R16783 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R16784 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R16785 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R16786 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R16787 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R16788 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R16789 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R16790 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R16791 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R16792 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R16793 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R16794 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R16795 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R16796 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R16797 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R16798 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R16799 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R16800 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R16801 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R16802 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R16803 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R16804 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R16805 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R16806 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R16807 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R16808 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R16809 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R16810 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R16811 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R16812 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R16813 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R16814 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R16815 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R16816 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R16817 XThC.XTBN.Y.n192 XThC.XTBN.Y.n191 208.964
R16818 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R16819 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R16820 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R16821 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R16822 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R16823 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R16824 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R16825 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R16826 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R16827 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R16828 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R16829 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R16830 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R16831 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R16832 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R16833 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R16834 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R16835 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R16836 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R16837 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R16838 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R16839 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R16840 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R16841 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R16842 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R16843 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R16844 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R16845 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R16846 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R16847 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R16848 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R16849 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R16850 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R16851 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R16852 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R16853 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R16854 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R16855 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R16856 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R16857 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R16858 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R16859 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R16860 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R16861 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R16862 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R16863 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R16864 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R16865 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R16866 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R16867 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R16868 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R16869 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R16870 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R16871 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R16872 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R16873 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R16874 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R16875 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R16876 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R16877 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R16878 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R16879 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R16880 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R16881 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R16882 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R16883 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R16884 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R16885 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R16886 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R16887 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R16888 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R16889 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R16890 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R16891 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R16892 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R16893 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R16894 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R16895 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R16896 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R16897 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R16898 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R16899 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R16900 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R16901 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R16902 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R16903 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R16904 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R16905 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R16906 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R16907 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R16908 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R16909 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R16910 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R16911 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R16912 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R16913 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R16914 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R16915 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R16916 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R16917 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R16918 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R16919 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R16920 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R16921 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R16922 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R16923 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R16924 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R16925 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R16926 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R16927 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R16928 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R16929 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R16930 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R16931 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R16932 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R16933 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R16934 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R16935 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R16936 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R16937 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R16938 XThC.XTBN.Y XThC.XTBN.Y.n188 96.8352
R16939 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R16940 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R16941 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R16942 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R16943 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R16944 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R16945 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R16946 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R16947 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R16948 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R16949 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R16950 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R16951 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R16952 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R16953 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R16954 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R16955 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R16956 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R16957 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R16958 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R16959 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R16960 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R16961 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R16962 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R16963 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R16964 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R16965 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R16966 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R16967 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R16968 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R16969 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R16970 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R16971 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R16972 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R16973 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R16974 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R16975 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R16976 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R16977 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R16978 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R16979 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R16980 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R16981 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R16982 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R16983 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R16984 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R16985 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R16986 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R16987 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R16988 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R16989 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R16990 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R16991 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R16992 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R16993 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R16994 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R16995 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R16996 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R16997 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R16998 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R16999 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R17000 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R17001 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R17002 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R17003 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R17004 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R17005 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R17006 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R17007 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R17008 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R17009 XThC.XTBN.Y.n191 XThC.XTBN.Y.t0 26.5955
R17010 XThC.XTBN.Y.n191 XThC.XTBN.Y.t1 26.5955
R17011 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 24.9236
R17012 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 24.9236
R17013 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R17014 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R17015 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R17016 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R17017 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R17018 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R17019 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R17020 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R17021 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R17022 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R17023 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R17024 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R17025 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R17026 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R17027 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R17028 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R17029 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R17030 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R17031 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R17032 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R17033 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R17034 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R17035 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R17036 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R17037 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R17038 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R17039 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R17040 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R17041 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R17042 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R17043 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R17044 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R17045 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R17046 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R17047 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R17048 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R17049 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R17050 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R17051 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R17052 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R17053 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R17054 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R17055 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R17056 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R17057 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R17058 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R17059 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R17060 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R17061 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R17062 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R17063 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R17064 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R17065 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R17066 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R17067 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R17068 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R17069 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R17070 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R17071 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R17072 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R17073 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R17074 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R17075 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R17076 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R17077 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R17078 XThC.XTBN.Y XThC.XTBN.Y.n190 12.5445
R17079 XThC.XTBN.Y XThC.XTBN.Y.n189 11.2645
R17080 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R17081 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R17082 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R17083 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R17084 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R17085 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R17086 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R17087 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R17088 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R17089 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R17090 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R17091 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R17092 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R17093 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R17094 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R17095 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R17096 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R17097 XThC.XTBN.Y.n189 XThC.XTBN.Y 6.1445
R17098 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R17099 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R17100 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R17101 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R17102 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R17103 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R17104 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R17105 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R17106 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R17107 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R17108 XThC.XTBN.Y.n190 XThC.XTBN.Y 4.8645
R17109 XThC.XTBN.Y.n189 XThC.XTBN.Y 4.65505
R17110 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R17111 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R17112 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R17113 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R17114 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R17115 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R17116 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R17117 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R17118 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R17119 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R17120 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R17121 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R17122 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R17123 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R17124 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R17125 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R17126 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R17127 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R17128 XThC.XTBN.Y.n192 XThC.XTBN.Y 2.0485
R17129 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R17130 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R17131 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R17132 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R17133 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R17134 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R17135 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R17136 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R17137 XThC.XTBN.Y XThC.XTBN.Y.n192 1.55202
R17138 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R17139 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R17140 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R17141 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R17142 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R17143 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R17144 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R17145 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R17146 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R17147 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R17148 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R17149 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R17150 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R17151 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R17152 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R17153 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R17154 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R17155 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R17156 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R17157 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R17158 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R17159 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R17160 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R17161 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R17162 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R17163 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R17164 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R17165 XThC.Tn[6].n71 XThC.Tn[6].n69 161.365
R17166 XThC.Tn[6].n67 XThC.Tn[6].n65 161.365
R17167 XThC.Tn[6].n63 XThC.Tn[6].n61 161.365
R17168 XThC.Tn[6].n59 XThC.Tn[6].n57 161.365
R17169 XThC.Tn[6].n55 XThC.Tn[6].n53 161.365
R17170 XThC.Tn[6].n51 XThC.Tn[6].n49 161.365
R17171 XThC.Tn[6].n47 XThC.Tn[6].n45 161.365
R17172 XThC.Tn[6].n43 XThC.Tn[6].n41 161.365
R17173 XThC.Tn[6].n39 XThC.Tn[6].n37 161.365
R17174 XThC.Tn[6].n35 XThC.Tn[6].n33 161.365
R17175 XThC.Tn[6].n31 XThC.Tn[6].n29 161.365
R17176 XThC.Tn[6].n27 XThC.Tn[6].n25 161.365
R17177 XThC.Tn[6].n23 XThC.Tn[6].n21 161.365
R17178 XThC.Tn[6].n19 XThC.Tn[6].n17 161.365
R17179 XThC.Tn[6].n15 XThC.Tn[6].n13 161.365
R17180 XThC.Tn[6].n12 XThC.Tn[6].n10 161.365
R17181 XThC.Tn[6].n69 XThC.Tn[6].t21 161.106
R17182 XThC.Tn[6].n65 XThC.Tn[6].t33 161.106
R17183 XThC.Tn[6].n61 XThC.Tn[6].t31 161.106
R17184 XThC.Tn[6].n57 XThC.Tn[6].t29 161.106
R17185 XThC.Tn[6].n53 XThC.Tn[6].t43 161.106
R17186 XThC.Tn[6].n49 XThC.Tn[6].t40 161.106
R17187 XThC.Tn[6].n45 XThC.Tn[6].t28 161.106
R17188 XThC.Tn[6].n41 XThC.Tn[6].t19 161.106
R17189 XThC.Tn[6].n37 XThC.Tn[6].t17 161.106
R17190 XThC.Tn[6].n33 XThC.Tn[6].t38 161.106
R17191 XThC.Tn[6].n29 XThC.Tn[6].t27 161.106
R17192 XThC.Tn[6].n25 XThC.Tn[6].t16 161.106
R17193 XThC.Tn[6].n21 XThC.Tn[6].t37 161.106
R17194 XThC.Tn[6].n17 XThC.Tn[6].t36 161.106
R17195 XThC.Tn[6].n13 XThC.Tn[6].t23 161.106
R17196 XThC.Tn[6].n10 XThC.Tn[6].t13 161.106
R17197 XThC.Tn[6].n69 XThC.Tn[6].t41 154.679
R17198 XThC.Tn[6].n65 XThC.Tn[6].t20 154.679
R17199 XThC.Tn[6].n61 XThC.Tn[6].t18 154.679
R17200 XThC.Tn[6].n57 XThC.Tn[6].t15 154.679
R17201 XThC.Tn[6].n53 XThC.Tn[6].t30 154.679
R17202 XThC.Tn[6].n49 XThC.Tn[6].t26 154.679
R17203 XThC.Tn[6].n45 XThC.Tn[6].t14 154.679
R17204 XThC.Tn[6].n41 XThC.Tn[6].t39 154.679
R17205 XThC.Tn[6].n37 XThC.Tn[6].t35 154.679
R17206 XThC.Tn[6].n33 XThC.Tn[6].t25 154.679
R17207 XThC.Tn[6].n29 XThC.Tn[6].t12 154.679
R17208 XThC.Tn[6].n25 XThC.Tn[6].t34 154.679
R17209 XThC.Tn[6].n21 XThC.Tn[6].t24 154.679
R17210 XThC.Tn[6].n17 XThC.Tn[6].t22 154.679
R17211 XThC.Tn[6].n13 XThC.Tn[6].t42 154.679
R17212 XThC.Tn[6].n10 XThC.Tn[6].t32 154.679
R17213 XThC.Tn[6].n7 XThC.Tn[6].n6 135.248
R17214 XThC.Tn[6].n9 XThC.Tn[6].n3 98.982
R17215 XThC.Tn[6].n8 XThC.Tn[6].n4 98.982
R17216 XThC.Tn[6].n7 XThC.Tn[6].n5 98.982
R17217 XThC.Tn[6].n9 XThC.Tn[6].n8 36.2672
R17218 XThC.Tn[6].n8 XThC.Tn[6].n7 36.2672
R17219 XThC.Tn[6].n73 XThC.Tn[6].n9 32.6405
R17220 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R17221 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R17222 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R17223 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R17224 XThC.Tn[6].n3 XThC.Tn[6].t8 24.9236
R17225 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R17226 XThC.Tn[6].n4 XThC.Tn[6].t10 24.9236
R17227 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R17228 XThC.Tn[6].n5 XThC.Tn[6].t1 24.9236
R17229 XThC.Tn[6].n5 XThC.Tn[6].t0 24.9236
R17230 XThC.Tn[6].n6 XThC.Tn[6].t3 24.9236
R17231 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R17232 XThC.Tn[6].n74 XThC.Tn[6].n2 18.5605
R17233 XThC.Tn[6].n74 XThC.Tn[6].n73 11.5205
R17234 XThC.Tn[6] XThC.Tn[6].n12 8.0245
R17235 XThC.Tn[6].n72 XThC.Tn[6].n71 7.9105
R17236 XThC.Tn[6].n68 XThC.Tn[6].n67 7.9105
R17237 XThC.Tn[6].n64 XThC.Tn[6].n63 7.9105
R17238 XThC.Tn[6].n60 XThC.Tn[6].n59 7.9105
R17239 XThC.Tn[6].n56 XThC.Tn[6].n55 7.9105
R17240 XThC.Tn[6].n52 XThC.Tn[6].n51 7.9105
R17241 XThC.Tn[6].n48 XThC.Tn[6].n47 7.9105
R17242 XThC.Tn[6].n44 XThC.Tn[6].n43 7.9105
R17243 XThC.Tn[6].n40 XThC.Tn[6].n39 7.9105
R17244 XThC.Tn[6].n36 XThC.Tn[6].n35 7.9105
R17245 XThC.Tn[6].n32 XThC.Tn[6].n31 7.9105
R17246 XThC.Tn[6].n28 XThC.Tn[6].n27 7.9105
R17247 XThC.Tn[6].n24 XThC.Tn[6].n23 7.9105
R17248 XThC.Tn[6].n20 XThC.Tn[6].n19 7.9105
R17249 XThC.Tn[6].n16 XThC.Tn[6].n15 7.9105
R17250 XThC.Tn[6].n73 XThC.Tn[6] 5.42203
R17251 XThC.Tn[6] XThC.Tn[6].n74 0.6405
R17252 XThC.Tn[6].n16 XThC.Tn[6] 0.235138
R17253 XThC.Tn[6].n20 XThC.Tn[6] 0.235138
R17254 XThC.Tn[6].n24 XThC.Tn[6] 0.235138
R17255 XThC.Tn[6].n28 XThC.Tn[6] 0.235138
R17256 XThC.Tn[6].n32 XThC.Tn[6] 0.235138
R17257 XThC.Tn[6].n36 XThC.Tn[6] 0.235138
R17258 XThC.Tn[6].n40 XThC.Tn[6] 0.235138
R17259 XThC.Tn[6].n44 XThC.Tn[6] 0.235138
R17260 XThC.Tn[6].n48 XThC.Tn[6] 0.235138
R17261 XThC.Tn[6].n52 XThC.Tn[6] 0.235138
R17262 XThC.Tn[6].n56 XThC.Tn[6] 0.235138
R17263 XThC.Tn[6].n60 XThC.Tn[6] 0.235138
R17264 XThC.Tn[6].n64 XThC.Tn[6] 0.235138
R17265 XThC.Tn[6].n68 XThC.Tn[6] 0.235138
R17266 XThC.Tn[6].n72 XThC.Tn[6] 0.235138
R17267 XThC.Tn[6] XThC.Tn[6].n16 0.114505
R17268 XThC.Tn[6] XThC.Tn[6].n20 0.114505
R17269 XThC.Tn[6] XThC.Tn[6].n24 0.114505
R17270 XThC.Tn[6] XThC.Tn[6].n28 0.114505
R17271 XThC.Tn[6] XThC.Tn[6].n32 0.114505
R17272 XThC.Tn[6] XThC.Tn[6].n36 0.114505
R17273 XThC.Tn[6] XThC.Tn[6].n40 0.114505
R17274 XThC.Tn[6] XThC.Tn[6].n44 0.114505
R17275 XThC.Tn[6] XThC.Tn[6].n48 0.114505
R17276 XThC.Tn[6] XThC.Tn[6].n52 0.114505
R17277 XThC.Tn[6] XThC.Tn[6].n56 0.114505
R17278 XThC.Tn[6] XThC.Tn[6].n60 0.114505
R17279 XThC.Tn[6] XThC.Tn[6].n64 0.114505
R17280 XThC.Tn[6] XThC.Tn[6].n68 0.114505
R17281 XThC.Tn[6] XThC.Tn[6].n72 0.114505
R17282 XThC.Tn[6].n71 XThC.Tn[6].n70 0.0599512
R17283 XThC.Tn[6].n67 XThC.Tn[6].n66 0.0599512
R17284 XThC.Tn[6].n63 XThC.Tn[6].n62 0.0599512
R17285 XThC.Tn[6].n59 XThC.Tn[6].n58 0.0599512
R17286 XThC.Tn[6].n55 XThC.Tn[6].n54 0.0599512
R17287 XThC.Tn[6].n51 XThC.Tn[6].n50 0.0599512
R17288 XThC.Tn[6].n47 XThC.Tn[6].n46 0.0599512
R17289 XThC.Tn[6].n43 XThC.Tn[6].n42 0.0599512
R17290 XThC.Tn[6].n39 XThC.Tn[6].n38 0.0599512
R17291 XThC.Tn[6].n35 XThC.Tn[6].n34 0.0599512
R17292 XThC.Tn[6].n31 XThC.Tn[6].n30 0.0599512
R17293 XThC.Tn[6].n27 XThC.Tn[6].n26 0.0599512
R17294 XThC.Tn[6].n23 XThC.Tn[6].n22 0.0599512
R17295 XThC.Tn[6].n19 XThC.Tn[6].n18 0.0599512
R17296 XThC.Tn[6].n15 XThC.Tn[6].n14 0.0599512
R17297 XThC.Tn[6].n12 XThC.Tn[6].n11 0.0599512
R17298 XThC.Tn[6].n70 XThC.Tn[6] 0.0469286
R17299 XThC.Tn[6].n66 XThC.Tn[6] 0.0469286
R17300 XThC.Tn[6].n62 XThC.Tn[6] 0.0469286
R17301 XThC.Tn[6].n58 XThC.Tn[6] 0.0469286
R17302 XThC.Tn[6].n54 XThC.Tn[6] 0.0469286
R17303 XThC.Tn[6].n50 XThC.Tn[6] 0.0469286
R17304 XThC.Tn[6].n46 XThC.Tn[6] 0.0469286
R17305 XThC.Tn[6].n42 XThC.Tn[6] 0.0469286
R17306 XThC.Tn[6].n38 XThC.Tn[6] 0.0469286
R17307 XThC.Tn[6].n34 XThC.Tn[6] 0.0469286
R17308 XThC.Tn[6].n30 XThC.Tn[6] 0.0469286
R17309 XThC.Tn[6].n26 XThC.Tn[6] 0.0469286
R17310 XThC.Tn[6].n22 XThC.Tn[6] 0.0469286
R17311 XThC.Tn[6].n18 XThC.Tn[6] 0.0469286
R17312 XThC.Tn[6].n14 XThC.Tn[6] 0.0469286
R17313 XThC.Tn[6].n11 XThC.Tn[6] 0.0469286
R17314 XThC.Tn[6].n70 XThC.Tn[6] 0.0401341
R17315 XThC.Tn[6].n66 XThC.Tn[6] 0.0401341
R17316 XThC.Tn[6].n62 XThC.Tn[6] 0.0401341
R17317 XThC.Tn[6].n58 XThC.Tn[6] 0.0401341
R17318 XThC.Tn[6].n54 XThC.Tn[6] 0.0401341
R17319 XThC.Tn[6].n50 XThC.Tn[6] 0.0401341
R17320 XThC.Tn[6].n46 XThC.Tn[6] 0.0401341
R17321 XThC.Tn[6].n42 XThC.Tn[6] 0.0401341
R17322 XThC.Tn[6].n38 XThC.Tn[6] 0.0401341
R17323 XThC.Tn[6].n34 XThC.Tn[6] 0.0401341
R17324 XThC.Tn[6].n30 XThC.Tn[6] 0.0401341
R17325 XThC.Tn[6].n26 XThC.Tn[6] 0.0401341
R17326 XThC.Tn[6].n22 XThC.Tn[6] 0.0401341
R17327 XThC.Tn[6].n18 XThC.Tn[6] 0.0401341
R17328 XThC.Tn[6].n14 XThC.Tn[6] 0.0401341
R17329 XThC.Tn[6].n11 XThC.Tn[6] 0.0401341
R17330 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R17331 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R17332 XThC.Tn[4].n71 XThC.Tn[4].n69 161.365
R17333 XThC.Tn[4].n67 XThC.Tn[4].n65 161.365
R17334 XThC.Tn[4].n63 XThC.Tn[4].n61 161.365
R17335 XThC.Tn[4].n59 XThC.Tn[4].n57 161.365
R17336 XThC.Tn[4].n55 XThC.Tn[4].n53 161.365
R17337 XThC.Tn[4].n51 XThC.Tn[4].n49 161.365
R17338 XThC.Tn[4].n47 XThC.Tn[4].n45 161.365
R17339 XThC.Tn[4].n43 XThC.Tn[4].n41 161.365
R17340 XThC.Tn[4].n39 XThC.Tn[4].n37 161.365
R17341 XThC.Tn[4].n35 XThC.Tn[4].n33 161.365
R17342 XThC.Tn[4].n31 XThC.Tn[4].n29 161.365
R17343 XThC.Tn[4].n27 XThC.Tn[4].n25 161.365
R17344 XThC.Tn[4].n23 XThC.Tn[4].n21 161.365
R17345 XThC.Tn[4].n19 XThC.Tn[4].n17 161.365
R17346 XThC.Tn[4].n15 XThC.Tn[4].n13 161.365
R17347 XThC.Tn[4].n12 XThC.Tn[4].n10 161.365
R17348 XThC.Tn[4].n69 XThC.Tn[4].t18 161.106
R17349 XThC.Tn[4].n65 XThC.Tn[4].t32 161.106
R17350 XThC.Tn[4].n61 XThC.Tn[4].t29 161.106
R17351 XThC.Tn[4].n57 XThC.Tn[4].t27 161.106
R17352 XThC.Tn[4].n53 XThC.Tn[4].t40 161.106
R17353 XThC.Tn[4].n49 XThC.Tn[4].t38 161.106
R17354 XThC.Tn[4].n45 XThC.Tn[4].t26 161.106
R17355 XThC.Tn[4].n41 XThC.Tn[4].t17 161.106
R17356 XThC.Tn[4].n37 XThC.Tn[4].t15 161.106
R17357 XThC.Tn[4].n33 XThC.Tn[4].t37 161.106
R17358 XThC.Tn[4].n29 XThC.Tn[4].t24 161.106
R17359 XThC.Tn[4].n25 XThC.Tn[4].t13 161.106
R17360 XThC.Tn[4].n21 XThC.Tn[4].t36 161.106
R17361 XThC.Tn[4].n17 XThC.Tn[4].t34 161.106
R17362 XThC.Tn[4].n13 XThC.Tn[4].t21 161.106
R17363 XThC.Tn[4].n10 XThC.Tn[4].t12 161.106
R17364 XThC.Tn[4].n69 XThC.Tn[4].t14 154.679
R17365 XThC.Tn[4].n65 XThC.Tn[4].t25 154.679
R17366 XThC.Tn[4].n61 XThC.Tn[4].t23 154.679
R17367 XThC.Tn[4].n57 XThC.Tn[4].t22 154.679
R17368 XThC.Tn[4].n53 XThC.Tn[4].t35 154.679
R17369 XThC.Tn[4].n49 XThC.Tn[4].t33 154.679
R17370 XThC.Tn[4].n45 XThC.Tn[4].t20 154.679
R17371 XThC.Tn[4].n41 XThC.Tn[4].t43 154.679
R17372 XThC.Tn[4].n37 XThC.Tn[4].t42 154.679
R17373 XThC.Tn[4].n33 XThC.Tn[4].t31 154.679
R17374 XThC.Tn[4].n29 XThC.Tn[4].t19 154.679
R17375 XThC.Tn[4].n25 XThC.Tn[4].t41 154.679
R17376 XThC.Tn[4].n21 XThC.Tn[4].t30 154.679
R17377 XThC.Tn[4].n17 XThC.Tn[4].t28 154.679
R17378 XThC.Tn[4].n13 XThC.Tn[4].t16 154.679
R17379 XThC.Tn[4].n10 XThC.Tn[4].t39 154.679
R17380 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R17381 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R17382 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R17383 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R17384 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R17385 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R17386 XThC.Tn[4].n73 XThC.Tn[4].n9 32.6405
R17387 XThC.Tn[4].n1 XThC.Tn[4].t7 26.5955
R17388 XThC.Tn[4].n1 XThC.Tn[4].t6 26.5955
R17389 XThC.Tn[4].n0 XThC.Tn[4].t5 26.5955
R17390 XThC.Tn[4].n0 XThC.Tn[4].t4 26.5955
R17391 XThC.Tn[4].n3 XThC.Tn[4].t9 24.9236
R17392 XThC.Tn[4].n3 XThC.Tn[4].t8 24.9236
R17393 XThC.Tn[4].n4 XThC.Tn[4].t11 24.9236
R17394 XThC.Tn[4].n4 XThC.Tn[4].t10 24.9236
R17395 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R17396 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R17397 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R17398 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R17399 XThC.Tn[4].n74 XThC.Tn[4].n2 18.5605
R17400 XThC.Tn[4].n74 XThC.Tn[4].n73 11.5205
R17401 XThC.Tn[4] XThC.Tn[4].n12 8.0245
R17402 XThC.Tn[4].n72 XThC.Tn[4].n71 7.9105
R17403 XThC.Tn[4].n68 XThC.Tn[4].n67 7.9105
R17404 XThC.Tn[4].n64 XThC.Tn[4].n63 7.9105
R17405 XThC.Tn[4].n60 XThC.Tn[4].n59 7.9105
R17406 XThC.Tn[4].n56 XThC.Tn[4].n55 7.9105
R17407 XThC.Tn[4].n52 XThC.Tn[4].n51 7.9105
R17408 XThC.Tn[4].n48 XThC.Tn[4].n47 7.9105
R17409 XThC.Tn[4].n44 XThC.Tn[4].n43 7.9105
R17410 XThC.Tn[4].n40 XThC.Tn[4].n39 7.9105
R17411 XThC.Tn[4].n36 XThC.Tn[4].n35 7.9105
R17412 XThC.Tn[4].n32 XThC.Tn[4].n31 7.9105
R17413 XThC.Tn[4].n28 XThC.Tn[4].n27 7.9105
R17414 XThC.Tn[4].n24 XThC.Tn[4].n23 7.9105
R17415 XThC.Tn[4].n20 XThC.Tn[4].n19 7.9105
R17416 XThC.Tn[4].n16 XThC.Tn[4].n15 7.9105
R17417 XThC.Tn[4].n73 XThC.Tn[4] 5.77342
R17418 XThC.Tn[4] XThC.Tn[4].n74 0.6405
R17419 XThC.Tn[4].n16 XThC.Tn[4] 0.235138
R17420 XThC.Tn[4].n20 XThC.Tn[4] 0.235138
R17421 XThC.Tn[4].n24 XThC.Tn[4] 0.235138
R17422 XThC.Tn[4].n28 XThC.Tn[4] 0.235138
R17423 XThC.Tn[4].n32 XThC.Tn[4] 0.235138
R17424 XThC.Tn[4].n36 XThC.Tn[4] 0.235138
R17425 XThC.Tn[4].n40 XThC.Tn[4] 0.235138
R17426 XThC.Tn[4].n44 XThC.Tn[4] 0.235138
R17427 XThC.Tn[4].n48 XThC.Tn[4] 0.235138
R17428 XThC.Tn[4].n52 XThC.Tn[4] 0.235138
R17429 XThC.Tn[4].n56 XThC.Tn[4] 0.235138
R17430 XThC.Tn[4].n60 XThC.Tn[4] 0.235138
R17431 XThC.Tn[4].n64 XThC.Tn[4] 0.235138
R17432 XThC.Tn[4].n68 XThC.Tn[4] 0.235138
R17433 XThC.Tn[4].n72 XThC.Tn[4] 0.235138
R17434 XThC.Tn[4] XThC.Tn[4].n16 0.114505
R17435 XThC.Tn[4] XThC.Tn[4].n20 0.114505
R17436 XThC.Tn[4] XThC.Tn[4].n24 0.114505
R17437 XThC.Tn[4] XThC.Tn[4].n28 0.114505
R17438 XThC.Tn[4] XThC.Tn[4].n32 0.114505
R17439 XThC.Tn[4] XThC.Tn[4].n36 0.114505
R17440 XThC.Tn[4] XThC.Tn[4].n40 0.114505
R17441 XThC.Tn[4] XThC.Tn[4].n44 0.114505
R17442 XThC.Tn[4] XThC.Tn[4].n48 0.114505
R17443 XThC.Tn[4] XThC.Tn[4].n52 0.114505
R17444 XThC.Tn[4] XThC.Tn[4].n56 0.114505
R17445 XThC.Tn[4] XThC.Tn[4].n60 0.114505
R17446 XThC.Tn[4] XThC.Tn[4].n64 0.114505
R17447 XThC.Tn[4] XThC.Tn[4].n68 0.114505
R17448 XThC.Tn[4] XThC.Tn[4].n72 0.114505
R17449 XThC.Tn[4].n71 XThC.Tn[4].n70 0.0599512
R17450 XThC.Tn[4].n67 XThC.Tn[4].n66 0.0599512
R17451 XThC.Tn[4].n63 XThC.Tn[4].n62 0.0599512
R17452 XThC.Tn[4].n59 XThC.Tn[4].n58 0.0599512
R17453 XThC.Tn[4].n55 XThC.Tn[4].n54 0.0599512
R17454 XThC.Tn[4].n51 XThC.Tn[4].n50 0.0599512
R17455 XThC.Tn[4].n47 XThC.Tn[4].n46 0.0599512
R17456 XThC.Tn[4].n43 XThC.Tn[4].n42 0.0599512
R17457 XThC.Tn[4].n39 XThC.Tn[4].n38 0.0599512
R17458 XThC.Tn[4].n35 XThC.Tn[4].n34 0.0599512
R17459 XThC.Tn[4].n31 XThC.Tn[4].n30 0.0599512
R17460 XThC.Tn[4].n27 XThC.Tn[4].n26 0.0599512
R17461 XThC.Tn[4].n23 XThC.Tn[4].n22 0.0599512
R17462 XThC.Tn[4].n19 XThC.Tn[4].n18 0.0599512
R17463 XThC.Tn[4].n15 XThC.Tn[4].n14 0.0599512
R17464 XThC.Tn[4].n12 XThC.Tn[4].n11 0.0599512
R17465 XThC.Tn[4].n70 XThC.Tn[4] 0.0469286
R17466 XThC.Tn[4].n66 XThC.Tn[4] 0.0469286
R17467 XThC.Tn[4].n62 XThC.Tn[4] 0.0469286
R17468 XThC.Tn[4].n58 XThC.Tn[4] 0.0469286
R17469 XThC.Tn[4].n54 XThC.Tn[4] 0.0469286
R17470 XThC.Tn[4].n50 XThC.Tn[4] 0.0469286
R17471 XThC.Tn[4].n46 XThC.Tn[4] 0.0469286
R17472 XThC.Tn[4].n42 XThC.Tn[4] 0.0469286
R17473 XThC.Tn[4].n38 XThC.Tn[4] 0.0469286
R17474 XThC.Tn[4].n34 XThC.Tn[4] 0.0469286
R17475 XThC.Tn[4].n30 XThC.Tn[4] 0.0469286
R17476 XThC.Tn[4].n26 XThC.Tn[4] 0.0469286
R17477 XThC.Tn[4].n22 XThC.Tn[4] 0.0469286
R17478 XThC.Tn[4].n18 XThC.Tn[4] 0.0469286
R17479 XThC.Tn[4].n14 XThC.Tn[4] 0.0469286
R17480 XThC.Tn[4].n11 XThC.Tn[4] 0.0469286
R17481 XThC.Tn[4].n70 XThC.Tn[4] 0.0401341
R17482 XThC.Tn[4].n66 XThC.Tn[4] 0.0401341
R17483 XThC.Tn[4].n62 XThC.Tn[4] 0.0401341
R17484 XThC.Tn[4].n58 XThC.Tn[4] 0.0401341
R17485 XThC.Tn[4].n54 XThC.Tn[4] 0.0401341
R17486 XThC.Tn[4].n50 XThC.Tn[4] 0.0401341
R17487 XThC.Tn[4].n46 XThC.Tn[4] 0.0401341
R17488 XThC.Tn[4].n42 XThC.Tn[4] 0.0401341
R17489 XThC.Tn[4].n38 XThC.Tn[4] 0.0401341
R17490 XThC.Tn[4].n34 XThC.Tn[4] 0.0401341
R17491 XThC.Tn[4].n30 XThC.Tn[4] 0.0401341
R17492 XThC.Tn[4].n26 XThC.Tn[4] 0.0401341
R17493 XThC.Tn[4].n22 XThC.Tn[4] 0.0401341
R17494 XThC.Tn[4].n18 XThC.Tn[4] 0.0401341
R17495 XThC.Tn[4].n14 XThC.Tn[4] 0.0401341
R17496 XThC.Tn[4].n11 XThC.Tn[4] 0.0401341
R17497 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R17498 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R17499 XThC.Tn[5].n71 XThC.Tn[5].n69 161.365
R17500 XThC.Tn[5].n67 XThC.Tn[5].n65 161.365
R17501 XThC.Tn[5].n63 XThC.Tn[5].n61 161.365
R17502 XThC.Tn[5].n59 XThC.Tn[5].n57 161.365
R17503 XThC.Tn[5].n55 XThC.Tn[5].n53 161.365
R17504 XThC.Tn[5].n51 XThC.Tn[5].n49 161.365
R17505 XThC.Tn[5].n47 XThC.Tn[5].n45 161.365
R17506 XThC.Tn[5].n43 XThC.Tn[5].n41 161.365
R17507 XThC.Tn[5].n39 XThC.Tn[5].n37 161.365
R17508 XThC.Tn[5].n35 XThC.Tn[5].n33 161.365
R17509 XThC.Tn[5].n31 XThC.Tn[5].n29 161.365
R17510 XThC.Tn[5].n27 XThC.Tn[5].n25 161.365
R17511 XThC.Tn[5].n23 XThC.Tn[5].n21 161.365
R17512 XThC.Tn[5].n19 XThC.Tn[5].n17 161.365
R17513 XThC.Tn[5].n15 XThC.Tn[5].n13 161.365
R17514 XThC.Tn[5].n12 XThC.Tn[5].n10 161.365
R17515 XThC.Tn[5].n69 XThC.Tn[5].t31 161.106
R17516 XThC.Tn[5].n65 XThC.Tn[5].t43 161.106
R17517 XThC.Tn[5].n61 XThC.Tn[5].t41 161.106
R17518 XThC.Tn[5].n57 XThC.Tn[5].t38 161.106
R17519 XThC.Tn[5].n53 XThC.Tn[5].t20 161.106
R17520 XThC.Tn[5].n49 XThC.Tn[5].t18 161.106
R17521 XThC.Tn[5].n45 XThC.Tn[5].t37 161.106
R17522 XThC.Tn[5].n41 XThC.Tn[5].t29 161.106
R17523 XThC.Tn[5].n37 XThC.Tn[5].t26 161.106
R17524 XThC.Tn[5].n33 XThC.Tn[5].t17 161.106
R17525 XThC.Tn[5].n29 XThC.Tn[5].t36 161.106
R17526 XThC.Tn[5].n25 XThC.Tn[5].t25 161.106
R17527 XThC.Tn[5].n21 XThC.Tn[5].t16 161.106
R17528 XThC.Tn[5].n17 XThC.Tn[5].t14 161.106
R17529 XThC.Tn[5].n13 XThC.Tn[5].t32 161.106
R17530 XThC.Tn[5].n10 XThC.Tn[5].t24 161.106
R17531 XThC.Tn[5].n69 XThC.Tn[5].t28 154.679
R17532 XThC.Tn[5].n65 XThC.Tn[5].t40 154.679
R17533 XThC.Tn[5].n61 XThC.Tn[5].t39 154.679
R17534 XThC.Tn[5].n57 XThC.Tn[5].t35 154.679
R17535 XThC.Tn[5].n53 XThC.Tn[5].t19 154.679
R17536 XThC.Tn[5].n49 XThC.Tn[5].t15 154.679
R17537 XThC.Tn[5].n45 XThC.Tn[5].t34 154.679
R17538 XThC.Tn[5].n41 XThC.Tn[5].t27 154.679
R17539 XThC.Tn[5].n37 XThC.Tn[5].t23 154.679
R17540 XThC.Tn[5].n33 XThC.Tn[5].t13 154.679
R17541 XThC.Tn[5].n29 XThC.Tn[5].t33 154.679
R17542 XThC.Tn[5].n25 XThC.Tn[5].t22 154.679
R17543 XThC.Tn[5].n21 XThC.Tn[5].t12 154.679
R17544 XThC.Tn[5].n17 XThC.Tn[5].t42 154.679
R17545 XThC.Tn[5].n13 XThC.Tn[5].t30 154.679
R17546 XThC.Tn[5].n10 XThC.Tn[5].t21 154.679
R17547 XThC.Tn[5].n7 XThC.Tn[5].n6 135.249
R17548 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R17549 XThC.Tn[5].n8 XThC.Tn[5].n4 98.981
R17550 XThC.Tn[5].n7 XThC.Tn[5].n5 98.981
R17551 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R17552 XThC.Tn[5].n8 XThC.Tn[5].n7 36.2672
R17553 XThC.Tn[5].n73 XThC.Tn[5].n9 32.6405
R17554 XThC.Tn[5].n1 XThC.Tn[5].t9 26.5955
R17555 XThC.Tn[5].n1 XThC.Tn[5].t8 26.5955
R17556 XThC.Tn[5].n0 XThC.Tn[5].t11 26.5955
R17557 XThC.Tn[5].n0 XThC.Tn[5].t10 26.5955
R17558 XThC.Tn[5].n3 XThC.Tn[5].t5 24.9236
R17559 XThC.Tn[5].n3 XThC.Tn[5].t4 24.9236
R17560 XThC.Tn[5].n4 XThC.Tn[5].t7 24.9236
R17561 XThC.Tn[5].n4 XThC.Tn[5].t6 24.9236
R17562 XThC.Tn[5].n5 XThC.Tn[5].t2 24.9236
R17563 XThC.Tn[5].n5 XThC.Tn[5].t1 24.9236
R17564 XThC.Tn[5].n6 XThC.Tn[5].t0 24.9236
R17565 XThC.Tn[5].n6 XThC.Tn[5].t3 24.9236
R17566 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R17567 XThC.Tn[5] XThC.Tn[5].n12 8.0245
R17568 XThC.Tn[5].n72 XThC.Tn[5].n71 7.9105
R17569 XThC.Tn[5].n68 XThC.Tn[5].n67 7.9105
R17570 XThC.Tn[5].n64 XThC.Tn[5].n63 7.9105
R17571 XThC.Tn[5].n60 XThC.Tn[5].n59 7.9105
R17572 XThC.Tn[5].n56 XThC.Tn[5].n55 7.9105
R17573 XThC.Tn[5].n52 XThC.Tn[5].n51 7.9105
R17574 XThC.Tn[5].n48 XThC.Tn[5].n47 7.9105
R17575 XThC.Tn[5].n44 XThC.Tn[5].n43 7.9105
R17576 XThC.Tn[5].n40 XThC.Tn[5].n39 7.9105
R17577 XThC.Tn[5].n36 XThC.Tn[5].n35 7.9105
R17578 XThC.Tn[5].n32 XThC.Tn[5].n31 7.9105
R17579 XThC.Tn[5].n28 XThC.Tn[5].n27 7.9105
R17580 XThC.Tn[5].n24 XThC.Tn[5].n23 7.9105
R17581 XThC.Tn[5].n20 XThC.Tn[5].n19 7.9105
R17582 XThC.Tn[5].n16 XThC.Tn[5].n15 7.9105
R17583 XThC.Tn[5] XThC.Tn[5].n73 6.7205
R17584 XThC.Tn[5].n73 XThC.Tn[5] 5.69842
R17585 XThC.Tn[5].n16 XThC.Tn[5] 0.235138
R17586 XThC.Tn[5].n20 XThC.Tn[5] 0.235138
R17587 XThC.Tn[5].n24 XThC.Tn[5] 0.235138
R17588 XThC.Tn[5].n28 XThC.Tn[5] 0.235138
R17589 XThC.Tn[5].n32 XThC.Tn[5] 0.235138
R17590 XThC.Tn[5].n36 XThC.Tn[5] 0.235138
R17591 XThC.Tn[5].n40 XThC.Tn[5] 0.235138
R17592 XThC.Tn[5].n44 XThC.Tn[5] 0.235138
R17593 XThC.Tn[5].n48 XThC.Tn[5] 0.235138
R17594 XThC.Tn[5].n52 XThC.Tn[5] 0.235138
R17595 XThC.Tn[5].n56 XThC.Tn[5] 0.235138
R17596 XThC.Tn[5].n60 XThC.Tn[5] 0.235138
R17597 XThC.Tn[5].n64 XThC.Tn[5] 0.235138
R17598 XThC.Tn[5].n68 XThC.Tn[5] 0.235138
R17599 XThC.Tn[5].n72 XThC.Tn[5] 0.235138
R17600 XThC.Tn[5] XThC.Tn[5].n16 0.114505
R17601 XThC.Tn[5] XThC.Tn[5].n20 0.114505
R17602 XThC.Tn[5] XThC.Tn[5].n24 0.114505
R17603 XThC.Tn[5] XThC.Tn[5].n28 0.114505
R17604 XThC.Tn[5] XThC.Tn[5].n32 0.114505
R17605 XThC.Tn[5] XThC.Tn[5].n36 0.114505
R17606 XThC.Tn[5] XThC.Tn[5].n40 0.114505
R17607 XThC.Tn[5] XThC.Tn[5].n44 0.114505
R17608 XThC.Tn[5] XThC.Tn[5].n48 0.114505
R17609 XThC.Tn[5] XThC.Tn[5].n52 0.114505
R17610 XThC.Tn[5] XThC.Tn[5].n56 0.114505
R17611 XThC.Tn[5] XThC.Tn[5].n60 0.114505
R17612 XThC.Tn[5] XThC.Tn[5].n64 0.114505
R17613 XThC.Tn[5] XThC.Tn[5].n68 0.114505
R17614 XThC.Tn[5] XThC.Tn[5].n72 0.114505
R17615 XThC.Tn[5].n71 XThC.Tn[5].n70 0.0599512
R17616 XThC.Tn[5].n67 XThC.Tn[5].n66 0.0599512
R17617 XThC.Tn[5].n63 XThC.Tn[5].n62 0.0599512
R17618 XThC.Tn[5].n59 XThC.Tn[5].n58 0.0599512
R17619 XThC.Tn[5].n55 XThC.Tn[5].n54 0.0599512
R17620 XThC.Tn[5].n51 XThC.Tn[5].n50 0.0599512
R17621 XThC.Tn[5].n47 XThC.Tn[5].n46 0.0599512
R17622 XThC.Tn[5].n43 XThC.Tn[5].n42 0.0599512
R17623 XThC.Tn[5].n39 XThC.Tn[5].n38 0.0599512
R17624 XThC.Tn[5].n35 XThC.Tn[5].n34 0.0599512
R17625 XThC.Tn[5].n31 XThC.Tn[5].n30 0.0599512
R17626 XThC.Tn[5].n27 XThC.Tn[5].n26 0.0599512
R17627 XThC.Tn[5].n23 XThC.Tn[5].n22 0.0599512
R17628 XThC.Tn[5].n19 XThC.Tn[5].n18 0.0599512
R17629 XThC.Tn[5].n15 XThC.Tn[5].n14 0.0599512
R17630 XThC.Tn[5].n12 XThC.Tn[5].n11 0.0599512
R17631 XThC.Tn[5].n70 XThC.Tn[5] 0.0469286
R17632 XThC.Tn[5].n66 XThC.Tn[5] 0.0469286
R17633 XThC.Tn[5].n62 XThC.Tn[5] 0.0469286
R17634 XThC.Tn[5].n58 XThC.Tn[5] 0.0469286
R17635 XThC.Tn[5].n54 XThC.Tn[5] 0.0469286
R17636 XThC.Tn[5].n50 XThC.Tn[5] 0.0469286
R17637 XThC.Tn[5].n46 XThC.Tn[5] 0.0469286
R17638 XThC.Tn[5].n42 XThC.Tn[5] 0.0469286
R17639 XThC.Tn[5].n38 XThC.Tn[5] 0.0469286
R17640 XThC.Tn[5].n34 XThC.Tn[5] 0.0469286
R17641 XThC.Tn[5].n30 XThC.Tn[5] 0.0469286
R17642 XThC.Tn[5].n26 XThC.Tn[5] 0.0469286
R17643 XThC.Tn[5].n22 XThC.Tn[5] 0.0469286
R17644 XThC.Tn[5].n18 XThC.Tn[5] 0.0469286
R17645 XThC.Tn[5].n14 XThC.Tn[5] 0.0469286
R17646 XThC.Tn[5].n11 XThC.Tn[5] 0.0469286
R17647 XThC.Tn[5].n70 XThC.Tn[5] 0.0401341
R17648 XThC.Tn[5].n66 XThC.Tn[5] 0.0401341
R17649 XThC.Tn[5].n62 XThC.Tn[5] 0.0401341
R17650 XThC.Tn[5].n58 XThC.Tn[5] 0.0401341
R17651 XThC.Tn[5].n54 XThC.Tn[5] 0.0401341
R17652 XThC.Tn[5].n50 XThC.Tn[5] 0.0401341
R17653 XThC.Tn[5].n46 XThC.Tn[5] 0.0401341
R17654 XThC.Tn[5].n42 XThC.Tn[5] 0.0401341
R17655 XThC.Tn[5].n38 XThC.Tn[5] 0.0401341
R17656 XThC.Tn[5].n34 XThC.Tn[5] 0.0401341
R17657 XThC.Tn[5].n30 XThC.Tn[5] 0.0401341
R17658 XThC.Tn[5].n26 XThC.Tn[5] 0.0401341
R17659 XThC.Tn[5].n22 XThC.Tn[5] 0.0401341
R17660 XThC.Tn[5].n18 XThC.Tn[5] 0.0401341
R17661 XThC.Tn[5].n14 XThC.Tn[5] 0.0401341
R17662 XThC.Tn[5].n11 XThC.Tn[5] 0.0401341
R17663 XThR.Tn[7].n5 XThR.Tn[7].n3 244.067
R17664 XThR.Tn[7].n2 XThR.Tn[7].n0 236.589
R17665 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R17666 XThR.Tn[7].n2 XThR.Tn[7].n1 200.321
R17667 XThR.Tn[7] XThR.Tn[7].n79 161.363
R17668 XThR.Tn[7] XThR.Tn[7].n74 161.363
R17669 XThR.Tn[7] XThR.Tn[7].n69 161.363
R17670 XThR.Tn[7] XThR.Tn[7].n64 161.363
R17671 XThR.Tn[7] XThR.Tn[7].n59 161.363
R17672 XThR.Tn[7] XThR.Tn[7].n54 161.363
R17673 XThR.Tn[7] XThR.Tn[7].n49 161.363
R17674 XThR.Tn[7] XThR.Tn[7].n44 161.363
R17675 XThR.Tn[7] XThR.Tn[7].n39 161.363
R17676 XThR.Tn[7] XThR.Tn[7].n34 161.363
R17677 XThR.Tn[7] XThR.Tn[7].n29 161.363
R17678 XThR.Tn[7] XThR.Tn[7].n24 161.363
R17679 XThR.Tn[7] XThR.Tn[7].n19 161.363
R17680 XThR.Tn[7] XThR.Tn[7].n14 161.363
R17681 XThR.Tn[7] XThR.Tn[7].n9 161.363
R17682 XThR.Tn[7] XThR.Tn[7].n7 161.363
R17683 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R17684 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R17685 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R17686 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R17687 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R17688 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R17689 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R17690 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R17691 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R17692 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R17693 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R17694 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R17695 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R17696 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R17697 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R17698 XThR.Tn[7].n80 XThR.Tn[7].t12 161.106
R17699 XThR.Tn[7].n79 XThR.Tn[7].t14 161.106
R17700 XThR.Tn[7].n75 XThR.Tn[7].t18 161.106
R17701 XThR.Tn[7].n74 XThR.Tn[7].t23 161.106
R17702 XThR.Tn[7].n70 XThR.Tn[7].t62 161.106
R17703 XThR.Tn[7].n69 XThR.Tn[7].t67 161.106
R17704 XThR.Tn[7].n65 XThR.Tn[7].t45 161.106
R17705 XThR.Tn[7].n64 XThR.Tn[7].t47 161.106
R17706 XThR.Tn[7].n60 XThR.Tn[7].t11 161.106
R17707 XThR.Tn[7].n59 XThR.Tn[7].t13 161.106
R17708 XThR.Tn[7].n55 XThR.Tn[7].t35 161.106
R17709 XThR.Tn[7].n54 XThR.Tn[7].t40 161.106
R17710 XThR.Tn[7].n50 XThR.Tn[7].t16 161.106
R17711 XThR.Tn[7].n49 XThR.Tn[7].t21 161.106
R17712 XThR.Tn[7].n45 XThR.Tn[7].t59 161.106
R17713 XThR.Tn[7].n44 XThR.Tn[7].t64 161.106
R17714 XThR.Tn[7].n40 XThR.Tn[7].t44 161.106
R17715 XThR.Tn[7].n39 XThR.Tn[7].t46 161.106
R17716 XThR.Tn[7].n35 XThR.Tn[7].t49 161.106
R17717 XThR.Tn[7].n34 XThR.Tn[7].t54 161.106
R17718 XThR.Tn[7].n30 XThR.Tn[7].t34 161.106
R17719 XThR.Tn[7].n29 XThR.Tn[7].t39 161.106
R17720 XThR.Tn[7].n25 XThR.Tn[7].t61 161.106
R17721 XThR.Tn[7].n24 XThR.Tn[7].t66 161.106
R17722 XThR.Tn[7].n20 XThR.Tn[7].t31 161.106
R17723 XThR.Tn[7].n19 XThR.Tn[7].t37 161.106
R17724 XThR.Tn[7].n15 XThR.Tn[7].t15 161.106
R17725 XThR.Tn[7].n14 XThR.Tn[7].t19 161.106
R17726 XThR.Tn[7].n10 XThR.Tn[7].t42 161.106
R17727 XThR.Tn[7].n9 XThR.Tn[7].t43 161.106
R17728 XThR.Tn[7].n7 XThR.Tn[7].t26 161.106
R17729 XThR.Tn[7].n80 XThR.Tn[7].t29 154.679
R17730 XThR.Tn[7].n79 XThR.Tn[7].t33 154.679
R17731 XThR.Tn[7].n75 XThR.Tn[7].t8 154.679
R17732 XThR.Tn[7].n74 XThR.Tn[7].t10 154.679
R17733 XThR.Tn[7].n70 XThR.Tn[7].t51 154.679
R17734 XThR.Tn[7].n69 XThR.Tn[7].t56 154.679
R17735 XThR.Tn[7].n65 XThR.Tn[7].t20 154.679
R17736 XThR.Tn[7].n64 XThR.Tn[7].t24 154.679
R17737 XThR.Tn[7].n60 XThR.Tn[7].t63 154.679
R17738 XThR.Tn[7].n59 XThR.Tn[7].t68 154.679
R17739 XThR.Tn[7].n55 XThR.Tn[7].t28 154.679
R17740 XThR.Tn[7].n54 XThR.Tn[7].t30 154.679
R17741 XThR.Tn[7].n50 XThR.Tn[7].t52 154.679
R17742 XThR.Tn[7].n49 XThR.Tn[7].t57 154.679
R17743 XThR.Tn[7].n45 XThR.Tn[7].t36 154.679
R17744 XThR.Tn[7].n44 XThR.Tn[7].t41 154.679
R17745 XThR.Tn[7].n40 XThR.Tn[7].t17 154.679
R17746 XThR.Tn[7].n39 XThR.Tn[7].t22 154.679
R17747 XThR.Tn[7].n35 XThR.Tn[7].t60 154.679
R17748 XThR.Tn[7].n34 XThR.Tn[7].t65 154.679
R17749 XThR.Tn[7].n30 XThR.Tn[7].t69 154.679
R17750 XThR.Tn[7].n29 XThR.Tn[7].t9 154.679
R17751 XThR.Tn[7].n25 XThR.Tn[7].t50 154.679
R17752 XThR.Tn[7].n24 XThR.Tn[7].t55 154.679
R17753 XThR.Tn[7].n20 XThR.Tn[7].t25 154.679
R17754 XThR.Tn[7].n19 XThR.Tn[7].t27 154.679
R17755 XThR.Tn[7].n15 XThR.Tn[7].t48 154.679
R17756 XThR.Tn[7].n14 XThR.Tn[7].t53 154.679
R17757 XThR.Tn[7].n10 XThR.Tn[7].t32 154.679
R17758 XThR.Tn[7].n9 XThR.Tn[7].t38 154.679
R17759 XThR.Tn[7].n7 XThR.Tn[7].t58 154.679
R17760 XThR.Tn[7].n4 XThR.Tn[7].t1 26.5955
R17761 XThR.Tn[7].n4 XThR.Tn[7].t0 26.5955
R17762 XThR.Tn[7].n3 XThR.Tn[7].t2 26.5955
R17763 XThR.Tn[7].n3 XThR.Tn[7].t3 26.5955
R17764 XThR.Tn[7].n0 XThR.Tn[7].t7 24.9236
R17765 XThR.Tn[7].n0 XThR.Tn[7].t4 24.9236
R17766 XThR.Tn[7].n1 XThR.Tn[7].t6 24.9236
R17767 XThR.Tn[7].n1 XThR.Tn[7].t5 24.9236
R17768 XThR.Tn[7] XThR.Tn[7].n2 16.079
R17769 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R17770 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R17771 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R17772 XThR.Tn[7] XThR.Tn[7].n8 5.34871
R17773 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R17774 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R17775 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R17776 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R17777 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R17778 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R17779 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R17780 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R17781 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R17782 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R17783 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R17784 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R17785 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R17786 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R17787 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R17788 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R17789 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R17790 XThR.Tn[7].n13 XThR.Tn[7] 2.51836
R17791 XThR.Tn[7].n18 XThR.Tn[7] 2.51836
R17792 XThR.Tn[7].n23 XThR.Tn[7] 2.51836
R17793 XThR.Tn[7].n28 XThR.Tn[7] 2.51836
R17794 XThR.Tn[7].n33 XThR.Tn[7] 2.51836
R17795 XThR.Tn[7].n38 XThR.Tn[7] 2.51836
R17796 XThR.Tn[7].n43 XThR.Tn[7] 2.51836
R17797 XThR.Tn[7].n48 XThR.Tn[7] 2.51836
R17798 XThR.Tn[7].n53 XThR.Tn[7] 2.51836
R17799 XThR.Tn[7].n58 XThR.Tn[7] 2.51836
R17800 XThR.Tn[7].n63 XThR.Tn[7] 2.51836
R17801 XThR.Tn[7].n68 XThR.Tn[7] 2.51836
R17802 XThR.Tn[7].n73 XThR.Tn[7] 2.51836
R17803 XThR.Tn[7].n78 XThR.Tn[7] 2.51836
R17804 XThR.Tn[7].n83 XThR.Tn[7] 2.51836
R17805 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R17806 XThR.Tn[7] XThR.Tn[7].n13 0.848714
R17807 XThR.Tn[7] XThR.Tn[7].n18 0.848714
R17808 XThR.Tn[7] XThR.Tn[7].n23 0.848714
R17809 XThR.Tn[7] XThR.Tn[7].n28 0.848714
R17810 XThR.Tn[7] XThR.Tn[7].n33 0.848714
R17811 XThR.Tn[7] XThR.Tn[7].n38 0.848714
R17812 XThR.Tn[7] XThR.Tn[7].n43 0.848714
R17813 XThR.Tn[7] XThR.Tn[7].n48 0.848714
R17814 XThR.Tn[7] XThR.Tn[7].n53 0.848714
R17815 XThR.Tn[7] XThR.Tn[7].n58 0.848714
R17816 XThR.Tn[7] XThR.Tn[7].n63 0.848714
R17817 XThR.Tn[7] XThR.Tn[7].n68 0.848714
R17818 XThR.Tn[7] XThR.Tn[7].n73 0.848714
R17819 XThR.Tn[7] XThR.Tn[7].n78 0.848714
R17820 XThR.Tn[7] XThR.Tn[7].n83 0.848714
R17821 XThR.Tn[7].n6 XThR.Tn[7] 0.830612
R17822 XThR.Tn[7].n8 XThR.Tn[7] 0.485653
R17823 XThR.Tn[7].n81 XThR.Tn[7] 0.21482
R17824 XThR.Tn[7].n76 XThR.Tn[7] 0.21482
R17825 XThR.Tn[7].n71 XThR.Tn[7] 0.21482
R17826 XThR.Tn[7].n66 XThR.Tn[7] 0.21482
R17827 XThR.Tn[7].n61 XThR.Tn[7] 0.21482
R17828 XThR.Tn[7].n56 XThR.Tn[7] 0.21482
R17829 XThR.Tn[7].n51 XThR.Tn[7] 0.21482
R17830 XThR.Tn[7].n46 XThR.Tn[7] 0.21482
R17831 XThR.Tn[7].n41 XThR.Tn[7] 0.21482
R17832 XThR.Tn[7].n36 XThR.Tn[7] 0.21482
R17833 XThR.Tn[7].n31 XThR.Tn[7] 0.21482
R17834 XThR.Tn[7].n26 XThR.Tn[7] 0.21482
R17835 XThR.Tn[7].n21 XThR.Tn[7] 0.21482
R17836 XThR.Tn[7].n16 XThR.Tn[7] 0.21482
R17837 XThR.Tn[7].n11 XThR.Tn[7] 0.21482
R17838 XThR.Tn[7].n82 XThR.Tn[7] 0.0608448
R17839 XThR.Tn[7].n77 XThR.Tn[7] 0.0608448
R17840 XThR.Tn[7].n72 XThR.Tn[7] 0.0608448
R17841 XThR.Tn[7].n67 XThR.Tn[7] 0.0608448
R17842 XThR.Tn[7].n62 XThR.Tn[7] 0.0608448
R17843 XThR.Tn[7].n57 XThR.Tn[7] 0.0608448
R17844 XThR.Tn[7].n52 XThR.Tn[7] 0.0608448
R17845 XThR.Tn[7].n47 XThR.Tn[7] 0.0608448
R17846 XThR.Tn[7].n42 XThR.Tn[7] 0.0608448
R17847 XThR.Tn[7].n37 XThR.Tn[7] 0.0608448
R17848 XThR.Tn[7].n32 XThR.Tn[7] 0.0608448
R17849 XThR.Tn[7].n27 XThR.Tn[7] 0.0608448
R17850 XThR.Tn[7].n22 XThR.Tn[7] 0.0608448
R17851 XThR.Tn[7].n17 XThR.Tn[7] 0.0608448
R17852 XThR.Tn[7].n12 XThR.Tn[7] 0.0608448
R17853 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R17854 XThR.Tn[7] XThR.Tn[7].n84 0.038
R17855 XThR.Tn[7].n8 XThR.Tn[7] 0.00744444
R17856 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00265517
R17857 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00265517
R17858 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00265517
R17859 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00265517
R17860 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00265517
R17861 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00265517
R17862 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00265517
R17863 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00265517
R17864 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00265517
R17865 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00265517
R17866 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00265517
R17867 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00265517
R17868 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00265517
R17869 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00265517
R17870 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00265517
R17871 XThC.Tn[12].n70 XThC.Tn[12].n69 256.103
R17872 XThC.Tn[12].n74 XThC.Tn[12].n72 243.68
R17873 XThC.Tn[12].n2 XThC.Tn[12].n0 241.847
R17874 XThC.Tn[12].n74 XThC.Tn[12].n73 205.28
R17875 XThC.Tn[12].n70 XThC.Tn[12].n68 202.095
R17876 XThC.Tn[12].n2 XThC.Tn[12].n1 185
R17877 XThC.Tn[12].n64 XThC.Tn[12].n62 161.365
R17878 XThC.Tn[12].n60 XThC.Tn[12].n58 161.365
R17879 XThC.Tn[12].n56 XThC.Tn[12].n54 161.365
R17880 XThC.Tn[12].n52 XThC.Tn[12].n50 161.365
R17881 XThC.Tn[12].n48 XThC.Tn[12].n46 161.365
R17882 XThC.Tn[12].n44 XThC.Tn[12].n42 161.365
R17883 XThC.Tn[12].n40 XThC.Tn[12].n38 161.365
R17884 XThC.Tn[12].n36 XThC.Tn[12].n34 161.365
R17885 XThC.Tn[12].n32 XThC.Tn[12].n30 161.365
R17886 XThC.Tn[12].n28 XThC.Tn[12].n26 161.365
R17887 XThC.Tn[12].n24 XThC.Tn[12].n22 161.365
R17888 XThC.Tn[12].n20 XThC.Tn[12].n18 161.365
R17889 XThC.Tn[12].n16 XThC.Tn[12].n14 161.365
R17890 XThC.Tn[12].n12 XThC.Tn[12].n10 161.365
R17891 XThC.Tn[12].n8 XThC.Tn[12].n6 161.365
R17892 XThC.Tn[12].n5 XThC.Tn[12].n3 161.365
R17893 XThC.Tn[12].n62 XThC.Tn[12].t28 161.106
R17894 XThC.Tn[12].n58 XThC.Tn[12].t42 161.106
R17895 XThC.Tn[12].n54 XThC.Tn[12].t39 161.106
R17896 XThC.Tn[12].n50 XThC.Tn[12].t37 161.106
R17897 XThC.Tn[12].n46 XThC.Tn[12].t18 161.106
R17898 XThC.Tn[12].n42 XThC.Tn[12].t16 161.106
R17899 XThC.Tn[12].n38 XThC.Tn[12].t36 161.106
R17900 XThC.Tn[12].n34 XThC.Tn[12].t27 161.106
R17901 XThC.Tn[12].n30 XThC.Tn[12].t25 161.106
R17902 XThC.Tn[12].n26 XThC.Tn[12].t15 161.106
R17903 XThC.Tn[12].n22 XThC.Tn[12].t34 161.106
R17904 XThC.Tn[12].n18 XThC.Tn[12].t23 161.106
R17905 XThC.Tn[12].n14 XThC.Tn[12].t14 161.106
R17906 XThC.Tn[12].n10 XThC.Tn[12].t12 161.106
R17907 XThC.Tn[12].n6 XThC.Tn[12].t31 161.106
R17908 XThC.Tn[12].n3 XThC.Tn[12].t22 161.106
R17909 XThC.Tn[12].n62 XThC.Tn[12].t24 154.679
R17910 XThC.Tn[12].n58 XThC.Tn[12].t35 154.679
R17911 XThC.Tn[12].n54 XThC.Tn[12].t33 154.679
R17912 XThC.Tn[12].n50 XThC.Tn[12].t32 154.679
R17913 XThC.Tn[12].n46 XThC.Tn[12].t13 154.679
R17914 XThC.Tn[12].n42 XThC.Tn[12].t43 154.679
R17915 XThC.Tn[12].n38 XThC.Tn[12].t30 154.679
R17916 XThC.Tn[12].n34 XThC.Tn[12].t21 154.679
R17917 XThC.Tn[12].n30 XThC.Tn[12].t20 154.679
R17918 XThC.Tn[12].n26 XThC.Tn[12].t41 154.679
R17919 XThC.Tn[12].n22 XThC.Tn[12].t29 154.679
R17920 XThC.Tn[12].n18 XThC.Tn[12].t19 154.679
R17921 XThC.Tn[12].n14 XThC.Tn[12].t40 154.679
R17922 XThC.Tn[12].n10 XThC.Tn[12].t38 154.679
R17923 XThC.Tn[12].n6 XThC.Tn[12].t26 154.679
R17924 XThC.Tn[12].n3 XThC.Tn[12].t17 154.679
R17925 XThC.Tn[12].n68 XThC.Tn[12].t1 26.5955
R17926 XThC.Tn[12].n68 XThC.Tn[12].t2 26.5955
R17927 XThC.Tn[12].n72 XThC.Tn[12].t9 26.5955
R17928 XThC.Tn[12].n72 XThC.Tn[12].t8 26.5955
R17929 XThC.Tn[12].n73 XThC.Tn[12].t11 26.5955
R17930 XThC.Tn[12].n73 XThC.Tn[12].t10 26.5955
R17931 XThC.Tn[12].n69 XThC.Tn[12].t0 26.5955
R17932 XThC.Tn[12].n69 XThC.Tn[12].t3 26.5955
R17933 XThC.Tn[12].n1 XThC.Tn[12].t5 24.9236
R17934 XThC.Tn[12].n1 XThC.Tn[12].t4 24.9236
R17935 XThC.Tn[12].n0 XThC.Tn[12].t7 24.9236
R17936 XThC.Tn[12].n0 XThC.Tn[12].t6 24.9236
R17937 XThC.Tn[12] XThC.Tn[12].n74 22.9652
R17938 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R17939 XThC.Tn[12].n71 XThC.Tn[12].n70 13.9299
R17940 XThC.Tn[12] XThC.Tn[12].n71 13.9299
R17941 XThC.Tn[12] XThC.Tn[12].n5 8.0245
R17942 XThC.Tn[12].n65 XThC.Tn[12].n64 7.9105
R17943 XThC.Tn[12].n61 XThC.Tn[12].n60 7.9105
R17944 XThC.Tn[12].n57 XThC.Tn[12].n56 7.9105
R17945 XThC.Tn[12].n53 XThC.Tn[12].n52 7.9105
R17946 XThC.Tn[12].n49 XThC.Tn[12].n48 7.9105
R17947 XThC.Tn[12].n45 XThC.Tn[12].n44 7.9105
R17948 XThC.Tn[12].n41 XThC.Tn[12].n40 7.9105
R17949 XThC.Tn[12].n37 XThC.Tn[12].n36 7.9105
R17950 XThC.Tn[12].n33 XThC.Tn[12].n32 7.9105
R17951 XThC.Tn[12].n29 XThC.Tn[12].n28 7.9105
R17952 XThC.Tn[12].n25 XThC.Tn[12].n24 7.9105
R17953 XThC.Tn[12].n21 XThC.Tn[12].n20 7.9105
R17954 XThC.Tn[12].n17 XThC.Tn[12].n16 7.9105
R17955 XThC.Tn[12].n13 XThC.Tn[12].n12 7.9105
R17956 XThC.Tn[12].n9 XThC.Tn[12].n8 7.9105
R17957 XThC.Tn[12].n67 XThC.Tn[12].n66 7.4309
R17958 XThC.Tn[12].n66 XThC.Tn[12] 4.71945
R17959 XThC.Tn[12].n71 XThC.Tn[12].n67 2.99115
R17960 XThC.Tn[12].n71 XThC.Tn[12] 2.87153
R17961 XThC.Tn[12].n67 XThC.Tn[12] 2.2734
R17962 XThC.Tn[12].n66 XThC.Tn[12] 0.88175
R17963 XThC.Tn[12].n9 XThC.Tn[12] 0.235138
R17964 XThC.Tn[12].n13 XThC.Tn[12] 0.235138
R17965 XThC.Tn[12].n17 XThC.Tn[12] 0.235138
R17966 XThC.Tn[12].n21 XThC.Tn[12] 0.235138
R17967 XThC.Tn[12].n25 XThC.Tn[12] 0.235138
R17968 XThC.Tn[12].n29 XThC.Tn[12] 0.235138
R17969 XThC.Tn[12].n33 XThC.Tn[12] 0.235138
R17970 XThC.Tn[12].n37 XThC.Tn[12] 0.235138
R17971 XThC.Tn[12].n41 XThC.Tn[12] 0.235138
R17972 XThC.Tn[12].n45 XThC.Tn[12] 0.235138
R17973 XThC.Tn[12].n49 XThC.Tn[12] 0.235138
R17974 XThC.Tn[12].n53 XThC.Tn[12] 0.235138
R17975 XThC.Tn[12].n57 XThC.Tn[12] 0.235138
R17976 XThC.Tn[12].n61 XThC.Tn[12] 0.235138
R17977 XThC.Tn[12].n65 XThC.Tn[12] 0.235138
R17978 XThC.Tn[12] XThC.Tn[12].n9 0.114505
R17979 XThC.Tn[12] XThC.Tn[12].n13 0.114505
R17980 XThC.Tn[12] XThC.Tn[12].n17 0.114505
R17981 XThC.Tn[12] XThC.Tn[12].n21 0.114505
R17982 XThC.Tn[12] XThC.Tn[12].n25 0.114505
R17983 XThC.Tn[12] XThC.Tn[12].n29 0.114505
R17984 XThC.Tn[12] XThC.Tn[12].n33 0.114505
R17985 XThC.Tn[12] XThC.Tn[12].n37 0.114505
R17986 XThC.Tn[12] XThC.Tn[12].n41 0.114505
R17987 XThC.Tn[12] XThC.Tn[12].n45 0.114505
R17988 XThC.Tn[12] XThC.Tn[12].n49 0.114505
R17989 XThC.Tn[12] XThC.Tn[12].n53 0.114505
R17990 XThC.Tn[12] XThC.Tn[12].n57 0.114505
R17991 XThC.Tn[12] XThC.Tn[12].n61 0.114505
R17992 XThC.Tn[12] XThC.Tn[12].n65 0.114505
R17993 XThC.Tn[12].n64 XThC.Tn[12].n63 0.0599512
R17994 XThC.Tn[12].n60 XThC.Tn[12].n59 0.0599512
R17995 XThC.Tn[12].n56 XThC.Tn[12].n55 0.0599512
R17996 XThC.Tn[12].n52 XThC.Tn[12].n51 0.0599512
R17997 XThC.Tn[12].n48 XThC.Tn[12].n47 0.0599512
R17998 XThC.Tn[12].n44 XThC.Tn[12].n43 0.0599512
R17999 XThC.Tn[12].n40 XThC.Tn[12].n39 0.0599512
R18000 XThC.Tn[12].n36 XThC.Tn[12].n35 0.0599512
R18001 XThC.Tn[12].n32 XThC.Tn[12].n31 0.0599512
R18002 XThC.Tn[12].n28 XThC.Tn[12].n27 0.0599512
R18003 XThC.Tn[12].n24 XThC.Tn[12].n23 0.0599512
R18004 XThC.Tn[12].n20 XThC.Tn[12].n19 0.0599512
R18005 XThC.Tn[12].n16 XThC.Tn[12].n15 0.0599512
R18006 XThC.Tn[12].n12 XThC.Tn[12].n11 0.0599512
R18007 XThC.Tn[12].n8 XThC.Tn[12].n7 0.0599512
R18008 XThC.Tn[12].n5 XThC.Tn[12].n4 0.0599512
R18009 XThC.Tn[12].n63 XThC.Tn[12] 0.0469286
R18010 XThC.Tn[12].n59 XThC.Tn[12] 0.0469286
R18011 XThC.Tn[12].n55 XThC.Tn[12] 0.0469286
R18012 XThC.Tn[12].n51 XThC.Tn[12] 0.0469286
R18013 XThC.Tn[12].n47 XThC.Tn[12] 0.0469286
R18014 XThC.Tn[12].n43 XThC.Tn[12] 0.0469286
R18015 XThC.Tn[12].n39 XThC.Tn[12] 0.0469286
R18016 XThC.Tn[12].n35 XThC.Tn[12] 0.0469286
R18017 XThC.Tn[12].n31 XThC.Tn[12] 0.0469286
R18018 XThC.Tn[12].n27 XThC.Tn[12] 0.0469286
R18019 XThC.Tn[12].n23 XThC.Tn[12] 0.0469286
R18020 XThC.Tn[12].n19 XThC.Tn[12] 0.0469286
R18021 XThC.Tn[12].n15 XThC.Tn[12] 0.0469286
R18022 XThC.Tn[12].n11 XThC.Tn[12] 0.0469286
R18023 XThC.Tn[12].n7 XThC.Tn[12] 0.0469286
R18024 XThC.Tn[12].n4 XThC.Tn[12] 0.0469286
R18025 XThC.Tn[12].n63 XThC.Tn[12] 0.0401341
R18026 XThC.Tn[12].n59 XThC.Tn[12] 0.0401341
R18027 XThC.Tn[12].n55 XThC.Tn[12] 0.0401341
R18028 XThC.Tn[12].n51 XThC.Tn[12] 0.0401341
R18029 XThC.Tn[12].n47 XThC.Tn[12] 0.0401341
R18030 XThC.Tn[12].n43 XThC.Tn[12] 0.0401341
R18031 XThC.Tn[12].n39 XThC.Tn[12] 0.0401341
R18032 XThC.Tn[12].n35 XThC.Tn[12] 0.0401341
R18033 XThC.Tn[12].n31 XThC.Tn[12] 0.0401341
R18034 XThC.Tn[12].n27 XThC.Tn[12] 0.0401341
R18035 XThC.Tn[12].n23 XThC.Tn[12] 0.0401341
R18036 XThC.Tn[12].n19 XThC.Tn[12] 0.0401341
R18037 XThC.Tn[12].n15 XThC.Tn[12] 0.0401341
R18038 XThC.Tn[12].n11 XThC.Tn[12] 0.0401341
R18039 XThC.Tn[12].n7 XThC.Tn[12] 0.0401341
R18040 XThC.Tn[12].n4 XThC.Tn[12] 0.0401341
R18041 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R18042 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R18043 XThC.Tn[1].n71 XThC.Tn[1].n69 161.365
R18044 XThC.Tn[1].n67 XThC.Tn[1].n65 161.365
R18045 XThC.Tn[1].n63 XThC.Tn[1].n61 161.365
R18046 XThC.Tn[1].n59 XThC.Tn[1].n57 161.365
R18047 XThC.Tn[1].n55 XThC.Tn[1].n53 161.365
R18048 XThC.Tn[1].n51 XThC.Tn[1].n49 161.365
R18049 XThC.Tn[1].n47 XThC.Tn[1].n45 161.365
R18050 XThC.Tn[1].n43 XThC.Tn[1].n41 161.365
R18051 XThC.Tn[1].n39 XThC.Tn[1].n37 161.365
R18052 XThC.Tn[1].n35 XThC.Tn[1].n33 161.365
R18053 XThC.Tn[1].n31 XThC.Tn[1].n29 161.365
R18054 XThC.Tn[1].n27 XThC.Tn[1].n25 161.365
R18055 XThC.Tn[1].n23 XThC.Tn[1].n21 161.365
R18056 XThC.Tn[1].n19 XThC.Tn[1].n17 161.365
R18057 XThC.Tn[1].n15 XThC.Tn[1].n13 161.365
R18058 XThC.Tn[1].n12 XThC.Tn[1].n10 161.365
R18059 XThC.Tn[1].n69 XThC.Tn[1].t20 161.106
R18060 XThC.Tn[1].n65 XThC.Tn[1].t34 161.106
R18061 XThC.Tn[1].n61 XThC.Tn[1].t31 161.106
R18062 XThC.Tn[1].n57 XThC.Tn[1].t29 161.106
R18063 XThC.Tn[1].n53 XThC.Tn[1].t42 161.106
R18064 XThC.Tn[1].n49 XThC.Tn[1].t40 161.106
R18065 XThC.Tn[1].n45 XThC.Tn[1].t28 161.106
R18066 XThC.Tn[1].n41 XThC.Tn[1].t19 161.106
R18067 XThC.Tn[1].n37 XThC.Tn[1].t17 161.106
R18068 XThC.Tn[1].n33 XThC.Tn[1].t39 161.106
R18069 XThC.Tn[1].n29 XThC.Tn[1].t26 161.106
R18070 XThC.Tn[1].n25 XThC.Tn[1].t15 161.106
R18071 XThC.Tn[1].n21 XThC.Tn[1].t38 161.106
R18072 XThC.Tn[1].n17 XThC.Tn[1].t36 161.106
R18073 XThC.Tn[1].n13 XThC.Tn[1].t23 161.106
R18074 XThC.Tn[1].n10 XThC.Tn[1].t14 161.106
R18075 XThC.Tn[1].n69 XThC.Tn[1].t16 154.679
R18076 XThC.Tn[1].n65 XThC.Tn[1].t27 154.679
R18077 XThC.Tn[1].n61 XThC.Tn[1].t25 154.679
R18078 XThC.Tn[1].n57 XThC.Tn[1].t24 154.679
R18079 XThC.Tn[1].n53 XThC.Tn[1].t37 154.679
R18080 XThC.Tn[1].n49 XThC.Tn[1].t35 154.679
R18081 XThC.Tn[1].n45 XThC.Tn[1].t22 154.679
R18082 XThC.Tn[1].n41 XThC.Tn[1].t13 154.679
R18083 XThC.Tn[1].n37 XThC.Tn[1].t12 154.679
R18084 XThC.Tn[1].n33 XThC.Tn[1].t33 154.679
R18085 XThC.Tn[1].n29 XThC.Tn[1].t21 154.679
R18086 XThC.Tn[1].n25 XThC.Tn[1].t43 154.679
R18087 XThC.Tn[1].n21 XThC.Tn[1].t32 154.679
R18088 XThC.Tn[1].n17 XThC.Tn[1].t30 154.679
R18089 XThC.Tn[1].n13 XThC.Tn[1].t18 154.679
R18090 XThC.Tn[1].n10 XThC.Tn[1].t41 154.679
R18091 XThC.Tn[1].n7 XThC.Tn[1].n6 135.249
R18092 XThC.Tn[1].n9 XThC.Tn[1].n3 98.981
R18093 XThC.Tn[1].n8 XThC.Tn[1].n4 98.981
R18094 XThC.Tn[1].n7 XThC.Tn[1].n5 98.981
R18095 XThC.Tn[1].n9 XThC.Tn[1].n8 36.2672
R18096 XThC.Tn[1].n8 XThC.Tn[1].n7 36.2672
R18097 XThC.Tn[1].n74 XThC.Tn[1].n9 32.6405
R18098 XThC.Tn[1].n1 XThC.Tn[1].t5 26.5955
R18099 XThC.Tn[1].n1 XThC.Tn[1].t4 26.5955
R18100 XThC.Tn[1].n0 XThC.Tn[1].t7 26.5955
R18101 XThC.Tn[1].n0 XThC.Tn[1].t6 26.5955
R18102 XThC.Tn[1].n3 XThC.Tn[1].t9 24.9236
R18103 XThC.Tn[1].n3 XThC.Tn[1].t8 24.9236
R18104 XThC.Tn[1].n4 XThC.Tn[1].t11 24.9236
R18105 XThC.Tn[1].n4 XThC.Tn[1].t10 24.9236
R18106 XThC.Tn[1].n5 XThC.Tn[1].t1 24.9236
R18107 XThC.Tn[1].n5 XThC.Tn[1].t0 24.9236
R18108 XThC.Tn[1].n6 XThC.Tn[1].t3 24.9236
R18109 XThC.Tn[1].n6 XThC.Tn[1].t2 24.9236
R18110 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R18111 XThC.Tn[1] XThC.Tn[1].n12 8.0245
R18112 XThC.Tn[1].n72 XThC.Tn[1].n71 7.9105
R18113 XThC.Tn[1].n68 XThC.Tn[1].n67 7.9105
R18114 XThC.Tn[1].n64 XThC.Tn[1].n63 7.9105
R18115 XThC.Tn[1].n60 XThC.Tn[1].n59 7.9105
R18116 XThC.Tn[1].n56 XThC.Tn[1].n55 7.9105
R18117 XThC.Tn[1].n52 XThC.Tn[1].n51 7.9105
R18118 XThC.Tn[1].n48 XThC.Tn[1].n47 7.9105
R18119 XThC.Tn[1].n44 XThC.Tn[1].n43 7.9105
R18120 XThC.Tn[1].n40 XThC.Tn[1].n39 7.9105
R18121 XThC.Tn[1].n36 XThC.Tn[1].n35 7.9105
R18122 XThC.Tn[1].n32 XThC.Tn[1].n31 7.9105
R18123 XThC.Tn[1].n28 XThC.Tn[1].n27 7.9105
R18124 XThC.Tn[1].n24 XThC.Tn[1].n23 7.9105
R18125 XThC.Tn[1].n20 XThC.Tn[1].n19 7.9105
R18126 XThC.Tn[1].n16 XThC.Tn[1].n15 7.9105
R18127 XThC.Tn[1] XThC.Tn[1].n74 6.7205
R18128 XThC.Tn[1].n73 XThC.Tn[1] 6.08068
R18129 XThC.Tn[1].n74 XThC.Tn[1].n73 4.65249
R18130 XThC.Tn[1].n73 XThC.Tn[1] 1.8942
R18131 XThC.Tn[1].n16 XThC.Tn[1] 0.235138
R18132 XThC.Tn[1].n20 XThC.Tn[1] 0.235138
R18133 XThC.Tn[1].n24 XThC.Tn[1] 0.235138
R18134 XThC.Tn[1].n28 XThC.Tn[1] 0.235138
R18135 XThC.Tn[1].n32 XThC.Tn[1] 0.235138
R18136 XThC.Tn[1].n36 XThC.Tn[1] 0.235138
R18137 XThC.Tn[1].n40 XThC.Tn[1] 0.235138
R18138 XThC.Tn[1].n44 XThC.Tn[1] 0.235138
R18139 XThC.Tn[1].n48 XThC.Tn[1] 0.235138
R18140 XThC.Tn[1].n52 XThC.Tn[1] 0.235138
R18141 XThC.Tn[1].n56 XThC.Tn[1] 0.235138
R18142 XThC.Tn[1].n60 XThC.Tn[1] 0.235138
R18143 XThC.Tn[1].n64 XThC.Tn[1] 0.235138
R18144 XThC.Tn[1].n68 XThC.Tn[1] 0.235138
R18145 XThC.Tn[1].n72 XThC.Tn[1] 0.235138
R18146 XThC.Tn[1] XThC.Tn[1].n16 0.114505
R18147 XThC.Tn[1] XThC.Tn[1].n20 0.114505
R18148 XThC.Tn[1] XThC.Tn[1].n24 0.114505
R18149 XThC.Tn[1] XThC.Tn[1].n28 0.114505
R18150 XThC.Tn[1] XThC.Tn[1].n32 0.114505
R18151 XThC.Tn[1] XThC.Tn[1].n36 0.114505
R18152 XThC.Tn[1] XThC.Tn[1].n40 0.114505
R18153 XThC.Tn[1] XThC.Tn[1].n44 0.114505
R18154 XThC.Tn[1] XThC.Tn[1].n48 0.114505
R18155 XThC.Tn[1] XThC.Tn[1].n52 0.114505
R18156 XThC.Tn[1] XThC.Tn[1].n56 0.114505
R18157 XThC.Tn[1] XThC.Tn[1].n60 0.114505
R18158 XThC.Tn[1] XThC.Tn[1].n64 0.114505
R18159 XThC.Tn[1] XThC.Tn[1].n68 0.114505
R18160 XThC.Tn[1] XThC.Tn[1].n72 0.114505
R18161 XThC.Tn[1].n71 XThC.Tn[1].n70 0.0599512
R18162 XThC.Tn[1].n67 XThC.Tn[1].n66 0.0599512
R18163 XThC.Tn[1].n63 XThC.Tn[1].n62 0.0599512
R18164 XThC.Tn[1].n59 XThC.Tn[1].n58 0.0599512
R18165 XThC.Tn[1].n55 XThC.Tn[1].n54 0.0599512
R18166 XThC.Tn[1].n51 XThC.Tn[1].n50 0.0599512
R18167 XThC.Tn[1].n47 XThC.Tn[1].n46 0.0599512
R18168 XThC.Tn[1].n43 XThC.Tn[1].n42 0.0599512
R18169 XThC.Tn[1].n39 XThC.Tn[1].n38 0.0599512
R18170 XThC.Tn[1].n35 XThC.Tn[1].n34 0.0599512
R18171 XThC.Tn[1].n31 XThC.Tn[1].n30 0.0599512
R18172 XThC.Tn[1].n27 XThC.Tn[1].n26 0.0599512
R18173 XThC.Tn[1].n23 XThC.Tn[1].n22 0.0599512
R18174 XThC.Tn[1].n19 XThC.Tn[1].n18 0.0599512
R18175 XThC.Tn[1].n15 XThC.Tn[1].n14 0.0599512
R18176 XThC.Tn[1].n12 XThC.Tn[1].n11 0.0599512
R18177 XThC.Tn[1].n70 XThC.Tn[1] 0.0469286
R18178 XThC.Tn[1].n66 XThC.Tn[1] 0.0469286
R18179 XThC.Tn[1].n62 XThC.Tn[1] 0.0469286
R18180 XThC.Tn[1].n58 XThC.Tn[1] 0.0469286
R18181 XThC.Tn[1].n54 XThC.Tn[1] 0.0469286
R18182 XThC.Tn[1].n50 XThC.Tn[1] 0.0469286
R18183 XThC.Tn[1].n46 XThC.Tn[1] 0.0469286
R18184 XThC.Tn[1].n42 XThC.Tn[1] 0.0469286
R18185 XThC.Tn[1].n38 XThC.Tn[1] 0.0469286
R18186 XThC.Tn[1].n34 XThC.Tn[1] 0.0469286
R18187 XThC.Tn[1].n30 XThC.Tn[1] 0.0469286
R18188 XThC.Tn[1].n26 XThC.Tn[1] 0.0469286
R18189 XThC.Tn[1].n22 XThC.Tn[1] 0.0469286
R18190 XThC.Tn[1].n18 XThC.Tn[1] 0.0469286
R18191 XThC.Tn[1].n14 XThC.Tn[1] 0.0469286
R18192 XThC.Tn[1].n11 XThC.Tn[1] 0.0469286
R18193 XThC.Tn[1].n70 XThC.Tn[1] 0.0401341
R18194 XThC.Tn[1].n66 XThC.Tn[1] 0.0401341
R18195 XThC.Tn[1].n62 XThC.Tn[1] 0.0401341
R18196 XThC.Tn[1].n58 XThC.Tn[1] 0.0401341
R18197 XThC.Tn[1].n54 XThC.Tn[1] 0.0401341
R18198 XThC.Tn[1].n50 XThC.Tn[1] 0.0401341
R18199 XThC.Tn[1].n46 XThC.Tn[1] 0.0401341
R18200 XThC.Tn[1].n42 XThC.Tn[1] 0.0401341
R18201 XThC.Tn[1].n38 XThC.Tn[1] 0.0401341
R18202 XThC.Tn[1].n34 XThC.Tn[1] 0.0401341
R18203 XThC.Tn[1].n30 XThC.Tn[1] 0.0401341
R18204 XThC.Tn[1].n26 XThC.Tn[1] 0.0401341
R18205 XThC.Tn[1].n22 XThC.Tn[1] 0.0401341
R18206 XThC.Tn[1].n18 XThC.Tn[1] 0.0401341
R18207 XThC.Tn[1].n14 XThC.Tn[1] 0.0401341
R18208 XThC.Tn[1].n11 XThC.Tn[1] 0.0401341
R18209 XThC.Tn[0].n2 XThC.Tn[0].n1 332.332
R18210 XThC.Tn[0].n2 XThC.Tn[0].n0 296.493
R18211 XThC.Tn[0].n71 XThC.Tn[0].n69 161.365
R18212 XThC.Tn[0].n67 XThC.Tn[0].n65 161.365
R18213 XThC.Tn[0].n63 XThC.Tn[0].n61 161.365
R18214 XThC.Tn[0].n59 XThC.Tn[0].n57 161.365
R18215 XThC.Tn[0].n55 XThC.Tn[0].n53 161.365
R18216 XThC.Tn[0].n51 XThC.Tn[0].n49 161.365
R18217 XThC.Tn[0].n47 XThC.Tn[0].n45 161.365
R18218 XThC.Tn[0].n43 XThC.Tn[0].n41 161.365
R18219 XThC.Tn[0].n39 XThC.Tn[0].n37 161.365
R18220 XThC.Tn[0].n35 XThC.Tn[0].n33 161.365
R18221 XThC.Tn[0].n31 XThC.Tn[0].n29 161.365
R18222 XThC.Tn[0].n27 XThC.Tn[0].n25 161.365
R18223 XThC.Tn[0].n23 XThC.Tn[0].n21 161.365
R18224 XThC.Tn[0].n19 XThC.Tn[0].n17 161.365
R18225 XThC.Tn[0].n15 XThC.Tn[0].n13 161.365
R18226 XThC.Tn[0].n12 XThC.Tn[0].n10 161.365
R18227 XThC.Tn[0].n69 XThC.Tn[0].t20 161.106
R18228 XThC.Tn[0].n65 XThC.Tn[0].t32 161.106
R18229 XThC.Tn[0].n61 XThC.Tn[0].t30 161.106
R18230 XThC.Tn[0].n57 XThC.Tn[0].t28 161.106
R18231 XThC.Tn[0].n53 XThC.Tn[0].t41 161.106
R18232 XThC.Tn[0].n49 XThC.Tn[0].t39 161.106
R18233 XThC.Tn[0].n45 XThC.Tn[0].t26 161.106
R18234 XThC.Tn[0].n41 XThC.Tn[0].t18 161.106
R18235 XThC.Tn[0].n37 XThC.Tn[0].t16 161.106
R18236 XThC.Tn[0].n33 XThC.Tn[0].t36 161.106
R18237 XThC.Tn[0].n29 XThC.Tn[0].t25 161.106
R18238 XThC.Tn[0].n25 XThC.Tn[0].t15 161.106
R18239 XThC.Tn[0].n21 XThC.Tn[0].t35 161.106
R18240 XThC.Tn[0].n17 XThC.Tn[0].t33 161.106
R18241 XThC.Tn[0].n13 XThC.Tn[0].t21 161.106
R18242 XThC.Tn[0].n10 XThC.Tn[0].t12 161.106
R18243 XThC.Tn[0].n69 XThC.Tn[0].t29 154.679
R18244 XThC.Tn[0].n65 XThC.Tn[0].t42 154.679
R18245 XThC.Tn[0].n61 XThC.Tn[0].t40 154.679
R18246 XThC.Tn[0].n57 XThC.Tn[0].t38 154.679
R18247 XThC.Tn[0].n53 XThC.Tn[0].t19 154.679
R18248 XThC.Tn[0].n49 XThC.Tn[0].t17 154.679
R18249 XThC.Tn[0].n45 XThC.Tn[0].t37 154.679
R18250 XThC.Tn[0].n41 XThC.Tn[0].t27 154.679
R18251 XThC.Tn[0].n37 XThC.Tn[0].t24 154.679
R18252 XThC.Tn[0].n33 XThC.Tn[0].t14 154.679
R18253 XThC.Tn[0].n29 XThC.Tn[0].t34 154.679
R18254 XThC.Tn[0].n25 XThC.Tn[0].t23 154.679
R18255 XThC.Tn[0].n21 XThC.Tn[0].t13 154.679
R18256 XThC.Tn[0].n17 XThC.Tn[0].t43 154.679
R18257 XThC.Tn[0].n13 XThC.Tn[0].t31 154.679
R18258 XThC.Tn[0].n10 XThC.Tn[0].t22 154.679
R18259 XThC.Tn[0].n7 XThC.Tn[0].n6 135.248
R18260 XThC.Tn[0].n9 XThC.Tn[0].n3 98.982
R18261 XThC.Tn[0].n8 XThC.Tn[0].n4 98.982
R18262 XThC.Tn[0].n7 XThC.Tn[0].n5 98.982
R18263 XThC.Tn[0].n9 XThC.Tn[0].n8 36.2672
R18264 XThC.Tn[0].n8 XThC.Tn[0].n7 36.2672
R18265 XThC.Tn[0].n74 XThC.Tn[0].n9 32.6405
R18266 XThC.Tn[0].n1 XThC.Tn[0].t10 26.5955
R18267 XThC.Tn[0].n1 XThC.Tn[0].t9 26.5955
R18268 XThC.Tn[0].n0 XThC.Tn[0].t8 26.5955
R18269 XThC.Tn[0].n0 XThC.Tn[0].t7 26.5955
R18270 XThC.Tn[0].n3 XThC.Tn[0].t4 24.9236
R18271 XThC.Tn[0].n3 XThC.Tn[0].t3 24.9236
R18272 XThC.Tn[0].n4 XThC.Tn[0].t6 24.9236
R18273 XThC.Tn[0].n4 XThC.Tn[0].t5 24.9236
R18274 XThC.Tn[0].n5 XThC.Tn[0].t1 24.9236
R18275 XThC.Tn[0].n5 XThC.Tn[0].t2 24.9236
R18276 XThC.Tn[0].n6 XThC.Tn[0].t11 24.9236
R18277 XThC.Tn[0].n6 XThC.Tn[0].t0 24.9236
R18278 XThC.Tn[0].n75 XThC.Tn[0].n2 18.5605
R18279 XThC.Tn[0].n75 XThC.Tn[0].n74 11.5205
R18280 XThC.Tn[0] XThC.Tn[0].n12 8.0245
R18281 XThC.Tn[0].n72 XThC.Tn[0].n71 7.9105
R18282 XThC.Tn[0].n68 XThC.Tn[0].n67 7.9105
R18283 XThC.Tn[0].n64 XThC.Tn[0].n63 7.9105
R18284 XThC.Tn[0].n60 XThC.Tn[0].n59 7.9105
R18285 XThC.Tn[0].n56 XThC.Tn[0].n55 7.9105
R18286 XThC.Tn[0].n52 XThC.Tn[0].n51 7.9105
R18287 XThC.Tn[0].n48 XThC.Tn[0].n47 7.9105
R18288 XThC.Tn[0].n44 XThC.Tn[0].n43 7.9105
R18289 XThC.Tn[0].n40 XThC.Tn[0].n39 7.9105
R18290 XThC.Tn[0].n36 XThC.Tn[0].n35 7.9105
R18291 XThC.Tn[0].n32 XThC.Tn[0].n31 7.9105
R18292 XThC.Tn[0].n28 XThC.Tn[0].n27 7.9105
R18293 XThC.Tn[0].n24 XThC.Tn[0].n23 7.9105
R18294 XThC.Tn[0].n20 XThC.Tn[0].n19 7.9105
R18295 XThC.Tn[0].n16 XThC.Tn[0].n15 7.9105
R18296 XThC.Tn[0].n73 XThC.Tn[0] 5.95611
R18297 XThC.Tn[0].n74 XThC.Tn[0].n73 4.6005
R18298 XThC.Tn[0].n73 XThC.Tn[0] 1.89022
R18299 XThC.Tn[0] XThC.Tn[0].n75 0.6405
R18300 XThC.Tn[0].n16 XThC.Tn[0] 0.235138
R18301 XThC.Tn[0].n20 XThC.Tn[0] 0.235138
R18302 XThC.Tn[0].n24 XThC.Tn[0] 0.235138
R18303 XThC.Tn[0].n28 XThC.Tn[0] 0.235138
R18304 XThC.Tn[0].n32 XThC.Tn[0] 0.235138
R18305 XThC.Tn[0].n36 XThC.Tn[0] 0.235138
R18306 XThC.Tn[0].n40 XThC.Tn[0] 0.235138
R18307 XThC.Tn[0].n44 XThC.Tn[0] 0.235138
R18308 XThC.Tn[0].n48 XThC.Tn[0] 0.235138
R18309 XThC.Tn[0].n52 XThC.Tn[0] 0.235138
R18310 XThC.Tn[0].n56 XThC.Tn[0] 0.235138
R18311 XThC.Tn[0].n60 XThC.Tn[0] 0.235138
R18312 XThC.Tn[0].n64 XThC.Tn[0] 0.235138
R18313 XThC.Tn[0].n68 XThC.Tn[0] 0.235138
R18314 XThC.Tn[0].n72 XThC.Tn[0] 0.235138
R18315 XThC.Tn[0] XThC.Tn[0].n16 0.114505
R18316 XThC.Tn[0] XThC.Tn[0].n20 0.114505
R18317 XThC.Tn[0] XThC.Tn[0].n24 0.114505
R18318 XThC.Tn[0] XThC.Tn[0].n28 0.114505
R18319 XThC.Tn[0] XThC.Tn[0].n32 0.114505
R18320 XThC.Tn[0] XThC.Tn[0].n36 0.114505
R18321 XThC.Tn[0] XThC.Tn[0].n40 0.114505
R18322 XThC.Tn[0] XThC.Tn[0].n44 0.114505
R18323 XThC.Tn[0] XThC.Tn[0].n48 0.114505
R18324 XThC.Tn[0] XThC.Tn[0].n52 0.114505
R18325 XThC.Tn[0] XThC.Tn[0].n56 0.114505
R18326 XThC.Tn[0] XThC.Tn[0].n60 0.114505
R18327 XThC.Tn[0] XThC.Tn[0].n64 0.114505
R18328 XThC.Tn[0] XThC.Tn[0].n68 0.114505
R18329 XThC.Tn[0] XThC.Tn[0].n72 0.114505
R18330 XThC.Tn[0].n71 XThC.Tn[0].n70 0.0599512
R18331 XThC.Tn[0].n67 XThC.Tn[0].n66 0.0599512
R18332 XThC.Tn[0].n63 XThC.Tn[0].n62 0.0599512
R18333 XThC.Tn[0].n59 XThC.Tn[0].n58 0.0599512
R18334 XThC.Tn[0].n55 XThC.Tn[0].n54 0.0599512
R18335 XThC.Tn[0].n51 XThC.Tn[0].n50 0.0599512
R18336 XThC.Tn[0].n47 XThC.Tn[0].n46 0.0599512
R18337 XThC.Tn[0].n43 XThC.Tn[0].n42 0.0599512
R18338 XThC.Tn[0].n39 XThC.Tn[0].n38 0.0599512
R18339 XThC.Tn[0].n35 XThC.Tn[0].n34 0.0599512
R18340 XThC.Tn[0].n31 XThC.Tn[0].n30 0.0599512
R18341 XThC.Tn[0].n27 XThC.Tn[0].n26 0.0599512
R18342 XThC.Tn[0].n23 XThC.Tn[0].n22 0.0599512
R18343 XThC.Tn[0].n19 XThC.Tn[0].n18 0.0599512
R18344 XThC.Tn[0].n15 XThC.Tn[0].n14 0.0599512
R18345 XThC.Tn[0].n12 XThC.Tn[0].n11 0.0599512
R18346 XThC.Tn[0].n70 XThC.Tn[0] 0.0469286
R18347 XThC.Tn[0].n66 XThC.Tn[0] 0.0469286
R18348 XThC.Tn[0].n62 XThC.Tn[0] 0.0469286
R18349 XThC.Tn[0].n58 XThC.Tn[0] 0.0469286
R18350 XThC.Tn[0].n54 XThC.Tn[0] 0.0469286
R18351 XThC.Tn[0].n50 XThC.Tn[0] 0.0469286
R18352 XThC.Tn[0].n46 XThC.Tn[0] 0.0469286
R18353 XThC.Tn[0].n42 XThC.Tn[0] 0.0469286
R18354 XThC.Tn[0].n38 XThC.Tn[0] 0.0469286
R18355 XThC.Tn[0].n34 XThC.Tn[0] 0.0469286
R18356 XThC.Tn[0].n30 XThC.Tn[0] 0.0469286
R18357 XThC.Tn[0].n26 XThC.Tn[0] 0.0469286
R18358 XThC.Tn[0].n22 XThC.Tn[0] 0.0469286
R18359 XThC.Tn[0].n18 XThC.Tn[0] 0.0469286
R18360 XThC.Tn[0].n14 XThC.Tn[0] 0.0469286
R18361 XThC.Tn[0].n11 XThC.Tn[0] 0.0469286
R18362 XThC.Tn[0].n70 XThC.Tn[0] 0.0401341
R18363 XThC.Tn[0].n66 XThC.Tn[0] 0.0401341
R18364 XThC.Tn[0].n62 XThC.Tn[0] 0.0401341
R18365 XThC.Tn[0].n58 XThC.Tn[0] 0.0401341
R18366 XThC.Tn[0].n54 XThC.Tn[0] 0.0401341
R18367 XThC.Tn[0].n50 XThC.Tn[0] 0.0401341
R18368 XThC.Tn[0].n46 XThC.Tn[0] 0.0401341
R18369 XThC.Tn[0].n42 XThC.Tn[0] 0.0401341
R18370 XThC.Tn[0].n38 XThC.Tn[0] 0.0401341
R18371 XThC.Tn[0].n34 XThC.Tn[0] 0.0401341
R18372 XThC.Tn[0].n30 XThC.Tn[0] 0.0401341
R18373 XThC.Tn[0].n26 XThC.Tn[0] 0.0401341
R18374 XThC.Tn[0].n22 XThC.Tn[0] 0.0401341
R18375 XThC.Tn[0].n18 XThC.Tn[0] 0.0401341
R18376 XThC.Tn[0].n14 XThC.Tn[0] 0.0401341
R18377 XThC.Tn[0].n11 XThC.Tn[0] 0.0401341
R18378 XThC.XTB4.Y.n21 XThC.XTB4.Y.t0 235.56
R18379 XThC.XTB4.Y.n3 XThC.XTB4.Y.t3 212.081
R18380 XThC.XTB4.Y.n2 XThC.XTB4.Y.t2 212.081
R18381 XThC.XTB4.Y.n8 XThC.XTB4.Y.t17 212.081
R18382 XThC.XTB4.Y.n0 XThC.XTB4.Y.t13 212.081
R18383 XThC.XTB4.Y.n12 XThC.XTB4.Y.t8 212.081
R18384 XThC.XTB4.Y.n13 XThC.XTB4.Y.t12 212.081
R18385 XThC.XTB4.Y.n15 XThC.XTB4.Y.t6 212.081
R18386 XThC.XTB4.Y.n11 XThC.XTB4.Y.t16 212.081
R18387 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 173.761
R18388 XThC.XTB4.Y.n14 XThC.XTB4.Y 158.656
R18389 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 152
R18390 XThC.XTB4.Y.n5 XThC.XTB4.Y.n1 152
R18391 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 152
R18392 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 152
R18393 XThC.XTB4.Y.n3 XThC.XTB4.Y.t14 139.78
R18394 XThC.XTB4.Y.n2 XThC.XTB4.Y.t10 139.78
R18395 XThC.XTB4.Y.n8 XThC.XTB4.Y.t7 139.78
R18396 XThC.XTB4.Y.n0 XThC.XTB4.Y.t4 139.78
R18397 XThC.XTB4.Y.n12 XThC.XTB4.Y.t11 139.78
R18398 XThC.XTB4.Y.n13 XThC.XTB4.Y.t15 139.78
R18399 XThC.XTB4.Y.n15 XThC.XTB4.Y.t9 139.78
R18400 XThC.XTB4.Y.n11 XThC.XTB4.Y.t5 139.78
R18401 XThC.XTB4.Y.n20 XThC.XTB4.Y.t1 133.386
R18402 XThC.XTB4.Y.n19 XThC.XTB4.Y.n10 72.9296
R18403 XThC.XTB4.Y.n13 XThC.XTB4.Y.n12 61.346
R18404 XThC.XTB4.Y.n7 XThC.XTB4.Y.n1 49.6611
R18405 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 45.2793
R18406 XThC.XTB4.Y.n4 XThC.XTB4.Y.n2 42.3581
R18407 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 38.1854
R18408 XThC.XTB4.Y.n16 XThC.XTB4.Y.n11 30.6732
R18409 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R18410 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R18411 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 30.6732
R18412 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 21.7605
R18413 XThC.XTB4.Y XThC.XTB4.Y.n20 19.5051
R18414 XThC.XTB4.Y.n4 XThC.XTB4.Y.n3 18.9884
R18415 XThC.XTB4.Y.n9 XThC.XTB4.Y.n0 16.0672
R18416 XThC.XTB4.Y.n17 XThC.XTB4.Y 14.7905
R18417 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 11.994
R18418 XThC.XTB4.Y.n10 XThC.XTB4.Y 11.5205
R18419 XThC.XTB4.Y.n6 XThC.XTB4.Y 10.2405
R18420 XThC.XTB4.Y.n2 XThC.XTB4.Y.n1 7.30353
R18421 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 7.24578
R18422 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 4.38232
R18423 XThC.XTB4.Y.n21 XThC.XTB4.Y 2.22659
R18424 XThC.XTB4.Y XThC.XTB4.Y.n21 1.55202
R18425 XThC.XTB4.Y.n18 XThC.XTB4.Y 0.966538
R18426 XThR.Tn[5].n88 XThR.Tn[5].n87 332.332
R18427 XThR.Tn[5].n88 XThR.Tn[5].n86 296.493
R18428 XThR.Tn[5] XThR.Tn[5].n79 161.363
R18429 XThR.Tn[5] XThR.Tn[5].n74 161.363
R18430 XThR.Tn[5] XThR.Tn[5].n69 161.363
R18431 XThR.Tn[5] XThR.Tn[5].n64 161.363
R18432 XThR.Tn[5] XThR.Tn[5].n59 161.363
R18433 XThR.Tn[5] XThR.Tn[5].n54 161.363
R18434 XThR.Tn[5] XThR.Tn[5].n49 161.363
R18435 XThR.Tn[5] XThR.Tn[5].n44 161.363
R18436 XThR.Tn[5] XThR.Tn[5].n39 161.363
R18437 XThR.Tn[5] XThR.Tn[5].n34 161.363
R18438 XThR.Tn[5] XThR.Tn[5].n29 161.363
R18439 XThR.Tn[5] XThR.Tn[5].n24 161.363
R18440 XThR.Tn[5] XThR.Tn[5].n19 161.363
R18441 XThR.Tn[5] XThR.Tn[5].n14 161.363
R18442 XThR.Tn[5] XThR.Tn[5].n9 161.363
R18443 XThR.Tn[5] XThR.Tn[5].n7 161.363
R18444 XThR.Tn[5].n81 XThR.Tn[5].n80 161.3
R18445 XThR.Tn[5].n76 XThR.Tn[5].n75 161.3
R18446 XThR.Tn[5].n71 XThR.Tn[5].n70 161.3
R18447 XThR.Tn[5].n66 XThR.Tn[5].n65 161.3
R18448 XThR.Tn[5].n61 XThR.Tn[5].n60 161.3
R18449 XThR.Tn[5].n56 XThR.Tn[5].n55 161.3
R18450 XThR.Tn[5].n51 XThR.Tn[5].n50 161.3
R18451 XThR.Tn[5].n46 XThR.Tn[5].n45 161.3
R18452 XThR.Tn[5].n41 XThR.Tn[5].n40 161.3
R18453 XThR.Tn[5].n36 XThR.Tn[5].n35 161.3
R18454 XThR.Tn[5].n31 XThR.Tn[5].n30 161.3
R18455 XThR.Tn[5].n26 XThR.Tn[5].n25 161.3
R18456 XThR.Tn[5].n21 XThR.Tn[5].n20 161.3
R18457 XThR.Tn[5].n16 XThR.Tn[5].n15 161.3
R18458 XThR.Tn[5].n11 XThR.Tn[5].n10 161.3
R18459 XThR.Tn[5].n80 XThR.Tn[5].t39 161.106
R18460 XThR.Tn[5].n79 XThR.Tn[5].t60 161.106
R18461 XThR.Tn[5].n75 XThR.Tn[5].t45 161.106
R18462 XThR.Tn[5].n74 XThR.Tn[5].t68 161.106
R18463 XThR.Tn[5].n70 XThR.Tn[5].t28 161.106
R18464 XThR.Tn[5].n69 XThR.Tn[5].t50 161.106
R18465 XThR.Tn[5].n65 XThR.Tn[5].t73 161.106
R18466 XThR.Tn[5].n64 XThR.Tn[5].t31 161.106
R18467 XThR.Tn[5].n60 XThR.Tn[5].t37 161.106
R18468 XThR.Tn[5].n59 XThR.Tn[5].t57 161.106
R18469 XThR.Tn[5].n55 XThR.Tn[5].t62 161.106
R18470 XThR.Tn[5].n54 XThR.Tn[5].t22 161.106
R18471 XThR.Tn[5].n50 XThR.Tn[5].t43 161.106
R18472 XThR.Tn[5].n49 XThR.Tn[5].t65 161.106
R18473 XThR.Tn[5].n45 XThR.Tn[5].t25 161.106
R18474 XThR.Tn[5].n44 XThR.Tn[5].t47 161.106
R18475 XThR.Tn[5].n40 XThR.Tn[5].t71 161.106
R18476 XThR.Tn[5].n39 XThR.Tn[5].t30 161.106
R18477 XThR.Tn[5].n35 XThR.Tn[5].t14 161.106
R18478 XThR.Tn[5].n34 XThR.Tn[5].t35 161.106
R18479 XThR.Tn[5].n30 XThR.Tn[5].t61 161.106
R18480 XThR.Tn[5].n29 XThR.Tn[5].t21 161.106
R18481 XThR.Tn[5].n25 XThR.Tn[5].t27 161.106
R18482 XThR.Tn[5].n24 XThR.Tn[5].t49 161.106
R18483 XThR.Tn[5].n20 XThR.Tn[5].t58 161.106
R18484 XThR.Tn[5].n19 XThR.Tn[5].t19 161.106
R18485 XThR.Tn[5].n15 XThR.Tn[5].t41 161.106
R18486 XThR.Tn[5].n14 XThR.Tn[5].t64 161.106
R18487 XThR.Tn[5].n10 XThR.Tn[5].t66 161.106
R18488 XThR.Tn[5].n9 XThR.Tn[5].t24 161.106
R18489 XThR.Tn[5].n7 XThR.Tn[5].t70 161.106
R18490 XThR.Tn[5].n80 XThR.Tn[5].t56 154.679
R18491 XThR.Tn[5].n79 XThR.Tn[5].t16 154.679
R18492 XThR.Tn[5].n75 XThR.Tn[5].t33 154.679
R18493 XThR.Tn[5].n74 XThR.Tn[5].t54 154.679
R18494 XThR.Tn[5].n70 XThR.Tn[5].t17 154.679
R18495 XThR.Tn[5].n69 XThR.Tn[5].t38 154.679
R18496 XThR.Tn[5].n65 XThR.Tn[5].t46 154.679
R18497 XThR.Tn[5].n64 XThR.Tn[5].t69 154.679
R18498 XThR.Tn[5].n60 XThR.Tn[5].t29 154.679
R18499 XThR.Tn[5].n59 XThR.Tn[5].t51 154.679
R18500 XThR.Tn[5].n55 XThR.Tn[5].t55 154.679
R18501 XThR.Tn[5].n54 XThR.Tn[5].t12 154.679
R18502 XThR.Tn[5].n50 XThR.Tn[5].t18 154.679
R18503 XThR.Tn[5].n49 XThR.Tn[5].t40 154.679
R18504 XThR.Tn[5].n45 XThR.Tn[5].t63 154.679
R18505 XThR.Tn[5].n44 XThR.Tn[5].t23 154.679
R18506 XThR.Tn[5].n40 XThR.Tn[5].t44 154.679
R18507 XThR.Tn[5].n39 XThR.Tn[5].t67 154.679
R18508 XThR.Tn[5].n35 XThR.Tn[5].t26 154.679
R18509 XThR.Tn[5].n34 XThR.Tn[5].t48 154.679
R18510 XThR.Tn[5].n30 XThR.Tn[5].t32 154.679
R18511 XThR.Tn[5].n29 XThR.Tn[5].t53 154.679
R18512 XThR.Tn[5].n25 XThR.Tn[5].t15 154.679
R18513 XThR.Tn[5].n24 XThR.Tn[5].t36 154.679
R18514 XThR.Tn[5].n20 XThR.Tn[5].t52 154.679
R18515 XThR.Tn[5].n19 XThR.Tn[5].t72 154.679
R18516 XThR.Tn[5].n15 XThR.Tn[5].t13 154.679
R18517 XThR.Tn[5].n14 XThR.Tn[5].t34 154.679
R18518 XThR.Tn[5].n10 XThR.Tn[5].t59 154.679
R18519 XThR.Tn[5].n9 XThR.Tn[5].t20 154.679
R18520 XThR.Tn[5].n7 XThR.Tn[5].t42 154.679
R18521 XThR.Tn[5].n2 XThR.Tn[5].n0 135.249
R18522 XThR.Tn[5].n2 XThR.Tn[5].n1 98.981
R18523 XThR.Tn[5].n4 XThR.Tn[5].n3 98.981
R18524 XThR.Tn[5].n6 XThR.Tn[5].n5 98.981
R18525 XThR.Tn[5].n4 XThR.Tn[5].n2 36.2672
R18526 XThR.Tn[5].n6 XThR.Tn[5].n4 36.2672
R18527 XThR.Tn[5].n85 XThR.Tn[5].n6 32.6405
R18528 XThR.Tn[5].n87 XThR.Tn[5].t1 26.5955
R18529 XThR.Tn[5].n87 XThR.Tn[5].t0 26.5955
R18530 XThR.Tn[5].n86 XThR.Tn[5].t2 26.5955
R18531 XThR.Tn[5].n86 XThR.Tn[5].t3 26.5955
R18532 XThR.Tn[5].n0 XThR.Tn[5].t8 24.9236
R18533 XThR.Tn[5].n0 XThR.Tn[5].t9 24.9236
R18534 XThR.Tn[5].n1 XThR.Tn[5].t11 24.9236
R18535 XThR.Tn[5].n1 XThR.Tn[5].t10 24.9236
R18536 XThR.Tn[5].n3 XThR.Tn[5].t6 24.9236
R18537 XThR.Tn[5].n3 XThR.Tn[5].t5 24.9236
R18538 XThR.Tn[5].n5 XThR.Tn[5].t7 24.9236
R18539 XThR.Tn[5].n5 XThR.Tn[5].t4 24.9236
R18540 XThR.Tn[5].n89 XThR.Tn[5].n88 18.5605
R18541 XThR.Tn[5].n89 XThR.Tn[5].n85 11.5205
R18542 XThR.Tn[5].n85 XThR.Tn[5] 5.71508
R18543 XThR.Tn[5] XThR.Tn[5].n8 5.34871
R18544 XThR.Tn[5].n13 XThR.Tn[5].n12 4.5005
R18545 XThR.Tn[5].n18 XThR.Tn[5].n17 4.5005
R18546 XThR.Tn[5].n23 XThR.Tn[5].n22 4.5005
R18547 XThR.Tn[5].n28 XThR.Tn[5].n27 4.5005
R18548 XThR.Tn[5].n33 XThR.Tn[5].n32 4.5005
R18549 XThR.Tn[5].n38 XThR.Tn[5].n37 4.5005
R18550 XThR.Tn[5].n43 XThR.Tn[5].n42 4.5005
R18551 XThR.Tn[5].n48 XThR.Tn[5].n47 4.5005
R18552 XThR.Tn[5].n53 XThR.Tn[5].n52 4.5005
R18553 XThR.Tn[5].n58 XThR.Tn[5].n57 4.5005
R18554 XThR.Tn[5].n63 XThR.Tn[5].n62 4.5005
R18555 XThR.Tn[5].n68 XThR.Tn[5].n67 4.5005
R18556 XThR.Tn[5].n73 XThR.Tn[5].n72 4.5005
R18557 XThR.Tn[5].n78 XThR.Tn[5].n77 4.5005
R18558 XThR.Tn[5].n83 XThR.Tn[5].n82 4.5005
R18559 XThR.Tn[5].n84 XThR.Tn[5] 3.70586
R18560 XThR.Tn[5].n13 XThR.Tn[5] 2.51836
R18561 XThR.Tn[5].n18 XThR.Tn[5] 2.51836
R18562 XThR.Tn[5].n23 XThR.Tn[5] 2.51836
R18563 XThR.Tn[5].n28 XThR.Tn[5] 2.51836
R18564 XThR.Tn[5].n33 XThR.Tn[5] 2.51836
R18565 XThR.Tn[5].n38 XThR.Tn[5] 2.51836
R18566 XThR.Tn[5].n43 XThR.Tn[5] 2.51836
R18567 XThR.Tn[5].n48 XThR.Tn[5] 2.51836
R18568 XThR.Tn[5].n53 XThR.Tn[5] 2.51836
R18569 XThR.Tn[5].n58 XThR.Tn[5] 2.51836
R18570 XThR.Tn[5].n63 XThR.Tn[5] 2.51836
R18571 XThR.Tn[5].n68 XThR.Tn[5] 2.51836
R18572 XThR.Tn[5].n73 XThR.Tn[5] 2.51836
R18573 XThR.Tn[5].n78 XThR.Tn[5] 2.51836
R18574 XThR.Tn[5].n83 XThR.Tn[5] 2.51836
R18575 XThR.Tn[5] XThR.Tn[5].n13 0.848714
R18576 XThR.Tn[5] XThR.Tn[5].n18 0.848714
R18577 XThR.Tn[5] XThR.Tn[5].n23 0.848714
R18578 XThR.Tn[5] XThR.Tn[5].n28 0.848714
R18579 XThR.Tn[5] XThR.Tn[5].n33 0.848714
R18580 XThR.Tn[5] XThR.Tn[5].n38 0.848714
R18581 XThR.Tn[5] XThR.Tn[5].n43 0.848714
R18582 XThR.Tn[5] XThR.Tn[5].n48 0.848714
R18583 XThR.Tn[5] XThR.Tn[5].n53 0.848714
R18584 XThR.Tn[5] XThR.Tn[5].n58 0.848714
R18585 XThR.Tn[5] XThR.Tn[5].n63 0.848714
R18586 XThR.Tn[5] XThR.Tn[5].n68 0.848714
R18587 XThR.Tn[5] XThR.Tn[5].n73 0.848714
R18588 XThR.Tn[5] XThR.Tn[5].n78 0.848714
R18589 XThR.Tn[5] XThR.Tn[5].n83 0.848714
R18590 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R18591 XThR.Tn[5].n8 XThR.Tn[5] 0.485653
R18592 XThR.Tn[5].n81 XThR.Tn[5] 0.21482
R18593 XThR.Tn[5].n76 XThR.Tn[5] 0.21482
R18594 XThR.Tn[5].n71 XThR.Tn[5] 0.21482
R18595 XThR.Tn[5].n66 XThR.Tn[5] 0.21482
R18596 XThR.Tn[5].n61 XThR.Tn[5] 0.21482
R18597 XThR.Tn[5].n56 XThR.Tn[5] 0.21482
R18598 XThR.Tn[5].n51 XThR.Tn[5] 0.21482
R18599 XThR.Tn[5].n46 XThR.Tn[5] 0.21482
R18600 XThR.Tn[5].n41 XThR.Tn[5] 0.21482
R18601 XThR.Tn[5].n36 XThR.Tn[5] 0.21482
R18602 XThR.Tn[5].n31 XThR.Tn[5] 0.21482
R18603 XThR.Tn[5].n26 XThR.Tn[5] 0.21482
R18604 XThR.Tn[5].n21 XThR.Tn[5] 0.21482
R18605 XThR.Tn[5].n16 XThR.Tn[5] 0.21482
R18606 XThR.Tn[5].n11 XThR.Tn[5] 0.21482
R18607 XThR.Tn[5].n82 XThR.Tn[5] 0.0608448
R18608 XThR.Tn[5].n77 XThR.Tn[5] 0.0608448
R18609 XThR.Tn[5].n72 XThR.Tn[5] 0.0608448
R18610 XThR.Tn[5].n67 XThR.Tn[5] 0.0608448
R18611 XThR.Tn[5].n62 XThR.Tn[5] 0.0608448
R18612 XThR.Tn[5].n57 XThR.Tn[5] 0.0608448
R18613 XThR.Tn[5].n52 XThR.Tn[5] 0.0608448
R18614 XThR.Tn[5].n47 XThR.Tn[5] 0.0608448
R18615 XThR.Tn[5].n42 XThR.Tn[5] 0.0608448
R18616 XThR.Tn[5].n37 XThR.Tn[5] 0.0608448
R18617 XThR.Tn[5].n32 XThR.Tn[5] 0.0608448
R18618 XThR.Tn[5].n27 XThR.Tn[5] 0.0608448
R18619 XThR.Tn[5].n22 XThR.Tn[5] 0.0608448
R18620 XThR.Tn[5].n17 XThR.Tn[5] 0.0608448
R18621 XThR.Tn[5].n12 XThR.Tn[5] 0.0608448
R18622 XThR.Tn[5].n84 XThR.Tn[5] 0.0540714
R18623 XThR.Tn[5] XThR.Tn[5].n84 0.038
R18624 XThR.Tn[5].n8 XThR.Tn[5] 0.00744444
R18625 XThR.Tn[5].n82 XThR.Tn[5].n81 0.00265517
R18626 XThR.Tn[5].n77 XThR.Tn[5].n76 0.00265517
R18627 XThR.Tn[5].n72 XThR.Tn[5].n71 0.00265517
R18628 XThR.Tn[5].n67 XThR.Tn[5].n66 0.00265517
R18629 XThR.Tn[5].n62 XThR.Tn[5].n61 0.00265517
R18630 XThR.Tn[5].n57 XThR.Tn[5].n56 0.00265517
R18631 XThR.Tn[5].n52 XThR.Tn[5].n51 0.00265517
R18632 XThR.Tn[5].n47 XThR.Tn[5].n46 0.00265517
R18633 XThR.Tn[5].n42 XThR.Tn[5].n41 0.00265517
R18634 XThR.Tn[5].n37 XThR.Tn[5].n36 0.00265517
R18635 XThR.Tn[5].n32 XThR.Tn[5].n31 0.00265517
R18636 XThR.Tn[5].n27 XThR.Tn[5].n26 0.00265517
R18637 XThR.Tn[5].n22 XThR.Tn[5].n21 0.00265517
R18638 XThR.Tn[5].n17 XThR.Tn[5].n16 0.00265517
R18639 XThR.Tn[5].n12 XThR.Tn[5].n11 0.00265517
R18640 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R18641 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R18642 XThC.Tn[2].n71 XThC.Tn[2].n69 161.365
R18643 XThC.Tn[2].n67 XThC.Tn[2].n65 161.365
R18644 XThC.Tn[2].n63 XThC.Tn[2].n61 161.365
R18645 XThC.Tn[2].n59 XThC.Tn[2].n57 161.365
R18646 XThC.Tn[2].n55 XThC.Tn[2].n53 161.365
R18647 XThC.Tn[2].n51 XThC.Tn[2].n49 161.365
R18648 XThC.Tn[2].n47 XThC.Tn[2].n45 161.365
R18649 XThC.Tn[2].n43 XThC.Tn[2].n41 161.365
R18650 XThC.Tn[2].n39 XThC.Tn[2].n37 161.365
R18651 XThC.Tn[2].n35 XThC.Tn[2].n33 161.365
R18652 XThC.Tn[2].n31 XThC.Tn[2].n29 161.365
R18653 XThC.Tn[2].n27 XThC.Tn[2].n25 161.365
R18654 XThC.Tn[2].n23 XThC.Tn[2].n21 161.365
R18655 XThC.Tn[2].n19 XThC.Tn[2].n17 161.365
R18656 XThC.Tn[2].n15 XThC.Tn[2].n13 161.365
R18657 XThC.Tn[2].n12 XThC.Tn[2].n10 161.365
R18658 XThC.Tn[2].n69 XThC.Tn[2].t12 161.106
R18659 XThC.Tn[2].n65 XThC.Tn[2].t26 161.106
R18660 XThC.Tn[2].n61 XThC.Tn[2].t23 161.106
R18661 XThC.Tn[2].n57 XThC.Tn[2].t21 161.106
R18662 XThC.Tn[2].n53 XThC.Tn[2].t34 161.106
R18663 XThC.Tn[2].n49 XThC.Tn[2].t32 161.106
R18664 XThC.Tn[2].n45 XThC.Tn[2].t20 161.106
R18665 XThC.Tn[2].n41 XThC.Tn[2].t43 161.106
R18666 XThC.Tn[2].n37 XThC.Tn[2].t41 161.106
R18667 XThC.Tn[2].n33 XThC.Tn[2].t31 161.106
R18668 XThC.Tn[2].n29 XThC.Tn[2].t18 161.106
R18669 XThC.Tn[2].n25 XThC.Tn[2].t39 161.106
R18670 XThC.Tn[2].n21 XThC.Tn[2].t30 161.106
R18671 XThC.Tn[2].n17 XThC.Tn[2].t28 161.106
R18672 XThC.Tn[2].n13 XThC.Tn[2].t15 161.106
R18673 XThC.Tn[2].n10 XThC.Tn[2].t38 161.106
R18674 XThC.Tn[2].n69 XThC.Tn[2].t40 154.679
R18675 XThC.Tn[2].n65 XThC.Tn[2].t19 154.679
R18676 XThC.Tn[2].n61 XThC.Tn[2].t17 154.679
R18677 XThC.Tn[2].n57 XThC.Tn[2].t16 154.679
R18678 XThC.Tn[2].n53 XThC.Tn[2].t29 154.679
R18679 XThC.Tn[2].n49 XThC.Tn[2].t27 154.679
R18680 XThC.Tn[2].n45 XThC.Tn[2].t14 154.679
R18681 XThC.Tn[2].n41 XThC.Tn[2].t37 154.679
R18682 XThC.Tn[2].n37 XThC.Tn[2].t36 154.679
R18683 XThC.Tn[2].n33 XThC.Tn[2].t25 154.679
R18684 XThC.Tn[2].n29 XThC.Tn[2].t13 154.679
R18685 XThC.Tn[2].n25 XThC.Tn[2].t35 154.679
R18686 XThC.Tn[2].n21 XThC.Tn[2].t24 154.679
R18687 XThC.Tn[2].n17 XThC.Tn[2].t22 154.679
R18688 XThC.Tn[2].n13 XThC.Tn[2].t42 154.679
R18689 XThC.Tn[2].n10 XThC.Tn[2].t33 154.679
R18690 XThC.Tn[2].n7 XThC.Tn[2].n6 135.248
R18691 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R18692 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R18693 XThC.Tn[2].n7 XThC.Tn[2].n5 98.982
R18694 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R18695 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R18696 XThC.Tn[2].n74 XThC.Tn[2].n9 32.6405
R18697 XThC.Tn[2].n1 XThC.Tn[2].t5 26.5955
R18698 XThC.Tn[2].n1 XThC.Tn[2].t4 26.5955
R18699 XThC.Tn[2].n0 XThC.Tn[2].t7 26.5955
R18700 XThC.Tn[2].n0 XThC.Tn[2].t6 26.5955
R18701 XThC.Tn[2].n3 XThC.Tn[2].t11 24.9236
R18702 XThC.Tn[2].n3 XThC.Tn[2].t10 24.9236
R18703 XThC.Tn[2].n4 XThC.Tn[2].t9 24.9236
R18704 XThC.Tn[2].n4 XThC.Tn[2].t8 24.9236
R18705 XThC.Tn[2].n5 XThC.Tn[2].t1 24.9236
R18706 XThC.Tn[2].n5 XThC.Tn[2].t2 24.9236
R18707 XThC.Tn[2].n6 XThC.Tn[2].t3 24.9236
R18708 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R18709 XThC.Tn[2].n75 XThC.Tn[2].n2 18.5605
R18710 XThC.Tn[2].n75 XThC.Tn[2].n74 11.5205
R18711 XThC.Tn[2] XThC.Tn[2].n12 8.0245
R18712 XThC.Tn[2].n72 XThC.Tn[2].n71 7.9105
R18713 XThC.Tn[2].n68 XThC.Tn[2].n67 7.9105
R18714 XThC.Tn[2].n64 XThC.Tn[2].n63 7.9105
R18715 XThC.Tn[2].n60 XThC.Tn[2].n59 7.9105
R18716 XThC.Tn[2].n56 XThC.Tn[2].n55 7.9105
R18717 XThC.Tn[2].n52 XThC.Tn[2].n51 7.9105
R18718 XThC.Tn[2].n48 XThC.Tn[2].n47 7.9105
R18719 XThC.Tn[2].n44 XThC.Tn[2].n43 7.9105
R18720 XThC.Tn[2].n40 XThC.Tn[2].n39 7.9105
R18721 XThC.Tn[2].n36 XThC.Tn[2].n35 7.9105
R18722 XThC.Tn[2].n32 XThC.Tn[2].n31 7.9105
R18723 XThC.Tn[2].n28 XThC.Tn[2].n27 7.9105
R18724 XThC.Tn[2].n24 XThC.Tn[2].n23 7.9105
R18725 XThC.Tn[2].n20 XThC.Tn[2].n19 7.9105
R18726 XThC.Tn[2].n16 XThC.Tn[2].n15 7.9105
R18727 XThC.Tn[2].n73 XThC.Tn[2] 5.58686
R18728 XThC.Tn[2].n74 XThC.Tn[2].n73 4.6005
R18729 XThC.Tn[2].n73 XThC.Tn[2] 1.83383
R18730 XThC.Tn[2] XThC.Tn[2].n75 0.6405
R18731 XThC.Tn[2].n16 XThC.Tn[2] 0.235138
R18732 XThC.Tn[2].n20 XThC.Tn[2] 0.235138
R18733 XThC.Tn[2].n24 XThC.Tn[2] 0.235138
R18734 XThC.Tn[2].n28 XThC.Tn[2] 0.235138
R18735 XThC.Tn[2].n32 XThC.Tn[2] 0.235138
R18736 XThC.Tn[2].n36 XThC.Tn[2] 0.235138
R18737 XThC.Tn[2].n40 XThC.Tn[2] 0.235138
R18738 XThC.Tn[2].n44 XThC.Tn[2] 0.235138
R18739 XThC.Tn[2].n48 XThC.Tn[2] 0.235138
R18740 XThC.Tn[2].n52 XThC.Tn[2] 0.235138
R18741 XThC.Tn[2].n56 XThC.Tn[2] 0.235138
R18742 XThC.Tn[2].n60 XThC.Tn[2] 0.235138
R18743 XThC.Tn[2].n64 XThC.Tn[2] 0.235138
R18744 XThC.Tn[2].n68 XThC.Tn[2] 0.235138
R18745 XThC.Tn[2].n72 XThC.Tn[2] 0.235138
R18746 XThC.Tn[2] XThC.Tn[2].n16 0.114505
R18747 XThC.Tn[2] XThC.Tn[2].n20 0.114505
R18748 XThC.Tn[2] XThC.Tn[2].n24 0.114505
R18749 XThC.Tn[2] XThC.Tn[2].n28 0.114505
R18750 XThC.Tn[2] XThC.Tn[2].n32 0.114505
R18751 XThC.Tn[2] XThC.Tn[2].n36 0.114505
R18752 XThC.Tn[2] XThC.Tn[2].n40 0.114505
R18753 XThC.Tn[2] XThC.Tn[2].n44 0.114505
R18754 XThC.Tn[2] XThC.Tn[2].n48 0.114505
R18755 XThC.Tn[2] XThC.Tn[2].n52 0.114505
R18756 XThC.Tn[2] XThC.Tn[2].n56 0.114505
R18757 XThC.Tn[2] XThC.Tn[2].n60 0.114505
R18758 XThC.Tn[2] XThC.Tn[2].n64 0.114505
R18759 XThC.Tn[2] XThC.Tn[2].n68 0.114505
R18760 XThC.Tn[2] XThC.Tn[2].n72 0.114505
R18761 XThC.Tn[2].n71 XThC.Tn[2].n70 0.0599512
R18762 XThC.Tn[2].n67 XThC.Tn[2].n66 0.0599512
R18763 XThC.Tn[2].n63 XThC.Tn[2].n62 0.0599512
R18764 XThC.Tn[2].n59 XThC.Tn[2].n58 0.0599512
R18765 XThC.Tn[2].n55 XThC.Tn[2].n54 0.0599512
R18766 XThC.Tn[2].n51 XThC.Tn[2].n50 0.0599512
R18767 XThC.Tn[2].n47 XThC.Tn[2].n46 0.0599512
R18768 XThC.Tn[2].n43 XThC.Tn[2].n42 0.0599512
R18769 XThC.Tn[2].n39 XThC.Tn[2].n38 0.0599512
R18770 XThC.Tn[2].n35 XThC.Tn[2].n34 0.0599512
R18771 XThC.Tn[2].n31 XThC.Tn[2].n30 0.0599512
R18772 XThC.Tn[2].n27 XThC.Tn[2].n26 0.0599512
R18773 XThC.Tn[2].n23 XThC.Tn[2].n22 0.0599512
R18774 XThC.Tn[2].n19 XThC.Tn[2].n18 0.0599512
R18775 XThC.Tn[2].n15 XThC.Tn[2].n14 0.0599512
R18776 XThC.Tn[2].n12 XThC.Tn[2].n11 0.0599512
R18777 XThC.Tn[2].n70 XThC.Tn[2] 0.0469286
R18778 XThC.Tn[2].n66 XThC.Tn[2] 0.0469286
R18779 XThC.Tn[2].n62 XThC.Tn[2] 0.0469286
R18780 XThC.Tn[2].n58 XThC.Tn[2] 0.0469286
R18781 XThC.Tn[2].n54 XThC.Tn[2] 0.0469286
R18782 XThC.Tn[2].n50 XThC.Tn[2] 0.0469286
R18783 XThC.Tn[2].n46 XThC.Tn[2] 0.0469286
R18784 XThC.Tn[2].n42 XThC.Tn[2] 0.0469286
R18785 XThC.Tn[2].n38 XThC.Tn[2] 0.0469286
R18786 XThC.Tn[2].n34 XThC.Tn[2] 0.0469286
R18787 XThC.Tn[2].n30 XThC.Tn[2] 0.0469286
R18788 XThC.Tn[2].n26 XThC.Tn[2] 0.0469286
R18789 XThC.Tn[2].n22 XThC.Tn[2] 0.0469286
R18790 XThC.Tn[2].n18 XThC.Tn[2] 0.0469286
R18791 XThC.Tn[2].n14 XThC.Tn[2] 0.0469286
R18792 XThC.Tn[2].n11 XThC.Tn[2] 0.0469286
R18793 XThC.Tn[2].n70 XThC.Tn[2] 0.0401341
R18794 XThC.Tn[2].n66 XThC.Tn[2] 0.0401341
R18795 XThC.Tn[2].n62 XThC.Tn[2] 0.0401341
R18796 XThC.Tn[2].n58 XThC.Tn[2] 0.0401341
R18797 XThC.Tn[2].n54 XThC.Tn[2] 0.0401341
R18798 XThC.Tn[2].n50 XThC.Tn[2] 0.0401341
R18799 XThC.Tn[2].n46 XThC.Tn[2] 0.0401341
R18800 XThC.Tn[2].n42 XThC.Tn[2] 0.0401341
R18801 XThC.Tn[2].n38 XThC.Tn[2] 0.0401341
R18802 XThC.Tn[2].n34 XThC.Tn[2] 0.0401341
R18803 XThC.Tn[2].n30 XThC.Tn[2] 0.0401341
R18804 XThC.Tn[2].n26 XThC.Tn[2] 0.0401341
R18805 XThC.Tn[2].n22 XThC.Tn[2] 0.0401341
R18806 XThC.Tn[2].n18 XThC.Tn[2] 0.0401341
R18807 XThC.Tn[2].n14 XThC.Tn[2] 0.0401341
R18808 XThC.Tn[2].n11 XThC.Tn[2] 0.0401341
R18809 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R18810 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R18811 XThR.Tn[0] XThR.Tn[0].n82 161.363
R18812 XThR.Tn[0] XThR.Tn[0].n77 161.363
R18813 XThR.Tn[0] XThR.Tn[0].n72 161.363
R18814 XThR.Tn[0] XThR.Tn[0].n67 161.363
R18815 XThR.Tn[0] XThR.Tn[0].n62 161.363
R18816 XThR.Tn[0] XThR.Tn[0].n57 161.363
R18817 XThR.Tn[0] XThR.Tn[0].n52 161.363
R18818 XThR.Tn[0] XThR.Tn[0].n47 161.363
R18819 XThR.Tn[0] XThR.Tn[0].n42 161.363
R18820 XThR.Tn[0] XThR.Tn[0].n37 161.363
R18821 XThR.Tn[0] XThR.Tn[0].n32 161.363
R18822 XThR.Tn[0] XThR.Tn[0].n27 161.363
R18823 XThR.Tn[0] XThR.Tn[0].n22 161.363
R18824 XThR.Tn[0] XThR.Tn[0].n17 161.363
R18825 XThR.Tn[0] XThR.Tn[0].n12 161.363
R18826 XThR.Tn[0] XThR.Tn[0].n10 161.363
R18827 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R18828 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R18829 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R18830 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R18831 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R18832 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R18833 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R18834 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R18835 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R18836 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R18837 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R18838 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R18839 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R18840 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R18841 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R18842 XThR.Tn[0].n83 XThR.Tn[0].t62 161.106
R18843 XThR.Tn[0].n82 XThR.Tn[0].t28 161.106
R18844 XThR.Tn[0].n78 XThR.Tn[0].t71 161.106
R18845 XThR.Tn[0].n77 XThR.Tn[0].t33 161.106
R18846 XThR.Tn[0].n73 XThR.Tn[0].t54 161.106
R18847 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R18848 XThR.Tn[0].n68 XThR.Tn[0].t36 161.106
R18849 XThR.Tn[0].n67 XThR.Tn[0].t59 161.106
R18850 XThR.Tn[0].n63 XThR.Tn[0].t61 161.106
R18851 XThR.Tn[0].n62 XThR.Tn[0].t27 161.106
R18852 XThR.Tn[0].n58 XThR.Tn[0].t25 161.106
R18853 XThR.Tn[0].n57 XThR.Tn[0].t49 161.106
R18854 XThR.Tn[0].n53 XThR.Tn[0].t69 161.106
R18855 XThR.Tn[0].n52 XThR.Tn[0].t31 161.106
R18856 XThR.Tn[0].n48 XThR.Tn[0].t51 161.106
R18857 XThR.Tn[0].n47 XThR.Tn[0].t13 161.106
R18858 XThR.Tn[0].n43 XThR.Tn[0].t35 161.106
R18859 XThR.Tn[0].n42 XThR.Tn[0].t57 161.106
R18860 XThR.Tn[0].n38 XThR.Tn[0].t40 161.106
R18861 XThR.Tn[0].n37 XThR.Tn[0].t64 161.106
R18862 XThR.Tn[0].n33 XThR.Tn[0].t24 161.106
R18863 XThR.Tn[0].n32 XThR.Tn[0].t48 161.106
R18864 XThR.Tn[0].n28 XThR.Tn[0].t53 161.106
R18865 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R18866 XThR.Tn[0].n23 XThR.Tn[0].t22 161.106
R18867 XThR.Tn[0].n22 XThR.Tn[0].t46 161.106
R18868 XThR.Tn[0].n18 XThR.Tn[0].t68 161.106
R18869 XThR.Tn[0].n17 XThR.Tn[0].t30 161.106
R18870 XThR.Tn[0].n13 XThR.Tn[0].t29 161.106
R18871 XThR.Tn[0].n12 XThR.Tn[0].t55 161.106
R18872 XThR.Tn[0].n10 XThR.Tn[0].t37 161.106
R18873 XThR.Tn[0].n83 XThR.Tn[0].t19 154.679
R18874 XThR.Tn[0].n82 XThR.Tn[0].t45 154.679
R18875 XThR.Tn[0].n78 XThR.Tn[0].t60 154.679
R18876 XThR.Tn[0].n77 XThR.Tn[0].t21 154.679
R18877 XThR.Tn[0].n73 XThR.Tn[0].t42 154.679
R18878 XThR.Tn[0].n72 XThR.Tn[0].t66 154.679
R18879 XThR.Tn[0].n68 XThR.Tn[0].t72 154.679
R18880 XThR.Tn[0].n67 XThR.Tn[0].t34 154.679
R18881 XThR.Tn[0].n63 XThR.Tn[0].t56 154.679
R18882 XThR.Tn[0].n62 XThR.Tn[0].t17 154.679
R18883 XThR.Tn[0].n58 XThR.Tn[0].t18 154.679
R18884 XThR.Tn[0].n57 XThR.Tn[0].t44 154.679
R18885 XThR.Tn[0].n53 XThR.Tn[0].t43 154.679
R18886 XThR.Tn[0].n52 XThR.Tn[0].t67 154.679
R18887 XThR.Tn[0].n48 XThR.Tn[0].t26 154.679
R18888 XThR.Tn[0].n47 XThR.Tn[0].t50 154.679
R18889 XThR.Tn[0].n43 XThR.Tn[0].t70 154.679
R18890 XThR.Tn[0].n42 XThR.Tn[0].t32 154.679
R18891 XThR.Tn[0].n38 XThR.Tn[0].t52 154.679
R18892 XThR.Tn[0].n37 XThR.Tn[0].t14 154.679
R18893 XThR.Tn[0].n33 XThR.Tn[0].t58 154.679
R18894 XThR.Tn[0].n32 XThR.Tn[0].t20 154.679
R18895 XThR.Tn[0].n28 XThR.Tn[0].t41 154.679
R18896 XThR.Tn[0].n27 XThR.Tn[0].t65 154.679
R18897 XThR.Tn[0].n23 XThR.Tn[0].t12 154.679
R18898 XThR.Tn[0].n22 XThR.Tn[0].t38 154.679
R18899 XThR.Tn[0].n18 XThR.Tn[0].t39 154.679
R18900 XThR.Tn[0].n17 XThR.Tn[0].t63 154.679
R18901 XThR.Tn[0].n13 XThR.Tn[0].t23 154.679
R18902 XThR.Tn[0].n12 XThR.Tn[0].t47 154.679
R18903 XThR.Tn[0].n10 XThR.Tn[0].t73 154.679
R18904 XThR.Tn[0].n7 XThR.Tn[0].n6 135.249
R18905 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R18906 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R18907 XThR.Tn[0].n7 XThR.Tn[0].n5 98.982
R18908 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R18909 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R18910 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R18911 XThR.Tn[0].n1 XThR.Tn[0].t5 26.5955
R18912 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R18913 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R18914 XThR.Tn[0].n0 XThR.Tn[0].t7 26.5955
R18915 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R18916 XThR.Tn[0].n3 XThR.Tn[0].t10 24.9236
R18917 XThR.Tn[0].n4 XThR.Tn[0].t8 24.9236
R18918 XThR.Tn[0].n4 XThR.Tn[0].t11 24.9236
R18919 XThR.Tn[0].n5 XThR.Tn[0].t2 24.9236
R18920 XThR.Tn[0].n5 XThR.Tn[0].t3 24.9236
R18921 XThR.Tn[0].n6 XThR.Tn[0].t1 24.9236
R18922 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R18923 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R18924 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R18925 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R18926 XThR.Tn[0] XThR.Tn[0].n11 5.34871
R18927 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R18928 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R18929 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R18930 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R18931 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R18932 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R18933 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R18934 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R18935 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R18936 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R18937 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R18938 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R18939 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R18940 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R18941 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R18942 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R18943 XThR.Tn[0].n16 XThR.Tn[0] 2.51836
R18944 XThR.Tn[0].n21 XThR.Tn[0] 2.51836
R18945 XThR.Tn[0].n26 XThR.Tn[0] 2.51836
R18946 XThR.Tn[0].n31 XThR.Tn[0] 2.51836
R18947 XThR.Tn[0].n36 XThR.Tn[0] 2.51836
R18948 XThR.Tn[0].n41 XThR.Tn[0] 2.51836
R18949 XThR.Tn[0].n46 XThR.Tn[0] 2.51836
R18950 XThR.Tn[0].n51 XThR.Tn[0] 2.51836
R18951 XThR.Tn[0].n56 XThR.Tn[0] 2.51836
R18952 XThR.Tn[0].n61 XThR.Tn[0] 2.51836
R18953 XThR.Tn[0].n66 XThR.Tn[0] 2.51836
R18954 XThR.Tn[0].n71 XThR.Tn[0] 2.51836
R18955 XThR.Tn[0].n76 XThR.Tn[0] 2.51836
R18956 XThR.Tn[0].n81 XThR.Tn[0] 2.51836
R18957 XThR.Tn[0].n86 XThR.Tn[0] 2.51836
R18958 XThR.Tn[0] XThR.Tn[0].n16 0.848714
R18959 XThR.Tn[0] XThR.Tn[0].n21 0.848714
R18960 XThR.Tn[0] XThR.Tn[0].n26 0.848714
R18961 XThR.Tn[0] XThR.Tn[0].n31 0.848714
R18962 XThR.Tn[0] XThR.Tn[0].n36 0.848714
R18963 XThR.Tn[0] XThR.Tn[0].n41 0.848714
R18964 XThR.Tn[0] XThR.Tn[0].n46 0.848714
R18965 XThR.Tn[0] XThR.Tn[0].n51 0.848714
R18966 XThR.Tn[0] XThR.Tn[0].n56 0.848714
R18967 XThR.Tn[0] XThR.Tn[0].n61 0.848714
R18968 XThR.Tn[0] XThR.Tn[0].n66 0.848714
R18969 XThR.Tn[0] XThR.Tn[0].n71 0.848714
R18970 XThR.Tn[0] XThR.Tn[0].n76 0.848714
R18971 XThR.Tn[0] XThR.Tn[0].n81 0.848714
R18972 XThR.Tn[0] XThR.Tn[0].n86 0.848714
R18973 XThR.Tn[0].n11 XThR.Tn[0] 0.485653
R18974 XThR.Tn[0].n84 XThR.Tn[0] 0.21482
R18975 XThR.Tn[0].n79 XThR.Tn[0] 0.21482
R18976 XThR.Tn[0].n74 XThR.Tn[0] 0.21482
R18977 XThR.Tn[0].n69 XThR.Tn[0] 0.21482
R18978 XThR.Tn[0].n64 XThR.Tn[0] 0.21482
R18979 XThR.Tn[0].n59 XThR.Tn[0] 0.21482
R18980 XThR.Tn[0].n54 XThR.Tn[0] 0.21482
R18981 XThR.Tn[0].n49 XThR.Tn[0] 0.21482
R18982 XThR.Tn[0].n44 XThR.Tn[0] 0.21482
R18983 XThR.Tn[0].n39 XThR.Tn[0] 0.21482
R18984 XThR.Tn[0].n34 XThR.Tn[0] 0.21482
R18985 XThR.Tn[0].n29 XThR.Tn[0] 0.21482
R18986 XThR.Tn[0].n24 XThR.Tn[0] 0.21482
R18987 XThR.Tn[0].n19 XThR.Tn[0] 0.21482
R18988 XThR.Tn[0].n14 XThR.Tn[0] 0.21482
R18989 XThR.Tn[0].n85 XThR.Tn[0] 0.0608448
R18990 XThR.Tn[0].n80 XThR.Tn[0] 0.0608448
R18991 XThR.Tn[0].n75 XThR.Tn[0] 0.0608448
R18992 XThR.Tn[0].n70 XThR.Tn[0] 0.0608448
R18993 XThR.Tn[0].n65 XThR.Tn[0] 0.0608448
R18994 XThR.Tn[0].n60 XThR.Tn[0] 0.0608448
R18995 XThR.Tn[0].n55 XThR.Tn[0] 0.0608448
R18996 XThR.Tn[0].n50 XThR.Tn[0] 0.0608448
R18997 XThR.Tn[0].n45 XThR.Tn[0] 0.0608448
R18998 XThR.Tn[0].n40 XThR.Tn[0] 0.0608448
R18999 XThR.Tn[0].n35 XThR.Tn[0] 0.0608448
R19000 XThR.Tn[0].n30 XThR.Tn[0] 0.0608448
R19001 XThR.Tn[0].n25 XThR.Tn[0] 0.0608448
R19002 XThR.Tn[0].n20 XThR.Tn[0] 0.0608448
R19003 XThR.Tn[0].n15 XThR.Tn[0] 0.0608448
R19004 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R19005 XThR.Tn[0] XThR.Tn[0].n87 0.038
R19006 XThR.Tn[0].n11 XThR.Tn[0] 0.00744444
R19007 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00265517
R19008 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00265517
R19009 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00265517
R19010 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00265517
R19011 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00265517
R19012 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00265517
R19013 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00265517
R19014 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00265517
R19015 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00265517
R19016 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00265517
R19017 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00265517
R19018 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00265517
R19019 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00265517
R19020 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00265517
R19021 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00265517
R19022 XThR.Tn[9].n87 XThR.Tn[9].n86 256.103
R19023 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R19024 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R19025 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R19026 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R19027 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R19028 XThR.Tn[9] XThR.Tn[9].n78 161.363
R19029 XThR.Tn[9] XThR.Tn[9].n73 161.363
R19030 XThR.Tn[9] XThR.Tn[9].n68 161.363
R19031 XThR.Tn[9] XThR.Tn[9].n63 161.363
R19032 XThR.Tn[9] XThR.Tn[9].n58 161.363
R19033 XThR.Tn[9] XThR.Tn[9].n53 161.363
R19034 XThR.Tn[9] XThR.Tn[9].n48 161.363
R19035 XThR.Tn[9] XThR.Tn[9].n43 161.363
R19036 XThR.Tn[9] XThR.Tn[9].n38 161.363
R19037 XThR.Tn[9] XThR.Tn[9].n33 161.363
R19038 XThR.Tn[9] XThR.Tn[9].n28 161.363
R19039 XThR.Tn[9] XThR.Tn[9].n23 161.363
R19040 XThR.Tn[9] XThR.Tn[9].n18 161.363
R19041 XThR.Tn[9] XThR.Tn[9].n13 161.363
R19042 XThR.Tn[9] XThR.Tn[9].n8 161.363
R19043 XThR.Tn[9] XThR.Tn[9].n6 161.363
R19044 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R19045 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R19046 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R19047 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R19048 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R19049 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R19050 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R19051 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R19052 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R19053 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R19054 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R19055 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R19056 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R19057 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R19058 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R19059 XThR.Tn[9].n79 XThR.Tn[9].t38 161.106
R19060 XThR.Tn[9].n78 XThR.Tn[9].t46 161.106
R19061 XThR.Tn[9].n74 XThR.Tn[9].t45 161.106
R19062 XThR.Tn[9].n73 XThR.Tn[9].t52 161.106
R19063 XThR.Tn[9].n69 XThR.Tn[9].t28 161.106
R19064 XThR.Tn[9].n68 XThR.Tn[9].t33 161.106
R19065 XThR.Tn[9].n64 XThR.Tn[9].t73 161.106
R19066 XThR.Tn[9].n63 XThR.Tn[9].t13 161.106
R19067 XThR.Tn[9].n59 XThR.Tn[9].t37 161.106
R19068 XThR.Tn[9].n58 XThR.Tn[9].t43 161.106
R19069 XThR.Tn[9].n54 XThR.Tn[9].t61 161.106
R19070 XThR.Tn[9].n53 XThR.Tn[9].t69 161.106
R19071 XThR.Tn[9].n49 XThR.Tn[9].t42 161.106
R19072 XThR.Tn[9].n48 XThR.Tn[9].t50 161.106
R19073 XThR.Tn[9].n44 XThR.Tn[9].t24 161.106
R19074 XThR.Tn[9].n43 XThR.Tn[9].t30 161.106
R19075 XThR.Tn[9].n39 XThR.Tn[9].t71 161.106
R19076 XThR.Tn[9].n38 XThR.Tn[9].t12 161.106
R19077 XThR.Tn[9].n34 XThR.Tn[9].t15 161.106
R19078 XThR.Tn[9].n33 XThR.Tn[9].t20 161.106
R19079 XThR.Tn[9].n29 XThR.Tn[9].t60 161.106
R19080 XThR.Tn[9].n28 XThR.Tn[9].t68 161.106
R19081 XThR.Tn[9].n24 XThR.Tn[9].t26 161.106
R19082 XThR.Tn[9].n23 XThR.Tn[9].t32 161.106
R19083 XThR.Tn[9].n19 XThR.Tn[9].t58 161.106
R19084 XThR.Tn[9].n18 XThR.Tn[9].t66 161.106
R19085 XThR.Tn[9].n14 XThR.Tn[9].t41 161.106
R19086 XThR.Tn[9].n13 XThR.Tn[9].t48 161.106
R19087 XThR.Tn[9].n9 XThR.Tn[9].t65 161.106
R19088 XThR.Tn[9].n8 XThR.Tn[9].t72 161.106
R19089 XThR.Tn[9].n6 XThR.Tn[9].t54 161.106
R19090 XThR.Tn[9].n79 XThR.Tn[9].t57 154.679
R19091 XThR.Tn[9].n78 XThR.Tn[9].t64 154.679
R19092 XThR.Tn[9].n74 XThR.Tn[9].t36 154.679
R19093 XThR.Tn[9].n73 XThR.Tn[9].t40 154.679
R19094 XThR.Tn[9].n69 XThR.Tn[9].t17 154.679
R19095 XThR.Tn[9].n68 XThR.Tn[9].t22 154.679
R19096 XThR.Tn[9].n64 XThR.Tn[9].t47 154.679
R19097 XThR.Tn[9].n63 XThR.Tn[9].t53 154.679
R19098 XThR.Tn[9].n59 XThR.Tn[9].t29 154.679
R19099 XThR.Tn[9].n58 XThR.Tn[9].t34 154.679
R19100 XThR.Tn[9].n54 XThR.Tn[9].t56 154.679
R19101 XThR.Tn[9].n53 XThR.Tn[9].t63 154.679
R19102 XThR.Tn[9].n49 XThR.Tn[9].t18 154.679
R19103 XThR.Tn[9].n48 XThR.Tn[9].t23 154.679
R19104 XThR.Tn[9].n44 XThR.Tn[9].t62 154.679
R19105 XThR.Tn[9].n43 XThR.Tn[9].t70 154.679
R19106 XThR.Tn[9].n39 XThR.Tn[9].t44 154.679
R19107 XThR.Tn[9].n38 XThR.Tn[9].t51 154.679
R19108 XThR.Tn[9].n34 XThR.Tn[9].t25 154.679
R19109 XThR.Tn[9].n33 XThR.Tn[9].t31 154.679
R19110 XThR.Tn[9].n29 XThR.Tn[9].t35 154.679
R19111 XThR.Tn[9].n28 XThR.Tn[9].t39 154.679
R19112 XThR.Tn[9].n24 XThR.Tn[9].t16 154.679
R19113 XThR.Tn[9].n23 XThR.Tn[9].t21 154.679
R19114 XThR.Tn[9].n19 XThR.Tn[9].t49 154.679
R19115 XThR.Tn[9].n18 XThR.Tn[9].t55 154.679
R19116 XThR.Tn[9].n14 XThR.Tn[9].t14 154.679
R19117 XThR.Tn[9].n13 XThR.Tn[9].t19 154.679
R19118 XThR.Tn[9].n9 XThR.Tn[9].t59 154.679
R19119 XThR.Tn[9].n8 XThR.Tn[9].t67 154.679
R19120 XThR.Tn[9].n6 XThR.Tn[9].t27 154.679
R19121 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R19122 XThR.Tn[9].n85 XThR.Tn[9].t2 26.5955
R19123 XThR.Tn[9].n85 XThR.Tn[9].t0 26.5955
R19124 XThR.Tn[9].n0 XThR.Tn[9].t10 26.5955
R19125 XThR.Tn[9].n0 XThR.Tn[9].t8 26.5955
R19126 XThR.Tn[9].n1 XThR.Tn[9].t11 26.5955
R19127 XThR.Tn[9].n1 XThR.Tn[9].t9 26.5955
R19128 XThR.Tn[9].n86 XThR.Tn[9].t3 26.5955
R19129 XThR.Tn[9].n86 XThR.Tn[9].t1 26.5955
R19130 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R19131 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R19132 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R19133 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R19134 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R19135 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R19136 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R19137 XThR.Tn[9] XThR.Tn[9].n7 5.34871
R19138 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R19139 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R19140 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R19141 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R19142 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R19143 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R19144 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R19145 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R19146 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R19147 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R19148 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R19149 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R19150 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R19151 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R19152 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R19153 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R19154 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R19155 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R19156 XThR.Tn[9].n12 XThR.Tn[9] 2.51836
R19157 XThR.Tn[9].n17 XThR.Tn[9] 2.51836
R19158 XThR.Tn[9].n22 XThR.Tn[9] 2.51836
R19159 XThR.Tn[9].n27 XThR.Tn[9] 2.51836
R19160 XThR.Tn[9].n32 XThR.Tn[9] 2.51836
R19161 XThR.Tn[9].n37 XThR.Tn[9] 2.51836
R19162 XThR.Tn[9].n42 XThR.Tn[9] 2.51836
R19163 XThR.Tn[9].n47 XThR.Tn[9] 2.51836
R19164 XThR.Tn[9].n52 XThR.Tn[9] 2.51836
R19165 XThR.Tn[9].n57 XThR.Tn[9] 2.51836
R19166 XThR.Tn[9].n62 XThR.Tn[9] 2.51836
R19167 XThR.Tn[9].n67 XThR.Tn[9] 2.51836
R19168 XThR.Tn[9].n72 XThR.Tn[9] 2.51836
R19169 XThR.Tn[9].n77 XThR.Tn[9] 2.51836
R19170 XThR.Tn[9].n82 XThR.Tn[9] 2.51836
R19171 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R19172 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R19173 XThR.Tn[9] XThR.Tn[9].n12 0.848714
R19174 XThR.Tn[9] XThR.Tn[9].n17 0.848714
R19175 XThR.Tn[9] XThR.Tn[9].n22 0.848714
R19176 XThR.Tn[9] XThR.Tn[9].n27 0.848714
R19177 XThR.Tn[9] XThR.Tn[9].n32 0.848714
R19178 XThR.Tn[9] XThR.Tn[9].n37 0.848714
R19179 XThR.Tn[9] XThR.Tn[9].n42 0.848714
R19180 XThR.Tn[9] XThR.Tn[9].n47 0.848714
R19181 XThR.Tn[9] XThR.Tn[9].n52 0.848714
R19182 XThR.Tn[9] XThR.Tn[9].n57 0.848714
R19183 XThR.Tn[9] XThR.Tn[9].n62 0.848714
R19184 XThR.Tn[9] XThR.Tn[9].n67 0.848714
R19185 XThR.Tn[9] XThR.Tn[9].n72 0.848714
R19186 XThR.Tn[9] XThR.Tn[9].n77 0.848714
R19187 XThR.Tn[9] XThR.Tn[9].n82 0.848714
R19188 XThR.Tn[9].n7 XThR.Tn[9] 0.485653
R19189 XThR.Tn[9].n80 XThR.Tn[9] 0.21482
R19190 XThR.Tn[9].n75 XThR.Tn[9] 0.21482
R19191 XThR.Tn[9].n70 XThR.Tn[9] 0.21482
R19192 XThR.Tn[9].n65 XThR.Tn[9] 0.21482
R19193 XThR.Tn[9].n60 XThR.Tn[9] 0.21482
R19194 XThR.Tn[9].n55 XThR.Tn[9] 0.21482
R19195 XThR.Tn[9].n50 XThR.Tn[9] 0.21482
R19196 XThR.Tn[9].n45 XThR.Tn[9] 0.21482
R19197 XThR.Tn[9].n40 XThR.Tn[9] 0.21482
R19198 XThR.Tn[9].n35 XThR.Tn[9] 0.21482
R19199 XThR.Tn[9].n30 XThR.Tn[9] 0.21482
R19200 XThR.Tn[9].n25 XThR.Tn[9] 0.21482
R19201 XThR.Tn[9].n20 XThR.Tn[9] 0.21482
R19202 XThR.Tn[9].n15 XThR.Tn[9] 0.21482
R19203 XThR.Tn[9].n10 XThR.Tn[9] 0.21482
R19204 XThR.Tn[9].n81 XThR.Tn[9] 0.0608448
R19205 XThR.Tn[9].n76 XThR.Tn[9] 0.0608448
R19206 XThR.Tn[9].n71 XThR.Tn[9] 0.0608448
R19207 XThR.Tn[9].n66 XThR.Tn[9] 0.0608448
R19208 XThR.Tn[9].n61 XThR.Tn[9] 0.0608448
R19209 XThR.Tn[9].n56 XThR.Tn[9] 0.0608448
R19210 XThR.Tn[9].n51 XThR.Tn[9] 0.0608448
R19211 XThR.Tn[9].n46 XThR.Tn[9] 0.0608448
R19212 XThR.Tn[9].n41 XThR.Tn[9] 0.0608448
R19213 XThR.Tn[9].n36 XThR.Tn[9] 0.0608448
R19214 XThR.Tn[9].n31 XThR.Tn[9] 0.0608448
R19215 XThR.Tn[9].n26 XThR.Tn[9] 0.0608448
R19216 XThR.Tn[9].n21 XThR.Tn[9] 0.0608448
R19217 XThR.Tn[9].n16 XThR.Tn[9] 0.0608448
R19218 XThR.Tn[9].n11 XThR.Tn[9] 0.0608448
R19219 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R19220 XThR.Tn[9] XThR.Tn[9].n83 0.038
R19221 XThR.Tn[9].n7 XThR.Tn[9] 0.00744444
R19222 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00265517
R19223 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00265517
R19224 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00265517
R19225 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00265517
R19226 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00265517
R19227 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00265517
R19228 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00265517
R19229 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00265517
R19230 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00265517
R19231 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00265517
R19232 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00265517
R19233 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00265517
R19234 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00265517
R19235 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00265517
R19236 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00265517
R19237 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R19238 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R19239 XThR.Tn[4] XThR.Tn[4].n82 161.363
R19240 XThR.Tn[4] XThR.Tn[4].n77 161.363
R19241 XThR.Tn[4] XThR.Tn[4].n72 161.363
R19242 XThR.Tn[4] XThR.Tn[4].n67 161.363
R19243 XThR.Tn[4] XThR.Tn[4].n62 161.363
R19244 XThR.Tn[4] XThR.Tn[4].n57 161.363
R19245 XThR.Tn[4] XThR.Tn[4].n52 161.363
R19246 XThR.Tn[4] XThR.Tn[4].n47 161.363
R19247 XThR.Tn[4] XThR.Tn[4].n42 161.363
R19248 XThR.Tn[4] XThR.Tn[4].n37 161.363
R19249 XThR.Tn[4] XThR.Tn[4].n32 161.363
R19250 XThR.Tn[4] XThR.Tn[4].n27 161.363
R19251 XThR.Tn[4] XThR.Tn[4].n22 161.363
R19252 XThR.Tn[4] XThR.Tn[4].n17 161.363
R19253 XThR.Tn[4] XThR.Tn[4].n12 161.363
R19254 XThR.Tn[4] XThR.Tn[4].n10 161.363
R19255 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R19256 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R19257 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R19258 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R19259 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R19260 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R19261 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R19262 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R19263 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R19264 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R19265 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R19266 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R19267 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R19268 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R19269 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R19270 XThR.Tn[4].n83 XThR.Tn[4].t61 161.106
R19271 XThR.Tn[4].n82 XThR.Tn[4].t63 161.106
R19272 XThR.Tn[4].n78 XThR.Tn[4].t67 161.106
R19273 XThR.Tn[4].n77 XThR.Tn[4].t72 161.106
R19274 XThR.Tn[4].n73 XThR.Tn[4].t49 161.106
R19275 XThR.Tn[4].n72 XThR.Tn[4].t54 161.106
R19276 XThR.Tn[4].n68 XThR.Tn[4].t32 161.106
R19277 XThR.Tn[4].n67 XThR.Tn[4].t34 161.106
R19278 XThR.Tn[4].n63 XThR.Tn[4].t60 161.106
R19279 XThR.Tn[4].n62 XThR.Tn[4].t62 161.106
R19280 XThR.Tn[4].n58 XThR.Tn[4].t22 161.106
R19281 XThR.Tn[4].n57 XThR.Tn[4].t27 161.106
R19282 XThR.Tn[4].n53 XThR.Tn[4].t65 161.106
R19283 XThR.Tn[4].n52 XThR.Tn[4].t70 161.106
R19284 XThR.Tn[4].n48 XThR.Tn[4].t46 161.106
R19285 XThR.Tn[4].n47 XThR.Tn[4].t51 161.106
R19286 XThR.Tn[4].n43 XThR.Tn[4].t31 161.106
R19287 XThR.Tn[4].n42 XThR.Tn[4].t33 161.106
R19288 XThR.Tn[4].n38 XThR.Tn[4].t36 161.106
R19289 XThR.Tn[4].n37 XThR.Tn[4].t41 161.106
R19290 XThR.Tn[4].n33 XThR.Tn[4].t21 161.106
R19291 XThR.Tn[4].n32 XThR.Tn[4].t26 161.106
R19292 XThR.Tn[4].n28 XThR.Tn[4].t48 161.106
R19293 XThR.Tn[4].n27 XThR.Tn[4].t53 161.106
R19294 XThR.Tn[4].n23 XThR.Tn[4].t18 161.106
R19295 XThR.Tn[4].n22 XThR.Tn[4].t24 161.106
R19296 XThR.Tn[4].n18 XThR.Tn[4].t64 161.106
R19297 XThR.Tn[4].n17 XThR.Tn[4].t68 161.106
R19298 XThR.Tn[4].n13 XThR.Tn[4].t29 161.106
R19299 XThR.Tn[4].n12 XThR.Tn[4].t30 161.106
R19300 XThR.Tn[4].n10 XThR.Tn[4].t13 161.106
R19301 XThR.Tn[4].n83 XThR.Tn[4].t16 154.679
R19302 XThR.Tn[4].n82 XThR.Tn[4].t19 154.679
R19303 XThR.Tn[4].n78 XThR.Tn[4].t57 154.679
R19304 XThR.Tn[4].n77 XThR.Tn[4].t59 154.679
R19305 XThR.Tn[4].n73 XThR.Tn[4].t38 154.679
R19306 XThR.Tn[4].n72 XThR.Tn[4].t43 154.679
R19307 XThR.Tn[4].n68 XThR.Tn[4].t69 154.679
R19308 XThR.Tn[4].n67 XThR.Tn[4].t73 154.679
R19309 XThR.Tn[4].n63 XThR.Tn[4].t50 154.679
R19310 XThR.Tn[4].n62 XThR.Tn[4].t55 154.679
R19311 XThR.Tn[4].n58 XThR.Tn[4].t15 154.679
R19312 XThR.Tn[4].n57 XThR.Tn[4].t17 154.679
R19313 XThR.Tn[4].n53 XThR.Tn[4].t39 154.679
R19314 XThR.Tn[4].n52 XThR.Tn[4].t44 154.679
R19315 XThR.Tn[4].n48 XThR.Tn[4].t23 154.679
R19316 XThR.Tn[4].n47 XThR.Tn[4].t28 154.679
R19317 XThR.Tn[4].n43 XThR.Tn[4].t66 154.679
R19318 XThR.Tn[4].n42 XThR.Tn[4].t71 154.679
R19319 XThR.Tn[4].n38 XThR.Tn[4].t47 154.679
R19320 XThR.Tn[4].n37 XThR.Tn[4].t52 154.679
R19321 XThR.Tn[4].n33 XThR.Tn[4].t56 154.679
R19322 XThR.Tn[4].n32 XThR.Tn[4].t58 154.679
R19323 XThR.Tn[4].n28 XThR.Tn[4].t37 154.679
R19324 XThR.Tn[4].n27 XThR.Tn[4].t42 154.679
R19325 XThR.Tn[4].n23 XThR.Tn[4].t12 154.679
R19326 XThR.Tn[4].n22 XThR.Tn[4].t14 154.679
R19327 XThR.Tn[4].n18 XThR.Tn[4].t35 154.679
R19328 XThR.Tn[4].n17 XThR.Tn[4].t40 154.679
R19329 XThR.Tn[4].n13 XThR.Tn[4].t20 154.679
R19330 XThR.Tn[4].n12 XThR.Tn[4].t25 154.679
R19331 XThR.Tn[4].n10 XThR.Tn[4].t45 154.679
R19332 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R19333 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R19334 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R19335 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R19336 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R19337 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R19338 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R19339 XThR.Tn[4].n1 XThR.Tn[4].t8 26.5955
R19340 XThR.Tn[4].n1 XThR.Tn[4].t11 26.5955
R19341 XThR.Tn[4].n0 XThR.Tn[4].t9 26.5955
R19342 XThR.Tn[4].n0 XThR.Tn[4].t10 26.5955
R19343 XThR.Tn[4].n3 XThR.Tn[4].t7 24.9236
R19344 XThR.Tn[4].n3 XThR.Tn[4].t4 24.9236
R19345 XThR.Tn[4].n4 XThR.Tn[4].t6 24.9236
R19346 XThR.Tn[4].n4 XThR.Tn[4].t5 24.9236
R19347 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R19348 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R19349 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R19350 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R19351 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R19352 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R19353 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R19354 XThR.Tn[4] XThR.Tn[4].n11 5.34871
R19355 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R19356 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R19357 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R19358 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R19359 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R19360 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R19361 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R19362 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R19363 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R19364 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R19365 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R19366 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R19367 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R19368 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R19369 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R19370 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R19371 XThR.Tn[4].n16 XThR.Tn[4] 2.51836
R19372 XThR.Tn[4].n21 XThR.Tn[4] 2.51836
R19373 XThR.Tn[4].n26 XThR.Tn[4] 2.51836
R19374 XThR.Tn[4].n31 XThR.Tn[4] 2.51836
R19375 XThR.Tn[4].n36 XThR.Tn[4] 2.51836
R19376 XThR.Tn[4].n41 XThR.Tn[4] 2.51836
R19377 XThR.Tn[4].n46 XThR.Tn[4] 2.51836
R19378 XThR.Tn[4].n51 XThR.Tn[4] 2.51836
R19379 XThR.Tn[4].n56 XThR.Tn[4] 2.51836
R19380 XThR.Tn[4].n61 XThR.Tn[4] 2.51836
R19381 XThR.Tn[4].n66 XThR.Tn[4] 2.51836
R19382 XThR.Tn[4].n71 XThR.Tn[4] 2.51836
R19383 XThR.Tn[4].n76 XThR.Tn[4] 2.51836
R19384 XThR.Tn[4].n81 XThR.Tn[4] 2.51836
R19385 XThR.Tn[4].n86 XThR.Tn[4] 2.51836
R19386 XThR.Tn[4] XThR.Tn[4].n16 0.848714
R19387 XThR.Tn[4] XThR.Tn[4].n21 0.848714
R19388 XThR.Tn[4] XThR.Tn[4].n26 0.848714
R19389 XThR.Tn[4] XThR.Tn[4].n31 0.848714
R19390 XThR.Tn[4] XThR.Tn[4].n36 0.848714
R19391 XThR.Tn[4] XThR.Tn[4].n41 0.848714
R19392 XThR.Tn[4] XThR.Tn[4].n46 0.848714
R19393 XThR.Tn[4] XThR.Tn[4].n51 0.848714
R19394 XThR.Tn[4] XThR.Tn[4].n56 0.848714
R19395 XThR.Tn[4] XThR.Tn[4].n61 0.848714
R19396 XThR.Tn[4] XThR.Tn[4].n66 0.848714
R19397 XThR.Tn[4] XThR.Tn[4].n71 0.848714
R19398 XThR.Tn[4] XThR.Tn[4].n76 0.848714
R19399 XThR.Tn[4] XThR.Tn[4].n81 0.848714
R19400 XThR.Tn[4] XThR.Tn[4].n86 0.848714
R19401 XThR.Tn[4].n11 XThR.Tn[4] 0.485653
R19402 XThR.Tn[4].n84 XThR.Tn[4] 0.21482
R19403 XThR.Tn[4].n79 XThR.Tn[4] 0.21482
R19404 XThR.Tn[4].n74 XThR.Tn[4] 0.21482
R19405 XThR.Tn[4].n69 XThR.Tn[4] 0.21482
R19406 XThR.Tn[4].n64 XThR.Tn[4] 0.21482
R19407 XThR.Tn[4].n59 XThR.Tn[4] 0.21482
R19408 XThR.Tn[4].n54 XThR.Tn[4] 0.21482
R19409 XThR.Tn[4].n49 XThR.Tn[4] 0.21482
R19410 XThR.Tn[4].n44 XThR.Tn[4] 0.21482
R19411 XThR.Tn[4].n39 XThR.Tn[4] 0.21482
R19412 XThR.Tn[4].n34 XThR.Tn[4] 0.21482
R19413 XThR.Tn[4].n29 XThR.Tn[4] 0.21482
R19414 XThR.Tn[4].n24 XThR.Tn[4] 0.21482
R19415 XThR.Tn[4].n19 XThR.Tn[4] 0.21482
R19416 XThR.Tn[4].n14 XThR.Tn[4] 0.21482
R19417 XThR.Tn[4].n85 XThR.Tn[4] 0.0608448
R19418 XThR.Tn[4].n80 XThR.Tn[4] 0.0608448
R19419 XThR.Tn[4].n75 XThR.Tn[4] 0.0608448
R19420 XThR.Tn[4].n70 XThR.Tn[4] 0.0608448
R19421 XThR.Tn[4].n65 XThR.Tn[4] 0.0608448
R19422 XThR.Tn[4].n60 XThR.Tn[4] 0.0608448
R19423 XThR.Tn[4].n55 XThR.Tn[4] 0.0608448
R19424 XThR.Tn[4].n50 XThR.Tn[4] 0.0608448
R19425 XThR.Tn[4].n45 XThR.Tn[4] 0.0608448
R19426 XThR.Tn[4].n40 XThR.Tn[4] 0.0608448
R19427 XThR.Tn[4].n35 XThR.Tn[4] 0.0608448
R19428 XThR.Tn[4].n30 XThR.Tn[4] 0.0608448
R19429 XThR.Tn[4].n25 XThR.Tn[4] 0.0608448
R19430 XThR.Tn[4].n20 XThR.Tn[4] 0.0608448
R19431 XThR.Tn[4].n15 XThR.Tn[4] 0.0608448
R19432 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R19433 XThR.Tn[4] XThR.Tn[4].n87 0.038
R19434 XThR.Tn[4].n11 XThR.Tn[4] 0.00744444
R19435 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00265517
R19436 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00265517
R19437 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00265517
R19438 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00265517
R19439 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00265517
R19440 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00265517
R19441 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00265517
R19442 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00265517
R19443 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00265517
R19444 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00265517
R19445 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00265517
R19446 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00265517
R19447 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00265517
R19448 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00265517
R19449 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00265517
R19450 Vbias.n1 Vbias.t4 651.571
R19451 Vbias.n1 Vbias.t5 651.571
R19452 Vbias.n2 Vbias.t0 651.571
R19453 Vbias.n2 Vbias.t3 651.571
R19454 Vbias.n376 Vbias.t129 119.309
R19455 Vbias.n8 Vbias.t110 119.309
R19456 Vbias.n334 Vbias.t87 119.309
R19457 Vbias.n285 Vbias.t73 119.309
R19458 Vbias.n278 Vbias.t198 119.309
R19459 Vbias.n280 Vbias.t176 119.309
R19460 Vbias.n274 Vbias.t49 119.309
R19461 Vbias.n229 Vbias.t137 119.309
R19462 Vbias.n185 Vbias.t9 119.309
R19463 Vbias.n225 Vbias.t250 119.309
R19464 Vbias.n181 Vbias.t55 119.309
R19465 Vbias.n122 Vbias.t249 119.309
R19466 Vbias.n82 Vbias.t30 119.309
R19467 Vbias.n176 Vbias.t13 119.309
R19468 Vbias.n78 Vbias.t140 119.309
R19469 Vbias.n75 Vbias.t79 119.309
R19470 Vbias.n414 Vbias.t201 119.309
R19471 Vbias.n372 Vbias.t130 119.309
R19472 Vbias.n333 Vbias.t160 119.309
R19473 Vbias.n331 Vbias.t88 119.309
R19474 Vbias.n543 Vbias.t17 119.309
R19475 Vbias.n272 Vbias.t195 119.309
R19476 Vbias.n270 Vbias.t122 119.309
R19477 Vbias.n636 Vbias.t154 119.309
R19478 Vbias.n186 Vbias.t83 119.309
R19479 Vbias.n188 Vbias.t10 119.309
R19480 Vbias.n767 Vbias.t128 119.309
R19481 Vbias.n85 Vbias.t6 119.309
R19482 Vbias.n83 Vbias.t100 119.309
R19483 Vbias.n136 Vbias.t31 119.309
R19484 Vbias.n77 Vbias.t216 119.309
R19485 Vbias.n74 Vbias.t174 119.309
R19486 Vbias.n411 Vbias.t41 119.309
R19487 Vbias.n369 Vbias.t229 119.309
R19488 Vbias.n326 Vbias.t261 119.309
R19489 Vbias.n328 Vbias.t185 119.309
R19490 Vbias.n540 Vbias.t113 119.309
R19491 Vbias.n267 Vbias.t37 119.309
R19492 Vbias.n269 Vbias.t222 119.309
R19493 Vbias.n639 Vbias.t257 119.309
R19494 Vbias.n191 Vbias.t180 119.309
R19495 Vbias.n189 Vbias.t108 119.309
R19496 Vbias.n770 Vbias.t226 119.309
R19497 Vbias.n86 Vbias.t103 119.309
R19498 Vbias.n88 Vbias.t203 119.309
R19499 Vbias.n139 Vbias.t132 119.309
R19500 Vbias.n72 Vbias.t59 119.309
R19501 Vbias.n69 Vbias.t182 119.309
R19502 Vbias.n408 Vbias.t56 119.309
R19503 Vbias.n366 Vbias.t242 119.309
R19504 Vbias.n325 Vbias.t14 119.309
R19505 Vbias.n323 Vbias.t196 119.309
R19506 Vbias.n537 Vbias.t124 119.309
R19507 Vbias.n266 Vbias.t48 119.309
R19508 Vbias.n264 Vbias.t235 119.309
R19509 Vbias.n642 Vbias.t8 119.309
R19510 Vbias.n192 Vbias.t188 119.309
R19511 Vbias.n194 Vbias.t117 119.309
R19512 Vbias.n773 Vbias.t241 119.309
R19513 Vbias.n91 Vbias.t115 119.309
R19514 Vbias.n89 Vbias.t214 119.309
R19515 Vbias.n142 Vbias.t139 119.309
R19516 Vbias.n71 Vbias.t67 119.309
R19517 Vbias.n68 Vbias.t15 119.309
R19518 Vbias.n405 Vbias.t141 119.309
R19519 Vbias.n363 Vbias.t69 119.309
R19520 Vbias.n320 Vbias.t99 119.309
R19521 Vbias.n322 Vbias.t29 119.309
R19522 Vbias.n534 Vbias.t213 119.309
R19523 Vbias.n261 Vbias.t135 119.309
R19524 Vbias.n263 Vbias.t63 119.309
R19525 Vbias.n645 Vbias.t93 119.309
R19526 Vbias.n197 Vbias.t23 119.309
R19527 Vbias.n195 Vbias.t208 119.309
R19528 Vbias.n776 Vbias.t66 119.309
R19529 Vbias.n92 Vbias.t206 119.309
R19530 Vbias.n94 Vbias.t38 119.309
R19531 Vbias.n145 Vbias.t224 119.309
R19532 Vbias.n66 Vbias.t152 119.309
R19533 Vbias.n63 Vbias.t101 119.309
R19534 Vbias.n402 Vbias.t227 119.309
R19535 Vbias.n360 Vbias.t156 119.309
R19536 Vbias.n319 Vbias.t183 119.309
R19537 Vbias.n317 Vbias.t112 119.309
R19538 Vbias.n531 Vbias.t40 119.309
R19539 Vbias.n260 Vbias.t221 119.309
R19540 Vbias.n258 Vbias.t150 119.309
R19541 Vbias.n648 Vbias.t179 119.309
R19542 Vbias.n198 Vbias.t107 119.309
R19543 Vbias.n200 Vbias.t36 119.309
R19544 Vbias.n779 Vbias.t155 119.309
R19545 Vbias.n97 Vbias.t34 119.309
R19546 Vbias.n95 Vbias.t131 119.309
R19547 Vbias.n148 Vbias.t58 119.309
R19548 Vbias.n65 Vbias.t245 119.309
R19549 Vbias.n62 Vbias.t184 119.309
R19550 Vbias.n399 Vbias.t60 119.309
R19551 Vbias.n357 Vbias.t247 119.309
R19552 Vbias.n314 Vbias.t18 119.309
R19553 Vbias.n316 Vbias.t200 119.309
R19554 Vbias.n528 Vbias.t127 119.309
R19555 Vbias.n255 Vbias.t50 119.309
R19556 Vbias.n257 Vbias.t237 119.309
R19557 Vbias.n651 Vbias.t11 119.309
R19558 Vbias.n203 Vbias.t192 119.309
R19559 Vbias.n201 Vbias.t120 119.309
R19560 Vbias.n782 Vbias.t244 119.309
R19561 Vbias.n98 Vbias.t116 119.309
R19562 Vbias.n100 Vbias.t218 119.309
R19563 Vbias.n151 Vbias.t145 119.309
R19564 Vbias.n60 Vbias.t72 119.309
R19565 Vbias.n57 Vbias.t19 119.309
R19566 Vbias.n396 Vbias.t147 119.309
R19567 Vbias.n354 Vbias.t76 119.309
R19568 Vbias.n313 Vbias.t102 119.309
R19569 Vbias.n311 Vbias.t33 119.309
R19570 Vbias.n525 Vbias.t219 119.309
R19571 Vbias.n254 Vbias.t138 119.309
R19572 Vbias.n252 Vbias.t68 119.309
R19573 Vbias.n654 Vbias.t98 119.309
R19574 Vbias.n204 Vbias.t28 119.309
R19575 Vbias.n206 Vbias.t212 119.309
R19576 Vbias.n785 Vbias.t74 119.309
R19577 Vbias.n103 Vbias.t209 119.309
R19578 Vbias.n101 Vbias.t42 119.309
R19579 Vbias.n154 Vbias.t230 119.309
R19580 Vbias.n59 Vbias.t158 119.309
R19581 Vbias.n56 Vbias.t39 119.309
R19582 Vbias.n393 Vbias.t169 119.309
R19583 Vbias.n351 Vbias.t96 119.309
R19584 Vbias.n308 Vbias.t125 119.309
R19585 Vbias.n310 Vbias.t53 119.309
R19586 Vbias.n522 Vbias.t240 119.309
R19587 Vbias.n249 Vbias.t163 119.309
R19588 Vbias.n251 Vbias.t91 119.309
R19589 Vbias.n657 Vbias.t118 119.309
R19590 Vbias.n209 Vbias.t45 119.309
R19591 Vbias.n207 Vbias.t234 119.309
R19592 Vbias.n788 Vbias.t94 119.309
R19593 Vbias.n104 Vbias.t231 119.309
R19594 Vbias.n106 Vbias.t70 119.309
R19595 Vbias.n157 Vbias.t253 119.309
R19596 Vbias.n54 Vbias.t178 119.309
R19597 Vbias.n51 Vbias.t111 119.309
R19598 Vbias.n390 Vbias.t246 119.309
R19599 Vbias.n348 Vbias.t171 119.309
R19600 Vbias.n307 Vbias.t199 119.309
R19601 Vbias.n305 Vbias.t126 119.309
R19602 Vbias.n519 Vbias.t54 119.309
R19603 Vbias.n248 Vbias.t236 119.309
R19604 Vbias.n246 Vbias.t164 119.309
R19605 Vbias.n660 Vbias.t190 119.309
R19606 Vbias.n210 Vbias.t119 119.309
R19607 Vbias.n212 Vbias.t46 119.309
R19608 Vbias.n791 Vbias.t167 119.309
R19609 Vbias.n109 Vbias.t43 119.309
R19610 Vbias.n107 Vbias.t143 119.309
R19611 Vbias.n160 Vbias.t71 119.309
R19612 Vbias.n53 Vbias.t254 119.309
R19613 Vbias.n50 Vbias.t202 119.309
R19614 Vbias.n387 Vbias.t75 119.309
R19615 Vbias.n345 Vbias.t258 119.309
R19616 Vbias.n302 Vbias.t32 119.309
R19617 Vbias.n304 Vbias.t217 119.309
R19618 Vbias.n516 Vbias.t144 119.309
R19619 Vbias.n243 Vbias.t65 119.309
R19620 Vbias.n245 Vbias.t251 119.309
R19621 Vbias.n663 Vbias.t27 119.309
R19622 Vbias.n215 Vbias.t211 119.309
R19623 Vbias.n213 Vbias.t136 119.309
R19624 Vbias.n794 Vbias.t256 119.309
R19625 Vbias.n110 Vbias.t134 119.309
R19626 Vbias.n112 Vbias.t228 119.309
R19627 Vbias.n163 Vbias.t157 119.309
R19628 Vbias.n48 Vbias.t84 119.309
R19629 Vbias.n45 Vbias.t223 119.309
R19630 Vbias.n384 Vbias.t95 119.309
R19631 Vbias.n342 Vbias.t25 119.309
R19632 Vbias.n301 Vbias.t52 119.309
R19633 Vbias.n299 Vbias.t239 119.309
R19634 Vbias.n513 Vbias.t166 119.309
R19635 Vbias.n242 Vbias.t90 119.309
R19636 Vbias.n240 Vbias.t21 119.309
R19637 Vbias.n666 Vbias.t44 119.309
R19638 Vbias.n216 Vbias.t233 119.309
R19639 Vbias.n218 Vbias.t162 119.309
R19640 Vbias.n797 Vbias.t22 119.309
R19641 Vbias.n115 Vbias.t159 119.309
R19642 Vbias.n113 Vbias.t252 119.309
R19643 Vbias.n166 Vbias.t177 119.309
R19644 Vbias.n47 Vbias.t106 119.309
R19645 Vbias.n44 Vbias.t114 119.309
R19646 Vbias.n381 Vbias.t248 119.309
R19647 Vbias.n339 Vbias.t173 119.309
R19648 Vbias.n296 Vbias.t205 119.309
R19649 Vbias.n298 Vbias.t133 119.309
R19650 Vbias.n510 Vbias.t62 119.309
R19651 Vbias.n237 Vbias.t243 119.309
R19652 Vbias.n239 Vbias.t168 119.309
R19653 Vbias.n669 Vbias.t197 119.309
R19654 Vbias.n221 Vbias.t123 119.309
R19655 Vbias.n219 Vbias.t51 119.309
R19656 Vbias.n800 Vbias.t172 119.309
R19657 Vbias.n116 Vbias.t47 119.309
R19658 Vbias.n118 Vbias.t148 119.309
R19659 Vbias.n169 Vbias.t77 119.309
R19660 Vbias.n42 Vbias.t259 119.309
R19661 Vbias.n39 Vbias.t142 119.309
R19662 Vbias.n378 Vbias.t12 119.309
R19663 Vbias.n336 Vbias.t193 119.309
R19664 Vbias.n288 Vbias.t225 119.309
R19665 Vbias.n286 Vbias.t153 119.309
R19666 Vbias.n507 Vbias.t81 119.309
R19667 Vbias.n236 Vbias.t7 119.309
R19668 Vbias.n234 Vbias.t187 119.309
R19669 Vbias.n672 Vbias.t220 119.309
R19670 Vbias.n222 Vbias.t149 119.309
R19671 Vbias.n224 Vbias.t80 119.309
R19672 Vbias.n803 Vbias.t191 119.309
R19673 Vbias.n121 Vbias.t78 119.309
R19674 Vbias.n119 Vbias.t170 119.309
R19675 Vbias.n172 Vbias.t97 119.309
R19676 Vbias.n41 Vbias.t26 119.309
R19677 Vbias.n38 Vbias.t151 119.309
R19678 Vbias.n10 Vbias.t24 119.309
R19679 Vbias.n9 Vbias.t210 119.309
R19680 Vbias.n12 Vbias.t238 119.309
R19681 Vbias.n14 Vbias.t165 119.309
R19682 Vbias.n16 Vbias.t92 119.309
R19683 Vbias.n18 Vbias.t20 119.309
R19684 Vbias.n20 Vbias.t204 119.309
R19685 Vbias.n22 Vbias.t232 119.309
R19686 Vbias.n24 Vbias.t161 119.309
R19687 Vbias.n26 Vbias.t89 119.309
R19688 Vbias.n28 Vbias.t207 119.309
R19689 Vbias.n30 Vbias.t85 119.309
R19690 Vbias.n32 Vbias.t175 119.309
R19691 Vbias.n34 Vbias.t104 119.309
R19692 Vbias.n36 Vbias.t35 119.309
R19693 Vbias.n129 Vbias.t61 119.309
R19694 Vbias.n904 Vbias.t260 119.309
R19695 Vbias.n128 Vbias.t194 119.309
R19696 Vbias.n79 Vbias.t215 119.309
R19697 Vbias.n125 Vbias.t86 119.309
R19698 Vbias.n893 Vbias.t186 119.309
R19699 Vbias.n807 Vbias.t109 119.309
R19700 Vbias.n182 Vbias.t189 119.309
R19701 Vbias.n226 Vbias.t64 119.309
R19702 Vbias.n634 Vbias.t82 119.309
R19703 Vbias.n629 Vbias.t105 119.309
R19704 Vbias.n273 Vbias.t121 119.309
R19705 Vbias.n279 Vbias.t255 119.309
R19706 Vbias.n329 Vbias.t16 119.309
R19707 Vbias.n292 Vbias.t146 119.309
R19708 Vbias.n6 Vbias.t181 119.309
R19709 Vbias.n335 Vbias.t57 119.309
R19710 Vbias.n0 Vbias.t1 77.1834
R19711 Vbias.n0 Vbias.t2 34.3787
R19712 Vbias.n3 Vbias.n1 4.78773
R19713 Vbias.n3 Vbias.n2 4.78773
R19714 Vbias.n415 Vbias.n414 4.5005
R19715 Vbias.n373 Vbias.n372 4.5005
R19716 Vbias.n422 Vbias.n333 4.5005
R19717 Vbias.n425 Vbias.n331 4.5005
R19718 Vbias.n544 Vbias.n543 4.5005
R19719 Vbias.n551 Vbias.n272 4.5005
R19720 Vbias.n554 Vbias.n270 4.5005
R19721 Vbias.n637 Vbias.n636 4.5005
R19722 Vbias.n760 Vbias.n186 4.5005
R19723 Vbias.n757 Vbias.n188 4.5005
R19724 Vbias.n768 Vbias.n767 4.5005
R19725 Vbias.n896 Vbias.n85 4.5005
R19726 Vbias.n899 Vbias.n83 4.5005
R19727 Vbias.n137 Vbias.n136 4.5005
R19728 Vbias.n909 Vbias.n77 4.5005
R19729 Vbias.n911 Vbias.n75 4.5005
R19730 Vbias.n412 Vbias.n411 4.5005
R19731 Vbias.n370 Vbias.n369 4.5005
R19732 Vbias.n431 Vbias.n326 4.5005
R19733 Vbias.n428 Vbias.n328 4.5005
R19734 Vbias.n541 Vbias.n540 4.5005
R19735 Vbias.n560 Vbias.n267 4.5005
R19736 Vbias.n557 Vbias.n269 4.5005
R19737 Vbias.n640 Vbias.n639 4.5005
R19738 Vbias.n751 Vbias.n191 4.5005
R19739 Vbias.n754 Vbias.n189 4.5005
R19740 Vbias.n771 Vbias.n770 4.5005
R19741 Vbias.n891 Vbias.n86 4.5005
R19742 Vbias.n888 Vbias.n88 4.5005
R19743 Vbias.n140 Vbias.n139 4.5005
R19744 Vbias.n916 Vbias.n72 4.5005
R19745 Vbias.n914 Vbias.n74 4.5005
R19746 Vbias.n409 Vbias.n408 4.5005
R19747 Vbias.n367 Vbias.n366 4.5005
R19748 Vbias.n434 Vbias.n325 4.5005
R19749 Vbias.n437 Vbias.n323 4.5005
R19750 Vbias.n538 Vbias.n537 4.5005
R19751 Vbias.n563 Vbias.n266 4.5005
R19752 Vbias.n566 Vbias.n264 4.5005
R19753 Vbias.n643 Vbias.n642 4.5005
R19754 Vbias.n748 Vbias.n192 4.5005
R19755 Vbias.n745 Vbias.n194 4.5005
R19756 Vbias.n774 Vbias.n773 4.5005
R19757 Vbias.n882 Vbias.n91 4.5005
R19758 Vbias.n885 Vbias.n89 4.5005
R19759 Vbias.n143 Vbias.n142 4.5005
R19760 Vbias.n919 Vbias.n71 4.5005
R19761 Vbias.n921 Vbias.n69 4.5005
R19762 Vbias.n406 Vbias.n405 4.5005
R19763 Vbias.n364 Vbias.n363 4.5005
R19764 Vbias.n443 Vbias.n320 4.5005
R19765 Vbias.n440 Vbias.n322 4.5005
R19766 Vbias.n535 Vbias.n534 4.5005
R19767 Vbias.n572 Vbias.n261 4.5005
R19768 Vbias.n569 Vbias.n263 4.5005
R19769 Vbias.n646 Vbias.n645 4.5005
R19770 Vbias.n739 Vbias.n197 4.5005
R19771 Vbias.n742 Vbias.n195 4.5005
R19772 Vbias.n777 Vbias.n776 4.5005
R19773 Vbias.n879 Vbias.n92 4.5005
R19774 Vbias.n876 Vbias.n94 4.5005
R19775 Vbias.n146 Vbias.n145 4.5005
R19776 Vbias.n926 Vbias.n66 4.5005
R19777 Vbias.n924 Vbias.n68 4.5005
R19778 Vbias.n403 Vbias.n402 4.5005
R19779 Vbias.n361 Vbias.n360 4.5005
R19780 Vbias.n446 Vbias.n319 4.5005
R19781 Vbias.n449 Vbias.n317 4.5005
R19782 Vbias.n532 Vbias.n531 4.5005
R19783 Vbias.n575 Vbias.n260 4.5005
R19784 Vbias.n578 Vbias.n258 4.5005
R19785 Vbias.n649 Vbias.n648 4.5005
R19786 Vbias.n736 Vbias.n198 4.5005
R19787 Vbias.n733 Vbias.n200 4.5005
R19788 Vbias.n780 Vbias.n779 4.5005
R19789 Vbias.n870 Vbias.n97 4.5005
R19790 Vbias.n873 Vbias.n95 4.5005
R19791 Vbias.n149 Vbias.n148 4.5005
R19792 Vbias.n929 Vbias.n65 4.5005
R19793 Vbias.n931 Vbias.n63 4.5005
R19794 Vbias.n400 Vbias.n399 4.5005
R19795 Vbias.n358 Vbias.n357 4.5005
R19796 Vbias.n455 Vbias.n314 4.5005
R19797 Vbias.n452 Vbias.n316 4.5005
R19798 Vbias.n529 Vbias.n528 4.5005
R19799 Vbias.n584 Vbias.n255 4.5005
R19800 Vbias.n581 Vbias.n257 4.5005
R19801 Vbias.n652 Vbias.n651 4.5005
R19802 Vbias.n727 Vbias.n203 4.5005
R19803 Vbias.n730 Vbias.n201 4.5005
R19804 Vbias.n783 Vbias.n782 4.5005
R19805 Vbias.n867 Vbias.n98 4.5005
R19806 Vbias.n864 Vbias.n100 4.5005
R19807 Vbias.n152 Vbias.n151 4.5005
R19808 Vbias.n936 Vbias.n60 4.5005
R19809 Vbias.n934 Vbias.n62 4.5005
R19810 Vbias.n397 Vbias.n396 4.5005
R19811 Vbias.n355 Vbias.n354 4.5005
R19812 Vbias.n458 Vbias.n313 4.5005
R19813 Vbias.n461 Vbias.n311 4.5005
R19814 Vbias.n526 Vbias.n525 4.5005
R19815 Vbias.n587 Vbias.n254 4.5005
R19816 Vbias.n590 Vbias.n252 4.5005
R19817 Vbias.n655 Vbias.n654 4.5005
R19818 Vbias.n724 Vbias.n204 4.5005
R19819 Vbias.n721 Vbias.n206 4.5005
R19820 Vbias.n786 Vbias.n785 4.5005
R19821 Vbias.n858 Vbias.n103 4.5005
R19822 Vbias.n861 Vbias.n101 4.5005
R19823 Vbias.n155 Vbias.n154 4.5005
R19824 Vbias.n939 Vbias.n59 4.5005
R19825 Vbias.n941 Vbias.n57 4.5005
R19826 Vbias.n394 Vbias.n393 4.5005
R19827 Vbias.n352 Vbias.n351 4.5005
R19828 Vbias.n467 Vbias.n308 4.5005
R19829 Vbias.n464 Vbias.n310 4.5005
R19830 Vbias.n523 Vbias.n522 4.5005
R19831 Vbias.n596 Vbias.n249 4.5005
R19832 Vbias.n593 Vbias.n251 4.5005
R19833 Vbias.n658 Vbias.n657 4.5005
R19834 Vbias.n715 Vbias.n209 4.5005
R19835 Vbias.n718 Vbias.n207 4.5005
R19836 Vbias.n789 Vbias.n788 4.5005
R19837 Vbias.n855 Vbias.n104 4.5005
R19838 Vbias.n852 Vbias.n106 4.5005
R19839 Vbias.n158 Vbias.n157 4.5005
R19840 Vbias.n946 Vbias.n54 4.5005
R19841 Vbias.n944 Vbias.n56 4.5005
R19842 Vbias.n391 Vbias.n390 4.5005
R19843 Vbias.n349 Vbias.n348 4.5005
R19844 Vbias.n470 Vbias.n307 4.5005
R19845 Vbias.n473 Vbias.n305 4.5005
R19846 Vbias.n520 Vbias.n519 4.5005
R19847 Vbias.n599 Vbias.n248 4.5005
R19848 Vbias.n602 Vbias.n246 4.5005
R19849 Vbias.n661 Vbias.n660 4.5005
R19850 Vbias.n712 Vbias.n210 4.5005
R19851 Vbias.n709 Vbias.n212 4.5005
R19852 Vbias.n792 Vbias.n791 4.5005
R19853 Vbias.n846 Vbias.n109 4.5005
R19854 Vbias.n849 Vbias.n107 4.5005
R19855 Vbias.n161 Vbias.n160 4.5005
R19856 Vbias.n949 Vbias.n53 4.5005
R19857 Vbias.n951 Vbias.n51 4.5005
R19858 Vbias.n388 Vbias.n387 4.5005
R19859 Vbias.n346 Vbias.n345 4.5005
R19860 Vbias.n479 Vbias.n302 4.5005
R19861 Vbias.n476 Vbias.n304 4.5005
R19862 Vbias.n517 Vbias.n516 4.5005
R19863 Vbias.n608 Vbias.n243 4.5005
R19864 Vbias.n605 Vbias.n245 4.5005
R19865 Vbias.n664 Vbias.n663 4.5005
R19866 Vbias.n703 Vbias.n215 4.5005
R19867 Vbias.n706 Vbias.n213 4.5005
R19868 Vbias.n795 Vbias.n794 4.5005
R19869 Vbias.n843 Vbias.n110 4.5005
R19870 Vbias.n840 Vbias.n112 4.5005
R19871 Vbias.n164 Vbias.n163 4.5005
R19872 Vbias.n956 Vbias.n48 4.5005
R19873 Vbias.n954 Vbias.n50 4.5005
R19874 Vbias.n385 Vbias.n384 4.5005
R19875 Vbias.n343 Vbias.n342 4.5005
R19876 Vbias.n482 Vbias.n301 4.5005
R19877 Vbias.n485 Vbias.n299 4.5005
R19878 Vbias.n514 Vbias.n513 4.5005
R19879 Vbias.n611 Vbias.n242 4.5005
R19880 Vbias.n614 Vbias.n240 4.5005
R19881 Vbias.n667 Vbias.n666 4.5005
R19882 Vbias.n700 Vbias.n216 4.5005
R19883 Vbias.n697 Vbias.n218 4.5005
R19884 Vbias.n798 Vbias.n797 4.5005
R19885 Vbias.n834 Vbias.n115 4.5005
R19886 Vbias.n837 Vbias.n113 4.5005
R19887 Vbias.n167 Vbias.n166 4.5005
R19888 Vbias.n959 Vbias.n47 4.5005
R19889 Vbias.n961 Vbias.n45 4.5005
R19890 Vbias.n382 Vbias.n381 4.5005
R19891 Vbias.n340 Vbias.n339 4.5005
R19892 Vbias.n491 Vbias.n296 4.5005
R19893 Vbias.n488 Vbias.n298 4.5005
R19894 Vbias.n511 Vbias.n510 4.5005
R19895 Vbias.n620 Vbias.n237 4.5005
R19896 Vbias.n617 Vbias.n239 4.5005
R19897 Vbias.n670 Vbias.n669 4.5005
R19898 Vbias.n691 Vbias.n221 4.5005
R19899 Vbias.n694 Vbias.n219 4.5005
R19900 Vbias.n801 Vbias.n800 4.5005
R19901 Vbias.n831 Vbias.n116 4.5005
R19902 Vbias.n828 Vbias.n118 4.5005
R19903 Vbias.n170 Vbias.n169 4.5005
R19904 Vbias.n966 Vbias.n42 4.5005
R19905 Vbias.n964 Vbias.n44 4.5005
R19906 Vbias.n379 Vbias.n378 4.5005
R19907 Vbias.n337 Vbias.n336 4.5005
R19908 Vbias.n494 Vbias.n288 4.5005
R19909 Vbias.n497 Vbias.n286 4.5005
R19910 Vbias.n508 Vbias.n507 4.5005
R19911 Vbias.n623 Vbias.n236 4.5005
R19912 Vbias.n626 Vbias.n234 4.5005
R19913 Vbias.n673 Vbias.n672 4.5005
R19914 Vbias.n688 Vbias.n222 4.5005
R19915 Vbias.n685 Vbias.n224 4.5005
R19916 Vbias.n804 Vbias.n803 4.5005
R19917 Vbias.n822 Vbias.n121 4.5005
R19918 Vbias.n825 Vbias.n119 4.5005
R19919 Vbias.n173 Vbias.n172 4.5005
R19920 Vbias.n969 Vbias.n41 4.5005
R19921 Vbias.n971 Vbias.n39 4.5005
R19922 Vbias.n11 Vbias.n10 4.5005
R19923 Vbias.n989 Vbias.n9 4.5005
R19924 Vbias.n13 Vbias.n12 4.5005
R19925 Vbias.n15 Vbias.n14 4.5005
R19926 Vbias.n17 Vbias.n16 4.5005
R19927 Vbias.n19 Vbias.n18 4.5005
R19928 Vbias.n21 Vbias.n20 4.5005
R19929 Vbias.n23 Vbias.n22 4.5005
R19930 Vbias.n25 Vbias.n24 4.5005
R19931 Vbias.n27 Vbias.n26 4.5005
R19932 Vbias.n29 Vbias.n28 4.5005
R19933 Vbias.n31 Vbias.n30 4.5005
R19934 Vbias.n33 Vbias.n32 4.5005
R19935 Vbias.n35 Vbias.n34 4.5005
R19936 Vbias.n37 Vbias.n36 4.5005
R19937 Vbias.n974 Vbias.n38 4.5005
R19938 Vbias.n131 Vbias.n129 4.5005
R19939 Vbias.n905 Vbias.n904 4.5005
R19940 Vbias.n907 Vbias.n78 4.5005
R19941 Vbias.n133 Vbias.n128 4.5005
R19942 Vbias.n177 Vbias.n176 4.5005
R19943 Vbias.n80 Vbias.n79 4.5005
R19944 Vbias.n901 Vbias.n82 4.5005
R19945 Vbias.n815 Vbias.n125 4.5005
R19946 Vbias.n818 Vbias.n122 4.5005
R19947 Vbias.n894 Vbias.n893 4.5005
R19948 Vbias.n766 Vbias.n181 4.5005
R19949 Vbias.n808 Vbias.n807 4.5005
R19950 Vbias.n681 Vbias.n225 4.5005
R19951 Vbias.n183 Vbias.n182 4.5005
R19952 Vbias.n762 Vbias.n185 4.5005
R19953 Vbias.n227 Vbias.n226 4.5005
R19954 Vbias.n677 Vbias.n229 4.5005
R19955 Vbias.n635 Vbias.n634 4.5005
R19956 Vbias.n275 Vbias.n274 4.5005
R19957 Vbias.n630 Vbias.n629 4.5005
R19958 Vbias.n283 Vbias.n280 4.5005
R19959 Vbias.n549 Vbias.n273 4.5005
R19960 Vbias.n546 Vbias.n278 4.5005
R19961 Vbias.n504 Vbias.n279 4.5005
R19962 Vbias.n501 Vbias.n285 4.5005
R19963 Vbias.n330 Vbias.n329 4.5005
R19964 Vbias.n420 Vbias.n334 4.5005
R19965 Vbias.n293 Vbias.n292 4.5005
R19966 Vbias.n994 Vbias.n6 4.5005
R19967 Vbias.n992 Vbias.n8 4.5005
R19968 Vbias.n375 Vbias.n335 4.5005
R19969 Vbias.n417 Vbias.n376 4.5005
R19970 Vbias Vbias.n291 3.95257
R19971 Vbias.n289 Vbias 3.95257
R19972 Vbias.n632 Vbias 3.95257
R19973 Vbias.n232 Vbias 3.95257
R19974 Vbias.n810 Vbias 3.95257
R19975 Vbias Vbias.n812 3.95257
R19976 Vbias.n135 Vbias 3.95257
R19977 Vbias Vbias.n126 3.95257
R19978 Vbias.n179 Vbias 3.95257
R19979 Vbias.n811 Vbias 3.95257
R19980 Vbias Vbias.n180 3.95257
R19981 Vbias Vbias.n633 3.95257
R19982 Vbias Vbias.n233 3.95257
R19983 Vbias.n290 Vbias 3.95257
R19984 Vbias Vbias.n5 3.95257
R19985 Vbias.n996 Vbias 3.95257
R19986 Vbias.n905 Vbias 3.50727
R19987 Vbias Vbias.n907 3.50727
R19988 Vbias Vbias.n80 3.50727
R19989 Vbias.n901 Vbias 3.50727
R19990 Vbias Vbias.n894 3.50727
R19991 Vbias Vbias.n766 3.50727
R19992 Vbias Vbias.n183 3.50727
R19993 Vbias.n762 Vbias 3.50727
R19994 Vbias Vbias.n635 3.50727
R19995 Vbias.n275 Vbias 3.50727
R19996 Vbias Vbias.n549 3.50727
R19997 Vbias.n546 Vbias 3.50727
R19998 Vbias Vbias.n330 3.50727
R19999 Vbias Vbias.n420 3.50727
R20000 Vbias.n375 Vbias 3.50727
R20001 Vbias.n417 Vbias 3.50727
R20002 Vbias.n131 Vbias.n130 3.4105
R20003 Vbias.n974 Vbias.n973 3.4105
R20004 Vbias.n972 Vbias.n971 3.4105
R20005 Vbias.n964 Vbias.n963 3.4105
R20006 Vbias.n962 Vbias.n961 3.4105
R20007 Vbias.n954 Vbias.n953 3.4105
R20008 Vbias.n952 Vbias.n951 3.4105
R20009 Vbias.n944 Vbias.n943 3.4105
R20010 Vbias.n942 Vbias.n941 3.4105
R20011 Vbias.n934 Vbias.n933 3.4105
R20012 Vbias.n932 Vbias.n931 3.4105
R20013 Vbias.n924 Vbias.n923 3.4105
R20014 Vbias.n922 Vbias.n921 3.4105
R20015 Vbias.n914 Vbias.n913 3.4105
R20016 Vbias.n912 Vbias.n911 3.4105
R20017 Vbias.n909 Vbias.n908 3.4105
R20018 Vbias.n917 Vbias.n916 3.4105
R20019 Vbias.n919 Vbias.n918 3.4105
R20020 Vbias.n927 Vbias.n926 3.4105
R20021 Vbias.n929 Vbias.n928 3.4105
R20022 Vbias.n937 Vbias.n936 3.4105
R20023 Vbias.n939 Vbias.n938 3.4105
R20024 Vbias.n947 Vbias.n946 3.4105
R20025 Vbias.n949 Vbias.n948 3.4105
R20026 Vbias.n957 Vbias.n956 3.4105
R20027 Vbias.n959 Vbias.n958 3.4105
R20028 Vbias.n967 Vbias.n966 3.4105
R20029 Vbias.n969 Vbias.n968 3.4105
R20030 Vbias.n127 Vbias.n37 3.4105
R20031 Vbias.n134 Vbias.n133 3.4105
R20032 Vbias.n178 Vbias.n177 3.4105
R20033 Vbias.n175 Vbias.n35 3.4105
R20034 Vbias.n174 Vbias.n173 3.4105
R20035 Vbias.n171 Vbias.n170 3.4105
R20036 Vbias.n168 Vbias.n167 3.4105
R20037 Vbias.n165 Vbias.n164 3.4105
R20038 Vbias.n162 Vbias.n161 3.4105
R20039 Vbias.n159 Vbias.n158 3.4105
R20040 Vbias.n156 Vbias.n155 3.4105
R20041 Vbias.n153 Vbias.n152 3.4105
R20042 Vbias.n150 Vbias.n149 3.4105
R20043 Vbias.n147 Vbias.n146 3.4105
R20044 Vbias.n144 Vbias.n143 3.4105
R20045 Vbias.n141 Vbias.n140 3.4105
R20046 Vbias.n138 Vbias.n137 3.4105
R20047 Vbias.n900 Vbias.n899 3.4105
R20048 Vbias.n888 Vbias.n887 3.4105
R20049 Vbias.n886 Vbias.n885 3.4105
R20050 Vbias.n876 Vbias.n875 3.4105
R20051 Vbias.n874 Vbias.n873 3.4105
R20052 Vbias.n864 Vbias.n863 3.4105
R20053 Vbias.n862 Vbias.n861 3.4105
R20054 Vbias.n852 Vbias.n851 3.4105
R20055 Vbias.n850 Vbias.n849 3.4105
R20056 Vbias.n840 Vbias.n839 3.4105
R20057 Vbias.n838 Vbias.n837 3.4105
R20058 Vbias.n828 Vbias.n827 3.4105
R20059 Vbias.n826 Vbias.n825 3.4105
R20060 Vbias.n813 Vbias.n33 3.4105
R20061 Vbias.n815 Vbias.n814 3.4105
R20062 Vbias.n819 Vbias.n818 3.4105
R20063 Vbias.n820 Vbias.n31 3.4105
R20064 Vbias.n822 Vbias.n821 3.4105
R20065 Vbias.n832 Vbias.n831 3.4105
R20066 Vbias.n834 Vbias.n833 3.4105
R20067 Vbias.n844 Vbias.n843 3.4105
R20068 Vbias.n846 Vbias.n845 3.4105
R20069 Vbias.n856 Vbias.n855 3.4105
R20070 Vbias.n858 Vbias.n857 3.4105
R20071 Vbias.n868 Vbias.n867 3.4105
R20072 Vbias.n870 Vbias.n869 3.4105
R20073 Vbias.n880 Vbias.n879 3.4105
R20074 Vbias.n882 Vbias.n881 3.4105
R20075 Vbias.n892 Vbias.n891 3.4105
R20076 Vbias.n896 Vbias.n895 3.4105
R20077 Vbias.n769 Vbias.n768 3.4105
R20078 Vbias.n772 Vbias.n771 3.4105
R20079 Vbias.n775 Vbias.n774 3.4105
R20080 Vbias.n778 Vbias.n777 3.4105
R20081 Vbias.n781 Vbias.n780 3.4105
R20082 Vbias.n784 Vbias.n783 3.4105
R20083 Vbias.n787 Vbias.n786 3.4105
R20084 Vbias.n790 Vbias.n789 3.4105
R20085 Vbias.n793 Vbias.n792 3.4105
R20086 Vbias.n796 Vbias.n795 3.4105
R20087 Vbias.n799 Vbias.n798 3.4105
R20088 Vbias.n802 Vbias.n801 3.4105
R20089 Vbias.n805 Vbias.n804 3.4105
R20090 Vbias.n806 Vbias.n29 3.4105
R20091 Vbias.n809 Vbias.n808 3.4105
R20092 Vbias.n682 Vbias.n681 3.4105
R20093 Vbias.n683 Vbias.n27 3.4105
R20094 Vbias.n685 Vbias.n684 3.4105
R20095 Vbias.n695 Vbias.n694 3.4105
R20096 Vbias.n697 Vbias.n696 3.4105
R20097 Vbias.n707 Vbias.n706 3.4105
R20098 Vbias.n709 Vbias.n708 3.4105
R20099 Vbias.n719 Vbias.n718 3.4105
R20100 Vbias.n721 Vbias.n720 3.4105
R20101 Vbias.n731 Vbias.n730 3.4105
R20102 Vbias.n733 Vbias.n732 3.4105
R20103 Vbias.n743 Vbias.n742 3.4105
R20104 Vbias.n745 Vbias.n744 3.4105
R20105 Vbias.n755 Vbias.n754 3.4105
R20106 Vbias.n757 Vbias.n756 3.4105
R20107 Vbias.n761 Vbias.n760 3.4105
R20108 Vbias.n751 Vbias.n750 3.4105
R20109 Vbias.n749 Vbias.n748 3.4105
R20110 Vbias.n739 Vbias.n738 3.4105
R20111 Vbias.n737 Vbias.n736 3.4105
R20112 Vbias.n727 Vbias.n726 3.4105
R20113 Vbias.n725 Vbias.n724 3.4105
R20114 Vbias.n715 Vbias.n714 3.4105
R20115 Vbias.n713 Vbias.n712 3.4105
R20116 Vbias.n703 Vbias.n702 3.4105
R20117 Vbias.n701 Vbias.n700 3.4105
R20118 Vbias.n691 Vbias.n690 3.4105
R20119 Vbias.n689 Vbias.n688 3.4105
R20120 Vbias.n230 Vbias.n25 3.4105
R20121 Vbias.n231 Vbias.n227 3.4105
R20122 Vbias.n677 Vbias.n676 3.4105
R20123 Vbias.n675 Vbias.n23 3.4105
R20124 Vbias.n674 Vbias.n673 3.4105
R20125 Vbias.n671 Vbias.n670 3.4105
R20126 Vbias.n668 Vbias.n667 3.4105
R20127 Vbias.n665 Vbias.n664 3.4105
R20128 Vbias.n662 Vbias.n661 3.4105
R20129 Vbias.n659 Vbias.n658 3.4105
R20130 Vbias.n656 Vbias.n655 3.4105
R20131 Vbias.n653 Vbias.n652 3.4105
R20132 Vbias.n650 Vbias.n649 3.4105
R20133 Vbias.n647 Vbias.n646 3.4105
R20134 Vbias.n644 Vbias.n643 3.4105
R20135 Vbias.n641 Vbias.n640 3.4105
R20136 Vbias.n638 Vbias.n637 3.4105
R20137 Vbias.n555 Vbias.n554 3.4105
R20138 Vbias.n557 Vbias.n556 3.4105
R20139 Vbias.n567 Vbias.n566 3.4105
R20140 Vbias.n569 Vbias.n568 3.4105
R20141 Vbias.n579 Vbias.n578 3.4105
R20142 Vbias.n581 Vbias.n580 3.4105
R20143 Vbias.n591 Vbias.n590 3.4105
R20144 Vbias.n593 Vbias.n592 3.4105
R20145 Vbias.n603 Vbias.n602 3.4105
R20146 Vbias.n605 Vbias.n604 3.4105
R20147 Vbias.n615 Vbias.n614 3.4105
R20148 Vbias.n617 Vbias.n616 3.4105
R20149 Vbias.n627 Vbias.n626 3.4105
R20150 Vbias.n628 Vbias.n21 3.4105
R20151 Vbias.n631 Vbias.n630 3.4105
R20152 Vbias.n283 Vbias.n282 3.4105
R20153 Vbias.n281 Vbias.n19 3.4105
R20154 Vbias.n623 Vbias.n622 3.4105
R20155 Vbias.n621 Vbias.n620 3.4105
R20156 Vbias.n611 Vbias.n610 3.4105
R20157 Vbias.n609 Vbias.n608 3.4105
R20158 Vbias.n599 Vbias.n598 3.4105
R20159 Vbias.n597 Vbias.n596 3.4105
R20160 Vbias.n587 Vbias.n586 3.4105
R20161 Vbias.n585 Vbias.n584 3.4105
R20162 Vbias.n575 Vbias.n574 3.4105
R20163 Vbias.n573 Vbias.n572 3.4105
R20164 Vbias.n563 Vbias.n562 3.4105
R20165 Vbias.n561 Vbias.n560 3.4105
R20166 Vbias.n551 Vbias.n550 3.4105
R20167 Vbias.n545 Vbias.n544 3.4105
R20168 Vbias.n542 Vbias.n541 3.4105
R20169 Vbias.n539 Vbias.n538 3.4105
R20170 Vbias.n536 Vbias.n535 3.4105
R20171 Vbias.n533 Vbias.n532 3.4105
R20172 Vbias.n530 Vbias.n529 3.4105
R20173 Vbias.n527 Vbias.n526 3.4105
R20174 Vbias.n524 Vbias.n523 3.4105
R20175 Vbias.n521 Vbias.n520 3.4105
R20176 Vbias.n518 Vbias.n517 3.4105
R20177 Vbias.n515 Vbias.n514 3.4105
R20178 Vbias.n512 Vbias.n511 3.4105
R20179 Vbias.n509 Vbias.n508 3.4105
R20180 Vbias.n506 Vbias.n17 3.4105
R20181 Vbias.n505 Vbias.n504 3.4105
R20182 Vbias.n501 Vbias.n500 3.4105
R20183 Vbias.n499 Vbias.n15 3.4105
R20184 Vbias.n498 Vbias.n497 3.4105
R20185 Vbias.n488 Vbias.n487 3.4105
R20186 Vbias.n486 Vbias.n485 3.4105
R20187 Vbias.n476 Vbias.n475 3.4105
R20188 Vbias.n474 Vbias.n473 3.4105
R20189 Vbias.n464 Vbias.n463 3.4105
R20190 Vbias.n462 Vbias.n461 3.4105
R20191 Vbias.n452 Vbias.n451 3.4105
R20192 Vbias.n450 Vbias.n449 3.4105
R20193 Vbias.n440 Vbias.n439 3.4105
R20194 Vbias.n438 Vbias.n437 3.4105
R20195 Vbias.n428 Vbias.n427 3.4105
R20196 Vbias.n426 Vbias.n425 3.4105
R20197 Vbias.n422 Vbias.n421 3.4105
R20198 Vbias.n432 Vbias.n431 3.4105
R20199 Vbias.n434 Vbias.n433 3.4105
R20200 Vbias.n444 Vbias.n443 3.4105
R20201 Vbias.n446 Vbias.n445 3.4105
R20202 Vbias.n456 Vbias.n455 3.4105
R20203 Vbias.n458 Vbias.n457 3.4105
R20204 Vbias.n468 Vbias.n467 3.4105
R20205 Vbias.n470 Vbias.n469 3.4105
R20206 Vbias.n480 Vbias.n479 3.4105
R20207 Vbias.n482 Vbias.n481 3.4105
R20208 Vbias.n492 Vbias.n491 3.4105
R20209 Vbias.n494 Vbias.n493 3.4105
R20210 Vbias.n295 Vbias.n13 3.4105
R20211 Vbias.n294 Vbias.n293 3.4105
R20212 Vbias.n992 Vbias.n991 3.4105
R20213 Vbias.n990 Vbias.n989 3.4105
R20214 Vbias.n338 Vbias.n337 3.4105
R20215 Vbias.n341 Vbias.n340 3.4105
R20216 Vbias.n344 Vbias.n343 3.4105
R20217 Vbias.n347 Vbias.n346 3.4105
R20218 Vbias.n350 Vbias.n349 3.4105
R20219 Vbias.n353 Vbias.n352 3.4105
R20220 Vbias.n356 Vbias.n355 3.4105
R20221 Vbias.n359 Vbias.n358 3.4105
R20222 Vbias.n362 Vbias.n361 3.4105
R20223 Vbias.n365 Vbias.n364 3.4105
R20224 Vbias.n368 Vbias.n367 3.4105
R20225 Vbias.n371 Vbias.n370 3.4105
R20226 Vbias.n374 Vbias.n373 3.4105
R20227 Vbias.n416 Vbias.n415 3.4105
R20228 Vbias.n413 Vbias.n412 3.4105
R20229 Vbias.n410 Vbias.n409 3.4105
R20230 Vbias.n407 Vbias.n406 3.4105
R20231 Vbias.n404 Vbias.n403 3.4105
R20232 Vbias.n401 Vbias.n400 3.4105
R20233 Vbias.n398 Vbias.n397 3.4105
R20234 Vbias.n395 Vbias.n394 3.4105
R20235 Vbias.n392 Vbias.n391 3.4105
R20236 Vbias.n389 Vbias.n388 3.4105
R20237 Vbias.n386 Vbias.n385 3.4105
R20238 Vbias.n383 Vbias.n382 3.4105
R20239 Vbias.n380 Vbias.n379 3.4105
R20240 Vbias.n377 Vbias.n11 3.4105
R20241 Vbias.n995 Vbias.n994 3.4105
R20242 Vbias.n415 Vbias.n332 2.9408
R20243 Vbias.n911 Vbias.n910 2.9408
R20244 Vbias.n412 Vbias.n327 2.9408
R20245 Vbias.n915 Vbias.n914 2.9408
R20246 Vbias.n409 Vbias.n324 2.9408
R20247 Vbias.n921 Vbias.n920 2.9408
R20248 Vbias.n406 Vbias.n321 2.9408
R20249 Vbias.n925 Vbias.n924 2.9408
R20250 Vbias.n403 Vbias.n318 2.9408
R20251 Vbias.n931 Vbias.n930 2.9408
R20252 Vbias.n400 Vbias.n315 2.9408
R20253 Vbias.n935 Vbias.n934 2.9408
R20254 Vbias.n397 Vbias.n312 2.9408
R20255 Vbias.n941 Vbias.n940 2.9408
R20256 Vbias.n394 Vbias.n309 2.9408
R20257 Vbias.n945 Vbias.n944 2.9408
R20258 Vbias.n391 Vbias.n306 2.9408
R20259 Vbias.n951 Vbias.n950 2.9408
R20260 Vbias.n388 Vbias.n303 2.9408
R20261 Vbias.n955 Vbias.n954 2.9408
R20262 Vbias.n385 Vbias.n300 2.9408
R20263 Vbias.n961 Vbias.n960 2.9408
R20264 Vbias.n382 Vbias.n297 2.9408
R20265 Vbias.n965 Vbias.n964 2.9408
R20266 Vbias.n379 Vbias.n287 2.9408
R20267 Vbias.n971 Vbias.n970 2.9408
R20268 Vbias.n988 Vbias.n11 2.9408
R20269 Vbias.n975 Vbias.n974 2.9408
R20270 Vbias.n132 Vbias.n131 2.9408
R20271 Vbias.n906 Vbias.n905 2.9408
R20272 Vbias.n994 Vbias.n993 2.9408
R20273 Vbias.n418 Vbias.n417 2.9408
R20274 Vbias.n423 Vbias.n332 2.76612
R20275 Vbias.n424 Vbias.n423 2.76612
R20276 Vbias.n424 Vbias.n271 2.76612
R20277 Vbias.n552 Vbias.n271 2.76612
R20278 Vbias.n553 Vbias.n552 2.76612
R20279 Vbias.n553 Vbias.n187 2.76612
R20280 Vbias.n759 Vbias.n187 2.76612
R20281 Vbias.n759 Vbias.n758 2.76612
R20282 Vbias.n758 Vbias.n84 2.76612
R20283 Vbias.n897 Vbias.n84 2.76612
R20284 Vbias.n898 Vbias.n897 2.76612
R20285 Vbias.n898 Vbias.n76 2.76612
R20286 Vbias.n910 Vbias.n76 2.76612
R20287 Vbias.n430 Vbias.n327 2.76612
R20288 Vbias.n430 Vbias.n429 2.76612
R20289 Vbias.n429 Vbias.n268 2.76612
R20290 Vbias.n559 Vbias.n268 2.76612
R20291 Vbias.n559 Vbias.n558 2.76612
R20292 Vbias.n558 Vbias.n190 2.76612
R20293 Vbias.n752 Vbias.n190 2.76612
R20294 Vbias.n753 Vbias.n752 2.76612
R20295 Vbias.n753 Vbias.n87 2.76612
R20296 Vbias.n890 Vbias.n87 2.76612
R20297 Vbias.n890 Vbias.n889 2.76612
R20298 Vbias.n889 Vbias.n73 2.76612
R20299 Vbias.n915 Vbias.n73 2.76612
R20300 Vbias.n435 Vbias.n324 2.76612
R20301 Vbias.n436 Vbias.n435 2.76612
R20302 Vbias.n436 Vbias.n265 2.76612
R20303 Vbias.n564 Vbias.n265 2.76612
R20304 Vbias.n565 Vbias.n564 2.76612
R20305 Vbias.n565 Vbias.n193 2.76612
R20306 Vbias.n747 Vbias.n193 2.76612
R20307 Vbias.n747 Vbias.n746 2.76612
R20308 Vbias.n746 Vbias.n90 2.76612
R20309 Vbias.n883 Vbias.n90 2.76612
R20310 Vbias.n884 Vbias.n883 2.76612
R20311 Vbias.n884 Vbias.n70 2.76612
R20312 Vbias.n920 Vbias.n70 2.76612
R20313 Vbias.n442 Vbias.n321 2.76612
R20314 Vbias.n442 Vbias.n441 2.76612
R20315 Vbias.n441 Vbias.n262 2.76612
R20316 Vbias.n571 Vbias.n262 2.76612
R20317 Vbias.n571 Vbias.n570 2.76612
R20318 Vbias.n570 Vbias.n196 2.76612
R20319 Vbias.n740 Vbias.n196 2.76612
R20320 Vbias.n741 Vbias.n740 2.76612
R20321 Vbias.n741 Vbias.n93 2.76612
R20322 Vbias.n878 Vbias.n93 2.76612
R20323 Vbias.n878 Vbias.n877 2.76612
R20324 Vbias.n877 Vbias.n67 2.76612
R20325 Vbias.n925 Vbias.n67 2.76612
R20326 Vbias.n447 Vbias.n318 2.76612
R20327 Vbias.n448 Vbias.n447 2.76612
R20328 Vbias.n448 Vbias.n259 2.76612
R20329 Vbias.n576 Vbias.n259 2.76612
R20330 Vbias.n577 Vbias.n576 2.76612
R20331 Vbias.n577 Vbias.n199 2.76612
R20332 Vbias.n735 Vbias.n199 2.76612
R20333 Vbias.n735 Vbias.n734 2.76612
R20334 Vbias.n734 Vbias.n96 2.76612
R20335 Vbias.n871 Vbias.n96 2.76612
R20336 Vbias.n872 Vbias.n871 2.76612
R20337 Vbias.n872 Vbias.n64 2.76612
R20338 Vbias.n930 Vbias.n64 2.76612
R20339 Vbias.n454 Vbias.n315 2.76612
R20340 Vbias.n454 Vbias.n453 2.76612
R20341 Vbias.n453 Vbias.n256 2.76612
R20342 Vbias.n583 Vbias.n256 2.76612
R20343 Vbias.n583 Vbias.n582 2.76612
R20344 Vbias.n582 Vbias.n202 2.76612
R20345 Vbias.n728 Vbias.n202 2.76612
R20346 Vbias.n729 Vbias.n728 2.76612
R20347 Vbias.n729 Vbias.n99 2.76612
R20348 Vbias.n866 Vbias.n99 2.76612
R20349 Vbias.n866 Vbias.n865 2.76612
R20350 Vbias.n865 Vbias.n61 2.76612
R20351 Vbias.n935 Vbias.n61 2.76612
R20352 Vbias.n459 Vbias.n312 2.76612
R20353 Vbias.n460 Vbias.n459 2.76612
R20354 Vbias.n460 Vbias.n253 2.76612
R20355 Vbias.n588 Vbias.n253 2.76612
R20356 Vbias.n589 Vbias.n588 2.76612
R20357 Vbias.n589 Vbias.n205 2.76612
R20358 Vbias.n723 Vbias.n205 2.76612
R20359 Vbias.n723 Vbias.n722 2.76612
R20360 Vbias.n722 Vbias.n102 2.76612
R20361 Vbias.n859 Vbias.n102 2.76612
R20362 Vbias.n860 Vbias.n859 2.76612
R20363 Vbias.n860 Vbias.n58 2.76612
R20364 Vbias.n940 Vbias.n58 2.76612
R20365 Vbias.n466 Vbias.n309 2.76612
R20366 Vbias.n466 Vbias.n465 2.76612
R20367 Vbias.n465 Vbias.n250 2.76612
R20368 Vbias.n595 Vbias.n250 2.76612
R20369 Vbias.n595 Vbias.n594 2.76612
R20370 Vbias.n594 Vbias.n208 2.76612
R20371 Vbias.n716 Vbias.n208 2.76612
R20372 Vbias.n717 Vbias.n716 2.76612
R20373 Vbias.n717 Vbias.n105 2.76612
R20374 Vbias.n854 Vbias.n105 2.76612
R20375 Vbias.n854 Vbias.n853 2.76612
R20376 Vbias.n853 Vbias.n55 2.76612
R20377 Vbias.n945 Vbias.n55 2.76612
R20378 Vbias.n471 Vbias.n306 2.76612
R20379 Vbias.n472 Vbias.n471 2.76612
R20380 Vbias.n472 Vbias.n247 2.76612
R20381 Vbias.n600 Vbias.n247 2.76612
R20382 Vbias.n601 Vbias.n600 2.76612
R20383 Vbias.n601 Vbias.n211 2.76612
R20384 Vbias.n711 Vbias.n211 2.76612
R20385 Vbias.n711 Vbias.n710 2.76612
R20386 Vbias.n710 Vbias.n108 2.76612
R20387 Vbias.n847 Vbias.n108 2.76612
R20388 Vbias.n848 Vbias.n847 2.76612
R20389 Vbias.n848 Vbias.n52 2.76612
R20390 Vbias.n950 Vbias.n52 2.76612
R20391 Vbias.n478 Vbias.n303 2.76612
R20392 Vbias.n478 Vbias.n477 2.76612
R20393 Vbias.n477 Vbias.n244 2.76612
R20394 Vbias.n607 Vbias.n244 2.76612
R20395 Vbias.n607 Vbias.n606 2.76612
R20396 Vbias.n606 Vbias.n214 2.76612
R20397 Vbias.n704 Vbias.n214 2.76612
R20398 Vbias.n705 Vbias.n704 2.76612
R20399 Vbias.n705 Vbias.n111 2.76612
R20400 Vbias.n842 Vbias.n111 2.76612
R20401 Vbias.n842 Vbias.n841 2.76612
R20402 Vbias.n841 Vbias.n49 2.76612
R20403 Vbias.n955 Vbias.n49 2.76612
R20404 Vbias.n483 Vbias.n300 2.76612
R20405 Vbias.n484 Vbias.n483 2.76612
R20406 Vbias.n484 Vbias.n241 2.76612
R20407 Vbias.n612 Vbias.n241 2.76612
R20408 Vbias.n613 Vbias.n612 2.76612
R20409 Vbias.n613 Vbias.n217 2.76612
R20410 Vbias.n699 Vbias.n217 2.76612
R20411 Vbias.n699 Vbias.n698 2.76612
R20412 Vbias.n698 Vbias.n114 2.76612
R20413 Vbias.n835 Vbias.n114 2.76612
R20414 Vbias.n836 Vbias.n835 2.76612
R20415 Vbias.n836 Vbias.n46 2.76612
R20416 Vbias.n960 Vbias.n46 2.76612
R20417 Vbias.n490 Vbias.n297 2.76612
R20418 Vbias.n490 Vbias.n489 2.76612
R20419 Vbias.n489 Vbias.n238 2.76612
R20420 Vbias.n619 Vbias.n238 2.76612
R20421 Vbias.n619 Vbias.n618 2.76612
R20422 Vbias.n618 Vbias.n220 2.76612
R20423 Vbias.n692 Vbias.n220 2.76612
R20424 Vbias.n693 Vbias.n692 2.76612
R20425 Vbias.n693 Vbias.n117 2.76612
R20426 Vbias.n830 Vbias.n117 2.76612
R20427 Vbias.n830 Vbias.n829 2.76612
R20428 Vbias.n829 Vbias.n43 2.76612
R20429 Vbias.n965 Vbias.n43 2.76612
R20430 Vbias.n495 Vbias.n287 2.76612
R20431 Vbias.n496 Vbias.n495 2.76612
R20432 Vbias.n496 Vbias.n235 2.76612
R20433 Vbias.n624 Vbias.n235 2.76612
R20434 Vbias.n625 Vbias.n624 2.76612
R20435 Vbias.n625 Vbias.n223 2.76612
R20436 Vbias.n687 Vbias.n223 2.76612
R20437 Vbias.n687 Vbias.n686 2.76612
R20438 Vbias.n686 Vbias.n120 2.76612
R20439 Vbias.n823 Vbias.n120 2.76612
R20440 Vbias.n824 Vbias.n823 2.76612
R20441 Vbias.n824 Vbias.n40 2.76612
R20442 Vbias.n970 Vbias.n40 2.76612
R20443 Vbias.n988 Vbias.n987 2.76612
R20444 Vbias.n987 Vbias.n986 2.76612
R20445 Vbias.n986 Vbias.n985 2.76612
R20446 Vbias.n985 Vbias.n984 2.76612
R20447 Vbias.n984 Vbias.n983 2.76612
R20448 Vbias.n983 Vbias.n982 2.76612
R20449 Vbias.n982 Vbias.n981 2.76612
R20450 Vbias.n981 Vbias.n980 2.76612
R20451 Vbias.n980 Vbias.n979 2.76612
R20452 Vbias.n979 Vbias.n978 2.76612
R20453 Vbias.n978 Vbias.n977 2.76612
R20454 Vbias.n977 Vbias.n976 2.76612
R20455 Vbias.n976 Vbias.n975 2.76612
R20456 Vbias.n906 Vbias.n903 2.76612
R20457 Vbias.n816 Vbias.n124 2.76612
R20458 Vbias.n132 Vbias.n124 2.76612
R20459 Vbias.n902 Vbias.n81 2.76612
R20460 Vbias.n903 Vbias.n902 2.76612
R20461 Vbias.n817 Vbias.n123 2.76612
R20462 Vbias.n817 Vbias.n816 2.76612
R20463 Vbias.n765 Vbias.n764 2.76612
R20464 Vbias.n765 Vbias.n81 2.76612
R20465 Vbias.n680 Vbias.n679 2.76612
R20466 Vbias.n680 Vbias.n123 2.76612
R20467 Vbias.n763 Vbias.n184 2.76612
R20468 Vbias.n764 Vbias.n763 2.76612
R20469 Vbias.n678 Vbias.n228 2.76612
R20470 Vbias.n679 Vbias.n678 2.76612
R20471 Vbias.n548 Vbias.n276 2.76612
R20472 Vbias.n276 Vbias.n184 2.76612
R20473 Vbias.n503 Vbias.n284 2.76612
R20474 Vbias.n284 Vbias.n228 2.76612
R20475 Vbias.n547 Vbias.n277 2.76612
R20476 Vbias.n548 Vbias.n547 2.76612
R20477 Vbias.n502 Vbias.n7 2.76612
R20478 Vbias.n503 Vbias.n502 2.76612
R20479 Vbias.n419 Vbias.n418 2.76612
R20480 Vbias.n419 Vbias.n277 2.76612
R20481 Vbias.n993 Vbias.n7 2.76612
R20482 Vbias.n4 Vbias.n3 2.06591
R20483 Vbias Vbias.n997 1.58434
R20484 Vbias.n4 Vbias.n0 1.13456
R20485 Vbias Vbias.n4 0.782551
R20486 Vbias.n997 Vbias 0.617767
R20487 Vbias.n996 Vbias.n5 0.603667
R20488 Vbias.n291 Vbias.n5 0.603667
R20489 Vbias.n291 Vbias.n290 0.603667
R20490 Vbias.n290 Vbias.n289 0.603667
R20491 Vbias.n289 Vbias.n233 0.603667
R20492 Vbias.n632 Vbias.n233 0.603667
R20493 Vbias.n633 Vbias.n632 0.603667
R20494 Vbias.n633 Vbias.n232 0.603667
R20495 Vbias.n232 Vbias.n180 0.603667
R20496 Vbias.n810 Vbias.n180 0.603667
R20497 Vbias.n811 Vbias.n810 0.603667
R20498 Vbias.n812 Vbias.n811 0.603667
R20499 Vbias.n812 Vbias.n179 0.603667
R20500 Vbias.n179 Vbias.n135 0.603667
R20501 Vbias.n135 Vbias.n126 0.603667
R20502 Vbias.n126 Vbias 0.5692
R20503 Vbias.n997 Vbias.n996 0.492433
R20504 Vbias.n130 Vbias 0.252372
R20505 Vbias.n973 Vbias 0.252372
R20506 Vbias.n972 Vbias 0.252372
R20507 Vbias.n963 Vbias 0.252372
R20508 Vbias.n962 Vbias 0.252372
R20509 Vbias.n953 Vbias 0.252372
R20510 Vbias.n952 Vbias 0.252372
R20511 Vbias.n943 Vbias 0.252372
R20512 Vbias.n942 Vbias 0.252372
R20513 Vbias.n933 Vbias 0.252372
R20514 Vbias.n932 Vbias 0.252372
R20515 Vbias.n923 Vbias 0.252372
R20516 Vbias.n922 Vbias 0.252372
R20517 Vbias.n913 Vbias 0.252372
R20518 Vbias.n912 Vbias 0.252372
R20519 Vbias.n908 Vbias 0.252372
R20520 Vbias.n917 Vbias 0.252372
R20521 Vbias.n918 Vbias 0.252372
R20522 Vbias.n927 Vbias 0.252372
R20523 Vbias.n928 Vbias 0.252372
R20524 Vbias.n937 Vbias 0.252372
R20525 Vbias.n938 Vbias 0.252372
R20526 Vbias.n947 Vbias 0.252372
R20527 Vbias.n948 Vbias 0.252372
R20528 Vbias.n957 Vbias 0.252372
R20529 Vbias.n958 Vbias 0.252372
R20530 Vbias.n967 Vbias 0.252372
R20531 Vbias.n968 Vbias 0.252372
R20532 Vbias.n127 Vbias 0.252372
R20533 Vbias.n134 Vbias 0.252372
R20534 Vbias.n178 Vbias 0.252372
R20535 Vbias.n175 Vbias 0.252372
R20536 Vbias.n174 Vbias 0.252372
R20537 Vbias.n171 Vbias 0.252372
R20538 Vbias.n168 Vbias 0.252372
R20539 Vbias.n165 Vbias 0.252372
R20540 Vbias.n162 Vbias 0.252372
R20541 Vbias.n159 Vbias 0.252372
R20542 Vbias.n156 Vbias 0.252372
R20543 Vbias.n153 Vbias 0.252372
R20544 Vbias.n150 Vbias 0.252372
R20545 Vbias.n147 Vbias 0.252372
R20546 Vbias.n144 Vbias 0.252372
R20547 Vbias.n141 Vbias 0.252372
R20548 Vbias.n138 Vbias 0.252372
R20549 Vbias Vbias.n900 0.252372
R20550 Vbias.n887 Vbias 0.252372
R20551 Vbias Vbias.n886 0.252372
R20552 Vbias.n875 Vbias 0.252372
R20553 Vbias Vbias.n874 0.252372
R20554 Vbias.n863 Vbias 0.252372
R20555 Vbias Vbias.n862 0.252372
R20556 Vbias.n851 Vbias 0.252372
R20557 Vbias Vbias.n850 0.252372
R20558 Vbias.n839 Vbias 0.252372
R20559 Vbias Vbias.n838 0.252372
R20560 Vbias.n827 Vbias 0.252372
R20561 Vbias Vbias.n826 0.252372
R20562 Vbias.n813 Vbias 0.252372
R20563 Vbias.n814 Vbias 0.252372
R20564 Vbias Vbias.n819 0.252372
R20565 Vbias Vbias.n820 0.252372
R20566 Vbias.n821 Vbias 0.252372
R20567 Vbias Vbias.n832 0.252372
R20568 Vbias.n833 Vbias 0.252372
R20569 Vbias Vbias.n844 0.252372
R20570 Vbias.n845 Vbias 0.252372
R20571 Vbias Vbias.n856 0.252372
R20572 Vbias.n857 Vbias 0.252372
R20573 Vbias Vbias.n868 0.252372
R20574 Vbias.n869 Vbias 0.252372
R20575 Vbias Vbias.n880 0.252372
R20576 Vbias.n881 Vbias 0.252372
R20577 Vbias Vbias.n892 0.252372
R20578 Vbias.n895 Vbias 0.252372
R20579 Vbias.n769 Vbias 0.252372
R20580 Vbias.n772 Vbias 0.252372
R20581 Vbias.n775 Vbias 0.252372
R20582 Vbias.n778 Vbias 0.252372
R20583 Vbias.n781 Vbias 0.252372
R20584 Vbias.n784 Vbias 0.252372
R20585 Vbias.n787 Vbias 0.252372
R20586 Vbias.n790 Vbias 0.252372
R20587 Vbias.n793 Vbias 0.252372
R20588 Vbias.n796 Vbias 0.252372
R20589 Vbias.n799 Vbias 0.252372
R20590 Vbias.n802 Vbias 0.252372
R20591 Vbias.n805 Vbias 0.252372
R20592 Vbias.n806 Vbias 0.252372
R20593 Vbias.n809 Vbias 0.252372
R20594 Vbias Vbias.n682 0.252372
R20595 Vbias Vbias.n683 0.252372
R20596 Vbias.n684 Vbias 0.252372
R20597 Vbias Vbias.n695 0.252372
R20598 Vbias.n696 Vbias 0.252372
R20599 Vbias Vbias.n707 0.252372
R20600 Vbias.n708 Vbias 0.252372
R20601 Vbias Vbias.n719 0.252372
R20602 Vbias.n720 Vbias 0.252372
R20603 Vbias Vbias.n731 0.252372
R20604 Vbias.n732 Vbias 0.252372
R20605 Vbias Vbias.n743 0.252372
R20606 Vbias.n744 Vbias 0.252372
R20607 Vbias Vbias.n755 0.252372
R20608 Vbias.n756 Vbias 0.252372
R20609 Vbias Vbias.n761 0.252372
R20610 Vbias.n750 Vbias 0.252372
R20611 Vbias Vbias.n749 0.252372
R20612 Vbias.n738 Vbias 0.252372
R20613 Vbias Vbias.n737 0.252372
R20614 Vbias.n726 Vbias 0.252372
R20615 Vbias Vbias.n725 0.252372
R20616 Vbias.n714 Vbias 0.252372
R20617 Vbias Vbias.n713 0.252372
R20618 Vbias.n702 Vbias 0.252372
R20619 Vbias Vbias.n701 0.252372
R20620 Vbias.n690 Vbias 0.252372
R20621 Vbias Vbias.n689 0.252372
R20622 Vbias.n230 Vbias 0.252372
R20623 Vbias.n231 Vbias 0.252372
R20624 Vbias.n676 Vbias 0.252372
R20625 Vbias.n675 Vbias 0.252372
R20626 Vbias.n674 Vbias 0.252372
R20627 Vbias.n671 Vbias 0.252372
R20628 Vbias.n668 Vbias 0.252372
R20629 Vbias.n665 Vbias 0.252372
R20630 Vbias.n662 Vbias 0.252372
R20631 Vbias.n659 Vbias 0.252372
R20632 Vbias.n656 Vbias 0.252372
R20633 Vbias.n653 Vbias 0.252372
R20634 Vbias.n650 Vbias 0.252372
R20635 Vbias.n647 Vbias 0.252372
R20636 Vbias.n644 Vbias 0.252372
R20637 Vbias.n641 Vbias 0.252372
R20638 Vbias.n638 Vbias 0.252372
R20639 Vbias.n555 Vbias 0.252372
R20640 Vbias.n556 Vbias 0.252372
R20641 Vbias.n567 Vbias 0.252372
R20642 Vbias.n568 Vbias 0.252372
R20643 Vbias.n579 Vbias 0.252372
R20644 Vbias.n580 Vbias 0.252372
R20645 Vbias.n591 Vbias 0.252372
R20646 Vbias.n592 Vbias 0.252372
R20647 Vbias.n603 Vbias 0.252372
R20648 Vbias.n604 Vbias 0.252372
R20649 Vbias.n615 Vbias 0.252372
R20650 Vbias.n616 Vbias 0.252372
R20651 Vbias.n627 Vbias 0.252372
R20652 Vbias.n628 Vbias 0.252372
R20653 Vbias.n631 Vbias 0.252372
R20654 Vbias.n282 Vbias 0.252372
R20655 Vbias.n281 Vbias 0.252372
R20656 Vbias.n622 Vbias 0.252372
R20657 Vbias.n621 Vbias 0.252372
R20658 Vbias.n610 Vbias 0.252372
R20659 Vbias.n609 Vbias 0.252372
R20660 Vbias.n598 Vbias 0.252372
R20661 Vbias.n597 Vbias 0.252372
R20662 Vbias.n586 Vbias 0.252372
R20663 Vbias.n585 Vbias 0.252372
R20664 Vbias.n574 Vbias 0.252372
R20665 Vbias.n573 Vbias 0.252372
R20666 Vbias.n562 Vbias 0.252372
R20667 Vbias.n561 Vbias 0.252372
R20668 Vbias.n550 Vbias 0.252372
R20669 Vbias Vbias.n545 0.252372
R20670 Vbias Vbias.n542 0.252372
R20671 Vbias Vbias.n539 0.252372
R20672 Vbias Vbias.n536 0.252372
R20673 Vbias Vbias.n533 0.252372
R20674 Vbias Vbias.n530 0.252372
R20675 Vbias Vbias.n527 0.252372
R20676 Vbias Vbias.n524 0.252372
R20677 Vbias Vbias.n521 0.252372
R20678 Vbias Vbias.n518 0.252372
R20679 Vbias Vbias.n515 0.252372
R20680 Vbias Vbias.n512 0.252372
R20681 Vbias Vbias.n509 0.252372
R20682 Vbias Vbias.n506 0.252372
R20683 Vbias Vbias.n505 0.252372
R20684 Vbias.n500 Vbias 0.252372
R20685 Vbias.n499 Vbias 0.252372
R20686 Vbias.n498 Vbias 0.252372
R20687 Vbias.n487 Vbias 0.252372
R20688 Vbias.n486 Vbias 0.252372
R20689 Vbias.n475 Vbias 0.252372
R20690 Vbias.n474 Vbias 0.252372
R20691 Vbias.n463 Vbias 0.252372
R20692 Vbias.n462 Vbias 0.252372
R20693 Vbias.n451 Vbias 0.252372
R20694 Vbias.n450 Vbias 0.252372
R20695 Vbias.n439 Vbias 0.252372
R20696 Vbias.n438 Vbias 0.252372
R20697 Vbias.n427 Vbias 0.252372
R20698 Vbias.n426 Vbias 0.252372
R20699 Vbias.n421 Vbias 0.252372
R20700 Vbias.n432 Vbias 0.252372
R20701 Vbias.n433 Vbias 0.252372
R20702 Vbias.n444 Vbias 0.252372
R20703 Vbias.n445 Vbias 0.252372
R20704 Vbias.n456 Vbias 0.252372
R20705 Vbias.n457 Vbias 0.252372
R20706 Vbias.n468 Vbias 0.252372
R20707 Vbias.n469 Vbias 0.252372
R20708 Vbias.n480 Vbias 0.252372
R20709 Vbias.n481 Vbias 0.252372
R20710 Vbias.n492 Vbias 0.252372
R20711 Vbias.n493 Vbias 0.252372
R20712 Vbias Vbias.n295 0.252372
R20713 Vbias Vbias.n294 0.252372
R20714 Vbias.n991 Vbias 0.252372
R20715 Vbias.n990 Vbias 0.252372
R20716 Vbias Vbias.n338 0.252372
R20717 Vbias Vbias.n341 0.252372
R20718 Vbias Vbias.n344 0.252372
R20719 Vbias Vbias.n347 0.252372
R20720 Vbias Vbias.n350 0.252372
R20721 Vbias Vbias.n353 0.252372
R20722 Vbias Vbias.n356 0.252372
R20723 Vbias Vbias.n359 0.252372
R20724 Vbias Vbias.n362 0.252372
R20725 Vbias Vbias.n365 0.252372
R20726 Vbias Vbias.n368 0.252372
R20727 Vbias Vbias.n371 0.252372
R20728 Vbias Vbias.n374 0.252372
R20729 Vbias Vbias.n416 0.252372
R20730 Vbias Vbias.n413 0.252372
R20731 Vbias Vbias.n410 0.252372
R20732 Vbias Vbias.n407 0.252372
R20733 Vbias Vbias.n404 0.252372
R20734 Vbias Vbias.n401 0.252372
R20735 Vbias Vbias.n398 0.252372
R20736 Vbias Vbias.n395 0.252372
R20737 Vbias Vbias.n392 0.252372
R20738 Vbias Vbias.n389 0.252372
R20739 Vbias Vbias.n386 0.252372
R20740 Vbias Vbias.n383 0.252372
R20741 Vbias Vbias.n380 0.252372
R20742 Vbias Vbias.n377 0.252372
R20743 Vbias.n995 Vbias 0.252372
R20744 Vbias.n373 Vbias.n332 0.175179
R20745 Vbias.n423 Vbias.n422 0.175179
R20746 Vbias.n425 Vbias.n424 0.175179
R20747 Vbias.n544 Vbias.n271 0.175179
R20748 Vbias.n552 Vbias.n551 0.175179
R20749 Vbias.n554 Vbias.n553 0.175179
R20750 Vbias.n637 Vbias.n187 0.175179
R20751 Vbias.n760 Vbias.n759 0.175179
R20752 Vbias.n758 Vbias.n757 0.175179
R20753 Vbias.n768 Vbias.n84 0.175179
R20754 Vbias.n897 Vbias.n896 0.175179
R20755 Vbias.n899 Vbias.n898 0.175179
R20756 Vbias.n137 Vbias.n76 0.175179
R20757 Vbias.n910 Vbias.n909 0.175179
R20758 Vbias.n370 Vbias.n327 0.175179
R20759 Vbias.n431 Vbias.n430 0.175179
R20760 Vbias.n429 Vbias.n428 0.175179
R20761 Vbias.n541 Vbias.n268 0.175179
R20762 Vbias.n560 Vbias.n559 0.175179
R20763 Vbias.n558 Vbias.n557 0.175179
R20764 Vbias.n640 Vbias.n190 0.175179
R20765 Vbias.n752 Vbias.n751 0.175179
R20766 Vbias.n754 Vbias.n753 0.175179
R20767 Vbias.n771 Vbias.n87 0.175179
R20768 Vbias.n891 Vbias.n890 0.175179
R20769 Vbias.n889 Vbias.n888 0.175179
R20770 Vbias.n140 Vbias.n73 0.175179
R20771 Vbias.n916 Vbias.n915 0.175179
R20772 Vbias.n367 Vbias.n324 0.175179
R20773 Vbias.n435 Vbias.n434 0.175179
R20774 Vbias.n437 Vbias.n436 0.175179
R20775 Vbias.n538 Vbias.n265 0.175179
R20776 Vbias.n564 Vbias.n563 0.175179
R20777 Vbias.n566 Vbias.n565 0.175179
R20778 Vbias.n643 Vbias.n193 0.175179
R20779 Vbias.n748 Vbias.n747 0.175179
R20780 Vbias.n746 Vbias.n745 0.175179
R20781 Vbias.n774 Vbias.n90 0.175179
R20782 Vbias.n883 Vbias.n882 0.175179
R20783 Vbias.n885 Vbias.n884 0.175179
R20784 Vbias.n143 Vbias.n70 0.175179
R20785 Vbias.n920 Vbias.n919 0.175179
R20786 Vbias.n364 Vbias.n321 0.175179
R20787 Vbias.n443 Vbias.n442 0.175179
R20788 Vbias.n441 Vbias.n440 0.175179
R20789 Vbias.n535 Vbias.n262 0.175179
R20790 Vbias.n572 Vbias.n571 0.175179
R20791 Vbias.n570 Vbias.n569 0.175179
R20792 Vbias.n646 Vbias.n196 0.175179
R20793 Vbias.n740 Vbias.n739 0.175179
R20794 Vbias.n742 Vbias.n741 0.175179
R20795 Vbias.n777 Vbias.n93 0.175179
R20796 Vbias.n879 Vbias.n878 0.175179
R20797 Vbias.n877 Vbias.n876 0.175179
R20798 Vbias.n146 Vbias.n67 0.175179
R20799 Vbias.n926 Vbias.n925 0.175179
R20800 Vbias.n361 Vbias.n318 0.175179
R20801 Vbias.n447 Vbias.n446 0.175179
R20802 Vbias.n449 Vbias.n448 0.175179
R20803 Vbias.n532 Vbias.n259 0.175179
R20804 Vbias.n576 Vbias.n575 0.175179
R20805 Vbias.n578 Vbias.n577 0.175179
R20806 Vbias.n649 Vbias.n199 0.175179
R20807 Vbias.n736 Vbias.n735 0.175179
R20808 Vbias.n734 Vbias.n733 0.175179
R20809 Vbias.n780 Vbias.n96 0.175179
R20810 Vbias.n871 Vbias.n870 0.175179
R20811 Vbias.n873 Vbias.n872 0.175179
R20812 Vbias.n149 Vbias.n64 0.175179
R20813 Vbias.n930 Vbias.n929 0.175179
R20814 Vbias.n358 Vbias.n315 0.175179
R20815 Vbias.n455 Vbias.n454 0.175179
R20816 Vbias.n453 Vbias.n452 0.175179
R20817 Vbias.n529 Vbias.n256 0.175179
R20818 Vbias.n584 Vbias.n583 0.175179
R20819 Vbias.n582 Vbias.n581 0.175179
R20820 Vbias.n652 Vbias.n202 0.175179
R20821 Vbias.n728 Vbias.n727 0.175179
R20822 Vbias.n730 Vbias.n729 0.175179
R20823 Vbias.n783 Vbias.n99 0.175179
R20824 Vbias.n867 Vbias.n866 0.175179
R20825 Vbias.n865 Vbias.n864 0.175179
R20826 Vbias.n152 Vbias.n61 0.175179
R20827 Vbias.n936 Vbias.n935 0.175179
R20828 Vbias.n355 Vbias.n312 0.175179
R20829 Vbias.n459 Vbias.n458 0.175179
R20830 Vbias.n461 Vbias.n460 0.175179
R20831 Vbias.n526 Vbias.n253 0.175179
R20832 Vbias.n588 Vbias.n587 0.175179
R20833 Vbias.n590 Vbias.n589 0.175179
R20834 Vbias.n655 Vbias.n205 0.175179
R20835 Vbias.n724 Vbias.n723 0.175179
R20836 Vbias.n722 Vbias.n721 0.175179
R20837 Vbias.n786 Vbias.n102 0.175179
R20838 Vbias.n859 Vbias.n858 0.175179
R20839 Vbias.n861 Vbias.n860 0.175179
R20840 Vbias.n155 Vbias.n58 0.175179
R20841 Vbias.n940 Vbias.n939 0.175179
R20842 Vbias.n352 Vbias.n309 0.175179
R20843 Vbias.n467 Vbias.n466 0.175179
R20844 Vbias.n465 Vbias.n464 0.175179
R20845 Vbias.n523 Vbias.n250 0.175179
R20846 Vbias.n596 Vbias.n595 0.175179
R20847 Vbias.n594 Vbias.n593 0.175179
R20848 Vbias.n658 Vbias.n208 0.175179
R20849 Vbias.n716 Vbias.n715 0.175179
R20850 Vbias.n718 Vbias.n717 0.175179
R20851 Vbias.n789 Vbias.n105 0.175179
R20852 Vbias.n855 Vbias.n854 0.175179
R20853 Vbias.n853 Vbias.n852 0.175179
R20854 Vbias.n158 Vbias.n55 0.175179
R20855 Vbias.n946 Vbias.n945 0.175179
R20856 Vbias.n349 Vbias.n306 0.175179
R20857 Vbias.n471 Vbias.n470 0.175179
R20858 Vbias.n473 Vbias.n472 0.175179
R20859 Vbias.n520 Vbias.n247 0.175179
R20860 Vbias.n600 Vbias.n599 0.175179
R20861 Vbias.n602 Vbias.n601 0.175179
R20862 Vbias.n661 Vbias.n211 0.175179
R20863 Vbias.n712 Vbias.n711 0.175179
R20864 Vbias.n710 Vbias.n709 0.175179
R20865 Vbias.n792 Vbias.n108 0.175179
R20866 Vbias.n847 Vbias.n846 0.175179
R20867 Vbias.n849 Vbias.n848 0.175179
R20868 Vbias.n161 Vbias.n52 0.175179
R20869 Vbias.n950 Vbias.n949 0.175179
R20870 Vbias.n346 Vbias.n303 0.175179
R20871 Vbias.n479 Vbias.n478 0.175179
R20872 Vbias.n477 Vbias.n476 0.175179
R20873 Vbias.n517 Vbias.n244 0.175179
R20874 Vbias.n608 Vbias.n607 0.175179
R20875 Vbias.n606 Vbias.n605 0.175179
R20876 Vbias.n664 Vbias.n214 0.175179
R20877 Vbias.n704 Vbias.n703 0.175179
R20878 Vbias.n706 Vbias.n705 0.175179
R20879 Vbias.n795 Vbias.n111 0.175179
R20880 Vbias.n843 Vbias.n842 0.175179
R20881 Vbias.n841 Vbias.n840 0.175179
R20882 Vbias.n164 Vbias.n49 0.175179
R20883 Vbias.n956 Vbias.n955 0.175179
R20884 Vbias.n343 Vbias.n300 0.175179
R20885 Vbias.n483 Vbias.n482 0.175179
R20886 Vbias.n485 Vbias.n484 0.175179
R20887 Vbias.n514 Vbias.n241 0.175179
R20888 Vbias.n612 Vbias.n611 0.175179
R20889 Vbias.n614 Vbias.n613 0.175179
R20890 Vbias.n667 Vbias.n217 0.175179
R20891 Vbias.n700 Vbias.n699 0.175179
R20892 Vbias.n698 Vbias.n697 0.175179
R20893 Vbias.n798 Vbias.n114 0.175179
R20894 Vbias.n835 Vbias.n834 0.175179
R20895 Vbias.n837 Vbias.n836 0.175179
R20896 Vbias.n167 Vbias.n46 0.175179
R20897 Vbias.n960 Vbias.n959 0.175179
R20898 Vbias.n340 Vbias.n297 0.175179
R20899 Vbias.n491 Vbias.n490 0.175179
R20900 Vbias.n489 Vbias.n488 0.175179
R20901 Vbias.n511 Vbias.n238 0.175179
R20902 Vbias.n620 Vbias.n619 0.175179
R20903 Vbias.n618 Vbias.n617 0.175179
R20904 Vbias.n670 Vbias.n220 0.175179
R20905 Vbias.n692 Vbias.n691 0.175179
R20906 Vbias.n694 Vbias.n693 0.175179
R20907 Vbias.n801 Vbias.n117 0.175179
R20908 Vbias.n831 Vbias.n830 0.175179
R20909 Vbias.n829 Vbias.n828 0.175179
R20910 Vbias.n170 Vbias.n43 0.175179
R20911 Vbias.n966 Vbias.n965 0.175179
R20912 Vbias.n337 Vbias.n287 0.175179
R20913 Vbias.n495 Vbias.n494 0.175179
R20914 Vbias.n497 Vbias.n496 0.175179
R20915 Vbias.n508 Vbias.n235 0.175179
R20916 Vbias.n624 Vbias.n623 0.175179
R20917 Vbias.n626 Vbias.n625 0.175179
R20918 Vbias.n673 Vbias.n223 0.175179
R20919 Vbias.n688 Vbias.n687 0.175179
R20920 Vbias.n686 Vbias.n685 0.175179
R20921 Vbias.n804 Vbias.n120 0.175179
R20922 Vbias.n823 Vbias.n822 0.175179
R20923 Vbias.n825 Vbias.n824 0.175179
R20924 Vbias.n173 Vbias.n40 0.175179
R20925 Vbias.n970 Vbias.n969 0.175179
R20926 Vbias.n989 Vbias.n988 0.175179
R20927 Vbias.n987 Vbias.n13 0.175179
R20928 Vbias.n986 Vbias.n15 0.175179
R20929 Vbias.n985 Vbias.n17 0.175179
R20930 Vbias.n984 Vbias.n19 0.175179
R20931 Vbias.n983 Vbias.n21 0.175179
R20932 Vbias.n982 Vbias.n23 0.175179
R20933 Vbias.n981 Vbias.n25 0.175179
R20934 Vbias.n980 Vbias.n27 0.175179
R20935 Vbias.n979 Vbias.n29 0.175179
R20936 Vbias.n978 Vbias.n31 0.175179
R20937 Vbias.n977 Vbias.n33 0.175179
R20938 Vbias.n976 Vbias.n35 0.175179
R20939 Vbias.n975 Vbias.n37 0.175179
R20940 Vbias.n907 Vbias.n906 0.175179
R20941 Vbias.n133 Vbias.n132 0.175179
R20942 Vbias.n177 Vbias.n124 0.175179
R20943 Vbias.n903 Vbias.n80 0.175179
R20944 Vbias.n902 Vbias.n901 0.175179
R20945 Vbias.n816 Vbias.n815 0.175179
R20946 Vbias.n818 Vbias.n817 0.175179
R20947 Vbias.n894 Vbias.n81 0.175179
R20948 Vbias.n766 Vbias.n765 0.175179
R20949 Vbias.n808 Vbias.n123 0.175179
R20950 Vbias.n681 Vbias.n680 0.175179
R20951 Vbias.n764 Vbias.n183 0.175179
R20952 Vbias.n763 Vbias.n762 0.175179
R20953 Vbias.n679 Vbias.n227 0.175179
R20954 Vbias.n678 Vbias.n677 0.175179
R20955 Vbias.n635 Vbias.n184 0.175179
R20956 Vbias.n276 Vbias.n275 0.175179
R20957 Vbias.n630 Vbias.n228 0.175179
R20958 Vbias.n284 Vbias.n283 0.175179
R20959 Vbias.n549 Vbias.n548 0.175179
R20960 Vbias.n547 Vbias.n546 0.175179
R20961 Vbias.n504 Vbias.n503 0.175179
R20962 Vbias.n502 Vbias.n501 0.175179
R20963 Vbias.n330 Vbias.n277 0.175179
R20964 Vbias.n420 Vbias.n419 0.175179
R20965 Vbias.n293 Vbias.n7 0.175179
R20966 Vbias.n993 Vbias.n992 0.175179
R20967 Vbias.n418 Vbias.n375 0.175179
R20968 Vbias.n294 Vbias 0.0972718
R20969 Vbias.n505 Vbias 0.0972718
R20970 Vbias Vbias.n631 0.0972718
R20971 Vbias Vbias.n231 0.0972718
R20972 Vbias Vbias.n809 0.0972718
R20973 Vbias.n814 Vbias 0.0972718
R20974 Vbias Vbias.n134 0.0972718
R20975 Vbias.n130 Vbias 0.0972718
R20976 Vbias.n973 Vbias 0.0972718
R20977 Vbias Vbias.n972 0.0972718
R20978 Vbias.n963 Vbias 0.0972718
R20979 Vbias Vbias.n962 0.0972718
R20980 Vbias.n953 Vbias 0.0972718
R20981 Vbias Vbias.n952 0.0972718
R20982 Vbias.n943 Vbias 0.0972718
R20983 Vbias Vbias.n942 0.0972718
R20984 Vbias.n933 Vbias 0.0972718
R20985 Vbias Vbias.n932 0.0972718
R20986 Vbias.n923 Vbias 0.0972718
R20987 Vbias Vbias.n922 0.0972718
R20988 Vbias.n913 Vbias 0.0972718
R20989 Vbias Vbias.n912 0.0972718
R20990 Vbias.n908 Vbias 0.0972718
R20991 Vbias Vbias.n917 0.0972718
R20992 Vbias.n918 Vbias 0.0972718
R20993 Vbias Vbias.n927 0.0972718
R20994 Vbias.n928 Vbias 0.0972718
R20995 Vbias Vbias.n937 0.0972718
R20996 Vbias.n938 Vbias 0.0972718
R20997 Vbias Vbias.n947 0.0972718
R20998 Vbias.n948 Vbias 0.0972718
R20999 Vbias Vbias.n957 0.0972718
R21000 Vbias.n958 Vbias 0.0972718
R21001 Vbias Vbias.n967 0.0972718
R21002 Vbias.n968 Vbias 0.0972718
R21003 Vbias Vbias.n127 0.0972718
R21004 Vbias Vbias.n178 0.0972718
R21005 Vbias Vbias.n175 0.0972718
R21006 Vbias Vbias.n174 0.0972718
R21007 Vbias Vbias.n171 0.0972718
R21008 Vbias Vbias.n168 0.0972718
R21009 Vbias Vbias.n165 0.0972718
R21010 Vbias Vbias.n162 0.0972718
R21011 Vbias Vbias.n159 0.0972718
R21012 Vbias Vbias.n156 0.0972718
R21013 Vbias Vbias.n153 0.0972718
R21014 Vbias Vbias.n150 0.0972718
R21015 Vbias Vbias.n147 0.0972718
R21016 Vbias Vbias.n144 0.0972718
R21017 Vbias Vbias.n141 0.0972718
R21018 Vbias Vbias.n138 0.0972718
R21019 Vbias.n900 Vbias 0.0972718
R21020 Vbias.n887 Vbias 0.0972718
R21021 Vbias.n886 Vbias 0.0972718
R21022 Vbias.n875 Vbias 0.0972718
R21023 Vbias.n874 Vbias 0.0972718
R21024 Vbias.n863 Vbias 0.0972718
R21025 Vbias.n862 Vbias 0.0972718
R21026 Vbias.n851 Vbias 0.0972718
R21027 Vbias.n850 Vbias 0.0972718
R21028 Vbias.n839 Vbias 0.0972718
R21029 Vbias.n838 Vbias 0.0972718
R21030 Vbias.n827 Vbias 0.0972718
R21031 Vbias.n826 Vbias 0.0972718
R21032 Vbias Vbias.n813 0.0972718
R21033 Vbias.n819 Vbias 0.0972718
R21034 Vbias.n820 Vbias 0.0972718
R21035 Vbias.n821 Vbias 0.0972718
R21036 Vbias.n832 Vbias 0.0972718
R21037 Vbias.n833 Vbias 0.0972718
R21038 Vbias.n844 Vbias 0.0972718
R21039 Vbias.n845 Vbias 0.0972718
R21040 Vbias.n856 Vbias 0.0972718
R21041 Vbias.n857 Vbias 0.0972718
R21042 Vbias.n868 Vbias 0.0972718
R21043 Vbias.n869 Vbias 0.0972718
R21044 Vbias.n880 Vbias 0.0972718
R21045 Vbias.n881 Vbias 0.0972718
R21046 Vbias.n892 Vbias 0.0972718
R21047 Vbias.n895 Vbias 0.0972718
R21048 Vbias Vbias.n769 0.0972718
R21049 Vbias Vbias.n772 0.0972718
R21050 Vbias Vbias.n775 0.0972718
R21051 Vbias Vbias.n778 0.0972718
R21052 Vbias Vbias.n781 0.0972718
R21053 Vbias Vbias.n784 0.0972718
R21054 Vbias Vbias.n787 0.0972718
R21055 Vbias Vbias.n790 0.0972718
R21056 Vbias Vbias.n793 0.0972718
R21057 Vbias Vbias.n796 0.0972718
R21058 Vbias Vbias.n799 0.0972718
R21059 Vbias Vbias.n802 0.0972718
R21060 Vbias Vbias.n805 0.0972718
R21061 Vbias Vbias.n806 0.0972718
R21062 Vbias.n682 Vbias 0.0972718
R21063 Vbias.n683 Vbias 0.0972718
R21064 Vbias.n684 Vbias 0.0972718
R21065 Vbias.n695 Vbias 0.0972718
R21066 Vbias.n696 Vbias 0.0972718
R21067 Vbias.n707 Vbias 0.0972718
R21068 Vbias.n708 Vbias 0.0972718
R21069 Vbias.n719 Vbias 0.0972718
R21070 Vbias.n720 Vbias 0.0972718
R21071 Vbias.n731 Vbias 0.0972718
R21072 Vbias.n732 Vbias 0.0972718
R21073 Vbias.n743 Vbias 0.0972718
R21074 Vbias.n744 Vbias 0.0972718
R21075 Vbias.n755 Vbias 0.0972718
R21076 Vbias.n756 Vbias 0.0972718
R21077 Vbias.n761 Vbias 0.0972718
R21078 Vbias.n750 Vbias 0.0972718
R21079 Vbias.n749 Vbias 0.0972718
R21080 Vbias.n738 Vbias 0.0972718
R21081 Vbias.n737 Vbias 0.0972718
R21082 Vbias.n726 Vbias 0.0972718
R21083 Vbias.n725 Vbias 0.0972718
R21084 Vbias.n714 Vbias 0.0972718
R21085 Vbias.n713 Vbias 0.0972718
R21086 Vbias.n702 Vbias 0.0972718
R21087 Vbias.n701 Vbias 0.0972718
R21088 Vbias.n690 Vbias 0.0972718
R21089 Vbias.n689 Vbias 0.0972718
R21090 Vbias Vbias.n230 0.0972718
R21091 Vbias.n676 Vbias 0.0972718
R21092 Vbias Vbias.n675 0.0972718
R21093 Vbias Vbias.n674 0.0972718
R21094 Vbias Vbias.n671 0.0972718
R21095 Vbias Vbias.n668 0.0972718
R21096 Vbias Vbias.n665 0.0972718
R21097 Vbias Vbias.n662 0.0972718
R21098 Vbias Vbias.n659 0.0972718
R21099 Vbias Vbias.n656 0.0972718
R21100 Vbias Vbias.n653 0.0972718
R21101 Vbias Vbias.n650 0.0972718
R21102 Vbias Vbias.n647 0.0972718
R21103 Vbias Vbias.n644 0.0972718
R21104 Vbias Vbias.n641 0.0972718
R21105 Vbias Vbias.n638 0.0972718
R21106 Vbias Vbias.n555 0.0972718
R21107 Vbias.n556 Vbias 0.0972718
R21108 Vbias Vbias.n567 0.0972718
R21109 Vbias.n568 Vbias 0.0972718
R21110 Vbias Vbias.n579 0.0972718
R21111 Vbias.n580 Vbias 0.0972718
R21112 Vbias Vbias.n591 0.0972718
R21113 Vbias.n592 Vbias 0.0972718
R21114 Vbias Vbias.n603 0.0972718
R21115 Vbias.n604 Vbias 0.0972718
R21116 Vbias Vbias.n615 0.0972718
R21117 Vbias.n616 Vbias 0.0972718
R21118 Vbias Vbias.n627 0.0972718
R21119 Vbias Vbias.n628 0.0972718
R21120 Vbias.n282 Vbias 0.0972718
R21121 Vbias Vbias.n281 0.0972718
R21122 Vbias.n622 Vbias 0.0972718
R21123 Vbias Vbias.n621 0.0972718
R21124 Vbias.n610 Vbias 0.0972718
R21125 Vbias Vbias.n609 0.0972718
R21126 Vbias.n598 Vbias 0.0972718
R21127 Vbias Vbias.n597 0.0972718
R21128 Vbias.n586 Vbias 0.0972718
R21129 Vbias Vbias.n585 0.0972718
R21130 Vbias.n574 Vbias 0.0972718
R21131 Vbias Vbias.n573 0.0972718
R21132 Vbias.n562 Vbias 0.0972718
R21133 Vbias Vbias.n561 0.0972718
R21134 Vbias.n550 Vbias 0.0972718
R21135 Vbias.n545 Vbias 0.0972718
R21136 Vbias.n542 Vbias 0.0972718
R21137 Vbias.n539 Vbias 0.0972718
R21138 Vbias.n536 Vbias 0.0972718
R21139 Vbias.n533 Vbias 0.0972718
R21140 Vbias.n530 Vbias 0.0972718
R21141 Vbias.n527 Vbias 0.0972718
R21142 Vbias.n524 Vbias 0.0972718
R21143 Vbias.n521 Vbias 0.0972718
R21144 Vbias.n518 Vbias 0.0972718
R21145 Vbias.n515 Vbias 0.0972718
R21146 Vbias.n512 Vbias 0.0972718
R21147 Vbias.n509 Vbias 0.0972718
R21148 Vbias.n506 Vbias 0.0972718
R21149 Vbias.n500 Vbias 0.0972718
R21150 Vbias Vbias.n499 0.0972718
R21151 Vbias Vbias.n498 0.0972718
R21152 Vbias.n487 Vbias 0.0972718
R21153 Vbias Vbias.n486 0.0972718
R21154 Vbias.n475 Vbias 0.0972718
R21155 Vbias Vbias.n474 0.0972718
R21156 Vbias.n463 Vbias 0.0972718
R21157 Vbias Vbias.n462 0.0972718
R21158 Vbias.n451 Vbias 0.0972718
R21159 Vbias Vbias.n450 0.0972718
R21160 Vbias.n439 Vbias 0.0972718
R21161 Vbias Vbias.n438 0.0972718
R21162 Vbias.n427 Vbias 0.0972718
R21163 Vbias Vbias.n426 0.0972718
R21164 Vbias.n421 Vbias 0.0972718
R21165 Vbias Vbias.n432 0.0972718
R21166 Vbias.n433 Vbias 0.0972718
R21167 Vbias Vbias.n444 0.0972718
R21168 Vbias.n445 Vbias 0.0972718
R21169 Vbias Vbias.n456 0.0972718
R21170 Vbias.n457 Vbias 0.0972718
R21171 Vbias Vbias.n468 0.0972718
R21172 Vbias.n469 Vbias 0.0972718
R21173 Vbias Vbias.n480 0.0972718
R21174 Vbias.n481 Vbias 0.0972718
R21175 Vbias Vbias.n492 0.0972718
R21176 Vbias.n493 Vbias 0.0972718
R21177 Vbias.n295 Vbias 0.0972718
R21178 Vbias.n991 Vbias 0.0972718
R21179 Vbias Vbias.n990 0.0972718
R21180 Vbias.n338 Vbias 0.0972718
R21181 Vbias.n341 Vbias 0.0972718
R21182 Vbias.n344 Vbias 0.0972718
R21183 Vbias.n347 Vbias 0.0972718
R21184 Vbias.n350 Vbias 0.0972718
R21185 Vbias.n353 Vbias 0.0972718
R21186 Vbias.n356 Vbias 0.0972718
R21187 Vbias.n359 Vbias 0.0972718
R21188 Vbias.n362 Vbias 0.0972718
R21189 Vbias.n365 Vbias 0.0972718
R21190 Vbias.n368 Vbias 0.0972718
R21191 Vbias.n371 Vbias 0.0972718
R21192 Vbias.n374 Vbias 0.0972718
R21193 Vbias.n416 Vbias 0.0972718
R21194 Vbias.n413 Vbias 0.0972718
R21195 Vbias.n410 Vbias 0.0972718
R21196 Vbias.n407 Vbias 0.0972718
R21197 Vbias.n404 Vbias 0.0972718
R21198 Vbias.n401 Vbias 0.0972718
R21199 Vbias.n398 Vbias 0.0972718
R21200 Vbias.n395 Vbias 0.0972718
R21201 Vbias.n392 Vbias 0.0972718
R21202 Vbias.n389 Vbias 0.0972718
R21203 Vbias.n386 Vbias 0.0972718
R21204 Vbias.n383 Vbias 0.0972718
R21205 Vbias.n380 Vbias 0.0972718
R21206 Vbias.n377 Vbias 0.0972718
R21207 Vbias Vbias.n995 0.0972718
R21208 Vbias.n376 Vbias 0.0489375
R21209 Vbias.n8 Vbias 0.0489375
R21210 Vbias.n334 Vbias 0.0489375
R21211 Vbias.n285 Vbias 0.0489375
R21212 Vbias.n278 Vbias 0.0489375
R21213 Vbias.n280 Vbias 0.0489375
R21214 Vbias.n274 Vbias 0.0489375
R21215 Vbias.n229 Vbias 0.0489375
R21216 Vbias.n185 Vbias 0.0489375
R21217 Vbias.n225 Vbias 0.0489375
R21218 Vbias.n181 Vbias 0.0489375
R21219 Vbias.n122 Vbias 0.0489375
R21220 Vbias.n82 Vbias 0.0489375
R21221 Vbias.n176 Vbias 0.0489375
R21222 Vbias.n78 Vbias 0.0489375
R21223 Vbias.n75 Vbias 0.0489375
R21224 Vbias.n414 Vbias 0.0489375
R21225 Vbias.n372 Vbias 0.0489375
R21226 Vbias.n333 Vbias 0.0489375
R21227 Vbias.n331 Vbias 0.0489375
R21228 Vbias.n543 Vbias 0.0489375
R21229 Vbias.n272 Vbias 0.0489375
R21230 Vbias.n270 Vbias 0.0489375
R21231 Vbias.n636 Vbias 0.0489375
R21232 Vbias.n186 Vbias 0.0489375
R21233 Vbias.n188 Vbias 0.0489375
R21234 Vbias.n767 Vbias 0.0489375
R21235 Vbias.n85 Vbias 0.0489375
R21236 Vbias.n83 Vbias 0.0489375
R21237 Vbias.n136 Vbias 0.0489375
R21238 Vbias.n77 Vbias 0.0489375
R21239 Vbias.n74 Vbias 0.0489375
R21240 Vbias.n411 Vbias 0.0489375
R21241 Vbias.n369 Vbias 0.0489375
R21242 Vbias.n326 Vbias 0.0489375
R21243 Vbias.n328 Vbias 0.0489375
R21244 Vbias.n540 Vbias 0.0489375
R21245 Vbias.n267 Vbias 0.0489375
R21246 Vbias.n269 Vbias 0.0489375
R21247 Vbias.n639 Vbias 0.0489375
R21248 Vbias.n191 Vbias 0.0489375
R21249 Vbias.n189 Vbias 0.0489375
R21250 Vbias.n770 Vbias 0.0489375
R21251 Vbias.n86 Vbias 0.0489375
R21252 Vbias.n88 Vbias 0.0489375
R21253 Vbias.n139 Vbias 0.0489375
R21254 Vbias.n72 Vbias 0.0489375
R21255 Vbias.n69 Vbias 0.0489375
R21256 Vbias.n408 Vbias 0.0489375
R21257 Vbias.n366 Vbias 0.0489375
R21258 Vbias.n325 Vbias 0.0489375
R21259 Vbias.n323 Vbias 0.0489375
R21260 Vbias.n537 Vbias 0.0489375
R21261 Vbias.n266 Vbias 0.0489375
R21262 Vbias.n264 Vbias 0.0489375
R21263 Vbias.n642 Vbias 0.0489375
R21264 Vbias.n192 Vbias 0.0489375
R21265 Vbias.n194 Vbias 0.0489375
R21266 Vbias.n773 Vbias 0.0489375
R21267 Vbias.n91 Vbias 0.0489375
R21268 Vbias.n89 Vbias 0.0489375
R21269 Vbias.n142 Vbias 0.0489375
R21270 Vbias.n71 Vbias 0.0489375
R21271 Vbias.n68 Vbias 0.0489375
R21272 Vbias.n405 Vbias 0.0489375
R21273 Vbias.n363 Vbias 0.0489375
R21274 Vbias.n320 Vbias 0.0489375
R21275 Vbias.n322 Vbias 0.0489375
R21276 Vbias.n534 Vbias 0.0489375
R21277 Vbias.n261 Vbias 0.0489375
R21278 Vbias.n263 Vbias 0.0489375
R21279 Vbias.n645 Vbias 0.0489375
R21280 Vbias.n197 Vbias 0.0489375
R21281 Vbias.n195 Vbias 0.0489375
R21282 Vbias.n776 Vbias 0.0489375
R21283 Vbias.n92 Vbias 0.0489375
R21284 Vbias.n94 Vbias 0.0489375
R21285 Vbias.n145 Vbias 0.0489375
R21286 Vbias.n66 Vbias 0.0489375
R21287 Vbias.n63 Vbias 0.0489375
R21288 Vbias.n402 Vbias 0.0489375
R21289 Vbias.n360 Vbias 0.0489375
R21290 Vbias.n319 Vbias 0.0489375
R21291 Vbias.n317 Vbias 0.0489375
R21292 Vbias.n531 Vbias 0.0489375
R21293 Vbias.n260 Vbias 0.0489375
R21294 Vbias.n258 Vbias 0.0489375
R21295 Vbias.n648 Vbias 0.0489375
R21296 Vbias.n198 Vbias 0.0489375
R21297 Vbias.n200 Vbias 0.0489375
R21298 Vbias.n779 Vbias 0.0489375
R21299 Vbias.n97 Vbias 0.0489375
R21300 Vbias.n95 Vbias 0.0489375
R21301 Vbias.n148 Vbias 0.0489375
R21302 Vbias.n65 Vbias 0.0489375
R21303 Vbias.n62 Vbias 0.0489375
R21304 Vbias.n399 Vbias 0.0489375
R21305 Vbias.n357 Vbias 0.0489375
R21306 Vbias.n314 Vbias 0.0489375
R21307 Vbias.n316 Vbias 0.0489375
R21308 Vbias.n528 Vbias 0.0489375
R21309 Vbias.n255 Vbias 0.0489375
R21310 Vbias.n257 Vbias 0.0489375
R21311 Vbias.n651 Vbias 0.0489375
R21312 Vbias.n203 Vbias 0.0489375
R21313 Vbias.n201 Vbias 0.0489375
R21314 Vbias.n782 Vbias 0.0489375
R21315 Vbias.n98 Vbias 0.0489375
R21316 Vbias.n100 Vbias 0.0489375
R21317 Vbias.n151 Vbias 0.0489375
R21318 Vbias.n60 Vbias 0.0489375
R21319 Vbias.n57 Vbias 0.0489375
R21320 Vbias.n396 Vbias 0.0489375
R21321 Vbias.n354 Vbias 0.0489375
R21322 Vbias.n313 Vbias 0.0489375
R21323 Vbias.n311 Vbias 0.0489375
R21324 Vbias.n525 Vbias 0.0489375
R21325 Vbias.n254 Vbias 0.0489375
R21326 Vbias.n252 Vbias 0.0489375
R21327 Vbias.n654 Vbias 0.0489375
R21328 Vbias.n204 Vbias 0.0489375
R21329 Vbias.n206 Vbias 0.0489375
R21330 Vbias.n785 Vbias 0.0489375
R21331 Vbias.n103 Vbias 0.0489375
R21332 Vbias.n101 Vbias 0.0489375
R21333 Vbias.n154 Vbias 0.0489375
R21334 Vbias.n59 Vbias 0.0489375
R21335 Vbias.n56 Vbias 0.0489375
R21336 Vbias.n393 Vbias 0.0489375
R21337 Vbias.n351 Vbias 0.0489375
R21338 Vbias.n308 Vbias 0.0489375
R21339 Vbias.n310 Vbias 0.0489375
R21340 Vbias.n522 Vbias 0.0489375
R21341 Vbias.n249 Vbias 0.0489375
R21342 Vbias.n251 Vbias 0.0489375
R21343 Vbias.n657 Vbias 0.0489375
R21344 Vbias.n209 Vbias 0.0489375
R21345 Vbias.n207 Vbias 0.0489375
R21346 Vbias.n788 Vbias 0.0489375
R21347 Vbias.n104 Vbias 0.0489375
R21348 Vbias.n106 Vbias 0.0489375
R21349 Vbias.n157 Vbias 0.0489375
R21350 Vbias.n54 Vbias 0.0489375
R21351 Vbias.n51 Vbias 0.0489375
R21352 Vbias.n390 Vbias 0.0489375
R21353 Vbias.n348 Vbias 0.0489375
R21354 Vbias.n307 Vbias 0.0489375
R21355 Vbias.n305 Vbias 0.0489375
R21356 Vbias.n519 Vbias 0.0489375
R21357 Vbias.n248 Vbias 0.0489375
R21358 Vbias.n246 Vbias 0.0489375
R21359 Vbias.n660 Vbias 0.0489375
R21360 Vbias.n210 Vbias 0.0489375
R21361 Vbias.n212 Vbias 0.0489375
R21362 Vbias.n791 Vbias 0.0489375
R21363 Vbias.n109 Vbias 0.0489375
R21364 Vbias.n107 Vbias 0.0489375
R21365 Vbias.n160 Vbias 0.0489375
R21366 Vbias.n53 Vbias 0.0489375
R21367 Vbias.n50 Vbias 0.0489375
R21368 Vbias.n387 Vbias 0.0489375
R21369 Vbias.n345 Vbias 0.0489375
R21370 Vbias.n302 Vbias 0.0489375
R21371 Vbias.n304 Vbias 0.0489375
R21372 Vbias.n516 Vbias 0.0489375
R21373 Vbias.n243 Vbias 0.0489375
R21374 Vbias.n245 Vbias 0.0489375
R21375 Vbias.n663 Vbias 0.0489375
R21376 Vbias.n215 Vbias 0.0489375
R21377 Vbias.n213 Vbias 0.0489375
R21378 Vbias.n794 Vbias 0.0489375
R21379 Vbias.n110 Vbias 0.0489375
R21380 Vbias.n112 Vbias 0.0489375
R21381 Vbias.n163 Vbias 0.0489375
R21382 Vbias.n48 Vbias 0.0489375
R21383 Vbias.n45 Vbias 0.0489375
R21384 Vbias.n384 Vbias 0.0489375
R21385 Vbias.n342 Vbias 0.0489375
R21386 Vbias.n301 Vbias 0.0489375
R21387 Vbias.n299 Vbias 0.0489375
R21388 Vbias.n513 Vbias 0.0489375
R21389 Vbias.n242 Vbias 0.0489375
R21390 Vbias.n240 Vbias 0.0489375
R21391 Vbias.n666 Vbias 0.0489375
R21392 Vbias.n216 Vbias 0.0489375
R21393 Vbias.n218 Vbias 0.0489375
R21394 Vbias.n797 Vbias 0.0489375
R21395 Vbias.n115 Vbias 0.0489375
R21396 Vbias.n113 Vbias 0.0489375
R21397 Vbias.n166 Vbias 0.0489375
R21398 Vbias.n47 Vbias 0.0489375
R21399 Vbias.n44 Vbias 0.0489375
R21400 Vbias.n381 Vbias 0.0489375
R21401 Vbias.n339 Vbias 0.0489375
R21402 Vbias.n296 Vbias 0.0489375
R21403 Vbias.n298 Vbias 0.0489375
R21404 Vbias.n510 Vbias 0.0489375
R21405 Vbias.n237 Vbias 0.0489375
R21406 Vbias.n239 Vbias 0.0489375
R21407 Vbias.n669 Vbias 0.0489375
R21408 Vbias.n221 Vbias 0.0489375
R21409 Vbias.n219 Vbias 0.0489375
R21410 Vbias.n800 Vbias 0.0489375
R21411 Vbias.n116 Vbias 0.0489375
R21412 Vbias.n118 Vbias 0.0489375
R21413 Vbias.n169 Vbias 0.0489375
R21414 Vbias.n42 Vbias 0.0489375
R21415 Vbias.n39 Vbias 0.0489375
R21416 Vbias.n378 Vbias 0.0489375
R21417 Vbias.n336 Vbias 0.0489375
R21418 Vbias.n288 Vbias 0.0489375
R21419 Vbias.n286 Vbias 0.0489375
R21420 Vbias.n507 Vbias 0.0489375
R21421 Vbias.n236 Vbias 0.0489375
R21422 Vbias.n234 Vbias 0.0489375
R21423 Vbias.n672 Vbias 0.0489375
R21424 Vbias.n222 Vbias 0.0489375
R21425 Vbias.n224 Vbias 0.0489375
R21426 Vbias.n803 Vbias 0.0489375
R21427 Vbias.n121 Vbias 0.0489375
R21428 Vbias.n119 Vbias 0.0489375
R21429 Vbias.n172 Vbias 0.0489375
R21430 Vbias.n41 Vbias 0.0489375
R21431 Vbias.n38 Vbias 0.0489375
R21432 Vbias.n10 Vbias 0.0489375
R21433 Vbias.n9 Vbias 0.0489375
R21434 Vbias.n12 Vbias 0.0489375
R21435 Vbias.n14 Vbias 0.0489375
R21436 Vbias.n16 Vbias 0.0489375
R21437 Vbias.n18 Vbias 0.0489375
R21438 Vbias.n20 Vbias 0.0489375
R21439 Vbias.n22 Vbias 0.0489375
R21440 Vbias.n24 Vbias 0.0489375
R21441 Vbias.n26 Vbias 0.0489375
R21442 Vbias.n28 Vbias 0.0489375
R21443 Vbias.n30 Vbias 0.0489375
R21444 Vbias.n32 Vbias 0.0489375
R21445 Vbias.n34 Vbias 0.0489375
R21446 Vbias.n36 Vbias 0.0489375
R21447 Vbias.n129 Vbias 0.0489375
R21448 Vbias.n904 Vbias 0.0489375
R21449 Vbias.n128 Vbias 0.0489375
R21450 Vbias.n79 Vbias 0.0489375
R21451 Vbias.n125 Vbias 0.0489375
R21452 Vbias.n893 Vbias 0.0489375
R21453 Vbias.n807 Vbias 0.0489375
R21454 Vbias.n182 Vbias 0.0489375
R21455 Vbias.n226 Vbias 0.0489375
R21456 Vbias.n634 Vbias 0.0489375
R21457 Vbias.n629 Vbias 0.0489375
R21458 Vbias.n273 Vbias 0.0489375
R21459 Vbias.n279 Vbias 0.0489375
R21460 Vbias.n329 Vbias 0.0489375
R21461 Vbias.n292 Vbias 0.0489375
R21462 Vbias.n6 Vbias 0.0489375
R21463 Vbias.n335 Vbias 0.0489375
R21464 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R21465 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R21466 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R21467 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R21468 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R21469 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R21470 XThR.Tn[12] XThR.Tn[12].n78 161.363
R21471 XThR.Tn[12] XThR.Tn[12].n73 161.363
R21472 XThR.Tn[12] XThR.Tn[12].n68 161.363
R21473 XThR.Tn[12] XThR.Tn[12].n63 161.363
R21474 XThR.Tn[12] XThR.Tn[12].n58 161.363
R21475 XThR.Tn[12] XThR.Tn[12].n53 161.363
R21476 XThR.Tn[12] XThR.Tn[12].n48 161.363
R21477 XThR.Tn[12] XThR.Tn[12].n43 161.363
R21478 XThR.Tn[12] XThR.Tn[12].n38 161.363
R21479 XThR.Tn[12] XThR.Tn[12].n33 161.363
R21480 XThR.Tn[12] XThR.Tn[12].n28 161.363
R21481 XThR.Tn[12] XThR.Tn[12].n23 161.363
R21482 XThR.Tn[12] XThR.Tn[12].n18 161.363
R21483 XThR.Tn[12] XThR.Tn[12].n13 161.363
R21484 XThR.Tn[12] XThR.Tn[12].n8 161.363
R21485 XThR.Tn[12] XThR.Tn[12].n6 161.363
R21486 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R21487 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R21488 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R21489 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R21490 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R21491 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R21492 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R21493 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R21494 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R21495 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R21496 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R21497 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R21498 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R21499 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R21500 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R21501 XThR.Tn[12].n79 XThR.Tn[12].t56 161.106
R21502 XThR.Tn[12].n78 XThR.Tn[12].t58 161.106
R21503 XThR.Tn[12].n74 XThR.Tn[12].t62 161.106
R21504 XThR.Tn[12].n73 XThR.Tn[12].t67 161.106
R21505 XThR.Tn[12].n69 XThR.Tn[12].t44 161.106
R21506 XThR.Tn[12].n68 XThR.Tn[12].t49 161.106
R21507 XThR.Tn[12].n64 XThR.Tn[12].t27 161.106
R21508 XThR.Tn[12].n63 XThR.Tn[12].t29 161.106
R21509 XThR.Tn[12].n59 XThR.Tn[12].t55 161.106
R21510 XThR.Tn[12].n58 XThR.Tn[12].t57 161.106
R21511 XThR.Tn[12].n54 XThR.Tn[12].t17 161.106
R21512 XThR.Tn[12].n53 XThR.Tn[12].t22 161.106
R21513 XThR.Tn[12].n49 XThR.Tn[12].t60 161.106
R21514 XThR.Tn[12].n48 XThR.Tn[12].t65 161.106
R21515 XThR.Tn[12].n44 XThR.Tn[12].t41 161.106
R21516 XThR.Tn[12].n43 XThR.Tn[12].t46 161.106
R21517 XThR.Tn[12].n39 XThR.Tn[12].t26 161.106
R21518 XThR.Tn[12].n38 XThR.Tn[12].t28 161.106
R21519 XThR.Tn[12].n34 XThR.Tn[12].t31 161.106
R21520 XThR.Tn[12].n33 XThR.Tn[12].t36 161.106
R21521 XThR.Tn[12].n29 XThR.Tn[12].t16 161.106
R21522 XThR.Tn[12].n28 XThR.Tn[12].t21 161.106
R21523 XThR.Tn[12].n24 XThR.Tn[12].t43 161.106
R21524 XThR.Tn[12].n23 XThR.Tn[12].t48 161.106
R21525 XThR.Tn[12].n19 XThR.Tn[12].t13 161.106
R21526 XThR.Tn[12].n18 XThR.Tn[12].t19 161.106
R21527 XThR.Tn[12].n14 XThR.Tn[12].t59 161.106
R21528 XThR.Tn[12].n13 XThR.Tn[12].t63 161.106
R21529 XThR.Tn[12].n9 XThR.Tn[12].t24 161.106
R21530 XThR.Tn[12].n8 XThR.Tn[12].t25 161.106
R21531 XThR.Tn[12].n6 XThR.Tn[12].t70 161.106
R21532 XThR.Tn[12].n79 XThR.Tn[12].t73 154.679
R21533 XThR.Tn[12].n78 XThR.Tn[12].t15 154.679
R21534 XThR.Tn[12].n74 XThR.Tn[12].t52 154.679
R21535 XThR.Tn[12].n73 XThR.Tn[12].t54 154.679
R21536 XThR.Tn[12].n69 XThR.Tn[12].t33 154.679
R21537 XThR.Tn[12].n68 XThR.Tn[12].t38 154.679
R21538 XThR.Tn[12].n64 XThR.Tn[12].t64 154.679
R21539 XThR.Tn[12].n63 XThR.Tn[12].t68 154.679
R21540 XThR.Tn[12].n59 XThR.Tn[12].t45 154.679
R21541 XThR.Tn[12].n58 XThR.Tn[12].t50 154.679
R21542 XThR.Tn[12].n54 XThR.Tn[12].t72 154.679
R21543 XThR.Tn[12].n53 XThR.Tn[12].t12 154.679
R21544 XThR.Tn[12].n49 XThR.Tn[12].t34 154.679
R21545 XThR.Tn[12].n48 XThR.Tn[12].t39 154.679
R21546 XThR.Tn[12].n44 XThR.Tn[12].t18 154.679
R21547 XThR.Tn[12].n43 XThR.Tn[12].t23 154.679
R21548 XThR.Tn[12].n39 XThR.Tn[12].t61 154.679
R21549 XThR.Tn[12].n38 XThR.Tn[12].t66 154.679
R21550 XThR.Tn[12].n34 XThR.Tn[12].t42 154.679
R21551 XThR.Tn[12].n33 XThR.Tn[12].t47 154.679
R21552 XThR.Tn[12].n29 XThR.Tn[12].t51 154.679
R21553 XThR.Tn[12].n28 XThR.Tn[12].t53 154.679
R21554 XThR.Tn[12].n24 XThR.Tn[12].t32 154.679
R21555 XThR.Tn[12].n23 XThR.Tn[12].t37 154.679
R21556 XThR.Tn[12].n19 XThR.Tn[12].t69 154.679
R21557 XThR.Tn[12].n18 XThR.Tn[12].t71 154.679
R21558 XThR.Tn[12].n14 XThR.Tn[12].t30 154.679
R21559 XThR.Tn[12].n13 XThR.Tn[12].t35 154.679
R21560 XThR.Tn[12].n9 XThR.Tn[12].t14 154.679
R21561 XThR.Tn[12].n8 XThR.Tn[12].t20 154.679
R21562 XThR.Tn[12].n6 XThR.Tn[12].t40 154.679
R21563 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R21564 XThR.Tn[12].n85 XThR.Tn[12].t2 26.5955
R21565 XThR.Tn[12].n85 XThR.Tn[12].t0 26.5955
R21566 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R21567 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R21568 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R21569 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R21570 XThR.Tn[12].n86 XThR.Tn[12].t3 26.5955
R21571 XThR.Tn[12].n86 XThR.Tn[12].t1 26.5955
R21572 XThR.Tn[12].n4 XThR.Tn[12].t6 24.9236
R21573 XThR.Tn[12].n4 XThR.Tn[12].t4 24.9236
R21574 XThR.Tn[12].n3 XThR.Tn[12].t7 24.9236
R21575 XThR.Tn[12].n3 XThR.Tn[12].t5 24.9236
R21576 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R21577 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R21578 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R21579 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R21580 XThR.Tn[12] XThR.Tn[12].n7 5.34871
R21581 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R21582 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R21583 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R21584 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R21585 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R21586 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R21587 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R21588 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R21589 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R21590 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R21591 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R21592 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R21593 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R21594 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R21595 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R21596 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R21597 XThR.Tn[12].n12 XThR.Tn[12] 2.51836
R21598 XThR.Tn[12].n17 XThR.Tn[12] 2.51836
R21599 XThR.Tn[12].n22 XThR.Tn[12] 2.51836
R21600 XThR.Tn[12].n27 XThR.Tn[12] 2.51836
R21601 XThR.Tn[12].n32 XThR.Tn[12] 2.51836
R21602 XThR.Tn[12].n37 XThR.Tn[12] 2.51836
R21603 XThR.Tn[12].n42 XThR.Tn[12] 2.51836
R21604 XThR.Tn[12].n47 XThR.Tn[12] 2.51836
R21605 XThR.Tn[12].n52 XThR.Tn[12] 2.51836
R21606 XThR.Tn[12].n57 XThR.Tn[12] 2.51836
R21607 XThR.Tn[12].n62 XThR.Tn[12] 2.51836
R21608 XThR.Tn[12].n67 XThR.Tn[12] 2.51836
R21609 XThR.Tn[12].n72 XThR.Tn[12] 2.51836
R21610 XThR.Tn[12].n77 XThR.Tn[12] 2.51836
R21611 XThR.Tn[12].n82 XThR.Tn[12] 2.51836
R21612 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R21613 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R21614 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R21615 XThR.Tn[12] XThR.Tn[12].n12 0.848714
R21616 XThR.Tn[12] XThR.Tn[12].n17 0.848714
R21617 XThR.Tn[12] XThR.Tn[12].n22 0.848714
R21618 XThR.Tn[12] XThR.Tn[12].n27 0.848714
R21619 XThR.Tn[12] XThR.Tn[12].n32 0.848714
R21620 XThR.Tn[12] XThR.Tn[12].n37 0.848714
R21621 XThR.Tn[12] XThR.Tn[12].n42 0.848714
R21622 XThR.Tn[12] XThR.Tn[12].n47 0.848714
R21623 XThR.Tn[12] XThR.Tn[12].n52 0.848714
R21624 XThR.Tn[12] XThR.Tn[12].n57 0.848714
R21625 XThR.Tn[12] XThR.Tn[12].n62 0.848714
R21626 XThR.Tn[12] XThR.Tn[12].n67 0.848714
R21627 XThR.Tn[12] XThR.Tn[12].n72 0.848714
R21628 XThR.Tn[12] XThR.Tn[12].n77 0.848714
R21629 XThR.Tn[12] XThR.Tn[12].n82 0.848714
R21630 XThR.Tn[12].n7 XThR.Tn[12] 0.485653
R21631 XThR.Tn[12].n80 XThR.Tn[12] 0.21482
R21632 XThR.Tn[12].n75 XThR.Tn[12] 0.21482
R21633 XThR.Tn[12].n70 XThR.Tn[12] 0.21482
R21634 XThR.Tn[12].n65 XThR.Tn[12] 0.21482
R21635 XThR.Tn[12].n60 XThR.Tn[12] 0.21482
R21636 XThR.Tn[12].n55 XThR.Tn[12] 0.21482
R21637 XThR.Tn[12].n50 XThR.Tn[12] 0.21482
R21638 XThR.Tn[12].n45 XThR.Tn[12] 0.21482
R21639 XThR.Tn[12].n40 XThR.Tn[12] 0.21482
R21640 XThR.Tn[12].n35 XThR.Tn[12] 0.21482
R21641 XThR.Tn[12].n30 XThR.Tn[12] 0.21482
R21642 XThR.Tn[12].n25 XThR.Tn[12] 0.21482
R21643 XThR.Tn[12].n20 XThR.Tn[12] 0.21482
R21644 XThR.Tn[12].n15 XThR.Tn[12] 0.21482
R21645 XThR.Tn[12].n10 XThR.Tn[12] 0.21482
R21646 XThR.Tn[12].n81 XThR.Tn[12] 0.0608448
R21647 XThR.Tn[12].n76 XThR.Tn[12] 0.0608448
R21648 XThR.Tn[12].n71 XThR.Tn[12] 0.0608448
R21649 XThR.Tn[12].n66 XThR.Tn[12] 0.0608448
R21650 XThR.Tn[12].n61 XThR.Tn[12] 0.0608448
R21651 XThR.Tn[12].n56 XThR.Tn[12] 0.0608448
R21652 XThR.Tn[12].n51 XThR.Tn[12] 0.0608448
R21653 XThR.Tn[12].n46 XThR.Tn[12] 0.0608448
R21654 XThR.Tn[12].n41 XThR.Tn[12] 0.0608448
R21655 XThR.Tn[12].n36 XThR.Tn[12] 0.0608448
R21656 XThR.Tn[12].n31 XThR.Tn[12] 0.0608448
R21657 XThR.Tn[12].n26 XThR.Tn[12] 0.0608448
R21658 XThR.Tn[12].n21 XThR.Tn[12] 0.0608448
R21659 XThR.Tn[12].n16 XThR.Tn[12] 0.0608448
R21660 XThR.Tn[12].n11 XThR.Tn[12] 0.0608448
R21661 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R21662 XThR.Tn[12] XThR.Tn[12].n83 0.038
R21663 XThR.Tn[12].n7 XThR.Tn[12] 0.00744444
R21664 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00265517
R21665 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00265517
R21666 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00265517
R21667 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00265517
R21668 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00265517
R21669 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00265517
R21670 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00265517
R21671 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00265517
R21672 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00265517
R21673 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00265517
R21674 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00265517
R21675 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00265517
R21676 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00265517
R21677 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00265517
R21678 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00265517
R21679 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R21680 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R21681 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R21682 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R21683 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R21684 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R21685 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R21686 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R21687 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R21688 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R21689 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R21690 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R21691 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R21692 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R21693 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R21694 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R21695 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R21696 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R21697 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R21698 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R21699 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R21700 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R21701 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R21702 XThC.XTB1.Y.n0 XThC.XTB1.Y.t1 132.067
R21703 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R21704 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R21705 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R21706 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R21707 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R21708 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R21709 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R21710 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R21711 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R21712 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R21713 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R21714 XThC.XTB1.Y.n2 XThC.XTB1.Y.t2 26.5955
R21715 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R21716 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R21717 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R21718 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R21719 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R21720 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R21721 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R21722 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R21723 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R21724 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R21725 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R21726 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R21727 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R21728 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R21729 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R21730 XThC.Tn[8].n71 XThC.Tn[8].n70 256.104
R21731 XThC.Tn[8].n75 XThC.Tn[8].n74 243.679
R21732 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R21733 XThC.Tn[8].n75 XThC.Tn[8].n73 205.28
R21734 XThC.Tn[8].n71 XThC.Tn[8].n69 202.095
R21735 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R21736 XThC.Tn[8].n65 XThC.Tn[8].n63 161.365
R21737 XThC.Tn[8].n61 XThC.Tn[8].n59 161.365
R21738 XThC.Tn[8].n57 XThC.Tn[8].n55 161.365
R21739 XThC.Tn[8].n53 XThC.Tn[8].n51 161.365
R21740 XThC.Tn[8].n49 XThC.Tn[8].n47 161.365
R21741 XThC.Tn[8].n45 XThC.Tn[8].n43 161.365
R21742 XThC.Tn[8].n41 XThC.Tn[8].n39 161.365
R21743 XThC.Tn[8].n37 XThC.Tn[8].n35 161.365
R21744 XThC.Tn[8].n33 XThC.Tn[8].n31 161.365
R21745 XThC.Tn[8].n29 XThC.Tn[8].n27 161.365
R21746 XThC.Tn[8].n25 XThC.Tn[8].n23 161.365
R21747 XThC.Tn[8].n21 XThC.Tn[8].n19 161.365
R21748 XThC.Tn[8].n17 XThC.Tn[8].n15 161.365
R21749 XThC.Tn[8].n13 XThC.Tn[8].n11 161.365
R21750 XThC.Tn[8].n9 XThC.Tn[8].n7 161.365
R21751 XThC.Tn[8].n6 XThC.Tn[8].n4 161.365
R21752 XThC.Tn[8].n63 XThC.Tn[8].t34 161.106
R21753 XThC.Tn[8].n59 XThC.Tn[8].t14 161.106
R21754 XThC.Tn[8].n55 XThC.Tn[8].t12 161.106
R21755 XThC.Tn[8].n51 XThC.Tn[8].t43 161.106
R21756 XThC.Tn[8].n47 XThC.Tn[8].t24 161.106
R21757 XThC.Tn[8].n43 XThC.Tn[8].t21 161.106
R21758 XThC.Tn[8].n39 XThC.Tn[8].t41 161.106
R21759 XThC.Tn[8].n35 XThC.Tn[8].t32 161.106
R21760 XThC.Tn[8].n31 XThC.Tn[8].t30 161.106
R21761 XThC.Tn[8].n27 XThC.Tn[8].t19 161.106
R21762 XThC.Tn[8].n23 XThC.Tn[8].t40 161.106
R21763 XThC.Tn[8].n19 XThC.Tn[8].t29 161.106
R21764 XThC.Tn[8].n15 XThC.Tn[8].t18 161.106
R21765 XThC.Tn[8].n11 XThC.Tn[8].t17 161.106
R21766 XThC.Tn[8].n7 XThC.Tn[8].t36 161.106
R21767 XThC.Tn[8].n4 XThC.Tn[8].t26 161.106
R21768 XThC.Tn[8].n63 XThC.Tn[8].t22 154.679
R21769 XThC.Tn[8].n59 XThC.Tn[8].t33 154.679
R21770 XThC.Tn[8].n55 XThC.Tn[8].t31 154.679
R21771 XThC.Tn[8].n51 XThC.Tn[8].t28 154.679
R21772 XThC.Tn[8].n47 XThC.Tn[8].t42 154.679
R21773 XThC.Tn[8].n43 XThC.Tn[8].t39 154.679
R21774 XThC.Tn[8].n39 XThC.Tn[8].t27 154.679
R21775 XThC.Tn[8].n35 XThC.Tn[8].t20 154.679
R21776 XThC.Tn[8].n31 XThC.Tn[8].t16 154.679
R21777 XThC.Tn[8].n27 XThC.Tn[8].t38 154.679
R21778 XThC.Tn[8].n23 XThC.Tn[8].t25 154.679
R21779 XThC.Tn[8].n19 XThC.Tn[8].t15 154.679
R21780 XThC.Tn[8].n15 XThC.Tn[8].t37 154.679
R21781 XThC.Tn[8].n11 XThC.Tn[8].t35 154.679
R21782 XThC.Tn[8].n7 XThC.Tn[8].t23 154.679
R21783 XThC.Tn[8].n4 XThC.Tn[8].t13 154.679
R21784 XThC.Tn[8].n69 XThC.Tn[8].t5 26.5955
R21785 XThC.Tn[8].n69 XThC.Tn[8].t6 26.5955
R21786 XThC.Tn[8].n70 XThC.Tn[8].t4 26.5955
R21787 XThC.Tn[8].n70 XThC.Tn[8].t7 26.5955
R21788 XThC.Tn[8].n73 XThC.Tn[8].t2 26.5955
R21789 XThC.Tn[8].n73 XThC.Tn[8].t1 26.5955
R21790 XThC.Tn[8].n74 XThC.Tn[8].t0 26.5955
R21791 XThC.Tn[8].n74 XThC.Tn[8].t3 26.5955
R21792 XThC.Tn[8].n1 XThC.Tn[8].t11 24.9236
R21793 XThC.Tn[8].n1 XThC.Tn[8].t10 24.9236
R21794 XThC.Tn[8].n0 XThC.Tn[8].t9 24.9236
R21795 XThC.Tn[8].n0 XThC.Tn[8].t8 24.9236
R21796 XThC.Tn[8] XThC.Tn[8].n75 22.9652
R21797 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R21798 XThC.Tn[8].n72 XThC.Tn[8].n71 13.9299
R21799 XThC.Tn[8] XThC.Tn[8].n72 13.9299
R21800 XThC.Tn[8] XThC.Tn[8].n6 8.0245
R21801 XThC.Tn[8].n66 XThC.Tn[8].n65 7.9105
R21802 XThC.Tn[8].n62 XThC.Tn[8].n61 7.9105
R21803 XThC.Tn[8].n58 XThC.Tn[8].n57 7.9105
R21804 XThC.Tn[8].n54 XThC.Tn[8].n53 7.9105
R21805 XThC.Tn[8].n50 XThC.Tn[8].n49 7.9105
R21806 XThC.Tn[8].n46 XThC.Tn[8].n45 7.9105
R21807 XThC.Tn[8].n42 XThC.Tn[8].n41 7.9105
R21808 XThC.Tn[8].n38 XThC.Tn[8].n37 7.9105
R21809 XThC.Tn[8].n34 XThC.Tn[8].n33 7.9105
R21810 XThC.Tn[8].n30 XThC.Tn[8].n29 7.9105
R21811 XThC.Tn[8].n26 XThC.Tn[8].n25 7.9105
R21812 XThC.Tn[8].n22 XThC.Tn[8].n21 7.9105
R21813 XThC.Tn[8].n18 XThC.Tn[8].n17 7.9105
R21814 XThC.Tn[8].n14 XThC.Tn[8].n13 7.9105
R21815 XThC.Tn[8].n10 XThC.Tn[8].n9 7.9105
R21816 XThC.Tn[8].n68 XThC.Tn[8].n67 7.42331
R21817 XThC.Tn[8].n67 XThC.Tn[8] 4.24005
R21818 XThC.Tn[8].n72 XThC.Tn[8].n68 2.99115
R21819 XThC.Tn[8].n72 XThC.Tn[8] 2.87153
R21820 XThC.Tn[8].n68 XThC.Tn[8] 2.2734
R21821 XThC.Tn[8].n3 XThC.Tn[8] 0.672375
R21822 XThC.Tn[8].n10 XThC.Tn[8] 0.235138
R21823 XThC.Tn[8].n14 XThC.Tn[8] 0.235138
R21824 XThC.Tn[8].n18 XThC.Tn[8] 0.235138
R21825 XThC.Tn[8].n22 XThC.Tn[8] 0.235138
R21826 XThC.Tn[8].n26 XThC.Tn[8] 0.235138
R21827 XThC.Tn[8].n30 XThC.Tn[8] 0.235138
R21828 XThC.Tn[8].n34 XThC.Tn[8] 0.235138
R21829 XThC.Tn[8].n38 XThC.Tn[8] 0.235138
R21830 XThC.Tn[8].n42 XThC.Tn[8] 0.235138
R21831 XThC.Tn[8].n46 XThC.Tn[8] 0.235138
R21832 XThC.Tn[8].n50 XThC.Tn[8] 0.235138
R21833 XThC.Tn[8].n54 XThC.Tn[8] 0.235138
R21834 XThC.Tn[8].n58 XThC.Tn[8] 0.235138
R21835 XThC.Tn[8].n62 XThC.Tn[8] 0.235138
R21836 XThC.Tn[8].n66 XThC.Tn[8] 0.235138
R21837 XThC.Tn[8].n67 XThC.Tn[8].n3 0.220435
R21838 XThC.Tn[8].n3 XThC.Tn[8] 0.168469
R21839 XThC.Tn[8] XThC.Tn[8].n10 0.114505
R21840 XThC.Tn[8] XThC.Tn[8].n14 0.114505
R21841 XThC.Tn[8] XThC.Tn[8].n18 0.114505
R21842 XThC.Tn[8] XThC.Tn[8].n22 0.114505
R21843 XThC.Tn[8] XThC.Tn[8].n26 0.114505
R21844 XThC.Tn[8] XThC.Tn[8].n30 0.114505
R21845 XThC.Tn[8] XThC.Tn[8].n34 0.114505
R21846 XThC.Tn[8] XThC.Tn[8].n38 0.114505
R21847 XThC.Tn[8] XThC.Tn[8].n42 0.114505
R21848 XThC.Tn[8] XThC.Tn[8].n46 0.114505
R21849 XThC.Tn[8] XThC.Tn[8].n50 0.114505
R21850 XThC.Tn[8] XThC.Tn[8].n54 0.114505
R21851 XThC.Tn[8] XThC.Tn[8].n58 0.114505
R21852 XThC.Tn[8] XThC.Tn[8].n62 0.114505
R21853 XThC.Tn[8] XThC.Tn[8].n66 0.114505
R21854 XThC.Tn[8].n65 XThC.Tn[8].n64 0.0599512
R21855 XThC.Tn[8].n61 XThC.Tn[8].n60 0.0599512
R21856 XThC.Tn[8].n57 XThC.Tn[8].n56 0.0599512
R21857 XThC.Tn[8].n53 XThC.Tn[8].n52 0.0599512
R21858 XThC.Tn[8].n49 XThC.Tn[8].n48 0.0599512
R21859 XThC.Tn[8].n45 XThC.Tn[8].n44 0.0599512
R21860 XThC.Tn[8].n41 XThC.Tn[8].n40 0.0599512
R21861 XThC.Tn[8].n37 XThC.Tn[8].n36 0.0599512
R21862 XThC.Tn[8].n33 XThC.Tn[8].n32 0.0599512
R21863 XThC.Tn[8].n29 XThC.Tn[8].n28 0.0599512
R21864 XThC.Tn[8].n25 XThC.Tn[8].n24 0.0599512
R21865 XThC.Tn[8].n21 XThC.Tn[8].n20 0.0599512
R21866 XThC.Tn[8].n17 XThC.Tn[8].n16 0.0599512
R21867 XThC.Tn[8].n13 XThC.Tn[8].n12 0.0599512
R21868 XThC.Tn[8].n9 XThC.Tn[8].n8 0.0599512
R21869 XThC.Tn[8].n6 XThC.Tn[8].n5 0.0599512
R21870 XThC.Tn[8].n64 XThC.Tn[8] 0.0469286
R21871 XThC.Tn[8].n60 XThC.Tn[8] 0.0469286
R21872 XThC.Tn[8].n56 XThC.Tn[8] 0.0469286
R21873 XThC.Tn[8].n52 XThC.Tn[8] 0.0469286
R21874 XThC.Tn[8].n48 XThC.Tn[8] 0.0469286
R21875 XThC.Tn[8].n44 XThC.Tn[8] 0.0469286
R21876 XThC.Tn[8].n40 XThC.Tn[8] 0.0469286
R21877 XThC.Tn[8].n36 XThC.Tn[8] 0.0469286
R21878 XThC.Tn[8].n32 XThC.Tn[8] 0.0469286
R21879 XThC.Tn[8].n28 XThC.Tn[8] 0.0469286
R21880 XThC.Tn[8].n24 XThC.Tn[8] 0.0469286
R21881 XThC.Tn[8].n20 XThC.Tn[8] 0.0469286
R21882 XThC.Tn[8].n16 XThC.Tn[8] 0.0469286
R21883 XThC.Tn[8].n12 XThC.Tn[8] 0.0469286
R21884 XThC.Tn[8].n8 XThC.Tn[8] 0.0469286
R21885 XThC.Tn[8].n5 XThC.Tn[8] 0.0469286
R21886 XThC.Tn[8].n64 XThC.Tn[8] 0.0401341
R21887 XThC.Tn[8].n60 XThC.Tn[8] 0.0401341
R21888 XThC.Tn[8].n56 XThC.Tn[8] 0.0401341
R21889 XThC.Tn[8].n52 XThC.Tn[8] 0.0401341
R21890 XThC.Tn[8].n48 XThC.Tn[8] 0.0401341
R21891 XThC.Tn[8].n44 XThC.Tn[8] 0.0401341
R21892 XThC.Tn[8].n40 XThC.Tn[8] 0.0401341
R21893 XThC.Tn[8].n36 XThC.Tn[8] 0.0401341
R21894 XThC.Tn[8].n32 XThC.Tn[8] 0.0401341
R21895 XThC.Tn[8].n28 XThC.Tn[8] 0.0401341
R21896 XThC.Tn[8].n24 XThC.Tn[8] 0.0401341
R21897 XThC.Tn[8].n20 XThC.Tn[8] 0.0401341
R21898 XThC.Tn[8].n16 XThC.Tn[8] 0.0401341
R21899 XThC.Tn[8].n12 XThC.Tn[8] 0.0401341
R21900 XThC.Tn[8].n8 XThC.Tn[8] 0.0401341
R21901 XThC.Tn[8].n5 XThC.Tn[8] 0.0401341
R21902 XThC.Tn[13].n2 XThC.Tn[13].n1 265.341
R21903 XThC.Tn[13].n5 XThC.Tn[13].n3 243.68
R21904 XThC.Tn[13].n74 XThC.Tn[13].n73 241.847
R21905 XThC.Tn[13].n5 XThC.Tn[13].n4 205.28
R21906 XThC.Tn[13].n2 XThC.Tn[13].n0 202.094
R21907 XThC.Tn[13].n74 XThC.Tn[13].n72 185
R21908 XThC.Tn[13].n68 XThC.Tn[13].n66 161.365
R21909 XThC.Tn[13].n64 XThC.Tn[13].n62 161.365
R21910 XThC.Tn[13].n60 XThC.Tn[13].n58 161.365
R21911 XThC.Tn[13].n56 XThC.Tn[13].n54 161.365
R21912 XThC.Tn[13].n52 XThC.Tn[13].n50 161.365
R21913 XThC.Tn[13].n48 XThC.Tn[13].n46 161.365
R21914 XThC.Tn[13].n44 XThC.Tn[13].n42 161.365
R21915 XThC.Tn[13].n40 XThC.Tn[13].n38 161.365
R21916 XThC.Tn[13].n36 XThC.Tn[13].n34 161.365
R21917 XThC.Tn[13].n32 XThC.Tn[13].n30 161.365
R21918 XThC.Tn[13].n28 XThC.Tn[13].n26 161.365
R21919 XThC.Tn[13].n24 XThC.Tn[13].n22 161.365
R21920 XThC.Tn[13].n20 XThC.Tn[13].n18 161.365
R21921 XThC.Tn[13].n16 XThC.Tn[13].n14 161.365
R21922 XThC.Tn[13].n12 XThC.Tn[13].n10 161.365
R21923 XThC.Tn[13].n9 XThC.Tn[13].n7 161.365
R21924 XThC.Tn[13].n66 XThC.Tn[13].t21 161.106
R21925 XThC.Tn[13].n62 XThC.Tn[13].t33 161.106
R21926 XThC.Tn[13].n58 XThC.Tn[13].t31 161.106
R21927 XThC.Tn[13].n54 XThC.Tn[13].t30 161.106
R21928 XThC.Tn[13].n50 XThC.Tn[13].t43 161.106
R21929 XThC.Tn[13].n46 XThC.Tn[13].t40 161.106
R21930 XThC.Tn[13].n42 XThC.Tn[13].t28 161.106
R21931 XThC.Tn[13].n38 XThC.Tn[13].t19 161.106
R21932 XThC.Tn[13].n34 XThC.Tn[13].t17 161.106
R21933 XThC.Tn[13].n30 XThC.Tn[13].t38 161.106
R21934 XThC.Tn[13].n26 XThC.Tn[13].t27 161.106
R21935 XThC.Tn[13].n22 XThC.Tn[13].t16 161.106
R21936 XThC.Tn[13].n18 XThC.Tn[13].t37 161.106
R21937 XThC.Tn[13].n14 XThC.Tn[13].t36 161.106
R21938 XThC.Tn[13].n10 XThC.Tn[13].t23 161.106
R21939 XThC.Tn[13].n7 XThC.Tn[13].t13 161.106
R21940 XThC.Tn[13].n66 XThC.Tn[13].t41 154.679
R21941 XThC.Tn[13].n62 XThC.Tn[13].t20 154.679
R21942 XThC.Tn[13].n58 XThC.Tn[13].t18 154.679
R21943 XThC.Tn[13].n54 XThC.Tn[13].t15 154.679
R21944 XThC.Tn[13].n50 XThC.Tn[13].t29 154.679
R21945 XThC.Tn[13].n46 XThC.Tn[13].t26 154.679
R21946 XThC.Tn[13].n42 XThC.Tn[13].t14 154.679
R21947 XThC.Tn[13].n38 XThC.Tn[13].t39 154.679
R21948 XThC.Tn[13].n34 XThC.Tn[13].t35 154.679
R21949 XThC.Tn[13].n30 XThC.Tn[13].t25 154.679
R21950 XThC.Tn[13].n26 XThC.Tn[13].t12 154.679
R21951 XThC.Tn[13].n22 XThC.Tn[13].t34 154.679
R21952 XThC.Tn[13].n18 XThC.Tn[13].t24 154.679
R21953 XThC.Tn[13].n14 XThC.Tn[13].t22 154.679
R21954 XThC.Tn[13].n10 XThC.Tn[13].t42 154.679
R21955 XThC.Tn[13].n7 XThC.Tn[13].t32 154.679
R21956 XThC.Tn[13].n1 XThC.Tn[13].t4 26.5955
R21957 XThC.Tn[13].n1 XThC.Tn[13].t7 26.5955
R21958 XThC.Tn[13].n0 XThC.Tn[13].t6 26.5955
R21959 XThC.Tn[13].n0 XThC.Tn[13].t5 26.5955
R21960 XThC.Tn[13].n3 XThC.Tn[13].t9 26.5955
R21961 XThC.Tn[13].n3 XThC.Tn[13].t8 26.5955
R21962 XThC.Tn[13].n4 XThC.Tn[13].t11 26.5955
R21963 XThC.Tn[13].n4 XThC.Tn[13].t10 26.5955
R21964 XThC.Tn[13].n72 XThC.Tn[13].t0 24.9236
R21965 XThC.Tn[13].n72 XThC.Tn[13].t2 24.9236
R21966 XThC.Tn[13].n73 XThC.Tn[13].t3 24.9236
R21967 XThC.Tn[13].n73 XThC.Tn[13].t1 24.9236
R21968 XThC.Tn[13] XThC.Tn[13].n5 22.9652
R21969 XThC.Tn[13] XThC.Tn[13].n74 18.8943
R21970 XThC.Tn[13].n6 XThC.Tn[13].n2 13.9299
R21971 XThC.Tn[13].n6 XThC.Tn[13] 13.9299
R21972 XThC.Tn[13] XThC.Tn[13].n9 8.0245
R21973 XThC.Tn[13].n69 XThC.Tn[13].n68 7.9105
R21974 XThC.Tn[13].n65 XThC.Tn[13].n64 7.9105
R21975 XThC.Tn[13].n61 XThC.Tn[13].n60 7.9105
R21976 XThC.Tn[13].n57 XThC.Tn[13].n56 7.9105
R21977 XThC.Tn[13].n53 XThC.Tn[13].n52 7.9105
R21978 XThC.Tn[13].n49 XThC.Tn[13].n48 7.9105
R21979 XThC.Tn[13].n45 XThC.Tn[13].n44 7.9105
R21980 XThC.Tn[13].n41 XThC.Tn[13].n40 7.9105
R21981 XThC.Tn[13].n37 XThC.Tn[13].n36 7.9105
R21982 XThC.Tn[13].n33 XThC.Tn[13].n32 7.9105
R21983 XThC.Tn[13].n29 XThC.Tn[13].n28 7.9105
R21984 XThC.Tn[13].n25 XThC.Tn[13].n24 7.9105
R21985 XThC.Tn[13].n21 XThC.Tn[13].n20 7.9105
R21986 XThC.Tn[13].n17 XThC.Tn[13].n16 7.9105
R21987 XThC.Tn[13].n13 XThC.Tn[13].n12 7.9105
R21988 XThC.Tn[13].n71 XThC.Tn[13].n70 7.46054
R21989 XThC.Tn[13] XThC.Tn[13].n71 6.34069
R21990 XThC.Tn[13].n70 XThC.Tn[13] 4.78838
R21991 XThC.Tn[13].n71 XThC.Tn[13] 1.79489
R21992 XThC.Tn[13].n70 XThC.Tn[13] 1.51436
R21993 XThC.Tn[13] XThC.Tn[13].n6 1.19676
R21994 XThC.Tn[13].n13 XThC.Tn[13] 0.235138
R21995 XThC.Tn[13].n17 XThC.Tn[13] 0.235138
R21996 XThC.Tn[13].n21 XThC.Tn[13] 0.235138
R21997 XThC.Tn[13].n25 XThC.Tn[13] 0.235138
R21998 XThC.Tn[13].n29 XThC.Tn[13] 0.235138
R21999 XThC.Tn[13].n33 XThC.Tn[13] 0.235138
R22000 XThC.Tn[13].n37 XThC.Tn[13] 0.235138
R22001 XThC.Tn[13].n41 XThC.Tn[13] 0.235138
R22002 XThC.Tn[13].n45 XThC.Tn[13] 0.235138
R22003 XThC.Tn[13].n49 XThC.Tn[13] 0.235138
R22004 XThC.Tn[13].n53 XThC.Tn[13] 0.235138
R22005 XThC.Tn[13].n57 XThC.Tn[13] 0.235138
R22006 XThC.Tn[13].n61 XThC.Tn[13] 0.235138
R22007 XThC.Tn[13].n65 XThC.Tn[13] 0.235138
R22008 XThC.Tn[13].n69 XThC.Tn[13] 0.235138
R22009 XThC.Tn[13] XThC.Tn[13].n13 0.114505
R22010 XThC.Tn[13] XThC.Tn[13].n17 0.114505
R22011 XThC.Tn[13] XThC.Tn[13].n21 0.114505
R22012 XThC.Tn[13] XThC.Tn[13].n25 0.114505
R22013 XThC.Tn[13] XThC.Tn[13].n29 0.114505
R22014 XThC.Tn[13] XThC.Tn[13].n33 0.114505
R22015 XThC.Tn[13] XThC.Tn[13].n37 0.114505
R22016 XThC.Tn[13] XThC.Tn[13].n41 0.114505
R22017 XThC.Tn[13] XThC.Tn[13].n45 0.114505
R22018 XThC.Tn[13] XThC.Tn[13].n49 0.114505
R22019 XThC.Tn[13] XThC.Tn[13].n53 0.114505
R22020 XThC.Tn[13] XThC.Tn[13].n57 0.114505
R22021 XThC.Tn[13] XThC.Tn[13].n61 0.114505
R22022 XThC.Tn[13] XThC.Tn[13].n65 0.114505
R22023 XThC.Tn[13] XThC.Tn[13].n69 0.114505
R22024 XThC.Tn[13].n68 XThC.Tn[13].n67 0.0599512
R22025 XThC.Tn[13].n64 XThC.Tn[13].n63 0.0599512
R22026 XThC.Tn[13].n60 XThC.Tn[13].n59 0.0599512
R22027 XThC.Tn[13].n56 XThC.Tn[13].n55 0.0599512
R22028 XThC.Tn[13].n52 XThC.Tn[13].n51 0.0599512
R22029 XThC.Tn[13].n48 XThC.Tn[13].n47 0.0599512
R22030 XThC.Tn[13].n44 XThC.Tn[13].n43 0.0599512
R22031 XThC.Tn[13].n40 XThC.Tn[13].n39 0.0599512
R22032 XThC.Tn[13].n36 XThC.Tn[13].n35 0.0599512
R22033 XThC.Tn[13].n32 XThC.Tn[13].n31 0.0599512
R22034 XThC.Tn[13].n28 XThC.Tn[13].n27 0.0599512
R22035 XThC.Tn[13].n24 XThC.Tn[13].n23 0.0599512
R22036 XThC.Tn[13].n20 XThC.Tn[13].n19 0.0599512
R22037 XThC.Tn[13].n16 XThC.Tn[13].n15 0.0599512
R22038 XThC.Tn[13].n12 XThC.Tn[13].n11 0.0599512
R22039 XThC.Tn[13].n9 XThC.Tn[13].n8 0.0599512
R22040 XThC.Tn[13].n67 XThC.Tn[13] 0.0469286
R22041 XThC.Tn[13].n63 XThC.Tn[13] 0.0469286
R22042 XThC.Tn[13].n59 XThC.Tn[13] 0.0469286
R22043 XThC.Tn[13].n55 XThC.Tn[13] 0.0469286
R22044 XThC.Tn[13].n51 XThC.Tn[13] 0.0469286
R22045 XThC.Tn[13].n47 XThC.Tn[13] 0.0469286
R22046 XThC.Tn[13].n43 XThC.Tn[13] 0.0469286
R22047 XThC.Tn[13].n39 XThC.Tn[13] 0.0469286
R22048 XThC.Tn[13].n35 XThC.Tn[13] 0.0469286
R22049 XThC.Tn[13].n31 XThC.Tn[13] 0.0469286
R22050 XThC.Tn[13].n27 XThC.Tn[13] 0.0469286
R22051 XThC.Tn[13].n23 XThC.Tn[13] 0.0469286
R22052 XThC.Tn[13].n19 XThC.Tn[13] 0.0469286
R22053 XThC.Tn[13].n15 XThC.Tn[13] 0.0469286
R22054 XThC.Tn[13].n11 XThC.Tn[13] 0.0469286
R22055 XThC.Tn[13].n8 XThC.Tn[13] 0.0469286
R22056 XThC.Tn[13].n67 XThC.Tn[13] 0.0401341
R22057 XThC.Tn[13].n63 XThC.Tn[13] 0.0401341
R22058 XThC.Tn[13].n59 XThC.Tn[13] 0.0401341
R22059 XThC.Tn[13].n55 XThC.Tn[13] 0.0401341
R22060 XThC.Tn[13].n51 XThC.Tn[13] 0.0401341
R22061 XThC.Tn[13].n47 XThC.Tn[13] 0.0401341
R22062 XThC.Tn[13].n43 XThC.Tn[13] 0.0401341
R22063 XThC.Tn[13].n39 XThC.Tn[13] 0.0401341
R22064 XThC.Tn[13].n35 XThC.Tn[13] 0.0401341
R22065 XThC.Tn[13].n31 XThC.Tn[13] 0.0401341
R22066 XThC.Tn[13].n27 XThC.Tn[13] 0.0401341
R22067 XThC.Tn[13].n23 XThC.Tn[13] 0.0401341
R22068 XThC.Tn[13].n19 XThC.Tn[13] 0.0401341
R22069 XThC.Tn[13].n15 XThC.Tn[13] 0.0401341
R22070 XThC.Tn[13].n11 XThC.Tn[13] 0.0401341
R22071 XThC.Tn[13].n8 XThC.Tn[13] 0.0401341
R22072 XThC.Tn[7].n5 XThC.Tn[7].n4 255.096
R22073 XThC.Tn[7].n2 XThC.Tn[7].n0 236.589
R22074 XThC.Tn[7].n5 XThC.Tn[7].n3 201.845
R22075 XThC.Tn[7].n2 XThC.Tn[7].n1 200.321
R22076 XThC.Tn[7].n67 XThC.Tn[7].n65 161.365
R22077 XThC.Tn[7].n63 XThC.Tn[7].n61 161.365
R22078 XThC.Tn[7].n59 XThC.Tn[7].n57 161.365
R22079 XThC.Tn[7].n55 XThC.Tn[7].n53 161.365
R22080 XThC.Tn[7].n51 XThC.Tn[7].n49 161.365
R22081 XThC.Tn[7].n47 XThC.Tn[7].n45 161.365
R22082 XThC.Tn[7].n43 XThC.Tn[7].n41 161.365
R22083 XThC.Tn[7].n39 XThC.Tn[7].n37 161.365
R22084 XThC.Tn[7].n35 XThC.Tn[7].n33 161.365
R22085 XThC.Tn[7].n31 XThC.Tn[7].n29 161.365
R22086 XThC.Tn[7].n27 XThC.Tn[7].n25 161.365
R22087 XThC.Tn[7].n23 XThC.Tn[7].n21 161.365
R22088 XThC.Tn[7].n19 XThC.Tn[7].n17 161.365
R22089 XThC.Tn[7].n15 XThC.Tn[7].n13 161.365
R22090 XThC.Tn[7].n11 XThC.Tn[7].n9 161.365
R22091 XThC.Tn[7].n8 XThC.Tn[7].n6 161.365
R22092 XThC.Tn[7].n65 XThC.Tn[7].t8 161.106
R22093 XThC.Tn[7].n61 XThC.Tn[7].t20 161.106
R22094 XThC.Tn[7].n57 XThC.Tn[7].t18 161.106
R22095 XThC.Tn[7].n53 XThC.Tn[7].t16 161.106
R22096 XThC.Tn[7].n49 XThC.Tn[7].t30 161.106
R22097 XThC.Tn[7].n45 XThC.Tn[7].t27 161.106
R22098 XThC.Tn[7].n41 XThC.Tn[7].t15 161.106
R22099 XThC.Tn[7].n37 XThC.Tn[7].t38 161.106
R22100 XThC.Tn[7].n33 XThC.Tn[7].t36 161.106
R22101 XThC.Tn[7].n29 XThC.Tn[7].t25 161.106
R22102 XThC.Tn[7].n25 XThC.Tn[7].t14 161.106
R22103 XThC.Tn[7].n21 XThC.Tn[7].t35 161.106
R22104 XThC.Tn[7].n17 XThC.Tn[7].t24 161.106
R22105 XThC.Tn[7].n13 XThC.Tn[7].t23 161.106
R22106 XThC.Tn[7].n9 XThC.Tn[7].t10 161.106
R22107 XThC.Tn[7].n6 XThC.Tn[7].t32 161.106
R22108 XThC.Tn[7].n65 XThC.Tn[7].t28 154.679
R22109 XThC.Tn[7].n61 XThC.Tn[7].t39 154.679
R22110 XThC.Tn[7].n57 XThC.Tn[7].t37 154.679
R22111 XThC.Tn[7].n53 XThC.Tn[7].t34 154.679
R22112 XThC.Tn[7].n49 XThC.Tn[7].t17 154.679
R22113 XThC.Tn[7].n45 XThC.Tn[7].t13 154.679
R22114 XThC.Tn[7].n41 XThC.Tn[7].t33 154.679
R22115 XThC.Tn[7].n37 XThC.Tn[7].t26 154.679
R22116 XThC.Tn[7].n33 XThC.Tn[7].t22 154.679
R22117 XThC.Tn[7].n29 XThC.Tn[7].t12 154.679
R22118 XThC.Tn[7].n25 XThC.Tn[7].t31 154.679
R22119 XThC.Tn[7].n21 XThC.Tn[7].t21 154.679
R22120 XThC.Tn[7].n17 XThC.Tn[7].t11 154.679
R22121 XThC.Tn[7].n13 XThC.Tn[7].t9 154.679
R22122 XThC.Tn[7].n9 XThC.Tn[7].t29 154.679
R22123 XThC.Tn[7].n6 XThC.Tn[7].t19 154.679
R22124 XThC.Tn[7].n4 XThC.Tn[7].t2 26.5955
R22125 XThC.Tn[7].n4 XThC.Tn[7].t1 26.5955
R22126 XThC.Tn[7].n3 XThC.Tn[7].t0 26.5955
R22127 XThC.Tn[7].n3 XThC.Tn[7].t3 26.5955
R22128 XThC.Tn[7] XThC.Tn[7].n5 26.4992
R22129 XThC.Tn[7].n0 XThC.Tn[7].t6 24.9236
R22130 XThC.Tn[7].n0 XThC.Tn[7].t5 24.9236
R22131 XThC.Tn[7].n1 XThC.Tn[7].t4 24.9236
R22132 XThC.Tn[7].n1 XThC.Tn[7].t7 24.9236
R22133 XThC.Tn[7].n70 XThC.Tn[7].n2 12.0894
R22134 XThC.Tn[7].n70 XThC.Tn[7] 9.64206
R22135 XThC.Tn[7].n69 XThC.Tn[7] 8.14595
R22136 XThC.Tn[7] XThC.Tn[7].n8 8.0245
R22137 XThC.Tn[7].n68 XThC.Tn[7].n67 7.9105
R22138 XThC.Tn[7].n64 XThC.Tn[7].n63 7.9105
R22139 XThC.Tn[7].n60 XThC.Tn[7].n59 7.9105
R22140 XThC.Tn[7].n56 XThC.Tn[7].n55 7.9105
R22141 XThC.Tn[7].n52 XThC.Tn[7].n51 7.9105
R22142 XThC.Tn[7].n48 XThC.Tn[7].n47 7.9105
R22143 XThC.Tn[7].n44 XThC.Tn[7].n43 7.9105
R22144 XThC.Tn[7].n40 XThC.Tn[7].n39 7.9105
R22145 XThC.Tn[7].n36 XThC.Tn[7].n35 7.9105
R22146 XThC.Tn[7].n32 XThC.Tn[7].n31 7.9105
R22147 XThC.Tn[7].n28 XThC.Tn[7].n27 7.9105
R22148 XThC.Tn[7].n24 XThC.Tn[7].n23 7.9105
R22149 XThC.Tn[7].n20 XThC.Tn[7].n19 7.9105
R22150 XThC.Tn[7].n16 XThC.Tn[7].n15 7.9105
R22151 XThC.Tn[7].n12 XThC.Tn[7].n11 7.9105
R22152 XThC.Tn[7].n69 XThC.Tn[7] 5.30358
R22153 XThC.Tn[7] XThC.Tn[7].n69 3.15894
R22154 XThC.Tn[7] XThC.Tn[7].n70 1.66284
R22155 XThC.Tn[7].n12 XThC.Tn[7] 0.235138
R22156 XThC.Tn[7].n16 XThC.Tn[7] 0.235138
R22157 XThC.Tn[7].n20 XThC.Tn[7] 0.235138
R22158 XThC.Tn[7].n24 XThC.Tn[7] 0.235138
R22159 XThC.Tn[7].n28 XThC.Tn[7] 0.235138
R22160 XThC.Tn[7].n32 XThC.Tn[7] 0.235138
R22161 XThC.Tn[7].n36 XThC.Tn[7] 0.235138
R22162 XThC.Tn[7].n40 XThC.Tn[7] 0.235138
R22163 XThC.Tn[7].n44 XThC.Tn[7] 0.235138
R22164 XThC.Tn[7].n48 XThC.Tn[7] 0.235138
R22165 XThC.Tn[7].n52 XThC.Tn[7] 0.235138
R22166 XThC.Tn[7].n56 XThC.Tn[7] 0.235138
R22167 XThC.Tn[7].n60 XThC.Tn[7] 0.235138
R22168 XThC.Tn[7].n64 XThC.Tn[7] 0.235138
R22169 XThC.Tn[7].n68 XThC.Tn[7] 0.235138
R22170 XThC.Tn[7] XThC.Tn[7].n12 0.114505
R22171 XThC.Tn[7] XThC.Tn[7].n16 0.114505
R22172 XThC.Tn[7] XThC.Tn[7].n20 0.114505
R22173 XThC.Tn[7] XThC.Tn[7].n24 0.114505
R22174 XThC.Tn[7] XThC.Tn[7].n28 0.114505
R22175 XThC.Tn[7] XThC.Tn[7].n32 0.114505
R22176 XThC.Tn[7] XThC.Tn[7].n36 0.114505
R22177 XThC.Tn[7] XThC.Tn[7].n40 0.114505
R22178 XThC.Tn[7] XThC.Tn[7].n44 0.114505
R22179 XThC.Tn[7] XThC.Tn[7].n48 0.114505
R22180 XThC.Tn[7] XThC.Tn[7].n52 0.114505
R22181 XThC.Tn[7] XThC.Tn[7].n56 0.114505
R22182 XThC.Tn[7] XThC.Tn[7].n60 0.114505
R22183 XThC.Tn[7] XThC.Tn[7].n64 0.114505
R22184 XThC.Tn[7] XThC.Tn[7].n68 0.114505
R22185 XThC.Tn[7].n67 XThC.Tn[7].n66 0.0599512
R22186 XThC.Tn[7].n63 XThC.Tn[7].n62 0.0599512
R22187 XThC.Tn[7].n59 XThC.Tn[7].n58 0.0599512
R22188 XThC.Tn[7].n55 XThC.Tn[7].n54 0.0599512
R22189 XThC.Tn[7].n51 XThC.Tn[7].n50 0.0599512
R22190 XThC.Tn[7].n47 XThC.Tn[7].n46 0.0599512
R22191 XThC.Tn[7].n43 XThC.Tn[7].n42 0.0599512
R22192 XThC.Tn[7].n39 XThC.Tn[7].n38 0.0599512
R22193 XThC.Tn[7].n35 XThC.Tn[7].n34 0.0599512
R22194 XThC.Tn[7].n31 XThC.Tn[7].n30 0.0599512
R22195 XThC.Tn[7].n27 XThC.Tn[7].n26 0.0599512
R22196 XThC.Tn[7].n23 XThC.Tn[7].n22 0.0599512
R22197 XThC.Tn[7].n19 XThC.Tn[7].n18 0.0599512
R22198 XThC.Tn[7].n15 XThC.Tn[7].n14 0.0599512
R22199 XThC.Tn[7].n11 XThC.Tn[7].n10 0.0599512
R22200 XThC.Tn[7].n8 XThC.Tn[7].n7 0.0599512
R22201 XThC.Tn[7].n66 XThC.Tn[7] 0.0469286
R22202 XThC.Tn[7].n62 XThC.Tn[7] 0.0469286
R22203 XThC.Tn[7].n58 XThC.Tn[7] 0.0469286
R22204 XThC.Tn[7].n54 XThC.Tn[7] 0.0469286
R22205 XThC.Tn[7].n50 XThC.Tn[7] 0.0469286
R22206 XThC.Tn[7].n46 XThC.Tn[7] 0.0469286
R22207 XThC.Tn[7].n42 XThC.Tn[7] 0.0469286
R22208 XThC.Tn[7].n38 XThC.Tn[7] 0.0469286
R22209 XThC.Tn[7].n34 XThC.Tn[7] 0.0469286
R22210 XThC.Tn[7].n30 XThC.Tn[7] 0.0469286
R22211 XThC.Tn[7].n26 XThC.Tn[7] 0.0469286
R22212 XThC.Tn[7].n22 XThC.Tn[7] 0.0469286
R22213 XThC.Tn[7].n18 XThC.Tn[7] 0.0469286
R22214 XThC.Tn[7].n14 XThC.Tn[7] 0.0469286
R22215 XThC.Tn[7].n10 XThC.Tn[7] 0.0469286
R22216 XThC.Tn[7].n7 XThC.Tn[7] 0.0469286
R22217 XThC.Tn[7].n66 XThC.Tn[7] 0.0401341
R22218 XThC.Tn[7].n62 XThC.Tn[7] 0.0401341
R22219 XThC.Tn[7].n58 XThC.Tn[7] 0.0401341
R22220 XThC.Tn[7].n54 XThC.Tn[7] 0.0401341
R22221 XThC.Tn[7].n50 XThC.Tn[7] 0.0401341
R22222 XThC.Tn[7].n46 XThC.Tn[7] 0.0401341
R22223 XThC.Tn[7].n42 XThC.Tn[7] 0.0401341
R22224 XThC.Tn[7].n38 XThC.Tn[7] 0.0401341
R22225 XThC.Tn[7].n34 XThC.Tn[7] 0.0401341
R22226 XThC.Tn[7].n30 XThC.Tn[7] 0.0401341
R22227 XThC.Tn[7].n26 XThC.Tn[7] 0.0401341
R22228 XThC.Tn[7].n22 XThC.Tn[7] 0.0401341
R22229 XThC.Tn[7].n18 XThC.Tn[7] 0.0401341
R22230 XThC.Tn[7].n14 XThC.Tn[7] 0.0401341
R22231 XThC.Tn[7].n10 XThC.Tn[7] 0.0401341
R22232 XThC.Tn[7].n7 XThC.Tn[7] 0.0401341
R22233 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R22234 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R22235 XThR.Tn[6] XThR.Tn[6].n82 161.363
R22236 XThR.Tn[6] XThR.Tn[6].n77 161.363
R22237 XThR.Tn[6] XThR.Tn[6].n72 161.363
R22238 XThR.Tn[6] XThR.Tn[6].n67 161.363
R22239 XThR.Tn[6] XThR.Tn[6].n62 161.363
R22240 XThR.Tn[6] XThR.Tn[6].n57 161.363
R22241 XThR.Tn[6] XThR.Tn[6].n52 161.363
R22242 XThR.Tn[6] XThR.Tn[6].n47 161.363
R22243 XThR.Tn[6] XThR.Tn[6].n42 161.363
R22244 XThR.Tn[6] XThR.Tn[6].n37 161.363
R22245 XThR.Tn[6] XThR.Tn[6].n32 161.363
R22246 XThR.Tn[6] XThR.Tn[6].n27 161.363
R22247 XThR.Tn[6] XThR.Tn[6].n22 161.363
R22248 XThR.Tn[6] XThR.Tn[6].n17 161.363
R22249 XThR.Tn[6] XThR.Tn[6].n12 161.363
R22250 XThR.Tn[6] XThR.Tn[6].n10 161.363
R22251 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R22252 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R22253 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R22254 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R22255 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R22256 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R22257 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R22258 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R22259 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R22260 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R22261 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R22262 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R22263 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R22264 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R22265 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R22266 XThR.Tn[6].n83 XThR.Tn[6].t21 161.106
R22267 XThR.Tn[6].n82 XThR.Tn[6].t37 161.106
R22268 XThR.Tn[6].n78 XThR.Tn[6].t28 161.106
R22269 XThR.Tn[6].n77 XThR.Tn[6].t47 161.106
R22270 XThR.Tn[6].n73 XThR.Tn[6].t71 161.106
R22271 XThR.Tn[6].n72 XThR.Tn[6].t29 161.106
R22272 XThR.Tn[6].n68 XThR.Tn[6].t53 161.106
R22273 XThR.Tn[6].n67 XThR.Tn[6].t72 161.106
R22274 XThR.Tn[6].n63 XThR.Tn[6].t19 161.106
R22275 XThR.Tn[6].n62 XThR.Tn[6].t35 161.106
R22276 XThR.Tn[6].n58 XThR.Tn[6].t44 161.106
R22277 XThR.Tn[6].n57 XThR.Tn[6].t63 161.106
R22278 XThR.Tn[6].n53 XThR.Tn[6].t23 161.106
R22279 XThR.Tn[6].n52 XThR.Tn[6].t43 161.106
R22280 XThR.Tn[6].n48 XThR.Tn[6].t67 161.106
R22281 XThR.Tn[6].n47 XThR.Tn[6].t24 161.106
R22282 XThR.Tn[6].n43 XThR.Tn[6].t52 161.106
R22283 XThR.Tn[6].n42 XThR.Tn[6].t68 161.106
R22284 XThR.Tn[6].n38 XThR.Tn[6].t58 161.106
R22285 XThR.Tn[6].n37 XThR.Tn[6].t13 161.106
R22286 XThR.Tn[6].n33 XThR.Tn[6].t42 161.106
R22287 XThR.Tn[6].n32 XThR.Tn[6].t60 161.106
R22288 XThR.Tn[6].n28 XThR.Tn[6].t70 161.106
R22289 XThR.Tn[6].n27 XThR.Tn[6].t27 161.106
R22290 XThR.Tn[6].n23 XThR.Tn[6].t39 161.106
R22291 XThR.Tn[6].n22 XThR.Tn[6].t56 161.106
R22292 XThR.Tn[6].n18 XThR.Tn[6].t22 161.106
R22293 XThR.Tn[6].n17 XThR.Tn[6].t40 161.106
R22294 XThR.Tn[6].n13 XThR.Tn[6].t49 161.106
R22295 XThR.Tn[6].n12 XThR.Tn[6].t66 161.106
R22296 XThR.Tn[6].n10 XThR.Tn[6].t50 161.106
R22297 XThR.Tn[6].n83 XThR.Tn[6].t38 154.679
R22298 XThR.Tn[6].n82 XThR.Tn[6].t55 154.679
R22299 XThR.Tn[6].n78 XThR.Tn[6].t16 154.679
R22300 XThR.Tn[6].n77 XThR.Tn[6].t34 154.679
R22301 XThR.Tn[6].n73 XThR.Tn[6].t62 154.679
R22302 XThR.Tn[6].n72 XThR.Tn[6].t17 154.679
R22303 XThR.Tn[6].n68 XThR.Tn[6].t30 154.679
R22304 XThR.Tn[6].n67 XThR.Tn[6].t48 154.679
R22305 XThR.Tn[6].n63 XThR.Tn[6].t73 154.679
R22306 XThR.Tn[6].n62 XThR.Tn[6].t31 154.679
R22307 XThR.Tn[6].n58 XThR.Tn[6].t36 154.679
R22308 XThR.Tn[6].n57 XThR.Tn[6].t54 154.679
R22309 XThR.Tn[6].n53 XThR.Tn[6].t64 154.679
R22310 XThR.Tn[6].n52 XThR.Tn[6].t18 154.679
R22311 XThR.Tn[6].n48 XThR.Tn[6].t46 154.679
R22312 XThR.Tn[6].n47 XThR.Tn[6].t65 154.679
R22313 XThR.Tn[6].n43 XThR.Tn[6].t25 154.679
R22314 XThR.Tn[6].n42 XThR.Tn[6].t45 154.679
R22315 XThR.Tn[6].n38 XThR.Tn[6].t69 154.679
R22316 XThR.Tn[6].n37 XThR.Tn[6].t26 154.679
R22317 XThR.Tn[6].n33 XThR.Tn[6].t14 154.679
R22318 XThR.Tn[6].n32 XThR.Tn[6].t33 154.679
R22319 XThR.Tn[6].n28 XThR.Tn[6].t61 154.679
R22320 XThR.Tn[6].n27 XThR.Tn[6].t15 154.679
R22321 XThR.Tn[6].n23 XThR.Tn[6].t32 154.679
R22322 XThR.Tn[6].n22 XThR.Tn[6].t51 154.679
R22323 XThR.Tn[6].n18 XThR.Tn[6].t57 154.679
R22324 XThR.Tn[6].n17 XThR.Tn[6].t12 154.679
R22325 XThR.Tn[6].n13 XThR.Tn[6].t41 154.679
R22326 XThR.Tn[6].n12 XThR.Tn[6].t59 154.679
R22327 XThR.Tn[6].n10 XThR.Tn[6].t20 154.679
R22328 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R22329 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R22330 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R22331 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R22332 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R22333 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R22334 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R22335 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R22336 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R22337 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R22338 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R22339 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R22340 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R22341 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R22342 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R22343 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R22344 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R22345 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R22346 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R22347 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R22348 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R22349 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R22350 XThR.Tn[6] XThR.Tn[6].n11 5.34871
R22351 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R22352 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R22353 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R22354 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R22355 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R22356 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R22357 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R22358 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R22359 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R22360 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R22361 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R22362 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R22363 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R22364 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R22365 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R22366 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R22367 XThR.Tn[6].n16 XThR.Tn[6] 2.51836
R22368 XThR.Tn[6].n21 XThR.Tn[6] 2.51836
R22369 XThR.Tn[6].n26 XThR.Tn[6] 2.51836
R22370 XThR.Tn[6].n31 XThR.Tn[6] 2.51836
R22371 XThR.Tn[6].n36 XThR.Tn[6] 2.51836
R22372 XThR.Tn[6].n41 XThR.Tn[6] 2.51836
R22373 XThR.Tn[6].n46 XThR.Tn[6] 2.51836
R22374 XThR.Tn[6].n51 XThR.Tn[6] 2.51836
R22375 XThR.Tn[6].n56 XThR.Tn[6] 2.51836
R22376 XThR.Tn[6].n61 XThR.Tn[6] 2.51836
R22377 XThR.Tn[6].n66 XThR.Tn[6] 2.51836
R22378 XThR.Tn[6].n71 XThR.Tn[6] 2.51836
R22379 XThR.Tn[6].n76 XThR.Tn[6] 2.51836
R22380 XThR.Tn[6].n81 XThR.Tn[6] 2.51836
R22381 XThR.Tn[6].n86 XThR.Tn[6] 2.51836
R22382 XThR.Tn[6] XThR.Tn[6].n16 0.848714
R22383 XThR.Tn[6] XThR.Tn[6].n21 0.848714
R22384 XThR.Tn[6] XThR.Tn[6].n26 0.848714
R22385 XThR.Tn[6] XThR.Tn[6].n31 0.848714
R22386 XThR.Tn[6] XThR.Tn[6].n36 0.848714
R22387 XThR.Tn[6] XThR.Tn[6].n41 0.848714
R22388 XThR.Tn[6] XThR.Tn[6].n46 0.848714
R22389 XThR.Tn[6] XThR.Tn[6].n51 0.848714
R22390 XThR.Tn[6] XThR.Tn[6].n56 0.848714
R22391 XThR.Tn[6] XThR.Tn[6].n61 0.848714
R22392 XThR.Tn[6] XThR.Tn[6].n66 0.848714
R22393 XThR.Tn[6] XThR.Tn[6].n71 0.848714
R22394 XThR.Tn[6] XThR.Tn[6].n76 0.848714
R22395 XThR.Tn[6] XThR.Tn[6].n81 0.848714
R22396 XThR.Tn[6] XThR.Tn[6].n86 0.848714
R22397 XThR.Tn[6].n11 XThR.Tn[6] 0.485653
R22398 XThR.Tn[6].n84 XThR.Tn[6] 0.21482
R22399 XThR.Tn[6].n79 XThR.Tn[6] 0.21482
R22400 XThR.Tn[6].n74 XThR.Tn[6] 0.21482
R22401 XThR.Tn[6].n69 XThR.Tn[6] 0.21482
R22402 XThR.Tn[6].n64 XThR.Tn[6] 0.21482
R22403 XThR.Tn[6].n59 XThR.Tn[6] 0.21482
R22404 XThR.Tn[6].n54 XThR.Tn[6] 0.21482
R22405 XThR.Tn[6].n49 XThR.Tn[6] 0.21482
R22406 XThR.Tn[6].n44 XThR.Tn[6] 0.21482
R22407 XThR.Tn[6].n39 XThR.Tn[6] 0.21482
R22408 XThR.Tn[6].n34 XThR.Tn[6] 0.21482
R22409 XThR.Tn[6].n29 XThR.Tn[6] 0.21482
R22410 XThR.Tn[6].n24 XThR.Tn[6] 0.21482
R22411 XThR.Tn[6].n19 XThR.Tn[6] 0.21482
R22412 XThR.Tn[6].n14 XThR.Tn[6] 0.21482
R22413 XThR.Tn[6].n85 XThR.Tn[6] 0.0608448
R22414 XThR.Tn[6].n80 XThR.Tn[6] 0.0608448
R22415 XThR.Tn[6].n75 XThR.Tn[6] 0.0608448
R22416 XThR.Tn[6].n70 XThR.Tn[6] 0.0608448
R22417 XThR.Tn[6].n65 XThR.Tn[6] 0.0608448
R22418 XThR.Tn[6].n60 XThR.Tn[6] 0.0608448
R22419 XThR.Tn[6].n55 XThR.Tn[6] 0.0608448
R22420 XThR.Tn[6].n50 XThR.Tn[6] 0.0608448
R22421 XThR.Tn[6].n45 XThR.Tn[6] 0.0608448
R22422 XThR.Tn[6].n40 XThR.Tn[6] 0.0608448
R22423 XThR.Tn[6].n35 XThR.Tn[6] 0.0608448
R22424 XThR.Tn[6].n30 XThR.Tn[6] 0.0608448
R22425 XThR.Tn[6].n25 XThR.Tn[6] 0.0608448
R22426 XThR.Tn[6].n20 XThR.Tn[6] 0.0608448
R22427 XThR.Tn[6].n15 XThR.Tn[6] 0.0608448
R22428 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R22429 XThR.Tn[6] XThR.Tn[6].n87 0.038
R22430 XThR.Tn[6].n11 XThR.Tn[6] 0.00744444
R22431 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00265517
R22432 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00265517
R22433 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00265517
R22434 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00265517
R22435 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00265517
R22436 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00265517
R22437 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00265517
R22438 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00265517
R22439 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00265517
R22440 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00265517
R22441 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00265517
R22442 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00265517
R22443 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00265517
R22444 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00265517
R22445 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00265517
R22446 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R22447 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R22448 XThR.Tn[11].n2 XThR.Tn[11].n0 241.847
R22449 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R22450 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R22451 XThR.Tn[11].n2 XThR.Tn[11].n1 185
R22452 XThR.Tn[11] XThR.Tn[11].n82 161.363
R22453 XThR.Tn[11] XThR.Tn[11].n77 161.363
R22454 XThR.Tn[11] XThR.Tn[11].n72 161.363
R22455 XThR.Tn[11] XThR.Tn[11].n67 161.363
R22456 XThR.Tn[11] XThR.Tn[11].n62 161.363
R22457 XThR.Tn[11] XThR.Tn[11].n57 161.363
R22458 XThR.Tn[11] XThR.Tn[11].n52 161.363
R22459 XThR.Tn[11] XThR.Tn[11].n47 161.363
R22460 XThR.Tn[11] XThR.Tn[11].n42 161.363
R22461 XThR.Tn[11] XThR.Tn[11].n37 161.363
R22462 XThR.Tn[11] XThR.Tn[11].n32 161.363
R22463 XThR.Tn[11] XThR.Tn[11].n27 161.363
R22464 XThR.Tn[11] XThR.Tn[11].n22 161.363
R22465 XThR.Tn[11] XThR.Tn[11].n17 161.363
R22466 XThR.Tn[11] XThR.Tn[11].n12 161.363
R22467 XThR.Tn[11] XThR.Tn[11].n10 161.363
R22468 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R22469 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R22470 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R22471 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R22472 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R22473 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R22474 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R22475 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R22476 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R22477 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R22478 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R22479 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R22480 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R22481 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R22482 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R22483 XThR.Tn[11].n83 XThR.Tn[11].t71 161.106
R22484 XThR.Tn[11].n82 XThR.Tn[11].t17 161.106
R22485 XThR.Tn[11].n78 XThR.Tn[11].t16 161.106
R22486 XThR.Tn[11].n77 XThR.Tn[11].t23 161.106
R22487 XThR.Tn[11].n73 XThR.Tn[11].t61 161.106
R22488 XThR.Tn[11].n72 XThR.Tn[11].t66 161.106
R22489 XThR.Tn[11].n68 XThR.Tn[11].t44 161.106
R22490 XThR.Tn[11].n67 XThR.Tn[11].t46 161.106
R22491 XThR.Tn[11].n63 XThR.Tn[11].t70 161.106
R22492 XThR.Tn[11].n62 XThR.Tn[11].t14 161.106
R22493 XThR.Tn[11].n58 XThR.Tn[11].t32 161.106
R22494 XThR.Tn[11].n57 XThR.Tn[11].t40 161.106
R22495 XThR.Tn[11].n53 XThR.Tn[11].t13 161.106
R22496 XThR.Tn[11].n52 XThR.Tn[11].t21 161.106
R22497 XThR.Tn[11].n48 XThR.Tn[11].t57 161.106
R22498 XThR.Tn[11].n47 XThR.Tn[11].t63 161.106
R22499 XThR.Tn[11].n43 XThR.Tn[11].t42 161.106
R22500 XThR.Tn[11].n42 XThR.Tn[11].t45 161.106
R22501 XThR.Tn[11].n38 XThR.Tn[11].t48 161.106
R22502 XThR.Tn[11].n37 XThR.Tn[11].t53 161.106
R22503 XThR.Tn[11].n33 XThR.Tn[11].t31 161.106
R22504 XThR.Tn[11].n32 XThR.Tn[11].t39 161.106
R22505 XThR.Tn[11].n28 XThR.Tn[11].t59 161.106
R22506 XThR.Tn[11].n27 XThR.Tn[11].t65 161.106
R22507 XThR.Tn[11].n23 XThR.Tn[11].t29 161.106
R22508 XThR.Tn[11].n22 XThR.Tn[11].t37 161.106
R22509 XThR.Tn[11].n18 XThR.Tn[11].t12 161.106
R22510 XThR.Tn[11].n17 XThR.Tn[11].t19 161.106
R22511 XThR.Tn[11].n13 XThR.Tn[11].t36 161.106
R22512 XThR.Tn[11].n12 XThR.Tn[11].t43 161.106
R22513 XThR.Tn[11].n10 XThR.Tn[11].t25 161.106
R22514 XThR.Tn[11].n83 XThR.Tn[11].t28 154.679
R22515 XThR.Tn[11].n82 XThR.Tn[11].t35 154.679
R22516 XThR.Tn[11].n78 XThR.Tn[11].t69 154.679
R22517 XThR.Tn[11].n77 XThR.Tn[11].t73 154.679
R22518 XThR.Tn[11].n73 XThR.Tn[11].t50 154.679
R22519 XThR.Tn[11].n72 XThR.Tn[11].t55 154.679
R22520 XThR.Tn[11].n68 XThR.Tn[11].t18 154.679
R22521 XThR.Tn[11].n67 XThR.Tn[11].t24 154.679
R22522 XThR.Tn[11].n63 XThR.Tn[11].t62 154.679
R22523 XThR.Tn[11].n62 XThR.Tn[11].t67 154.679
R22524 XThR.Tn[11].n58 XThR.Tn[11].t27 154.679
R22525 XThR.Tn[11].n57 XThR.Tn[11].t34 154.679
R22526 XThR.Tn[11].n53 XThR.Tn[11].t51 154.679
R22527 XThR.Tn[11].n52 XThR.Tn[11].t56 154.679
R22528 XThR.Tn[11].n48 XThR.Tn[11].t33 154.679
R22529 XThR.Tn[11].n47 XThR.Tn[11].t41 154.679
R22530 XThR.Tn[11].n43 XThR.Tn[11].t15 154.679
R22531 XThR.Tn[11].n42 XThR.Tn[11].t22 154.679
R22532 XThR.Tn[11].n38 XThR.Tn[11].t58 154.679
R22533 XThR.Tn[11].n37 XThR.Tn[11].t64 154.679
R22534 XThR.Tn[11].n33 XThR.Tn[11].t68 154.679
R22535 XThR.Tn[11].n32 XThR.Tn[11].t72 154.679
R22536 XThR.Tn[11].n28 XThR.Tn[11].t49 154.679
R22537 XThR.Tn[11].n27 XThR.Tn[11].t54 154.679
R22538 XThR.Tn[11].n23 XThR.Tn[11].t20 154.679
R22539 XThR.Tn[11].n22 XThR.Tn[11].t26 154.679
R22540 XThR.Tn[11].n18 XThR.Tn[11].t47 154.679
R22541 XThR.Tn[11].n17 XThR.Tn[11].t52 154.679
R22542 XThR.Tn[11].n13 XThR.Tn[11].t30 154.679
R22543 XThR.Tn[11].n12 XThR.Tn[11].t38 154.679
R22544 XThR.Tn[11].n10 XThR.Tn[11].t60 154.679
R22545 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R22546 XThR.Tn[11].n6 XThR.Tn[11].t4 26.5955
R22547 XThR.Tn[11].n6 XThR.Tn[11].t6 26.5955
R22548 XThR.Tn[11].n7 XThR.Tn[11].t2 26.5955
R22549 XThR.Tn[11].n7 XThR.Tn[11].t5 26.5955
R22550 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R22551 XThR.Tn[11].n3 XThR.Tn[11].t10 26.5955
R22552 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R22553 XThR.Tn[11].n4 XThR.Tn[11].t11 26.5955
R22554 XThR.Tn[11].n0 XThR.Tn[11].t7 24.9236
R22555 XThR.Tn[11].n0 XThR.Tn[11].t1 24.9236
R22556 XThR.Tn[11].n1 XThR.Tn[11].t0 24.9236
R22557 XThR.Tn[11].n1 XThR.Tn[11].t3 24.9236
R22558 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R22559 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R22560 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R22561 XThR.Tn[11] XThR.Tn[11].n11 5.34871
R22562 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R22563 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R22564 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R22565 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R22566 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R22567 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R22568 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R22569 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R22570 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R22571 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R22572 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R22573 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R22574 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R22575 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R22576 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R22577 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R22578 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R22579 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R22580 XThR.Tn[11].n16 XThR.Tn[11] 2.51836
R22581 XThR.Tn[11].n21 XThR.Tn[11] 2.51836
R22582 XThR.Tn[11].n26 XThR.Tn[11] 2.51836
R22583 XThR.Tn[11].n31 XThR.Tn[11] 2.51836
R22584 XThR.Tn[11].n36 XThR.Tn[11] 2.51836
R22585 XThR.Tn[11].n41 XThR.Tn[11] 2.51836
R22586 XThR.Tn[11].n46 XThR.Tn[11] 2.51836
R22587 XThR.Tn[11].n51 XThR.Tn[11] 2.51836
R22588 XThR.Tn[11].n56 XThR.Tn[11] 2.51836
R22589 XThR.Tn[11].n61 XThR.Tn[11] 2.51836
R22590 XThR.Tn[11].n66 XThR.Tn[11] 2.51836
R22591 XThR.Tn[11].n71 XThR.Tn[11] 2.51836
R22592 XThR.Tn[11].n76 XThR.Tn[11] 2.51836
R22593 XThR.Tn[11].n81 XThR.Tn[11] 2.51836
R22594 XThR.Tn[11].n86 XThR.Tn[11] 2.51836
R22595 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R22596 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R22597 XThR.Tn[11] XThR.Tn[11].n16 0.848714
R22598 XThR.Tn[11] XThR.Tn[11].n21 0.848714
R22599 XThR.Tn[11] XThR.Tn[11].n26 0.848714
R22600 XThR.Tn[11] XThR.Tn[11].n31 0.848714
R22601 XThR.Tn[11] XThR.Tn[11].n36 0.848714
R22602 XThR.Tn[11] XThR.Tn[11].n41 0.848714
R22603 XThR.Tn[11] XThR.Tn[11].n46 0.848714
R22604 XThR.Tn[11] XThR.Tn[11].n51 0.848714
R22605 XThR.Tn[11] XThR.Tn[11].n56 0.848714
R22606 XThR.Tn[11] XThR.Tn[11].n61 0.848714
R22607 XThR.Tn[11] XThR.Tn[11].n66 0.848714
R22608 XThR.Tn[11] XThR.Tn[11].n71 0.848714
R22609 XThR.Tn[11] XThR.Tn[11].n76 0.848714
R22610 XThR.Tn[11] XThR.Tn[11].n81 0.848714
R22611 XThR.Tn[11] XThR.Tn[11].n86 0.848714
R22612 XThR.Tn[11].n11 XThR.Tn[11] 0.485653
R22613 XThR.Tn[11].n84 XThR.Tn[11] 0.21482
R22614 XThR.Tn[11].n79 XThR.Tn[11] 0.21482
R22615 XThR.Tn[11].n74 XThR.Tn[11] 0.21482
R22616 XThR.Tn[11].n69 XThR.Tn[11] 0.21482
R22617 XThR.Tn[11].n64 XThR.Tn[11] 0.21482
R22618 XThR.Tn[11].n59 XThR.Tn[11] 0.21482
R22619 XThR.Tn[11].n54 XThR.Tn[11] 0.21482
R22620 XThR.Tn[11].n49 XThR.Tn[11] 0.21482
R22621 XThR.Tn[11].n44 XThR.Tn[11] 0.21482
R22622 XThR.Tn[11].n39 XThR.Tn[11] 0.21482
R22623 XThR.Tn[11].n34 XThR.Tn[11] 0.21482
R22624 XThR.Tn[11].n29 XThR.Tn[11] 0.21482
R22625 XThR.Tn[11].n24 XThR.Tn[11] 0.21482
R22626 XThR.Tn[11].n19 XThR.Tn[11] 0.21482
R22627 XThR.Tn[11].n14 XThR.Tn[11] 0.21482
R22628 XThR.Tn[11].n85 XThR.Tn[11] 0.0608448
R22629 XThR.Tn[11].n80 XThR.Tn[11] 0.0608448
R22630 XThR.Tn[11].n75 XThR.Tn[11] 0.0608448
R22631 XThR.Tn[11].n70 XThR.Tn[11] 0.0608448
R22632 XThR.Tn[11].n65 XThR.Tn[11] 0.0608448
R22633 XThR.Tn[11].n60 XThR.Tn[11] 0.0608448
R22634 XThR.Tn[11].n55 XThR.Tn[11] 0.0608448
R22635 XThR.Tn[11].n50 XThR.Tn[11] 0.0608448
R22636 XThR.Tn[11].n45 XThR.Tn[11] 0.0608448
R22637 XThR.Tn[11].n40 XThR.Tn[11] 0.0608448
R22638 XThR.Tn[11].n35 XThR.Tn[11] 0.0608448
R22639 XThR.Tn[11].n30 XThR.Tn[11] 0.0608448
R22640 XThR.Tn[11].n25 XThR.Tn[11] 0.0608448
R22641 XThR.Tn[11].n20 XThR.Tn[11] 0.0608448
R22642 XThR.Tn[11].n15 XThR.Tn[11] 0.0608448
R22643 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R22644 XThR.Tn[11] XThR.Tn[11].n87 0.038
R22645 XThR.Tn[11].n11 XThR.Tn[11] 0.00744444
R22646 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00265517
R22647 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00265517
R22648 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00265517
R22649 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00265517
R22650 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00265517
R22651 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00265517
R22652 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00265517
R22653 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00265517
R22654 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00265517
R22655 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00265517
R22656 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00265517
R22657 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00265517
R22658 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00265517
R22659 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00265517
R22660 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00265517
R22661 XThR.Tn[13].n87 XThR.Tn[13].n86 256.104
R22662 XThR.Tn[13].n2 XThR.Tn[13].n1 243.68
R22663 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R22664 XThR.Tn[13].n2 XThR.Tn[13].n0 205.28
R22665 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R22666 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R22667 XThR.Tn[13] XThR.Tn[13].n78 161.363
R22668 XThR.Tn[13] XThR.Tn[13].n73 161.363
R22669 XThR.Tn[13] XThR.Tn[13].n68 161.363
R22670 XThR.Tn[13] XThR.Tn[13].n63 161.363
R22671 XThR.Tn[13] XThR.Tn[13].n58 161.363
R22672 XThR.Tn[13] XThR.Tn[13].n53 161.363
R22673 XThR.Tn[13] XThR.Tn[13].n48 161.363
R22674 XThR.Tn[13] XThR.Tn[13].n43 161.363
R22675 XThR.Tn[13] XThR.Tn[13].n38 161.363
R22676 XThR.Tn[13] XThR.Tn[13].n33 161.363
R22677 XThR.Tn[13] XThR.Tn[13].n28 161.363
R22678 XThR.Tn[13] XThR.Tn[13].n23 161.363
R22679 XThR.Tn[13] XThR.Tn[13].n18 161.363
R22680 XThR.Tn[13] XThR.Tn[13].n13 161.363
R22681 XThR.Tn[13] XThR.Tn[13].n8 161.363
R22682 XThR.Tn[13] XThR.Tn[13].n6 161.363
R22683 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R22684 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R22685 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R22686 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R22687 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R22688 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R22689 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R22690 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R22691 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R22692 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R22693 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R22694 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R22695 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R22696 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R22697 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R22698 XThR.Tn[13].n79 XThR.Tn[13].t28 161.106
R22699 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R22700 XThR.Tn[13].n74 XThR.Tn[13].t37 161.106
R22701 XThR.Tn[13].n73 XThR.Tn[13].t61 161.106
R22702 XThR.Tn[13].n69 XThR.Tn[13].t20 161.106
R22703 XThR.Tn[13].n68 XThR.Tn[13].t44 161.106
R22704 XThR.Tn[13].n64 XThR.Tn[13].t64 161.106
R22705 XThR.Tn[13].n63 XThR.Tn[13].t25 161.106
R22706 XThR.Tn[13].n59 XThR.Tn[13].t27 161.106
R22707 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R22708 XThR.Tn[13].n54 XThR.Tn[13].t53 161.106
R22709 XThR.Tn[13].n53 XThR.Tn[13].t15 161.106
R22710 XThR.Tn[13].n49 XThR.Tn[13].t35 161.106
R22711 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R22712 XThR.Tn[13].n44 XThR.Tn[13].t17 161.106
R22713 XThR.Tn[13].n43 XThR.Tn[13].t41 161.106
R22714 XThR.Tn[13].n39 XThR.Tn[13].t63 161.106
R22715 XThR.Tn[13].n38 XThR.Tn[13].t23 161.106
R22716 XThR.Tn[13].n34 XThR.Tn[13].t68 161.106
R22717 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R22718 XThR.Tn[13].n29 XThR.Tn[13].t52 161.106
R22719 XThR.Tn[13].n28 XThR.Tn[13].t14 161.106
R22720 XThR.Tn[13].n24 XThR.Tn[13].t19 161.106
R22721 XThR.Tn[13].n23 XThR.Tn[13].t43 161.106
R22722 XThR.Tn[13].n19 XThR.Tn[13].t50 161.106
R22723 XThR.Tn[13].n18 XThR.Tn[13].t12 161.106
R22724 XThR.Tn[13].n14 XThR.Tn[13].t33 161.106
R22725 XThR.Tn[13].n13 XThR.Tn[13].t58 161.106
R22726 XThR.Tn[13].n9 XThR.Tn[13].t57 161.106
R22727 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R22728 XThR.Tn[13].n6 XThR.Tn[13].t65 161.106
R22729 XThR.Tn[13].n79 XThR.Tn[13].t47 154.679
R22730 XThR.Tn[13].n78 XThR.Tn[13].t73 154.679
R22731 XThR.Tn[13].n74 XThR.Tn[13].t26 154.679
R22732 XThR.Tn[13].n73 XThR.Tn[13].t49 154.679
R22733 XThR.Tn[13].n69 XThR.Tn[13].t70 154.679
R22734 XThR.Tn[13].n68 XThR.Tn[13].t32 154.679
R22735 XThR.Tn[13].n64 XThR.Tn[13].t38 154.679
R22736 XThR.Tn[13].n63 XThR.Tn[13].t62 154.679
R22737 XThR.Tn[13].n59 XThR.Tn[13].t22 154.679
R22738 XThR.Tn[13].n58 XThR.Tn[13].t45 154.679
R22739 XThR.Tn[13].n54 XThR.Tn[13].t46 154.679
R22740 XThR.Tn[13].n53 XThR.Tn[13].t72 154.679
R22741 XThR.Tn[13].n49 XThR.Tn[13].t71 154.679
R22742 XThR.Tn[13].n48 XThR.Tn[13].t34 154.679
R22743 XThR.Tn[13].n44 XThR.Tn[13].t54 154.679
R22744 XThR.Tn[13].n43 XThR.Tn[13].t16 154.679
R22745 XThR.Tn[13].n39 XThR.Tn[13].t36 154.679
R22746 XThR.Tn[13].n38 XThR.Tn[13].t60 154.679
R22747 XThR.Tn[13].n34 XThR.Tn[13].t18 154.679
R22748 XThR.Tn[13].n33 XThR.Tn[13].t42 154.679
R22749 XThR.Tn[13].n29 XThR.Tn[13].t24 154.679
R22750 XThR.Tn[13].n28 XThR.Tn[13].t48 154.679
R22751 XThR.Tn[13].n24 XThR.Tn[13].t69 154.679
R22752 XThR.Tn[13].n23 XThR.Tn[13].t31 154.679
R22753 XThR.Tn[13].n19 XThR.Tn[13].t40 154.679
R22754 XThR.Tn[13].n18 XThR.Tn[13].t66 154.679
R22755 XThR.Tn[13].n14 XThR.Tn[13].t67 154.679
R22756 XThR.Tn[13].n13 XThR.Tn[13].t29 154.679
R22757 XThR.Tn[13].n9 XThR.Tn[13].t51 154.679
R22758 XThR.Tn[13].n8 XThR.Tn[13].t13 154.679
R22759 XThR.Tn[13].n6 XThR.Tn[13].t39 154.679
R22760 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R22761 XThR.Tn[13].n85 XThR.Tn[13].t6 26.5955
R22762 XThR.Tn[13].n85 XThR.Tn[13].t4 26.5955
R22763 XThR.Tn[13].n86 XThR.Tn[13].t7 26.5955
R22764 XThR.Tn[13].n86 XThR.Tn[13].t5 26.5955
R22765 XThR.Tn[13].n0 XThR.Tn[13].t2 26.5955
R22766 XThR.Tn[13].n0 XThR.Tn[13].t0 26.5955
R22767 XThR.Tn[13].n1 XThR.Tn[13].t1 26.5955
R22768 XThR.Tn[13].n1 XThR.Tn[13].t3 26.5955
R22769 XThR.Tn[13].n4 XThR.Tn[13].t10 24.9236
R22770 XThR.Tn[13].n4 XThR.Tn[13].t8 24.9236
R22771 XThR.Tn[13].n3 XThR.Tn[13].t11 24.9236
R22772 XThR.Tn[13].n3 XThR.Tn[13].t9 24.9236
R22773 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R22774 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R22775 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R22776 XThR.Tn[13] XThR.Tn[13].n7 5.34871
R22777 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R22778 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R22779 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R22780 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R22781 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R22782 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R22783 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R22784 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R22785 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R22786 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R22787 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R22788 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R22789 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R22790 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R22791 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R22792 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R22793 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R22794 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R22795 XThR.Tn[13].n12 XThR.Tn[13] 2.51836
R22796 XThR.Tn[13].n17 XThR.Tn[13] 2.51836
R22797 XThR.Tn[13].n22 XThR.Tn[13] 2.51836
R22798 XThR.Tn[13].n27 XThR.Tn[13] 2.51836
R22799 XThR.Tn[13].n32 XThR.Tn[13] 2.51836
R22800 XThR.Tn[13].n37 XThR.Tn[13] 2.51836
R22801 XThR.Tn[13].n42 XThR.Tn[13] 2.51836
R22802 XThR.Tn[13].n47 XThR.Tn[13] 2.51836
R22803 XThR.Tn[13].n52 XThR.Tn[13] 2.51836
R22804 XThR.Tn[13].n57 XThR.Tn[13] 2.51836
R22805 XThR.Tn[13].n62 XThR.Tn[13] 2.51836
R22806 XThR.Tn[13].n67 XThR.Tn[13] 2.51836
R22807 XThR.Tn[13].n72 XThR.Tn[13] 2.51836
R22808 XThR.Tn[13].n77 XThR.Tn[13] 2.51836
R22809 XThR.Tn[13].n82 XThR.Tn[13] 2.51836
R22810 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R22811 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R22812 XThR.Tn[13] XThR.Tn[13].n12 0.848714
R22813 XThR.Tn[13] XThR.Tn[13].n17 0.848714
R22814 XThR.Tn[13] XThR.Tn[13].n22 0.848714
R22815 XThR.Tn[13] XThR.Tn[13].n27 0.848714
R22816 XThR.Tn[13] XThR.Tn[13].n32 0.848714
R22817 XThR.Tn[13] XThR.Tn[13].n37 0.848714
R22818 XThR.Tn[13] XThR.Tn[13].n42 0.848714
R22819 XThR.Tn[13] XThR.Tn[13].n47 0.848714
R22820 XThR.Tn[13] XThR.Tn[13].n52 0.848714
R22821 XThR.Tn[13] XThR.Tn[13].n57 0.848714
R22822 XThR.Tn[13] XThR.Tn[13].n62 0.848714
R22823 XThR.Tn[13] XThR.Tn[13].n67 0.848714
R22824 XThR.Tn[13] XThR.Tn[13].n72 0.848714
R22825 XThR.Tn[13] XThR.Tn[13].n77 0.848714
R22826 XThR.Tn[13] XThR.Tn[13].n82 0.848714
R22827 XThR.Tn[13].n7 XThR.Tn[13] 0.485653
R22828 XThR.Tn[13].n80 XThR.Tn[13] 0.21482
R22829 XThR.Tn[13].n75 XThR.Tn[13] 0.21482
R22830 XThR.Tn[13].n70 XThR.Tn[13] 0.21482
R22831 XThR.Tn[13].n65 XThR.Tn[13] 0.21482
R22832 XThR.Tn[13].n60 XThR.Tn[13] 0.21482
R22833 XThR.Tn[13].n55 XThR.Tn[13] 0.21482
R22834 XThR.Tn[13].n50 XThR.Tn[13] 0.21482
R22835 XThR.Tn[13].n45 XThR.Tn[13] 0.21482
R22836 XThR.Tn[13].n40 XThR.Tn[13] 0.21482
R22837 XThR.Tn[13].n35 XThR.Tn[13] 0.21482
R22838 XThR.Tn[13].n30 XThR.Tn[13] 0.21482
R22839 XThR.Tn[13].n25 XThR.Tn[13] 0.21482
R22840 XThR.Tn[13].n20 XThR.Tn[13] 0.21482
R22841 XThR.Tn[13].n15 XThR.Tn[13] 0.21482
R22842 XThR.Tn[13].n10 XThR.Tn[13] 0.21482
R22843 XThR.Tn[13].n81 XThR.Tn[13] 0.0608448
R22844 XThR.Tn[13].n76 XThR.Tn[13] 0.0608448
R22845 XThR.Tn[13].n71 XThR.Tn[13] 0.0608448
R22846 XThR.Tn[13].n66 XThR.Tn[13] 0.0608448
R22847 XThR.Tn[13].n61 XThR.Tn[13] 0.0608448
R22848 XThR.Tn[13].n56 XThR.Tn[13] 0.0608448
R22849 XThR.Tn[13].n51 XThR.Tn[13] 0.0608448
R22850 XThR.Tn[13].n46 XThR.Tn[13] 0.0608448
R22851 XThR.Tn[13].n41 XThR.Tn[13] 0.0608448
R22852 XThR.Tn[13].n36 XThR.Tn[13] 0.0608448
R22853 XThR.Tn[13].n31 XThR.Tn[13] 0.0608448
R22854 XThR.Tn[13].n26 XThR.Tn[13] 0.0608448
R22855 XThR.Tn[13].n21 XThR.Tn[13] 0.0608448
R22856 XThR.Tn[13].n16 XThR.Tn[13] 0.0608448
R22857 XThR.Tn[13].n11 XThR.Tn[13] 0.0608448
R22858 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R22859 XThR.Tn[13] XThR.Tn[13].n83 0.038
R22860 XThR.Tn[13].n7 XThR.Tn[13] 0.00744444
R22861 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00265517
R22862 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00265517
R22863 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00265517
R22864 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00265517
R22865 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00265517
R22866 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00265517
R22867 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00265517
R22868 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00265517
R22869 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00265517
R22870 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00265517
R22871 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00265517
R22872 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00265517
R22873 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00265517
R22874 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00265517
R22875 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00265517
R22876 XThC.Tn[14].n70 XThC.Tn[14].n69 256.103
R22877 XThC.Tn[14].n74 XThC.Tn[14].n72 243.68
R22878 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22879 XThC.Tn[14].n74 XThC.Tn[14].n73 205.28
R22880 XThC.Tn[14].n70 XThC.Tn[14].n68 202.095
R22881 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22882 XThC.Tn[14].n64 XThC.Tn[14].n62 161.365
R22883 XThC.Tn[14].n60 XThC.Tn[14].n58 161.365
R22884 XThC.Tn[14].n56 XThC.Tn[14].n54 161.365
R22885 XThC.Tn[14].n52 XThC.Tn[14].n50 161.365
R22886 XThC.Tn[14].n48 XThC.Tn[14].n46 161.365
R22887 XThC.Tn[14].n44 XThC.Tn[14].n42 161.365
R22888 XThC.Tn[14].n40 XThC.Tn[14].n38 161.365
R22889 XThC.Tn[14].n36 XThC.Tn[14].n34 161.365
R22890 XThC.Tn[14].n32 XThC.Tn[14].n30 161.365
R22891 XThC.Tn[14].n28 XThC.Tn[14].n26 161.365
R22892 XThC.Tn[14].n24 XThC.Tn[14].n22 161.365
R22893 XThC.Tn[14].n20 XThC.Tn[14].n18 161.365
R22894 XThC.Tn[14].n16 XThC.Tn[14].n14 161.365
R22895 XThC.Tn[14].n12 XThC.Tn[14].n10 161.365
R22896 XThC.Tn[14].n8 XThC.Tn[14].n6 161.365
R22897 XThC.Tn[14].n5 XThC.Tn[14].n3 161.365
R22898 XThC.Tn[14].n62 XThC.Tn[14].t33 161.106
R22899 XThC.Tn[14].n58 XThC.Tn[14].t12 161.106
R22900 XThC.Tn[14].n54 XThC.Tn[14].t43 161.106
R22901 XThC.Tn[14].n50 XThC.Tn[14].t40 161.106
R22902 XThC.Tn[14].n46 XThC.Tn[14].t22 161.106
R22903 XThC.Tn[14].n42 XThC.Tn[14].t20 161.106
R22904 XThC.Tn[14].n38 XThC.Tn[14].t39 161.106
R22905 XThC.Tn[14].n34 XThC.Tn[14].t31 161.106
R22906 XThC.Tn[14].n30 XThC.Tn[14].t28 161.106
R22907 XThC.Tn[14].n26 XThC.Tn[14].t19 161.106
R22908 XThC.Tn[14].n22 XThC.Tn[14].t38 161.106
R22909 XThC.Tn[14].n18 XThC.Tn[14].t27 161.106
R22910 XThC.Tn[14].n14 XThC.Tn[14].t18 161.106
R22911 XThC.Tn[14].n10 XThC.Tn[14].t16 161.106
R22912 XThC.Tn[14].n6 XThC.Tn[14].t34 161.106
R22913 XThC.Tn[14].n3 XThC.Tn[14].t26 161.106
R22914 XThC.Tn[14].n62 XThC.Tn[14].t30 154.679
R22915 XThC.Tn[14].n58 XThC.Tn[14].t42 154.679
R22916 XThC.Tn[14].n54 XThC.Tn[14].t41 154.679
R22917 XThC.Tn[14].n50 XThC.Tn[14].t37 154.679
R22918 XThC.Tn[14].n46 XThC.Tn[14].t21 154.679
R22919 XThC.Tn[14].n42 XThC.Tn[14].t17 154.679
R22920 XThC.Tn[14].n38 XThC.Tn[14].t36 154.679
R22921 XThC.Tn[14].n34 XThC.Tn[14].t29 154.679
R22922 XThC.Tn[14].n30 XThC.Tn[14].t25 154.679
R22923 XThC.Tn[14].n26 XThC.Tn[14].t15 154.679
R22924 XThC.Tn[14].n22 XThC.Tn[14].t35 154.679
R22925 XThC.Tn[14].n18 XThC.Tn[14].t24 154.679
R22926 XThC.Tn[14].n14 XThC.Tn[14].t14 154.679
R22927 XThC.Tn[14].n10 XThC.Tn[14].t13 154.679
R22928 XThC.Tn[14].n6 XThC.Tn[14].t32 154.679
R22929 XThC.Tn[14].n3 XThC.Tn[14].t23 154.679
R22930 XThC.Tn[14].n68 XThC.Tn[14].t0 26.5955
R22931 XThC.Tn[14].n68 XThC.Tn[14].t1 26.5955
R22932 XThC.Tn[14].n72 XThC.Tn[14].t11 26.5955
R22933 XThC.Tn[14].n72 XThC.Tn[14].t10 26.5955
R22934 XThC.Tn[14].n73 XThC.Tn[14].t9 26.5955
R22935 XThC.Tn[14].n73 XThC.Tn[14].t8 26.5955
R22936 XThC.Tn[14].n69 XThC.Tn[14].t3 26.5955
R22937 XThC.Tn[14].n69 XThC.Tn[14].t2 26.5955
R22938 XThC.Tn[14].n1 XThC.Tn[14].t5 24.9236
R22939 XThC.Tn[14].n1 XThC.Tn[14].t7 24.9236
R22940 XThC.Tn[14].n0 XThC.Tn[14].t4 24.9236
R22941 XThC.Tn[14].n0 XThC.Tn[14].t6 24.9236
R22942 XThC.Tn[14] XThC.Tn[14].n74 22.9652
R22943 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22944 XThC.Tn[14].n71 XThC.Tn[14].n70 13.9299
R22945 XThC.Tn[14] XThC.Tn[14].n71 13.9299
R22946 XThC.Tn[14] XThC.Tn[14].n5 8.0245
R22947 XThC.Tn[14].n65 XThC.Tn[14].n64 7.9105
R22948 XThC.Tn[14].n61 XThC.Tn[14].n60 7.9105
R22949 XThC.Tn[14].n57 XThC.Tn[14].n56 7.9105
R22950 XThC.Tn[14].n53 XThC.Tn[14].n52 7.9105
R22951 XThC.Tn[14].n49 XThC.Tn[14].n48 7.9105
R22952 XThC.Tn[14].n45 XThC.Tn[14].n44 7.9105
R22953 XThC.Tn[14].n41 XThC.Tn[14].n40 7.9105
R22954 XThC.Tn[14].n37 XThC.Tn[14].n36 7.9105
R22955 XThC.Tn[14].n33 XThC.Tn[14].n32 7.9105
R22956 XThC.Tn[14].n29 XThC.Tn[14].n28 7.9105
R22957 XThC.Tn[14].n25 XThC.Tn[14].n24 7.9105
R22958 XThC.Tn[14].n21 XThC.Tn[14].n20 7.9105
R22959 XThC.Tn[14].n17 XThC.Tn[14].n16 7.9105
R22960 XThC.Tn[14].n13 XThC.Tn[14].n12 7.9105
R22961 XThC.Tn[14].n9 XThC.Tn[14].n8 7.9105
R22962 XThC.Tn[14].n67 XThC.Tn[14].n66 7.51947
R22963 XThC.Tn[14].n66 XThC.Tn[14] 5.85107
R22964 XThC.Tn[14].n71 XThC.Tn[14].n67 2.99115
R22965 XThC.Tn[14].n71 XThC.Tn[14] 2.87153
R22966 XThC.Tn[14].n67 XThC.Tn[14] 2.2734
R22967 XThC.Tn[14].n66 XThC.Tn[14] 1.06164
R22968 XThC.Tn[14].n9 XThC.Tn[14] 0.235138
R22969 XThC.Tn[14].n13 XThC.Tn[14] 0.235138
R22970 XThC.Tn[14].n17 XThC.Tn[14] 0.235138
R22971 XThC.Tn[14].n21 XThC.Tn[14] 0.235138
R22972 XThC.Tn[14].n25 XThC.Tn[14] 0.235138
R22973 XThC.Tn[14].n29 XThC.Tn[14] 0.235138
R22974 XThC.Tn[14].n33 XThC.Tn[14] 0.235138
R22975 XThC.Tn[14].n37 XThC.Tn[14] 0.235138
R22976 XThC.Tn[14].n41 XThC.Tn[14] 0.235138
R22977 XThC.Tn[14].n45 XThC.Tn[14] 0.235138
R22978 XThC.Tn[14].n49 XThC.Tn[14] 0.235138
R22979 XThC.Tn[14].n53 XThC.Tn[14] 0.235138
R22980 XThC.Tn[14].n57 XThC.Tn[14] 0.235138
R22981 XThC.Tn[14].n61 XThC.Tn[14] 0.235138
R22982 XThC.Tn[14].n65 XThC.Tn[14] 0.235138
R22983 XThC.Tn[14] XThC.Tn[14].n9 0.114505
R22984 XThC.Tn[14] XThC.Tn[14].n13 0.114505
R22985 XThC.Tn[14] XThC.Tn[14].n17 0.114505
R22986 XThC.Tn[14] XThC.Tn[14].n21 0.114505
R22987 XThC.Tn[14] XThC.Tn[14].n25 0.114505
R22988 XThC.Tn[14] XThC.Tn[14].n29 0.114505
R22989 XThC.Tn[14] XThC.Tn[14].n33 0.114505
R22990 XThC.Tn[14] XThC.Tn[14].n37 0.114505
R22991 XThC.Tn[14] XThC.Tn[14].n41 0.114505
R22992 XThC.Tn[14] XThC.Tn[14].n45 0.114505
R22993 XThC.Tn[14] XThC.Tn[14].n49 0.114505
R22994 XThC.Tn[14] XThC.Tn[14].n53 0.114505
R22995 XThC.Tn[14] XThC.Tn[14].n57 0.114505
R22996 XThC.Tn[14] XThC.Tn[14].n61 0.114505
R22997 XThC.Tn[14] XThC.Tn[14].n65 0.114505
R22998 XThC.Tn[14].n64 XThC.Tn[14].n63 0.0599512
R22999 XThC.Tn[14].n60 XThC.Tn[14].n59 0.0599512
R23000 XThC.Tn[14].n56 XThC.Tn[14].n55 0.0599512
R23001 XThC.Tn[14].n52 XThC.Tn[14].n51 0.0599512
R23002 XThC.Tn[14].n48 XThC.Tn[14].n47 0.0599512
R23003 XThC.Tn[14].n44 XThC.Tn[14].n43 0.0599512
R23004 XThC.Tn[14].n40 XThC.Tn[14].n39 0.0599512
R23005 XThC.Tn[14].n36 XThC.Tn[14].n35 0.0599512
R23006 XThC.Tn[14].n32 XThC.Tn[14].n31 0.0599512
R23007 XThC.Tn[14].n28 XThC.Tn[14].n27 0.0599512
R23008 XThC.Tn[14].n24 XThC.Tn[14].n23 0.0599512
R23009 XThC.Tn[14].n20 XThC.Tn[14].n19 0.0599512
R23010 XThC.Tn[14].n16 XThC.Tn[14].n15 0.0599512
R23011 XThC.Tn[14].n12 XThC.Tn[14].n11 0.0599512
R23012 XThC.Tn[14].n8 XThC.Tn[14].n7 0.0599512
R23013 XThC.Tn[14].n5 XThC.Tn[14].n4 0.0599512
R23014 XThC.Tn[14].n63 XThC.Tn[14] 0.0469286
R23015 XThC.Tn[14].n59 XThC.Tn[14] 0.0469286
R23016 XThC.Tn[14].n55 XThC.Tn[14] 0.0469286
R23017 XThC.Tn[14].n51 XThC.Tn[14] 0.0469286
R23018 XThC.Tn[14].n47 XThC.Tn[14] 0.0469286
R23019 XThC.Tn[14].n43 XThC.Tn[14] 0.0469286
R23020 XThC.Tn[14].n39 XThC.Tn[14] 0.0469286
R23021 XThC.Tn[14].n35 XThC.Tn[14] 0.0469286
R23022 XThC.Tn[14].n31 XThC.Tn[14] 0.0469286
R23023 XThC.Tn[14].n27 XThC.Tn[14] 0.0469286
R23024 XThC.Tn[14].n23 XThC.Tn[14] 0.0469286
R23025 XThC.Tn[14].n19 XThC.Tn[14] 0.0469286
R23026 XThC.Tn[14].n15 XThC.Tn[14] 0.0469286
R23027 XThC.Tn[14].n11 XThC.Tn[14] 0.0469286
R23028 XThC.Tn[14].n7 XThC.Tn[14] 0.0469286
R23029 XThC.Tn[14].n4 XThC.Tn[14] 0.0469286
R23030 XThC.Tn[14].n63 XThC.Tn[14] 0.0401341
R23031 XThC.Tn[14].n59 XThC.Tn[14] 0.0401341
R23032 XThC.Tn[14].n55 XThC.Tn[14] 0.0401341
R23033 XThC.Tn[14].n51 XThC.Tn[14] 0.0401341
R23034 XThC.Tn[14].n47 XThC.Tn[14] 0.0401341
R23035 XThC.Tn[14].n43 XThC.Tn[14] 0.0401341
R23036 XThC.Tn[14].n39 XThC.Tn[14] 0.0401341
R23037 XThC.Tn[14].n35 XThC.Tn[14] 0.0401341
R23038 XThC.Tn[14].n31 XThC.Tn[14] 0.0401341
R23039 XThC.Tn[14].n27 XThC.Tn[14] 0.0401341
R23040 XThC.Tn[14].n23 XThC.Tn[14] 0.0401341
R23041 XThC.Tn[14].n19 XThC.Tn[14] 0.0401341
R23042 XThC.Tn[14].n15 XThC.Tn[14] 0.0401341
R23043 XThC.Tn[14].n11 XThC.Tn[14] 0.0401341
R23044 XThC.Tn[14].n7 XThC.Tn[14] 0.0401341
R23045 XThC.Tn[14].n4 XThC.Tn[14] 0.0401341
R23046 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R23047 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R23048 XThR.Tn[1] XThR.Tn[1].n82 161.363
R23049 XThR.Tn[1] XThR.Tn[1].n77 161.363
R23050 XThR.Tn[1] XThR.Tn[1].n72 161.363
R23051 XThR.Tn[1] XThR.Tn[1].n67 161.363
R23052 XThR.Tn[1] XThR.Tn[1].n62 161.363
R23053 XThR.Tn[1] XThR.Tn[1].n57 161.363
R23054 XThR.Tn[1] XThR.Tn[1].n52 161.363
R23055 XThR.Tn[1] XThR.Tn[1].n47 161.363
R23056 XThR.Tn[1] XThR.Tn[1].n42 161.363
R23057 XThR.Tn[1] XThR.Tn[1].n37 161.363
R23058 XThR.Tn[1] XThR.Tn[1].n32 161.363
R23059 XThR.Tn[1] XThR.Tn[1].n27 161.363
R23060 XThR.Tn[1] XThR.Tn[1].n22 161.363
R23061 XThR.Tn[1] XThR.Tn[1].n17 161.363
R23062 XThR.Tn[1] XThR.Tn[1].n12 161.363
R23063 XThR.Tn[1] XThR.Tn[1].n10 161.363
R23064 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R23065 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R23066 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R23067 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R23068 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R23069 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R23070 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R23071 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R23072 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R23073 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R23074 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R23075 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R23076 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R23077 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R23078 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R23079 XThR.Tn[1].n83 XThR.Tn[1].t43 161.106
R23080 XThR.Tn[1].n82 XThR.Tn[1].t45 161.106
R23081 XThR.Tn[1].n78 XThR.Tn[1].t49 161.106
R23082 XThR.Tn[1].n77 XThR.Tn[1].t54 161.106
R23083 XThR.Tn[1].n73 XThR.Tn[1].t31 161.106
R23084 XThR.Tn[1].n72 XThR.Tn[1].t36 161.106
R23085 XThR.Tn[1].n68 XThR.Tn[1].t14 161.106
R23086 XThR.Tn[1].n67 XThR.Tn[1].t16 161.106
R23087 XThR.Tn[1].n63 XThR.Tn[1].t42 161.106
R23088 XThR.Tn[1].n62 XThR.Tn[1].t44 161.106
R23089 XThR.Tn[1].n58 XThR.Tn[1].t66 161.106
R23090 XThR.Tn[1].n57 XThR.Tn[1].t71 161.106
R23091 XThR.Tn[1].n53 XThR.Tn[1].t47 161.106
R23092 XThR.Tn[1].n52 XThR.Tn[1].t52 161.106
R23093 XThR.Tn[1].n48 XThR.Tn[1].t28 161.106
R23094 XThR.Tn[1].n47 XThR.Tn[1].t33 161.106
R23095 XThR.Tn[1].n43 XThR.Tn[1].t13 161.106
R23096 XThR.Tn[1].n42 XThR.Tn[1].t15 161.106
R23097 XThR.Tn[1].n38 XThR.Tn[1].t18 161.106
R23098 XThR.Tn[1].n37 XThR.Tn[1].t23 161.106
R23099 XThR.Tn[1].n33 XThR.Tn[1].t65 161.106
R23100 XThR.Tn[1].n32 XThR.Tn[1].t70 161.106
R23101 XThR.Tn[1].n28 XThR.Tn[1].t30 161.106
R23102 XThR.Tn[1].n27 XThR.Tn[1].t35 161.106
R23103 XThR.Tn[1].n23 XThR.Tn[1].t62 161.106
R23104 XThR.Tn[1].n22 XThR.Tn[1].t68 161.106
R23105 XThR.Tn[1].n18 XThR.Tn[1].t46 161.106
R23106 XThR.Tn[1].n17 XThR.Tn[1].t50 161.106
R23107 XThR.Tn[1].n13 XThR.Tn[1].t73 161.106
R23108 XThR.Tn[1].n12 XThR.Tn[1].t12 161.106
R23109 XThR.Tn[1].n10 XThR.Tn[1].t57 161.106
R23110 XThR.Tn[1].n83 XThR.Tn[1].t60 154.679
R23111 XThR.Tn[1].n82 XThR.Tn[1].t63 154.679
R23112 XThR.Tn[1].n78 XThR.Tn[1].t39 154.679
R23113 XThR.Tn[1].n77 XThR.Tn[1].t41 154.679
R23114 XThR.Tn[1].n73 XThR.Tn[1].t20 154.679
R23115 XThR.Tn[1].n72 XThR.Tn[1].t25 154.679
R23116 XThR.Tn[1].n68 XThR.Tn[1].t51 154.679
R23117 XThR.Tn[1].n67 XThR.Tn[1].t55 154.679
R23118 XThR.Tn[1].n63 XThR.Tn[1].t32 154.679
R23119 XThR.Tn[1].n62 XThR.Tn[1].t37 154.679
R23120 XThR.Tn[1].n58 XThR.Tn[1].t59 154.679
R23121 XThR.Tn[1].n57 XThR.Tn[1].t61 154.679
R23122 XThR.Tn[1].n53 XThR.Tn[1].t21 154.679
R23123 XThR.Tn[1].n52 XThR.Tn[1].t26 154.679
R23124 XThR.Tn[1].n48 XThR.Tn[1].t67 154.679
R23125 XThR.Tn[1].n47 XThR.Tn[1].t72 154.679
R23126 XThR.Tn[1].n43 XThR.Tn[1].t48 154.679
R23127 XThR.Tn[1].n42 XThR.Tn[1].t53 154.679
R23128 XThR.Tn[1].n38 XThR.Tn[1].t29 154.679
R23129 XThR.Tn[1].n37 XThR.Tn[1].t34 154.679
R23130 XThR.Tn[1].n33 XThR.Tn[1].t38 154.679
R23131 XThR.Tn[1].n32 XThR.Tn[1].t40 154.679
R23132 XThR.Tn[1].n28 XThR.Tn[1].t19 154.679
R23133 XThR.Tn[1].n27 XThR.Tn[1].t24 154.679
R23134 XThR.Tn[1].n23 XThR.Tn[1].t56 154.679
R23135 XThR.Tn[1].n22 XThR.Tn[1].t58 154.679
R23136 XThR.Tn[1].n18 XThR.Tn[1].t17 154.679
R23137 XThR.Tn[1].n17 XThR.Tn[1].t22 154.679
R23138 XThR.Tn[1].n13 XThR.Tn[1].t64 154.679
R23139 XThR.Tn[1].n12 XThR.Tn[1].t69 154.679
R23140 XThR.Tn[1].n10 XThR.Tn[1].t27 154.679
R23141 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R23142 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R23143 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R23144 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R23145 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R23146 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R23147 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R23148 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R23149 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R23150 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R23151 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R23152 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R23153 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R23154 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R23155 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R23156 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R23157 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R23158 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R23159 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R23160 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R23161 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R23162 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R23163 XThR.Tn[1] XThR.Tn[1].n11 5.34871
R23164 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R23165 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R23166 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R23167 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R23168 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R23169 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R23170 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R23171 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R23172 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R23173 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R23174 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R23175 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R23176 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R23177 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R23178 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R23179 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R23180 XThR.Tn[1].n16 XThR.Tn[1] 2.51836
R23181 XThR.Tn[1].n21 XThR.Tn[1] 2.51836
R23182 XThR.Tn[1].n26 XThR.Tn[1] 2.51836
R23183 XThR.Tn[1].n31 XThR.Tn[1] 2.51836
R23184 XThR.Tn[1].n36 XThR.Tn[1] 2.51836
R23185 XThR.Tn[1].n41 XThR.Tn[1] 2.51836
R23186 XThR.Tn[1].n46 XThR.Tn[1] 2.51836
R23187 XThR.Tn[1].n51 XThR.Tn[1] 2.51836
R23188 XThR.Tn[1].n56 XThR.Tn[1] 2.51836
R23189 XThR.Tn[1].n61 XThR.Tn[1] 2.51836
R23190 XThR.Tn[1].n66 XThR.Tn[1] 2.51836
R23191 XThR.Tn[1].n71 XThR.Tn[1] 2.51836
R23192 XThR.Tn[1].n76 XThR.Tn[1] 2.51836
R23193 XThR.Tn[1].n81 XThR.Tn[1] 2.51836
R23194 XThR.Tn[1].n86 XThR.Tn[1] 2.51836
R23195 XThR.Tn[1] XThR.Tn[1].n16 0.848714
R23196 XThR.Tn[1] XThR.Tn[1].n21 0.848714
R23197 XThR.Tn[1] XThR.Tn[1].n26 0.848714
R23198 XThR.Tn[1] XThR.Tn[1].n31 0.848714
R23199 XThR.Tn[1] XThR.Tn[1].n36 0.848714
R23200 XThR.Tn[1] XThR.Tn[1].n41 0.848714
R23201 XThR.Tn[1] XThR.Tn[1].n46 0.848714
R23202 XThR.Tn[1] XThR.Tn[1].n51 0.848714
R23203 XThR.Tn[1] XThR.Tn[1].n56 0.848714
R23204 XThR.Tn[1] XThR.Tn[1].n61 0.848714
R23205 XThR.Tn[1] XThR.Tn[1].n66 0.848714
R23206 XThR.Tn[1] XThR.Tn[1].n71 0.848714
R23207 XThR.Tn[1] XThR.Tn[1].n76 0.848714
R23208 XThR.Tn[1] XThR.Tn[1].n81 0.848714
R23209 XThR.Tn[1] XThR.Tn[1].n86 0.848714
R23210 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R23211 XThR.Tn[1].n11 XThR.Tn[1] 0.485653
R23212 XThR.Tn[1].n84 XThR.Tn[1] 0.21482
R23213 XThR.Tn[1].n79 XThR.Tn[1] 0.21482
R23214 XThR.Tn[1].n74 XThR.Tn[1] 0.21482
R23215 XThR.Tn[1].n69 XThR.Tn[1] 0.21482
R23216 XThR.Tn[1].n64 XThR.Tn[1] 0.21482
R23217 XThR.Tn[1].n59 XThR.Tn[1] 0.21482
R23218 XThR.Tn[1].n54 XThR.Tn[1] 0.21482
R23219 XThR.Tn[1].n49 XThR.Tn[1] 0.21482
R23220 XThR.Tn[1].n44 XThR.Tn[1] 0.21482
R23221 XThR.Tn[1].n39 XThR.Tn[1] 0.21482
R23222 XThR.Tn[1].n34 XThR.Tn[1] 0.21482
R23223 XThR.Tn[1].n29 XThR.Tn[1] 0.21482
R23224 XThR.Tn[1].n24 XThR.Tn[1] 0.21482
R23225 XThR.Tn[1].n19 XThR.Tn[1] 0.21482
R23226 XThR.Tn[1].n14 XThR.Tn[1] 0.21482
R23227 XThR.Tn[1].n85 XThR.Tn[1] 0.0608448
R23228 XThR.Tn[1].n80 XThR.Tn[1] 0.0608448
R23229 XThR.Tn[1].n75 XThR.Tn[1] 0.0608448
R23230 XThR.Tn[1].n70 XThR.Tn[1] 0.0608448
R23231 XThR.Tn[1].n65 XThR.Tn[1] 0.0608448
R23232 XThR.Tn[1].n60 XThR.Tn[1] 0.0608448
R23233 XThR.Tn[1].n55 XThR.Tn[1] 0.0608448
R23234 XThR.Tn[1].n50 XThR.Tn[1] 0.0608448
R23235 XThR.Tn[1].n45 XThR.Tn[1] 0.0608448
R23236 XThR.Tn[1].n40 XThR.Tn[1] 0.0608448
R23237 XThR.Tn[1].n35 XThR.Tn[1] 0.0608448
R23238 XThR.Tn[1].n30 XThR.Tn[1] 0.0608448
R23239 XThR.Tn[1].n25 XThR.Tn[1] 0.0608448
R23240 XThR.Tn[1].n20 XThR.Tn[1] 0.0608448
R23241 XThR.Tn[1].n15 XThR.Tn[1] 0.0608448
R23242 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R23243 XThR.Tn[1] XThR.Tn[1].n87 0.038
R23244 XThR.Tn[1].n11 XThR.Tn[1] 0.00744444
R23245 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00265517
R23246 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00265517
R23247 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00265517
R23248 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00265517
R23249 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00265517
R23250 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00265517
R23251 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00265517
R23252 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00265517
R23253 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00265517
R23254 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00265517
R23255 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00265517
R23256 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00265517
R23257 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00265517
R23258 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00265517
R23259 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00265517
R23260 XThR.Tn[10].n5 XThR.Tn[10].n4 256.103
R23261 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R23262 XThR.Tn[10].n88 XThR.Tn[10].n86 241.847
R23263 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R23264 XThR.Tn[10].n5 XThR.Tn[10].n3 202.095
R23265 XThR.Tn[10].n88 XThR.Tn[10].n87 185
R23266 XThR.Tn[10] XThR.Tn[10].n79 161.363
R23267 XThR.Tn[10] XThR.Tn[10].n74 161.363
R23268 XThR.Tn[10] XThR.Tn[10].n69 161.363
R23269 XThR.Tn[10] XThR.Tn[10].n64 161.363
R23270 XThR.Tn[10] XThR.Tn[10].n59 161.363
R23271 XThR.Tn[10] XThR.Tn[10].n54 161.363
R23272 XThR.Tn[10] XThR.Tn[10].n49 161.363
R23273 XThR.Tn[10] XThR.Tn[10].n44 161.363
R23274 XThR.Tn[10] XThR.Tn[10].n39 161.363
R23275 XThR.Tn[10] XThR.Tn[10].n34 161.363
R23276 XThR.Tn[10] XThR.Tn[10].n29 161.363
R23277 XThR.Tn[10] XThR.Tn[10].n24 161.363
R23278 XThR.Tn[10] XThR.Tn[10].n19 161.363
R23279 XThR.Tn[10] XThR.Tn[10].n14 161.363
R23280 XThR.Tn[10] XThR.Tn[10].n9 161.363
R23281 XThR.Tn[10] XThR.Tn[10].n7 161.363
R23282 XThR.Tn[10].n81 XThR.Tn[10].n80 161.3
R23283 XThR.Tn[10].n76 XThR.Tn[10].n75 161.3
R23284 XThR.Tn[10].n71 XThR.Tn[10].n70 161.3
R23285 XThR.Tn[10].n66 XThR.Tn[10].n65 161.3
R23286 XThR.Tn[10].n61 XThR.Tn[10].n60 161.3
R23287 XThR.Tn[10].n56 XThR.Tn[10].n55 161.3
R23288 XThR.Tn[10].n51 XThR.Tn[10].n50 161.3
R23289 XThR.Tn[10].n46 XThR.Tn[10].n45 161.3
R23290 XThR.Tn[10].n41 XThR.Tn[10].n40 161.3
R23291 XThR.Tn[10].n36 XThR.Tn[10].n35 161.3
R23292 XThR.Tn[10].n31 XThR.Tn[10].n30 161.3
R23293 XThR.Tn[10].n26 XThR.Tn[10].n25 161.3
R23294 XThR.Tn[10].n21 XThR.Tn[10].n20 161.3
R23295 XThR.Tn[10].n16 XThR.Tn[10].n15 161.3
R23296 XThR.Tn[10].n11 XThR.Tn[10].n10 161.3
R23297 XThR.Tn[10].n80 XThR.Tn[10].t17 161.106
R23298 XThR.Tn[10].n79 XThR.Tn[10].t38 161.106
R23299 XThR.Tn[10].n75 XThR.Tn[10].t23 161.106
R23300 XThR.Tn[10].n74 XThR.Tn[10].t46 161.106
R23301 XThR.Tn[10].n70 XThR.Tn[10].t68 161.106
R23302 XThR.Tn[10].n69 XThR.Tn[10].t28 161.106
R23303 XThR.Tn[10].n65 XThR.Tn[10].t51 161.106
R23304 XThR.Tn[10].n64 XThR.Tn[10].t71 161.106
R23305 XThR.Tn[10].n60 XThR.Tn[10].t15 161.106
R23306 XThR.Tn[10].n59 XThR.Tn[10].t35 161.106
R23307 XThR.Tn[10].n55 XThR.Tn[10].t40 161.106
R23308 XThR.Tn[10].n54 XThR.Tn[10].t62 161.106
R23309 XThR.Tn[10].n50 XThR.Tn[10].t21 161.106
R23310 XThR.Tn[10].n49 XThR.Tn[10].t43 161.106
R23311 XThR.Tn[10].n45 XThR.Tn[10].t65 161.106
R23312 XThR.Tn[10].n44 XThR.Tn[10].t25 161.106
R23313 XThR.Tn[10].n40 XThR.Tn[10].t49 161.106
R23314 XThR.Tn[10].n39 XThR.Tn[10].t70 161.106
R23315 XThR.Tn[10].n35 XThR.Tn[10].t54 161.106
R23316 XThR.Tn[10].n34 XThR.Tn[10].t13 161.106
R23317 XThR.Tn[10].n30 XThR.Tn[10].t39 161.106
R23318 XThR.Tn[10].n29 XThR.Tn[10].t61 161.106
R23319 XThR.Tn[10].n25 XThR.Tn[10].t67 161.106
R23320 XThR.Tn[10].n24 XThR.Tn[10].t27 161.106
R23321 XThR.Tn[10].n20 XThR.Tn[10].t36 161.106
R23322 XThR.Tn[10].n19 XThR.Tn[10].t59 161.106
R23323 XThR.Tn[10].n15 XThR.Tn[10].t19 161.106
R23324 XThR.Tn[10].n14 XThR.Tn[10].t42 161.106
R23325 XThR.Tn[10].n10 XThR.Tn[10].t44 161.106
R23326 XThR.Tn[10].n9 XThR.Tn[10].t64 161.106
R23327 XThR.Tn[10].n7 XThR.Tn[10].t48 161.106
R23328 XThR.Tn[10].n80 XThR.Tn[10].t34 154.679
R23329 XThR.Tn[10].n79 XThR.Tn[10].t56 154.679
R23330 XThR.Tn[10].n75 XThR.Tn[10].t73 154.679
R23331 XThR.Tn[10].n74 XThR.Tn[10].t32 154.679
R23332 XThR.Tn[10].n70 XThR.Tn[10].t57 154.679
R23333 XThR.Tn[10].n69 XThR.Tn[10].t16 154.679
R23334 XThR.Tn[10].n65 XThR.Tn[10].t24 154.679
R23335 XThR.Tn[10].n64 XThR.Tn[10].t47 154.679
R23336 XThR.Tn[10].n60 XThR.Tn[10].t69 154.679
R23337 XThR.Tn[10].n59 XThR.Tn[10].t29 154.679
R23338 XThR.Tn[10].n55 XThR.Tn[10].t33 154.679
R23339 XThR.Tn[10].n54 XThR.Tn[10].t52 154.679
R23340 XThR.Tn[10].n50 XThR.Tn[10].t58 154.679
R23341 XThR.Tn[10].n49 XThR.Tn[10].t18 154.679
R23342 XThR.Tn[10].n45 XThR.Tn[10].t41 154.679
R23343 XThR.Tn[10].n44 XThR.Tn[10].t63 154.679
R23344 XThR.Tn[10].n40 XThR.Tn[10].t22 154.679
R23345 XThR.Tn[10].n39 XThR.Tn[10].t45 154.679
R23346 XThR.Tn[10].n35 XThR.Tn[10].t66 154.679
R23347 XThR.Tn[10].n34 XThR.Tn[10].t26 154.679
R23348 XThR.Tn[10].n30 XThR.Tn[10].t72 154.679
R23349 XThR.Tn[10].n29 XThR.Tn[10].t31 154.679
R23350 XThR.Tn[10].n25 XThR.Tn[10].t55 154.679
R23351 XThR.Tn[10].n24 XThR.Tn[10].t14 154.679
R23352 XThR.Tn[10].n20 XThR.Tn[10].t30 154.679
R23353 XThR.Tn[10].n19 XThR.Tn[10].t50 154.679
R23354 XThR.Tn[10].n15 XThR.Tn[10].t53 154.679
R23355 XThR.Tn[10].n14 XThR.Tn[10].t12 154.679
R23356 XThR.Tn[10].n10 XThR.Tn[10].t37 154.679
R23357 XThR.Tn[10].n9 XThR.Tn[10].t60 154.679
R23358 XThR.Tn[10].n7 XThR.Tn[10].t20 154.679
R23359 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R23360 XThR.Tn[10].n3 XThR.Tn[10].t9 26.5955
R23361 XThR.Tn[10].n3 XThR.Tn[10].t11 26.5955
R23362 XThR.Tn[10].n4 XThR.Tn[10].t1 26.5955
R23363 XThR.Tn[10].n4 XThR.Tn[10].t10 26.5955
R23364 XThR.Tn[10].n0 XThR.Tn[10].t7 26.5955
R23365 XThR.Tn[10].n0 XThR.Tn[10].t5 26.5955
R23366 XThR.Tn[10].n1 XThR.Tn[10].t8 26.5955
R23367 XThR.Tn[10].n1 XThR.Tn[10].t6 26.5955
R23368 XThR.Tn[10].n86 XThR.Tn[10].t2 24.9236
R23369 XThR.Tn[10].n86 XThR.Tn[10].t4 24.9236
R23370 XThR.Tn[10].n87 XThR.Tn[10].t3 24.9236
R23371 XThR.Tn[10].n87 XThR.Tn[10].t0 24.9236
R23372 XThR.Tn[10] XThR.Tn[10].n88 18.8943
R23373 XThR.Tn[10].n6 XThR.Tn[10].n5 13.5534
R23374 XThR.Tn[10].n85 XThR.Tn[10] 7.84567
R23375 XThR.Tn[10] XThR.Tn[10].n85 6.34069
R23376 XThR.Tn[10] XThR.Tn[10].n8 5.34871
R23377 XThR.Tn[10].n13 XThR.Tn[10].n12 4.5005
R23378 XThR.Tn[10].n18 XThR.Tn[10].n17 4.5005
R23379 XThR.Tn[10].n23 XThR.Tn[10].n22 4.5005
R23380 XThR.Tn[10].n28 XThR.Tn[10].n27 4.5005
R23381 XThR.Tn[10].n33 XThR.Tn[10].n32 4.5005
R23382 XThR.Tn[10].n38 XThR.Tn[10].n37 4.5005
R23383 XThR.Tn[10].n43 XThR.Tn[10].n42 4.5005
R23384 XThR.Tn[10].n48 XThR.Tn[10].n47 4.5005
R23385 XThR.Tn[10].n53 XThR.Tn[10].n52 4.5005
R23386 XThR.Tn[10].n58 XThR.Tn[10].n57 4.5005
R23387 XThR.Tn[10].n63 XThR.Tn[10].n62 4.5005
R23388 XThR.Tn[10].n68 XThR.Tn[10].n67 4.5005
R23389 XThR.Tn[10].n73 XThR.Tn[10].n72 4.5005
R23390 XThR.Tn[10].n78 XThR.Tn[10].n77 4.5005
R23391 XThR.Tn[10].n83 XThR.Tn[10].n82 4.5005
R23392 XThR.Tn[10].n84 XThR.Tn[10] 3.70586
R23393 XThR.Tn[10].n13 XThR.Tn[10] 2.51836
R23394 XThR.Tn[10].n18 XThR.Tn[10] 2.51836
R23395 XThR.Tn[10].n23 XThR.Tn[10] 2.51836
R23396 XThR.Tn[10].n28 XThR.Tn[10] 2.51836
R23397 XThR.Tn[10].n33 XThR.Tn[10] 2.51836
R23398 XThR.Tn[10].n38 XThR.Tn[10] 2.51836
R23399 XThR.Tn[10].n43 XThR.Tn[10] 2.51836
R23400 XThR.Tn[10].n48 XThR.Tn[10] 2.51836
R23401 XThR.Tn[10].n53 XThR.Tn[10] 2.51836
R23402 XThR.Tn[10].n58 XThR.Tn[10] 2.51836
R23403 XThR.Tn[10].n63 XThR.Tn[10] 2.51836
R23404 XThR.Tn[10].n68 XThR.Tn[10] 2.51836
R23405 XThR.Tn[10].n73 XThR.Tn[10] 2.51836
R23406 XThR.Tn[10].n78 XThR.Tn[10] 2.51836
R23407 XThR.Tn[10].n83 XThR.Tn[10] 2.51836
R23408 XThR.Tn[10].n85 XThR.Tn[10] 1.79489
R23409 XThR.Tn[10].n6 XThR.Tn[10] 1.50638
R23410 XThR.Tn[10] XThR.Tn[10].n6 1.19676
R23411 XThR.Tn[10] XThR.Tn[10].n13 0.848714
R23412 XThR.Tn[10] XThR.Tn[10].n18 0.848714
R23413 XThR.Tn[10] XThR.Tn[10].n23 0.848714
R23414 XThR.Tn[10] XThR.Tn[10].n28 0.848714
R23415 XThR.Tn[10] XThR.Tn[10].n33 0.848714
R23416 XThR.Tn[10] XThR.Tn[10].n38 0.848714
R23417 XThR.Tn[10] XThR.Tn[10].n43 0.848714
R23418 XThR.Tn[10] XThR.Tn[10].n48 0.848714
R23419 XThR.Tn[10] XThR.Tn[10].n53 0.848714
R23420 XThR.Tn[10] XThR.Tn[10].n58 0.848714
R23421 XThR.Tn[10] XThR.Tn[10].n63 0.848714
R23422 XThR.Tn[10] XThR.Tn[10].n68 0.848714
R23423 XThR.Tn[10] XThR.Tn[10].n73 0.848714
R23424 XThR.Tn[10] XThR.Tn[10].n78 0.848714
R23425 XThR.Tn[10] XThR.Tn[10].n83 0.848714
R23426 XThR.Tn[10].n8 XThR.Tn[10] 0.485653
R23427 XThR.Tn[10].n81 XThR.Tn[10] 0.21482
R23428 XThR.Tn[10].n76 XThR.Tn[10] 0.21482
R23429 XThR.Tn[10].n71 XThR.Tn[10] 0.21482
R23430 XThR.Tn[10].n66 XThR.Tn[10] 0.21482
R23431 XThR.Tn[10].n61 XThR.Tn[10] 0.21482
R23432 XThR.Tn[10].n56 XThR.Tn[10] 0.21482
R23433 XThR.Tn[10].n51 XThR.Tn[10] 0.21482
R23434 XThR.Tn[10].n46 XThR.Tn[10] 0.21482
R23435 XThR.Tn[10].n41 XThR.Tn[10] 0.21482
R23436 XThR.Tn[10].n36 XThR.Tn[10] 0.21482
R23437 XThR.Tn[10].n31 XThR.Tn[10] 0.21482
R23438 XThR.Tn[10].n26 XThR.Tn[10] 0.21482
R23439 XThR.Tn[10].n21 XThR.Tn[10] 0.21482
R23440 XThR.Tn[10].n16 XThR.Tn[10] 0.21482
R23441 XThR.Tn[10].n11 XThR.Tn[10] 0.21482
R23442 XThR.Tn[10].n82 XThR.Tn[10] 0.0608448
R23443 XThR.Tn[10].n77 XThR.Tn[10] 0.0608448
R23444 XThR.Tn[10].n72 XThR.Tn[10] 0.0608448
R23445 XThR.Tn[10].n67 XThR.Tn[10] 0.0608448
R23446 XThR.Tn[10].n62 XThR.Tn[10] 0.0608448
R23447 XThR.Tn[10].n57 XThR.Tn[10] 0.0608448
R23448 XThR.Tn[10].n52 XThR.Tn[10] 0.0608448
R23449 XThR.Tn[10].n47 XThR.Tn[10] 0.0608448
R23450 XThR.Tn[10].n42 XThR.Tn[10] 0.0608448
R23451 XThR.Tn[10].n37 XThR.Tn[10] 0.0608448
R23452 XThR.Tn[10].n32 XThR.Tn[10] 0.0608448
R23453 XThR.Tn[10].n27 XThR.Tn[10] 0.0608448
R23454 XThR.Tn[10].n22 XThR.Tn[10] 0.0608448
R23455 XThR.Tn[10].n17 XThR.Tn[10] 0.0608448
R23456 XThR.Tn[10].n12 XThR.Tn[10] 0.0608448
R23457 XThR.Tn[10].n84 XThR.Tn[10] 0.0540714
R23458 XThR.Tn[10] XThR.Tn[10].n84 0.038
R23459 XThR.Tn[10].n8 XThR.Tn[10] 0.00744444
R23460 XThR.Tn[10].n82 XThR.Tn[10].n81 0.00265517
R23461 XThR.Tn[10].n77 XThR.Tn[10].n76 0.00265517
R23462 XThR.Tn[10].n72 XThR.Tn[10].n71 0.00265517
R23463 XThR.Tn[10].n67 XThR.Tn[10].n66 0.00265517
R23464 XThR.Tn[10].n62 XThR.Tn[10].n61 0.00265517
R23465 XThR.Tn[10].n57 XThR.Tn[10].n56 0.00265517
R23466 XThR.Tn[10].n52 XThR.Tn[10].n51 0.00265517
R23467 XThR.Tn[10].n47 XThR.Tn[10].n46 0.00265517
R23468 XThR.Tn[10].n42 XThR.Tn[10].n41 0.00265517
R23469 XThR.Tn[10].n37 XThR.Tn[10].n36 0.00265517
R23470 XThR.Tn[10].n32 XThR.Tn[10].n31 0.00265517
R23471 XThR.Tn[10].n27 XThR.Tn[10].n26 0.00265517
R23472 XThR.Tn[10].n22 XThR.Tn[10].n21 0.00265517
R23473 XThR.Tn[10].n17 XThR.Tn[10].n16 0.00265517
R23474 XThR.Tn[10].n12 XThR.Tn[10].n11 0.00265517
R23475 XThC.Tn[9].n70 XThC.Tn[9].n69 265.341
R23476 XThC.Tn[9].n74 XThC.Tn[9].n72 243.68
R23477 XThC.Tn[9].n2 XThC.Tn[9].n0 241.847
R23478 XThC.Tn[9].n74 XThC.Tn[9].n73 205.28
R23479 XThC.Tn[9].n70 XThC.Tn[9].n68 202.094
R23480 XThC.Tn[9].n2 XThC.Tn[9].n1 185
R23481 XThC.Tn[9].n64 XThC.Tn[9].n62 161.365
R23482 XThC.Tn[9].n60 XThC.Tn[9].n58 161.365
R23483 XThC.Tn[9].n56 XThC.Tn[9].n54 161.365
R23484 XThC.Tn[9].n52 XThC.Tn[9].n50 161.365
R23485 XThC.Tn[9].n48 XThC.Tn[9].n46 161.365
R23486 XThC.Tn[9].n44 XThC.Tn[9].n42 161.365
R23487 XThC.Tn[9].n40 XThC.Tn[9].n38 161.365
R23488 XThC.Tn[9].n36 XThC.Tn[9].n34 161.365
R23489 XThC.Tn[9].n32 XThC.Tn[9].n30 161.365
R23490 XThC.Tn[9].n28 XThC.Tn[9].n26 161.365
R23491 XThC.Tn[9].n24 XThC.Tn[9].n22 161.365
R23492 XThC.Tn[9].n20 XThC.Tn[9].n18 161.365
R23493 XThC.Tn[9].n16 XThC.Tn[9].n14 161.365
R23494 XThC.Tn[9].n12 XThC.Tn[9].n10 161.365
R23495 XThC.Tn[9].n8 XThC.Tn[9].n6 161.365
R23496 XThC.Tn[9].n5 XThC.Tn[9].n3 161.365
R23497 XThC.Tn[9].n62 XThC.Tn[9].t39 161.106
R23498 XThC.Tn[9].n58 XThC.Tn[9].t19 161.106
R23499 XThC.Tn[9].n54 XThC.Tn[9].t17 161.106
R23500 XThC.Tn[9].n50 XThC.Tn[9].t15 161.106
R23501 XThC.Tn[9].n46 XThC.Tn[9].t29 161.106
R23502 XThC.Tn[9].n42 XThC.Tn[9].t27 161.106
R23503 XThC.Tn[9].n38 XThC.Tn[9].t14 161.106
R23504 XThC.Tn[9].n34 XThC.Tn[9].t37 161.106
R23505 XThC.Tn[9].n30 XThC.Tn[9].t36 161.106
R23506 XThC.Tn[9].n26 XThC.Tn[9].t25 161.106
R23507 XThC.Tn[9].n22 XThC.Tn[9].t12 161.106
R23508 XThC.Tn[9].n18 XThC.Tn[9].t35 161.106
R23509 XThC.Tn[9].n14 XThC.Tn[9].t23 161.106
R23510 XThC.Tn[9].n10 XThC.Tn[9].t22 161.106
R23511 XThC.Tn[9].n6 XThC.Tn[9].t42 161.106
R23512 XThC.Tn[9].n3 XThC.Tn[9].t33 161.106
R23513 XThC.Tn[9].n62 XThC.Tn[9].t13 154.679
R23514 XThC.Tn[9].n58 XThC.Tn[9].t26 154.679
R23515 XThC.Tn[9].n54 XThC.Tn[9].t24 154.679
R23516 XThC.Tn[9].n50 XThC.Tn[9].t21 154.679
R23517 XThC.Tn[9].n46 XThC.Tn[9].t34 154.679
R23518 XThC.Tn[9].n42 XThC.Tn[9].t32 154.679
R23519 XThC.Tn[9].n38 XThC.Tn[9].t20 154.679
R23520 XThC.Tn[9].n34 XThC.Tn[9].t43 154.679
R23521 XThC.Tn[9].n30 XThC.Tn[9].t41 154.679
R23522 XThC.Tn[9].n26 XThC.Tn[9].t31 154.679
R23523 XThC.Tn[9].n22 XThC.Tn[9].t18 154.679
R23524 XThC.Tn[9].n18 XThC.Tn[9].t40 154.679
R23525 XThC.Tn[9].n14 XThC.Tn[9].t30 154.679
R23526 XThC.Tn[9].n10 XThC.Tn[9].t28 154.679
R23527 XThC.Tn[9].n6 XThC.Tn[9].t16 154.679
R23528 XThC.Tn[9].n3 XThC.Tn[9].t38 154.679
R23529 XThC.Tn[9].n69 XThC.Tn[9].t2 26.5955
R23530 XThC.Tn[9].n69 XThC.Tn[9].t1 26.5955
R23531 XThC.Tn[9].n72 XThC.Tn[9].t9 26.5955
R23532 XThC.Tn[9].n72 XThC.Tn[9].t8 26.5955
R23533 XThC.Tn[9].n73 XThC.Tn[9].t11 26.5955
R23534 XThC.Tn[9].n73 XThC.Tn[9].t10 26.5955
R23535 XThC.Tn[9].n68 XThC.Tn[9].t0 26.5955
R23536 XThC.Tn[9].n68 XThC.Tn[9].t3 26.5955
R23537 XThC.Tn[9].n1 XThC.Tn[9].t6 24.9236
R23538 XThC.Tn[9].n1 XThC.Tn[9].t7 24.9236
R23539 XThC.Tn[9].n0 XThC.Tn[9].t5 24.9236
R23540 XThC.Tn[9].n0 XThC.Tn[9].t4 24.9236
R23541 XThC.Tn[9] XThC.Tn[9].n74 22.9652
R23542 XThC.Tn[9] XThC.Tn[9].n2 18.8943
R23543 XThC.Tn[9].n71 XThC.Tn[9].n70 13.9299
R23544 XThC.Tn[9] XThC.Tn[9].n71 13.9299
R23545 XThC.Tn[9] XThC.Tn[9].n5 8.0245
R23546 XThC.Tn[9].n65 XThC.Tn[9].n64 7.9105
R23547 XThC.Tn[9].n61 XThC.Tn[9].n60 7.9105
R23548 XThC.Tn[9].n57 XThC.Tn[9].n56 7.9105
R23549 XThC.Tn[9].n53 XThC.Tn[9].n52 7.9105
R23550 XThC.Tn[9].n49 XThC.Tn[9].n48 7.9105
R23551 XThC.Tn[9].n45 XThC.Tn[9].n44 7.9105
R23552 XThC.Tn[9].n41 XThC.Tn[9].n40 7.9105
R23553 XThC.Tn[9].n37 XThC.Tn[9].n36 7.9105
R23554 XThC.Tn[9].n33 XThC.Tn[9].n32 7.9105
R23555 XThC.Tn[9].n29 XThC.Tn[9].n28 7.9105
R23556 XThC.Tn[9].n25 XThC.Tn[9].n24 7.9105
R23557 XThC.Tn[9].n21 XThC.Tn[9].n20 7.9105
R23558 XThC.Tn[9].n17 XThC.Tn[9].n16 7.9105
R23559 XThC.Tn[9].n13 XThC.Tn[9].n12 7.9105
R23560 XThC.Tn[9].n9 XThC.Tn[9].n8 7.9105
R23561 XThC.Tn[9].n67 XThC.Tn[9].n66 7.44831
R23562 XThC.Tn[9].n67 XThC.Tn[9] 6.34069
R23563 XThC.Tn[9].n66 XThC.Tn[9] 4.25199
R23564 XThC.Tn[9] XThC.Tn[9].n67 1.79489
R23565 XThC.Tn[9].n71 XThC.Tn[9] 1.19676
R23566 XThC.Tn[9].n66 XThC.Tn[9] 0.657022
R23567 XThC.Tn[9].n9 XThC.Tn[9] 0.235138
R23568 XThC.Tn[9].n13 XThC.Tn[9] 0.235138
R23569 XThC.Tn[9].n17 XThC.Tn[9] 0.235138
R23570 XThC.Tn[9].n21 XThC.Tn[9] 0.235138
R23571 XThC.Tn[9].n25 XThC.Tn[9] 0.235138
R23572 XThC.Tn[9].n29 XThC.Tn[9] 0.235138
R23573 XThC.Tn[9].n33 XThC.Tn[9] 0.235138
R23574 XThC.Tn[9].n37 XThC.Tn[9] 0.235138
R23575 XThC.Tn[9].n41 XThC.Tn[9] 0.235138
R23576 XThC.Tn[9].n45 XThC.Tn[9] 0.235138
R23577 XThC.Tn[9].n49 XThC.Tn[9] 0.235138
R23578 XThC.Tn[9].n53 XThC.Tn[9] 0.235138
R23579 XThC.Tn[9].n57 XThC.Tn[9] 0.235138
R23580 XThC.Tn[9].n61 XThC.Tn[9] 0.235138
R23581 XThC.Tn[9].n65 XThC.Tn[9] 0.235138
R23582 XThC.Tn[9] XThC.Tn[9].n9 0.114505
R23583 XThC.Tn[9] XThC.Tn[9].n13 0.114505
R23584 XThC.Tn[9] XThC.Tn[9].n17 0.114505
R23585 XThC.Tn[9] XThC.Tn[9].n21 0.114505
R23586 XThC.Tn[9] XThC.Tn[9].n25 0.114505
R23587 XThC.Tn[9] XThC.Tn[9].n29 0.114505
R23588 XThC.Tn[9] XThC.Tn[9].n33 0.114505
R23589 XThC.Tn[9] XThC.Tn[9].n37 0.114505
R23590 XThC.Tn[9] XThC.Tn[9].n41 0.114505
R23591 XThC.Tn[9] XThC.Tn[9].n45 0.114505
R23592 XThC.Tn[9] XThC.Tn[9].n49 0.114505
R23593 XThC.Tn[9] XThC.Tn[9].n53 0.114505
R23594 XThC.Tn[9] XThC.Tn[9].n57 0.114505
R23595 XThC.Tn[9] XThC.Tn[9].n61 0.114505
R23596 XThC.Tn[9] XThC.Tn[9].n65 0.114505
R23597 XThC.Tn[9].n64 XThC.Tn[9].n63 0.0599512
R23598 XThC.Tn[9].n60 XThC.Tn[9].n59 0.0599512
R23599 XThC.Tn[9].n56 XThC.Tn[9].n55 0.0599512
R23600 XThC.Tn[9].n52 XThC.Tn[9].n51 0.0599512
R23601 XThC.Tn[9].n48 XThC.Tn[9].n47 0.0599512
R23602 XThC.Tn[9].n44 XThC.Tn[9].n43 0.0599512
R23603 XThC.Tn[9].n40 XThC.Tn[9].n39 0.0599512
R23604 XThC.Tn[9].n36 XThC.Tn[9].n35 0.0599512
R23605 XThC.Tn[9].n32 XThC.Tn[9].n31 0.0599512
R23606 XThC.Tn[9].n28 XThC.Tn[9].n27 0.0599512
R23607 XThC.Tn[9].n24 XThC.Tn[9].n23 0.0599512
R23608 XThC.Tn[9].n20 XThC.Tn[9].n19 0.0599512
R23609 XThC.Tn[9].n16 XThC.Tn[9].n15 0.0599512
R23610 XThC.Tn[9].n12 XThC.Tn[9].n11 0.0599512
R23611 XThC.Tn[9].n8 XThC.Tn[9].n7 0.0599512
R23612 XThC.Tn[9].n5 XThC.Tn[9].n4 0.0599512
R23613 XThC.Tn[9].n63 XThC.Tn[9] 0.0469286
R23614 XThC.Tn[9].n59 XThC.Tn[9] 0.0469286
R23615 XThC.Tn[9].n55 XThC.Tn[9] 0.0469286
R23616 XThC.Tn[9].n51 XThC.Tn[9] 0.0469286
R23617 XThC.Tn[9].n47 XThC.Tn[9] 0.0469286
R23618 XThC.Tn[9].n43 XThC.Tn[9] 0.0469286
R23619 XThC.Tn[9].n39 XThC.Tn[9] 0.0469286
R23620 XThC.Tn[9].n35 XThC.Tn[9] 0.0469286
R23621 XThC.Tn[9].n31 XThC.Tn[9] 0.0469286
R23622 XThC.Tn[9].n27 XThC.Tn[9] 0.0469286
R23623 XThC.Tn[9].n23 XThC.Tn[9] 0.0469286
R23624 XThC.Tn[9].n19 XThC.Tn[9] 0.0469286
R23625 XThC.Tn[9].n15 XThC.Tn[9] 0.0469286
R23626 XThC.Tn[9].n11 XThC.Tn[9] 0.0469286
R23627 XThC.Tn[9].n7 XThC.Tn[9] 0.0469286
R23628 XThC.Tn[9].n4 XThC.Tn[9] 0.0469286
R23629 XThC.Tn[9].n63 XThC.Tn[9] 0.0401341
R23630 XThC.Tn[9].n59 XThC.Tn[9] 0.0401341
R23631 XThC.Tn[9].n55 XThC.Tn[9] 0.0401341
R23632 XThC.Tn[9].n51 XThC.Tn[9] 0.0401341
R23633 XThC.Tn[9].n47 XThC.Tn[9] 0.0401341
R23634 XThC.Tn[9].n43 XThC.Tn[9] 0.0401341
R23635 XThC.Tn[9].n39 XThC.Tn[9] 0.0401341
R23636 XThC.Tn[9].n35 XThC.Tn[9] 0.0401341
R23637 XThC.Tn[9].n31 XThC.Tn[9] 0.0401341
R23638 XThC.Tn[9].n27 XThC.Tn[9] 0.0401341
R23639 XThC.Tn[9].n23 XThC.Tn[9] 0.0401341
R23640 XThC.Tn[9].n19 XThC.Tn[9] 0.0401341
R23641 XThC.Tn[9].n15 XThC.Tn[9] 0.0401341
R23642 XThC.Tn[9].n11 XThC.Tn[9] 0.0401341
R23643 XThC.Tn[9].n7 XThC.Tn[9] 0.0401341
R23644 XThC.Tn[9].n4 XThC.Tn[9] 0.0401341
R23645 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R23646 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R23647 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R23648 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R23649 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R23650 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R23651 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R23652 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R23653 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R23654 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R23655 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R23656 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R23657 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R23658 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R23659 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R23660 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R23661 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R23662 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R23663 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R23664 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R23665 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R23666 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R23667 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R23668 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R23669 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R23670 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R23671 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R23672 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R23673 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R23674 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R23675 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R23676 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R23677 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R23678 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R23679 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R23680 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R23681 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R23682 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R23683 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R23684 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R23685 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R23686 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R23687 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R23688 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R23689 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R23690 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R23691 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R23692 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R23693 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R23694 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R23695 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R23696 data[4].n3 data[4].t0 231.835
R23697 data[4].n0 data[4].t3 230.155
R23698 data[4].n0 data[4].t1 157.856
R23699 data[4].n3 data[4].t2 157.07
R23700 data[4].n1 data[4].n0 152
R23701 data[4].n4 data[4].n3 152
R23702 data[4].n2 data[4].n1 25.6681
R23703 data[4].n4 data[4].n2 10.7642
R23704 data[4].n2 data[4] 2.763
R23705 data[4].n1 data[4] 2.10199
R23706 data[4] data[4].n4 2.01193
R23707 XThC.Tn[11].n70 XThC.Tn[11].n69 265.341
R23708 XThC.Tn[11].n74 XThC.Tn[11].n72 243.68
R23709 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R23710 XThC.Tn[11].n74 XThC.Tn[11].n73 205.28
R23711 XThC.Tn[11].n70 XThC.Tn[11].n68 202.094
R23712 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R23713 XThC.Tn[11].n64 XThC.Tn[11].n62 161.365
R23714 XThC.Tn[11].n60 XThC.Tn[11].n58 161.365
R23715 XThC.Tn[11].n56 XThC.Tn[11].n54 161.365
R23716 XThC.Tn[11].n52 XThC.Tn[11].n50 161.365
R23717 XThC.Tn[11].n48 XThC.Tn[11].n46 161.365
R23718 XThC.Tn[11].n44 XThC.Tn[11].n42 161.365
R23719 XThC.Tn[11].n40 XThC.Tn[11].n38 161.365
R23720 XThC.Tn[11].n36 XThC.Tn[11].n34 161.365
R23721 XThC.Tn[11].n32 XThC.Tn[11].n30 161.365
R23722 XThC.Tn[11].n28 XThC.Tn[11].n26 161.365
R23723 XThC.Tn[11].n24 XThC.Tn[11].n22 161.365
R23724 XThC.Tn[11].n20 XThC.Tn[11].n18 161.365
R23725 XThC.Tn[11].n16 XThC.Tn[11].n14 161.365
R23726 XThC.Tn[11].n12 XThC.Tn[11].n10 161.365
R23727 XThC.Tn[11].n8 XThC.Tn[11].n6 161.365
R23728 XThC.Tn[11].n5 XThC.Tn[11].n3 161.365
R23729 XThC.Tn[11].n62 XThC.Tn[11].t12 161.106
R23730 XThC.Tn[11].n58 XThC.Tn[11].t26 161.106
R23731 XThC.Tn[11].n54 XThC.Tn[11].t23 161.106
R23732 XThC.Tn[11].n50 XThC.Tn[11].t21 161.106
R23733 XThC.Tn[11].n46 XThC.Tn[11].t34 161.106
R23734 XThC.Tn[11].n42 XThC.Tn[11].t32 161.106
R23735 XThC.Tn[11].n38 XThC.Tn[11].t20 161.106
R23736 XThC.Tn[11].n34 XThC.Tn[11].t43 161.106
R23737 XThC.Tn[11].n30 XThC.Tn[11].t41 161.106
R23738 XThC.Tn[11].n26 XThC.Tn[11].t31 161.106
R23739 XThC.Tn[11].n22 XThC.Tn[11].t18 161.106
R23740 XThC.Tn[11].n18 XThC.Tn[11].t39 161.106
R23741 XThC.Tn[11].n14 XThC.Tn[11].t30 161.106
R23742 XThC.Tn[11].n10 XThC.Tn[11].t28 161.106
R23743 XThC.Tn[11].n6 XThC.Tn[11].t15 161.106
R23744 XThC.Tn[11].n3 XThC.Tn[11].t38 161.106
R23745 XThC.Tn[11].n62 XThC.Tn[11].t40 154.679
R23746 XThC.Tn[11].n58 XThC.Tn[11].t19 154.679
R23747 XThC.Tn[11].n54 XThC.Tn[11].t17 154.679
R23748 XThC.Tn[11].n50 XThC.Tn[11].t16 154.679
R23749 XThC.Tn[11].n46 XThC.Tn[11].t29 154.679
R23750 XThC.Tn[11].n42 XThC.Tn[11].t27 154.679
R23751 XThC.Tn[11].n38 XThC.Tn[11].t14 154.679
R23752 XThC.Tn[11].n34 XThC.Tn[11].t37 154.679
R23753 XThC.Tn[11].n30 XThC.Tn[11].t36 154.679
R23754 XThC.Tn[11].n26 XThC.Tn[11].t25 154.679
R23755 XThC.Tn[11].n22 XThC.Tn[11].t13 154.679
R23756 XThC.Tn[11].n18 XThC.Tn[11].t35 154.679
R23757 XThC.Tn[11].n14 XThC.Tn[11].t24 154.679
R23758 XThC.Tn[11].n10 XThC.Tn[11].t22 154.679
R23759 XThC.Tn[11].n6 XThC.Tn[11].t42 154.679
R23760 XThC.Tn[11].n3 XThC.Tn[11].t33 154.679
R23761 XThC.Tn[11].n68 XThC.Tn[11].t1 26.5955
R23762 XThC.Tn[11].n68 XThC.Tn[11].t2 26.5955
R23763 XThC.Tn[11].n72 XThC.Tn[11].t8 26.5955
R23764 XThC.Tn[11].n72 XThC.Tn[11].t11 26.5955
R23765 XThC.Tn[11].n73 XThC.Tn[11].t10 26.5955
R23766 XThC.Tn[11].n73 XThC.Tn[11].t9 26.5955
R23767 XThC.Tn[11].n69 XThC.Tn[11].t0 26.5955
R23768 XThC.Tn[11].n69 XThC.Tn[11].t3 26.5955
R23769 XThC.Tn[11].n1 XThC.Tn[11].t4 24.9236
R23770 XThC.Tn[11].n1 XThC.Tn[11].t5 24.9236
R23771 XThC.Tn[11].n0 XThC.Tn[11].t7 24.9236
R23772 XThC.Tn[11].n0 XThC.Tn[11].t6 24.9236
R23773 XThC.Tn[11] XThC.Tn[11].n74 22.9652
R23774 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R23775 XThC.Tn[11].n71 XThC.Tn[11].n70 13.9299
R23776 XThC.Tn[11] XThC.Tn[11].n71 13.9299
R23777 XThC.Tn[11] XThC.Tn[11].n5 8.0245
R23778 XThC.Tn[11].n65 XThC.Tn[11].n64 7.9105
R23779 XThC.Tn[11].n61 XThC.Tn[11].n60 7.9105
R23780 XThC.Tn[11].n57 XThC.Tn[11].n56 7.9105
R23781 XThC.Tn[11].n53 XThC.Tn[11].n52 7.9105
R23782 XThC.Tn[11].n49 XThC.Tn[11].n48 7.9105
R23783 XThC.Tn[11].n45 XThC.Tn[11].n44 7.9105
R23784 XThC.Tn[11].n41 XThC.Tn[11].n40 7.9105
R23785 XThC.Tn[11].n37 XThC.Tn[11].n36 7.9105
R23786 XThC.Tn[11].n33 XThC.Tn[11].n32 7.9105
R23787 XThC.Tn[11].n29 XThC.Tn[11].n28 7.9105
R23788 XThC.Tn[11].n25 XThC.Tn[11].n24 7.9105
R23789 XThC.Tn[11].n21 XThC.Tn[11].n20 7.9105
R23790 XThC.Tn[11].n17 XThC.Tn[11].n16 7.9105
R23791 XThC.Tn[11].n13 XThC.Tn[11].n12 7.9105
R23792 XThC.Tn[11].n9 XThC.Tn[11].n8 7.9105
R23793 XThC.Tn[11].n67 XThC.Tn[11].n66 7.44831
R23794 XThC.Tn[11].n67 XThC.Tn[11] 6.34069
R23795 XThC.Tn[11].n66 XThC.Tn[11] 4.37928
R23796 XThC.Tn[11] XThC.Tn[11].n67 1.79489
R23797 XThC.Tn[11].n71 XThC.Tn[11] 1.19676
R23798 XThC.Tn[11].n66 XThC.Tn[11] 1.0918
R23799 XThC.Tn[11].n9 XThC.Tn[11] 0.235138
R23800 XThC.Tn[11].n13 XThC.Tn[11] 0.235138
R23801 XThC.Tn[11].n17 XThC.Tn[11] 0.235138
R23802 XThC.Tn[11].n21 XThC.Tn[11] 0.235138
R23803 XThC.Tn[11].n25 XThC.Tn[11] 0.235138
R23804 XThC.Tn[11].n29 XThC.Tn[11] 0.235138
R23805 XThC.Tn[11].n33 XThC.Tn[11] 0.235138
R23806 XThC.Tn[11].n37 XThC.Tn[11] 0.235138
R23807 XThC.Tn[11].n41 XThC.Tn[11] 0.235138
R23808 XThC.Tn[11].n45 XThC.Tn[11] 0.235138
R23809 XThC.Tn[11].n49 XThC.Tn[11] 0.235138
R23810 XThC.Tn[11].n53 XThC.Tn[11] 0.235138
R23811 XThC.Tn[11].n57 XThC.Tn[11] 0.235138
R23812 XThC.Tn[11].n61 XThC.Tn[11] 0.235138
R23813 XThC.Tn[11].n65 XThC.Tn[11] 0.235138
R23814 XThC.Tn[11] XThC.Tn[11].n9 0.114505
R23815 XThC.Tn[11] XThC.Tn[11].n13 0.114505
R23816 XThC.Tn[11] XThC.Tn[11].n17 0.114505
R23817 XThC.Tn[11] XThC.Tn[11].n21 0.114505
R23818 XThC.Tn[11] XThC.Tn[11].n25 0.114505
R23819 XThC.Tn[11] XThC.Tn[11].n29 0.114505
R23820 XThC.Tn[11] XThC.Tn[11].n33 0.114505
R23821 XThC.Tn[11] XThC.Tn[11].n37 0.114505
R23822 XThC.Tn[11] XThC.Tn[11].n41 0.114505
R23823 XThC.Tn[11] XThC.Tn[11].n45 0.114505
R23824 XThC.Tn[11] XThC.Tn[11].n49 0.114505
R23825 XThC.Tn[11] XThC.Tn[11].n53 0.114505
R23826 XThC.Tn[11] XThC.Tn[11].n57 0.114505
R23827 XThC.Tn[11] XThC.Tn[11].n61 0.114505
R23828 XThC.Tn[11] XThC.Tn[11].n65 0.114505
R23829 XThC.Tn[11].n64 XThC.Tn[11].n63 0.0599512
R23830 XThC.Tn[11].n60 XThC.Tn[11].n59 0.0599512
R23831 XThC.Tn[11].n56 XThC.Tn[11].n55 0.0599512
R23832 XThC.Tn[11].n52 XThC.Tn[11].n51 0.0599512
R23833 XThC.Tn[11].n48 XThC.Tn[11].n47 0.0599512
R23834 XThC.Tn[11].n44 XThC.Tn[11].n43 0.0599512
R23835 XThC.Tn[11].n40 XThC.Tn[11].n39 0.0599512
R23836 XThC.Tn[11].n36 XThC.Tn[11].n35 0.0599512
R23837 XThC.Tn[11].n32 XThC.Tn[11].n31 0.0599512
R23838 XThC.Tn[11].n28 XThC.Tn[11].n27 0.0599512
R23839 XThC.Tn[11].n24 XThC.Tn[11].n23 0.0599512
R23840 XThC.Tn[11].n20 XThC.Tn[11].n19 0.0599512
R23841 XThC.Tn[11].n16 XThC.Tn[11].n15 0.0599512
R23842 XThC.Tn[11].n12 XThC.Tn[11].n11 0.0599512
R23843 XThC.Tn[11].n8 XThC.Tn[11].n7 0.0599512
R23844 XThC.Tn[11].n5 XThC.Tn[11].n4 0.0599512
R23845 XThC.Tn[11].n63 XThC.Tn[11] 0.0469286
R23846 XThC.Tn[11].n59 XThC.Tn[11] 0.0469286
R23847 XThC.Tn[11].n55 XThC.Tn[11] 0.0469286
R23848 XThC.Tn[11].n51 XThC.Tn[11] 0.0469286
R23849 XThC.Tn[11].n47 XThC.Tn[11] 0.0469286
R23850 XThC.Tn[11].n43 XThC.Tn[11] 0.0469286
R23851 XThC.Tn[11].n39 XThC.Tn[11] 0.0469286
R23852 XThC.Tn[11].n35 XThC.Tn[11] 0.0469286
R23853 XThC.Tn[11].n31 XThC.Tn[11] 0.0469286
R23854 XThC.Tn[11].n27 XThC.Tn[11] 0.0469286
R23855 XThC.Tn[11].n23 XThC.Tn[11] 0.0469286
R23856 XThC.Tn[11].n19 XThC.Tn[11] 0.0469286
R23857 XThC.Tn[11].n15 XThC.Tn[11] 0.0469286
R23858 XThC.Tn[11].n11 XThC.Tn[11] 0.0469286
R23859 XThC.Tn[11].n7 XThC.Tn[11] 0.0469286
R23860 XThC.Tn[11].n4 XThC.Tn[11] 0.0469286
R23861 XThC.Tn[11].n63 XThC.Tn[11] 0.0401341
R23862 XThC.Tn[11].n59 XThC.Tn[11] 0.0401341
R23863 XThC.Tn[11].n55 XThC.Tn[11] 0.0401341
R23864 XThC.Tn[11].n51 XThC.Tn[11] 0.0401341
R23865 XThC.Tn[11].n47 XThC.Tn[11] 0.0401341
R23866 XThC.Tn[11].n43 XThC.Tn[11] 0.0401341
R23867 XThC.Tn[11].n39 XThC.Tn[11] 0.0401341
R23868 XThC.Tn[11].n35 XThC.Tn[11] 0.0401341
R23869 XThC.Tn[11].n31 XThC.Tn[11] 0.0401341
R23870 XThC.Tn[11].n27 XThC.Tn[11] 0.0401341
R23871 XThC.Tn[11].n23 XThC.Tn[11] 0.0401341
R23872 XThC.Tn[11].n19 XThC.Tn[11] 0.0401341
R23873 XThC.Tn[11].n15 XThC.Tn[11] 0.0401341
R23874 XThC.Tn[11].n11 XThC.Tn[11] 0.0401341
R23875 XThC.Tn[11].n7 XThC.Tn[11] 0.0401341
R23876 XThC.Tn[11].n4 XThC.Tn[11] 0.0401341
R23877 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R23878 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R23879 XThR.Tn[3] XThR.Tn[3].n82 161.363
R23880 XThR.Tn[3] XThR.Tn[3].n77 161.363
R23881 XThR.Tn[3] XThR.Tn[3].n72 161.363
R23882 XThR.Tn[3] XThR.Tn[3].n67 161.363
R23883 XThR.Tn[3] XThR.Tn[3].n62 161.363
R23884 XThR.Tn[3] XThR.Tn[3].n57 161.363
R23885 XThR.Tn[3] XThR.Tn[3].n52 161.363
R23886 XThR.Tn[3] XThR.Tn[3].n47 161.363
R23887 XThR.Tn[3] XThR.Tn[3].n42 161.363
R23888 XThR.Tn[3] XThR.Tn[3].n37 161.363
R23889 XThR.Tn[3] XThR.Tn[3].n32 161.363
R23890 XThR.Tn[3] XThR.Tn[3].n27 161.363
R23891 XThR.Tn[3] XThR.Tn[3].n22 161.363
R23892 XThR.Tn[3] XThR.Tn[3].n17 161.363
R23893 XThR.Tn[3] XThR.Tn[3].n12 161.363
R23894 XThR.Tn[3] XThR.Tn[3].n10 161.363
R23895 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R23896 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R23897 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R23898 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R23899 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R23900 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R23901 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R23902 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R23903 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R23904 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R23905 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R23906 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R23907 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R23908 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R23909 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R23910 XThR.Tn[3].n83 XThR.Tn[3].t65 161.106
R23911 XThR.Tn[3].n82 XThR.Tn[3].t37 161.106
R23912 XThR.Tn[3].n78 XThR.Tn[3].t70 161.106
R23913 XThR.Tn[3].n77 XThR.Tn[3].t46 161.106
R23914 XThR.Tn[3].n73 XThR.Tn[3].t53 161.106
R23915 XThR.Tn[3].n72 XThR.Tn[3].t29 161.106
R23916 XThR.Tn[3].n68 XThR.Tn[3].t35 161.106
R23917 XThR.Tn[3].n67 XThR.Tn[3].t73 161.106
R23918 XThR.Tn[3].n63 XThR.Tn[3].t64 161.106
R23919 XThR.Tn[3].n62 XThR.Tn[3].t36 161.106
R23920 XThR.Tn[3].n58 XThR.Tn[3].t24 161.106
R23921 XThR.Tn[3].n57 XThR.Tn[3].t62 161.106
R23922 XThR.Tn[3].n53 XThR.Tn[3].t68 161.106
R23923 XThR.Tn[3].n52 XThR.Tn[3].t44 161.106
R23924 XThR.Tn[3].n48 XThR.Tn[3].t50 161.106
R23925 XThR.Tn[3].n47 XThR.Tn[3].t26 161.106
R23926 XThR.Tn[3].n43 XThR.Tn[3].t33 161.106
R23927 XThR.Tn[3].n42 XThR.Tn[3].t71 161.106
R23928 XThR.Tn[3].n38 XThR.Tn[3].t39 161.106
R23929 XThR.Tn[3].n37 XThR.Tn[3].t14 161.106
R23930 XThR.Tn[3].n33 XThR.Tn[3].t23 161.106
R23931 XThR.Tn[3].n32 XThR.Tn[3].t61 161.106
R23932 XThR.Tn[3].n28 XThR.Tn[3].t52 161.106
R23933 XThR.Tn[3].n27 XThR.Tn[3].t28 161.106
R23934 XThR.Tn[3].n23 XThR.Tn[3].t21 161.106
R23935 XThR.Tn[3].n22 XThR.Tn[3].t57 161.106
R23936 XThR.Tn[3].n18 XThR.Tn[3].t67 161.106
R23937 XThR.Tn[3].n17 XThR.Tn[3].t40 161.106
R23938 XThR.Tn[3].n13 XThR.Tn[3].t31 161.106
R23939 XThR.Tn[3].n12 XThR.Tn[3].t66 161.106
R23940 XThR.Tn[3].n10 XThR.Tn[3].t48 161.106
R23941 XThR.Tn[3].n83 XThR.Tn[3].t19 154.679
R23942 XThR.Tn[3].n82 XThR.Tn[3].t56 154.679
R23943 XThR.Tn[3].n78 XThR.Tn[3].t59 154.679
R23944 XThR.Tn[3].n77 XThR.Tn[3].t34 154.679
R23945 XThR.Tn[3].n73 XThR.Tn[3].t42 154.679
R23946 XThR.Tn[3].n72 XThR.Tn[3].t16 154.679
R23947 XThR.Tn[3].n68 XThR.Tn[3].t72 154.679
R23948 XThR.Tn[3].n67 XThR.Tn[3].t47 154.679
R23949 XThR.Tn[3].n63 XThR.Tn[3].t54 154.679
R23950 XThR.Tn[3].n62 XThR.Tn[3].t30 154.679
R23951 XThR.Tn[3].n58 XThR.Tn[3].t18 154.679
R23952 XThR.Tn[3].n57 XThR.Tn[3].t55 154.679
R23953 XThR.Tn[3].n53 XThR.Tn[3].t43 154.679
R23954 XThR.Tn[3].n52 XThR.Tn[3].t17 154.679
R23955 XThR.Tn[3].n48 XThR.Tn[3].t25 154.679
R23956 XThR.Tn[3].n47 XThR.Tn[3].t63 154.679
R23957 XThR.Tn[3].n43 XThR.Tn[3].t69 154.679
R23958 XThR.Tn[3].n42 XThR.Tn[3].t45 154.679
R23959 XThR.Tn[3].n38 XThR.Tn[3].t51 154.679
R23960 XThR.Tn[3].n37 XThR.Tn[3].t27 154.679
R23961 XThR.Tn[3].n33 XThR.Tn[3].t58 154.679
R23962 XThR.Tn[3].n32 XThR.Tn[3].t32 154.679
R23963 XThR.Tn[3].n28 XThR.Tn[3].t41 154.679
R23964 XThR.Tn[3].n27 XThR.Tn[3].t15 154.679
R23965 XThR.Tn[3].n23 XThR.Tn[3].t12 154.679
R23966 XThR.Tn[3].n22 XThR.Tn[3].t49 154.679
R23967 XThR.Tn[3].n18 XThR.Tn[3].t38 154.679
R23968 XThR.Tn[3].n17 XThR.Tn[3].t13 154.679
R23969 XThR.Tn[3].n13 XThR.Tn[3].t22 154.679
R23970 XThR.Tn[3].n12 XThR.Tn[3].t60 154.679
R23971 XThR.Tn[3].n10 XThR.Tn[3].t20 154.679
R23972 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R23973 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R23974 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R23975 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R23976 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R23977 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R23978 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R23979 XThR.Tn[3].n1 XThR.Tn[3].t4 26.5955
R23980 XThR.Tn[3].n1 XThR.Tn[3].t7 26.5955
R23981 XThR.Tn[3].n0 XThR.Tn[3].t5 26.5955
R23982 XThR.Tn[3].n0 XThR.Tn[3].t6 26.5955
R23983 XThR.Tn[3].n3 XThR.Tn[3].t11 24.9236
R23984 XThR.Tn[3].n3 XThR.Tn[3].t8 24.9236
R23985 XThR.Tn[3].n4 XThR.Tn[3].t10 24.9236
R23986 XThR.Tn[3].n4 XThR.Tn[3].t9 24.9236
R23987 XThR.Tn[3].n5 XThR.Tn[3].t2 24.9236
R23988 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R23989 XThR.Tn[3].n6 XThR.Tn[3].t3 24.9236
R23990 XThR.Tn[3].n6 XThR.Tn[3].t0 24.9236
R23991 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R23992 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R23993 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R23994 XThR.Tn[3] XThR.Tn[3].n11 5.34871
R23995 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R23996 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R23997 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R23998 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R23999 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R24000 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R24001 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R24002 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R24003 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R24004 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R24005 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R24006 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R24007 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R24008 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R24009 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R24010 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R24011 XThR.Tn[3].n16 XThR.Tn[3] 2.51836
R24012 XThR.Tn[3].n21 XThR.Tn[3] 2.51836
R24013 XThR.Tn[3].n26 XThR.Tn[3] 2.51836
R24014 XThR.Tn[3].n31 XThR.Tn[3] 2.51836
R24015 XThR.Tn[3].n36 XThR.Tn[3] 2.51836
R24016 XThR.Tn[3].n41 XThR.Tn[3] 2.51836
R24017 XThR.Tn[3].n46 XThR.Tn[3] 2.51836
R24018 XThR.Tn[3].n51 XThR.Tn[3] 2.51836
R24019 XThR.Tn[3].n56 XThR.Tn[3] 2.51836
R24020 XThR.Tn[3].n61 XThR.Tn[3] 2.51836
R24021 XThR.Tn[3].n66 XThR.Tn[3] 2.51836
R24022 XThR.Tn[3].n71 XThR.Tn[3] 2.51836
R24023 XThR.Tn[3].n76 XThR.Tn[3] 2.51836
R24024 XThR.Tn[3].n81 XThR.Tn[3] 2.51836
R24025 XThR.Tn[3].n86 XThR.Tn[3] 2.51836
R24026 XThR.Tn[3] XThR.Tn[3].n16 0.848714
R24027 XThR.Tn[3] XThR.Tn[3].n21 0.848714
R24028 XThR.Tn[3] XThR.Tn[3].n26 0.848714
R24029 XThR.Tn[3] XThR.Tn[3].n31 0.848714
R24030 XThR.Tn[3] XThR.Tn[3].n36 0.848714
R24031 XThR.Tn[3] XThR.Tn[3].n41 0.848714
R24032 XThR.Tn[3] XThR.Tn[3].n46 0.848714
R24033 XThR.Tn[3] XThR.Tn[3].n51 0.848714
R24034 XThR.Tn[3] XThR.Tn[3].n56 0.848714
R24035 XThR.Tn[3] XThR.Tn[3].n61 0.848714
R24036 XThR.Tn[3] XThR.Tn[3].n66 0.848714
R24037 XThR.Tn[3] XThR.Tn[3].n71 0.848714
R24038 XThR.Tn[3] XThR.Tn[3].n76 0.848714
R24039 XThR.Tn[3] XThR.Tn[3].n81 0.848714
R24040 XThR.Tn[3] XThR.Tn[3].n86 0.848714
R24041 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R24042 XThR.Tn[3].n11 XThR.Tn[3] 0.485653
R24043 XThR.Tn[3].n84 XThR.Tn[3] 0.21482
R24044 XThR.Tn[3].n79 XThR.Tn[3] 0.21482
R24045 XThR.Tn[3].n74 XThR.Tn[3] 0.21482
R24046 XThR.Tn[3].n69 XThR.Tn[3] 0.21482
R24047 XThR.Tn[3].n64 XThR.Tn[3] 0.21482
R24048 XThR.Tn[3].n59 XThR.Tn[3] 0.21482
R24049 XThR.Tn[3].n54 XThR.Tn[3] 0.21482
R24050 XThR.Tn[3].n49 XThR.Tn[3] 0.21482
R24051 XThR.Tn[3].n44 XThR.Tn[3] 0.21482
R24052 XThR.Tn[3].n39 XThR.Tn[3] 0.21482
R24053 XThR.Tn[3].n34 XThR.Tn[3] 0.21482
R24054 XThR.Tn[3].n29 XThR.Tn[3] 0.21482
R24055 XThR.Tn[3].n24 XThR.Tn[3] 0.21482
R24056 XThR.Tn[3].n19 XThR.Tn[3] 0.21482
R24057 XThR.Tn[3].n14 XThR.Tn[3] 0.21482
R24058 XThR.Tn[3].n85 XThR.Tn[3] 0.0608448
R24059 XThR.Tn[3].n80 XThR.Tn[3] 0.0608448
R24060 XThR.Tn[3].n75 XThR.Tn[3] 0.0608448
R24061 XThR.Tn[3].n70 XThR.Tn[3] 0.0608448
R24062 XThR.Tn[3].n65 XThR.Tn[3] 0.0608448
R24063 XThR.Tn[3].n60 XThR.Tn[3] 0.0608448
R24064 XThR.Tn[3].n55 XThR.Tn[3] 0.0608448
R24065 XThR.Tn[3].n50 XThR.Tn[3] 0.0608448
R24066 XThR.Tn[3].n45 XThR.Tn[3] 0.0608448
R24067 XThR.Tn[3].n40 XThR.Tn[3] 0.0608448
R24068 XThR.Tn[3].n35 XThR.Tn[3] 0.0608448
R24069 XThR.Tn[3].n30 XThR.Tn[3] 0.0608448
R24070 XThR.Tn[3].n25 XThR.Tn[3] 0.0608448
R24071 XThR.Tn[3].n20 XThR.Tn[3] 0.0608448
R24072 XThR.Tn[3].n15 XThR.Tn[3] 0.0608448
R24073 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R24074 XThR.Tn[3] XThR.Tn[3].n87 0.038
R24075 XThR.Tn[3].n11 XThR.Tn[3] 0.00744444
R24076 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00265517
R24077 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00265517
R24078 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00265517
R24079 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00265517
R24080 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00265517
R24081 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00265517
R24082 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00265517
R24083 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00265517
R24084 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00265517
R24085 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00265517
R24086 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00265517
R24087 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00265517
R24088 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00265517
R24089 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00265517
R24090 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00265517
R24091 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R24092 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R24093 XThR.Tn[2] XThR.Tn[2].n82 161.363
R24094 XThR.Tn[2] XThR.Tn[2].n77 161.363
R24095 XThR.Tn[2] XThR.Tn[2].n72 161.363
R24096 XThR.Tn[2] XThR.Tn[2].n67 161.363
R24097 XThR.Tn[2] XThR.Tn[2].n62 161.363
R24098 XThR.Tn[2] XThR.Tn[2].n57 161.363
R24099 XThR.Tn[2] XThR.Tn[2].n52 161.363
R24100 XThR.Tn[2] XThR.Tn[2].n47 161.363
R24101 XThR.Tn[2] XThR.Tn[2].n42 161.363
R24102 XThR.Tn[2] XThR.Tn[2].n37 161.363
R24103 XThR.Tn[2] XThR.Tn[2].n32 161.363
R24104 XThR.Tn[2] XThR.Tn[2].n27 161.363
R24105 XThR.Tn[2] XThR.Tn[2].n22 161.363
R24106 XThR.Tn[2] XThR.Tn[2].n17 161.363
R24107 XThR.Tn[2] XThR.Tn[2].n12 161.363
R24108 XThR.Tn[2] XThR.Tn[2].n10 161.363
R24109 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R24110 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R24111 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R24112 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R24113 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R24114 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R24115 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R24116 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R24117 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R24118 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R24119 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R24120 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R24121 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R24122 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R24123 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R24124 XThR.Tn[2].n83 XThR.Tn[2].t38 161.106
R24125 XThR.Tn[2].n82 XThR.Tn[2].t46 161.106
R24126 XThR.Tn[2].n78 XThR.Tn[2].t45 161.106
R24127 XThR.Tn[2].n77 XThR.Tn[2].t52 161.106
R24128 XThR.Tn[2].n73 XThR.Tn[2].t28 161.106
R24129 XThR.Tn[2].n72 XThR.Tn[2].t33 161.106
R24130 XThR.Tn[2].n68 XThR.Tn[2].t73 161.106
R24131 XThR.Tn[2].n67 XThR.Tn[2].t13 161.106
R24132 XThR.Tn[2].n63 XThR.Tn[2].t37 161.106
R24133 XThR.Tn[2].n62 XThR.Tn[2].t43 161.106
R24134 XThR.Tn[2].n58 XThR.Tn[2].t61 161.106
R24135 XThR.Tn[2].n57 XThR.Tn[2].t69 161.106
R24136 XThR.Tn[2].n53 XThR.Tn[2].t42 161.106
R24137 XThR.Tn[2].n52 XThR.Tn[2].t50 161.106
R24138 XThR.Tn[2].n48 XThR.Tn[2].t24 161.106
R24139 XThR.Tn[2].n47 XThR.Tn[2].t30 161.106
R24140 XThR.Tn[2].n43 XThR.Tn[2].t71 161.106
R24141 XThR.Tn[2].n42 XThR.Tn[2].t12 161.106
R24142 XThR.Tn[2].n38 XThR.Tn[2].t15 161.106
R24143 XThR.Tn[2].n37 XThR.Tn[2].t20 161.106
R24144 XThR.Tn[2].n33 XThR.Tn[2].t60 161.106
R24145 XThR.Tn[2].n32 XThR.Tn[2].t68 161.106
R24146 XThR.Tn[2].n28 XThR.Tn[2].t26 161.106
R24147 XThR.Tn[2].n27 XThR.Tn[2].t32 161.106
R24148 XThR.Tn[2].n23 XThR.Tn[2].t58 161.106
R24149 XThR.Tn[2].n22 XThR.Tn[2].t66 161.106
R24150 XThR.Tn[2].n18 XThR.Tn[2].t41 161.106
R24151 XThR.Tn[2].n17 XThR.Tn[2].t48 161.106
R24152 XThR.Tn[2].n13 XThR.Tn[2].t65 161.106
R24153 XThR.Tn[2].n12 XThR.Tn[2].t72 161.106
R24154 XThR.Tn[2].n10 XThR.Tn[2].t54 161.106
R24155 XThR.Tn[2].n83 XThR.Tn[2].t57 154.679
R24156 XThR.Tn[2].n82 XThR.Tn[2].t64 154.679
R24157 XThR.Tn[2].n78 XThR.Tn[2].t36 154.679
R24158 XThR.Tn[2].n77 XThR.Tn[2].t40 154.679
R24159 XThR.Tn[2].n73 XThR.Tn[2].t17 154.679
R24160 XThR.Tn[2].n72 XThR.Tn[2].t22 154.679
R24161 XThR.Tn[2].n68 XThR.Tn[2].t47 154.679
R24162 XThR.Tn[2].n67 XThR.Tn[2].t53 154.679
R24163 XThR.Tn[2].n63 XThR.Tn[2].t29 154.679
R24164 XThR.Tn[2].n62 XThR.Tn[2].t34 154.679
R24165 XThR.Tn[2].n58 XThR.Tn[2].t56 154.679
R24166 XThR.Tn[2].n57 XThR.Tn[2].t62 154.679
R24167 XThR.Tn[2].n53 XThR.Tn[2].t18 154.679
R24168 XThR.Tn[2].n52 XThR.Tn[2].t23 154.679
R24169 XThR.Tn[2].n48 XThR.Tn[2].t63 154.679
R24170 XThR.Tn[2].n47 XThR.Tn[2].t70 154.679
R24171 XThR.Tn[2].n43 XThR.Tn[2].t44 154.679
R24172 XThR.Tn[2].n42 XThR.Tn[2].t51 154.679
R24173 XThR.Tn[2].n38 XThR.Tn[2].t25 154.679
R24174 XThR.Tn[2].n37 XThR.Tn[2].t31 154.679
R24175 XThR.Tn[2].n33 XThR.Tn[2].t35 154.679
R24176 XThR.Tn[2].n32 XThR.Tn[2].t39 154.679
R24177 XThR.Tn[2].n28 XThR.Tn[2].t16 154.679
R24178 XThR.Tn[2].n27 XThR.Tn[2].t21 154.679
R24179 XThR.Tn[2].n23 XThR.Tn[2].t49 154.679
R24180 XThR.Tn[2].n22 XThR.Tn[2].t55 154.679
R24181 XThR.Tn[2].n18 XThR.Tn[2].t14 154.679
R24182 XThR.Tn[2].n17 XThR.Tn[2].t19 154.679
R24183 XThR.Tn[2].n13 XThR.Tn[2].t59 154.679
R24184 XThR.Tn[2].n12 XThR.Tn[2].t67 154.679
R24185 XThR.Tn[2].n10 XThR.Tn[2].t27 154.679
R24186 XThR.Tn[2].n7 XThR.Tn[2].n6 135.249
R24187 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R24188 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R24189 XThR.Tn[2].n7 XThR.Tn[2].n5 98.982
R24190 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R24191 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R24192 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R24193 XThR.Tn[2].n1 XThR.Tn[2].t5 26.5955
R24194 XThR.Tn[2].n1 XThR.Tn[2].t4 26.5955
R24195 XThR.Tn[2].n0 XThR.Tn[2].t6 26.5955
R24196 XThR.Tn[2].n0 XThR.Tn[2].t3 26.5955
R24197 XThR.Tn[2].n3 XThR.Tn[2].t9 24.9236
R24198 XThR.Tn[2].n3 XThR.Tn[2].t10 24.9236
R24199 XThR.Tn[2].n4 XThR.Tn[2].t8 24.9236
R24200 XThR.Tn[2].n4 XThR.Tn[2].t7 24.9236
R24201 XThR.Tn[2].n5 XThR.Tn[2].t11 24.9236
R24202 XThR.Tn[2].n5 XThR.Tn[2].t1 24.9236
R24203 XThR.Tn[2].n6 XThR.Tn[2].t2 24.9236
R24204 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R24205 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R24206 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R24207 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R24208 XThR.Tn[2] XThR.Tn[2].n11 5.34871
R24209 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R24210 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R24211 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R24212 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R24213 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R24214 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R24215 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R24216 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R24217 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R24218 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R24219 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R24220 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R24221 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R24222 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R24223 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R24224 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R24225 XThR.Tn[2].n16 XThR.Tn[2] 2.51836
R24226 XThR.Tn[2].n21 XThR.Tn[2] 2.51836
R24227 XThR.Tn[2].n26 XThR.Tn[2] 2.51836
R24228 XThR.Tn[2].n31 XThR.Tn[2] 2.51836
R24229 XThR.Tn[2].n36 XThR.Tn[2] 2.51836
R24230 XThR.Tn[2].n41 XThR.Tn[2] 2.51836
R24231 XThR.Tn[2].n46 XThR.Tn[2] 2.51836
R24232 XThR.Tn[2].n51 XThR.Tn[2] 2.51836
R24233 XThR.Tn[2].n56 XThR.Tn[2] 2.51836
R24234 XThR.Tn[2].n61 XThR.Tn[2] 2.51836
R24235 XThR.Tn[2].n66 XThR.Tn[2] 2.51836
R24236 XThR.Tn[2].n71 XThR.Tn[2] 2.51836
R24237 XThR.Tn[2].n76 XThR.Tn[2] 2.51836
R24238 XThR.Tn[2].n81 XThR.Tn[2] 2.51836
R24239 XThR.Tn[2].n86 XThR.Tn[2] 2.51836
R24240 XThR.Tn[2] XThR.Tn[2].n16 0.848714
R24241 XThR.Tn[2] XThR.Tn[2].n21 0.848714
R24242 XThR.Tn[2] XThR.Tn[2].n26 0.848714
R24243 XThR.Tn[2] XThR.Tn[2].n31 0.848714
R24244 XThR.Tn[2] XThR.Tn[2].n36 0.848714
R24245 XThR.Tn[2] XThR.Tn[2].n41 0.848714
R24246 XThR.Tn[2] XThR.Tn[2].n46 0.848714
R24247 XThR.Tn[2] XThR.Tn[2].n51 0.848714
R24248 XThR.Tn[2] XThR.Tn[2].n56 0.848714
R24249 XThR.Tn[2] XThR.Tn[2].n61 0.848714
R24250 XThR.Tn[2] XThR.Tn[2].n66 0.848714
R24251 XThR.Tn[2] XThR.Tn[2].n71 0.848714
R24252 XThR.Tn[2] XThR.Tn[2].n76 0.848714
R24253 XThR.Tn[2] XThR.Tn[2].n81 0.848714
R24254 XThR.Tn[2] XThR.Tn[2].n86 0.848714
R24255 XThR.Tn[2].n11 XThR.Tn[2] 0.485653
R24256 XThR.Tn[2].n84 XThR.Tn[2] 0.21482
R24257 XThR.Tn[2].n79 XThR.Tn[2] 0.21482
R24258 XThR.Tn[2].n74 XThR.Tn[2] 0.21482
R24259 XThR.Tn[2].n69 XThR.Tn[2] 0.21482
R24260 XThR.Tn[2].n64 XThR.Tn[2] 0.21482
R24261 XThR.Tn[2].n59 XThR.Tn[2] 0.21482
R24262 XThR.Tn[2].n54 XThR.Tn[2] 0.21482
R24263 XThR.Tn[2].n49 XThR.Tn[2] 0.21482
R24264 XThR.Tn[2].n44 XThR.Tn[2] 0.21482
R24265 XThR.Tn[2].n39 XThR.Tn[2] 0.21482
R24266 XThR.Tn[2].n34 XThR.Tn[2] 0.21482
R24267 XThR.Tn[2].n29 XThR.Tn[2] 0.21482
R24268 XThR.Tn[2].n24 XThR.Tn[2] 0.21482
R24269 XThR.Tn[2].n19 XThR.Tn[2] 0.21482
R24270 XThR.Tn[2].n14 XThR.Tn[2] 0.21482
R24271 XThR.Tn[2].n85 XThR.Tn[2] 0.0608448
R24272 XThR.Tn[2].n80 XThR.Tn[2] 0.0608448
R24273 XThR.Tn[2].n75 XThR.Tn[2] 0.0608448
R24274 XThR.Tn[2].n70 XThR.Tn[2] 0.0608448
R24275 XThR.Tn[2].n65 XThR.Tn[2] 0.0608448
R24276 XThR.Tn[2].n60 XThR.Tn[2] 0.0608448
R24277 XThR.Tn[2].n55 XThR.Tn[2] 0.0608448
R24278 XThR.Tn[2].n50 XThR.Tn[2] 0.0608448
R24279 XThR.Tn[2].n45 XThR.Tn[2] 0.0608448
R24280 XThR.Tn[2].n40 XThR.Tn[2] 0.0608448
R24281 XThR.Tn[2].n35 XThR.Tn[2] 0.0608448
R24282 XThR.Tn[2].n30 XThR.Tn[2] 0.0608448
R24283 XThR.Tn[2].n25 XThR.Tn[2] 0.0608448
R24284 XThR.Tn[2].n20 XThR.Tn[2] 0.0608448
R24285 XThR.Tn[2].n15 XThR.Tn[2] 0.0608448
R24286 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R24287 XThR.Tn[2] XThR.Tn[2].n87 0.038
R24288 XThR.Tn[2].n11 XThR.Tn[2] 0.00744444
R24289 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00265517
R24290 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00265517
R24291 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00265517
R24292 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00265517
R24293 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00265517
R24294 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00265517
R24295 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00265517
R24296 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00265517
R24297 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00265517
R24298 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00265517
R24299 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00265517
R24300 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00265517
R24301 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00265517
R24302 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00265517
R24303 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00265517
R24304 data[0].n1 data[0].t0 230.155
R24305 data[0].n0 data[0].t2 228.463
R24306 data[0].n1 data[0].t1 157.856
R24307 data[0].n0 data[0].t3 157.07
R24308 data[0].n2 data[0].n1 152.768
R24309 data[0].n4 data[0].n0 152.256
R24310 data[0].n3 data[0].n2 24.1398
R24311 data[0].n4 data[0].n3 9.48418
R24312 data[0] data[0].n4 6.1445
R24313 data[0].n2 data[0] 5.6325
R24314 data[0].n3 data[0] 2.638
R24315 XThR.XTB4.Y XThR.XTB4.Y.t0 230.518
R24316 XThR.XTB4.Y.n10 XThR.XTB4.Y.t12 212.081
R24317 XThR.XTB4.Y.n11 XThR.XTB4.Y.t2 212.081
R24318 XThR.XTB4.Y.n16 XThR.XTB4.Y.t7 212.081
R24319 XThR.XTB4.Y.n17 XThR.XTB4.Y.t6 212.081
R24320 XThR.XTB4.Y.n0 XThR.XTB4.Y.t17 212.081
R24321 XThR.XTB4.Y.n1 XThR.XTB4.Y.t5 212.081
R24322 XThR.XTB4.Y.n3 XThR.XTB4.Y.t15 212.081
R24323 XThR.XTB4.Y.n4 XThR.XTB4.Y.t4 212.081
R24324 XThR.XTB4.Y.n13 XThR.XTB4.Y.n12 173.761
R24325 XThR.XTB4.Y.n2 XThR.XTB4.Y 167.361
R24326 XThR.XTB4.Y.n19 XThR.XTB4.Y.n18 152
R24327 XThR.XTB4.Y.n15 XThR.XTB4.Y.n14 152
R24328 XThR.XTB4.Y.n13 XThR.XTB4.Y.n9 152
R24329 XThR.XTB4.Y.n6 XThR.XTB4.Y.n5 152
R24330 XThR.XTB4.Y.n10 XThR.XTB4.Y.t3 139.78
R24331 XThR.XTB4.Y.n11 XThR.XTB4.Y.t9 139.78
R24332 XThR.XTB4.Y.n16 XThR.XTB4.Y.t14 139.78
R24333 XThR.XTB4.Y.n17 XThR.XTB4.Y.t11 139.78
R24334 XThR.XTB4.Y.n0 XThR.XTB4.Y.t10 139.78
R24335 XThR.XTB4.Y.n1 XThR.XTB4.Y.t16 139.78
R24336 XThR.XTB4.Y.n3 XThR.XTB4.Y.t8 139.78
R24337 XThR.XTB4.Y.n4 XThR.XTB4.Y.t13 139.78
R24338 XThR.XTB4.Y.n21 XThR.XTB4.Y.t1 133.386
R24339 XThR.XTB4.Y.n20 XThR.XTB4.Y.n19 72.9296
R24340 XThR.XTB4.Y.n1 XThR.XTB4.Y.n0 61.346
R24341 XThR.XTB4.Y.n15 XThR.XTB4.Y.n9 49.6611
R24342 XThR.XTB4.Y.n18 XThR.XTB4.Y.n16 45.2793
R24343 XThR.XTB4.Y.n12 XThR.XTB4.Y.n11 42.3581
R24344 XThR.XTB4.Y.n20 XThR.XTB4.Y.n8 38.1854
R24345 XThR.XTB4.Y.n2 XThR.XTB4.Y.n1 30.6732
R24346 XThR.XTB4.Y.n3 XThR.XTB4.Y.n2 30.6732
R24347 XThR.XTB4.Y.n5 XThR.XTB4.Y.n3 30.6732
R24348 XThR.XTB4.Y.n5 XThR.XTB4.Y.n4 30.6732
R24349 XThR.XTB4.Y XThR.XTB4.Y.n21 28.966
R24350 XThR.XTB4.Y.n14 XThR.XTB4.Y.n13 21.7605
R24351 XThR.XTB4.Y.n14 XThR.XTB4.Y 21.1205
R24352 XThR.XTB4.Y.n12 XThR.XTB4.Y.n10 18.9884
R24353 XThR.XTB4.Y.n18 XThR.XTB4.Y.n17 16.0672
R24354 XThR.XTB4.Y.n21 XThR.XTB4.Y.n20 11.994
R24355 XThR.XTB4.Y.n22 XThR.XTB4.Y 11.6875
R24356 XThR.XTB4.Y.n8 XThR.XTB4.Y.n7 8.21182
R24357 XThR.XTB4.Y.n11 XThR.XTB4.Y.n9 7.30353
R24358 XThR.XTB4.Y.n8 XThR.XTB4.Y.n6 7.24578
R24359 XThR.XTB4.Y.n22 XThR.XTB4.Y 7.23528
R24360 XThR.XTB4.Y.n6 XThR.XTB4.Y 6.08654
R24361 XThR.XTB4.Y XThR.XTB4.Y.n22 5.04292
R24362 XThR.XTB4.Y.n16 XThR.XTB4.Y.n15 4.38232
R24363 XThR.XTB4.Y.n7 XThR.XTB4.Y 1.79489
R24364 XThR.XTB4.Y.n7 XThR.XTB4.Y 0.966538
R24365 XThR.XTB4.Y.n19 XThR.XTB4.Y 0.6405
R24366 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R24367 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R24368 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R24369 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R24370 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R24371 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R24372 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R24373 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R24374 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24375 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24376 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24377 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24378 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24379 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24380 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24381 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24382 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24383 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24384 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24385 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24386 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24387 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24388 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24389 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24390 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24391 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24392 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24393 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24394 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24395 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24396 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24397 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24398 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24399 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24400 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24401 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24402 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24403 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24404 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24405 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24406 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24407 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24408 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24409 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24410 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24411 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24412 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24413 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24414 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24415 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24416 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24417 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24418 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R24419 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R24420 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R24421 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R24422 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R24423 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R24424 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R24425 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R24426 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R24427 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R24428 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R24429 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R24430 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R24431 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R24432 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R24433 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R24434 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R24435 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R24436 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R24437 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R24438 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R24439 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R24440 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R24441 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R24442 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R24443 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R24444 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R24445 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R24446 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R24447 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R24448 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R24449 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R24450 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R24451 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R24452 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R24453 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R24454 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R24455 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R24456 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R24457 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R24458 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R24459 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R24460 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R24461 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R24462 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R24463 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R24464 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R24465 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R24466 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R24467 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R24468 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R24469 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R24470 XThC.Tn[3].n2 XThC.Tn[3].n1 332.332
R24471 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R24472 XThC.Tn[3].n71 XThC.Tn[3].n69 161.365
R24473 XThC.Tn[3].n67 XThC.Tn[3].n65 161.365
R24474 XThC.Tn[3].n63 XThC.Tn[3].n61 161.365
R24475 XThC.Tn[3].n59 XThC.Tn[3].n57 161.365
R24476 XThC.Tn[3].n55 XThC.Tn[3].n53 161.365
R24477 XThC.Tn[3].n51 XThC.Tn[3].n49 161.365
R24478 XThC.Tn[3].n47 XThC.Tn[3].n45 161.365
R24479 XThC.Tn[3].n43 XThC.Tn[3].n41 161.365
R24480 XThC.Tn[3].n39 XThC.Tn[3].n37 161.365
R24481 XThC.Tn[3].n35 XThC.Tn[3].n33 161.365
R24482 XThC.Tn[3].n31 XThC.Tn[3].n29 161.365
R24483 XThC.Tn[3].n27 XThC.Tn[3].n25 161.365
R24484 XThC.Tn[3].n23 XThC.Tn[3].n21 161.365
R24485 XThC.Tn[3].n19 XThC.Tn[3].n17 161.365
R24486 XThC.Tn[3].n15 XThC.Tn[3].n13 161.365
R24487 XThC.Tn[3].n12 XThC.Tn[3].n10 161.365
R24488 XThC.Tn[3].n69 XThC.Tn[3].t34 161.106
R24489 XThC.Tn[3].n65 XThC.Tn[3].t14 161.106
R24490 XThC.Tn[3].n61 XThC.Tn[3].t12 161.106
R24491 XThC.Tn[3].n57 XThC.Tn[3].t43 161.106
R24492 XThC.Tn[3].n53 XThC.Tn[3].t24 161.106
R24493 XThC.Tn[3].n49 XThC.Tn[3].t21 161.106
R24494 XThC.Tn[3].n45 XThC.Tn[3].t41 161.106
R24495 XThC.Tn[3].n41 XThC.Tn[3].t32 161.106
R24496 XThC.Tn[3].n37 XThC.Tn[3].t30 161.106
R24497 XThC.Tn[3].n33 XThC.Tn[3].t19 161.106
R24498 XThC.Tn[3].n29 XThC.Tn[3].t40 161.106
R24499 XThC.Tn[3].n25 XThC.Tn[3].t29 161.106
R24500 XThC.Tn[3].n21 XThC.Tn[3].t18 161.106
R24501 XThC.Tn[3].n17 XThC.Tn[3].t17 161.106
R24502 XThC.Tn[3].n13 XThC.Tn[3].t36 161.106
R24503 XThC.Tn[3].n10 XThC.Tn[3].t26 161.106
R24504 XThC.Tn[3].n69 XThC.Tn[3].t22 154.679
R24505 XThC.Tn[3].n65 XThC.Tn[3].t33 154.679
R24506 XThC.Tn[3].n61 XThC.Tn[3].t31 154.679
R24507 XThC.Tn[3].n57 XThC.Tn[3].t28 154.679
R24508 XThC.Tn[3].n53 XThC.Tn[3].t42 154.679
R24509 XThC.Tn[3].n49 XThC.Tn[3].t39 154.679
R24510 XThC.Tn[3].n45 XThC.Tn[3].t27 154.679
R24511 XThC.Tn[3].n41 XThC.Tn[3].t20 154.679
R24512 XThC.Tn[3].n37 XThC.Tn[3].t16 154.679
R24513 XThC.Tn[3].n33 XThC.Tn[3].t38 154.679
R24514 XThC.Tn[3].n29 XThC.Tn[3].t25 154.679
R24515 XThC.Tn[3].n25 XThC.Tn[3].t15 154.679
R24516 XThC.Tn[3].n21 XThC.Tn[3].t37 154.679
R24517 XThC.Tn[3].n17 XThC.Tn[3].t35 154.679
R24518 XThC.Tn[3].n13 XThC.Tn[3].t23 154.679
R24519 XThC.Tn[3].n10 XThC.Tn[3].t13 154.679
R24520 XThC.Tn[3].n7 XThC.Tn[3].n6 135.249
R24521 XThC.Tn[3].n9 XThC.Tn[3].n3 98.981
R24522 XThC.Tn[3].n8 XThC.Tn[3].n4 98.981
R24523 XThC.Tn[3].n7 XThC.Tn[3].n5 98.981
R24524 XThC.Tn[3].n9 XThC.Tn[3].n8 36.2672
R24525 XThC.Tn[3].n8 XThC.Tn[3].n7 36.2672
R24526 XThC.Tn[3].n74 XThC.Tn[3].n9 32.6405
R24527 XThC.Tn[3].n1 XThC.Tn[3].t7 26.5955
R24528 XThC.Tn[3].n1 XThC.Tn[3].t6 26.5955
R24529 XThC.Tn[3].n0 XThC.Tn[3].t5 26.5955
R24530 XThC.Tn[3].n0 XThC.Tn[3].t4 26.5955
R24531 XThC.Tn[3].n3 XThC.Tn[3].t9 24.9236
R24532 XThC.Tn[3].n3 XThC.Tn[3].t8 24.9236
R24533 XThC.Tn[3].n4 XThC.Tn[3].t11 24.9236
R24534 XThC.Tn[3].n4 XThC.Tn[3].t10 24.9236
R24535 XThC.Tn[3].n5 XThC.Tn[3].t1 24.9236
R24536 XThC.Tn[3].n5 XThC.Tn[3].t0 24.9236
R24537 XThC.Tn[3].n6 XThC.Tn[3].t3 24.9236
R24538 XThC.Tn[3].n6 XThC.Tn[3].t2 24.9236
R24539 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R24540 XThC.Tn[3] XThC.Tn[3].n12 8.0245
R24541 XThC.Tn[3].n72 XThC.Tn[3].n71 7.9105
R24542 XThC.Tn[3].n68 XThC.Tn[3].n67 7.9105
R24543 XThC.Tn[3].n64 XThC.Tn[3].n63 7.9105
R24544 XThC.Tn[3].n60 XThC.Tn[3].n59 7.9105
R24545 XThC.Tn[3].n56 XThC.Tn[3].n55 7.9105
R24546 XThC.Tn[3].n52 XThC.Tn[3].n51 7.9105
R24547 XThC.Tn[3].n48 XThC.Tn[3].n47 7.9105
R24548 XThC.Tn[3].n44 XThC.Tn[3].n43 7.9105
R24549 XThC.Tn[3].n40 XThC.Tn[3].n39 7.9105
R24550 XThC.Tn[3].n36 XThC.Tn[3].n35 7.9105
R24551 XThC.Tn[3].n32 XThC.Tn[3].n31 7.9105
R24552 XThC.Tn[3].n28 XThC.Tn[3].n27 7.9105
R24553 XThC.Tn[3].n24 XThC.Tn[3].n23 7.9105
R24554 XThC.Tn[3].n20 XThC.Tn[3].n19 7.9105
R24555 XThC.Tn[3].n16 XThC.Tn[3].n15 7.9105
R24556 XThC.Tn[3].n73 XThC.Tn[3] 7.48718
R24557 XThC.Tn[3] XThC.Tn[3].n74 6.7205
R24558 XThC.Tn[3].n74 XThC.Tn[3].n73 5.06464
R24559 XThC.Tn[3].n73 XThC.Tn[3] 1.18175
R24560 XThC.Tn[3].n16 XThC.Tn[3] 0.235138
R24561 XThC.Tn[3].n20 XThC.Tn[3] 0.235138
R24562 XThC.Tn[3].n24 XThC.Tn[3] 0.235138
R24563 XThC.Tn[3].n28 XThC.Tn[3] 0.235138
R24564 XThC.Tn[3].n32 XThC.Tn[3] 0.235138
R24565 XThC.Tn[3].n36 XThC.Tn[3] 0.235138
R24566 XThC.Tn[3].n40 XThC.Tn[3] 0.235138
R24567 XThC.Tn[3].n44 XThC.Tn[3] 0.235138
R24568 XThC.Tn[3].n48 XThC.Tn[3] 0.235138
R24569 XThC.Tn[3].n52 XThC.Tn[3] 0.235138
R24570 XThC.Tn[3].n56 XThC.Tn[3] 0.235138
R24571 XThC.Tn[3].n60 XThC.Tn[3] 0.235138
R24572 XThC.Tn[3].n64 XThC.Tn[3] 0.235138
R24573 XThC.Tn[3].n68 XThC.Tn[3] 0.235138
R24574 XThC.Tn[3].n72 XThC.Tn[3] 0.235138
R24575 XThC.Tn[3] XThC.Tn[3].n16 0.114505
R24576 XThC.Tn[3] XThC.Tn[3].n20 0.114505
R24577 XThC.Tn[3] XThC.Tn[3].n24 0.114505
R24578 XThC.Tn[3] XThC.Tn[3].n28 0.114505
R24579 XThC.Tn[3] XThC.Tn[3].n32 0.114505
R24580 XThC.Tn[3] XThC.Tn[3].n36 0.114505
R24581 XThC.Tn[3] XThC.Tn[3].n40 0.114505
R24582 XThC.Tn[3] XThC.Tn[3].n44 0.114505
R24583 XThC.Tn[3] XThC.Tn[3].n48 0.114505
R24584 XThC.Tn[3] XThC.Tn[3].n52 0.114505
R24585 XThC.Tn[3] XThC.Tn[3].n56 0.114505
R24586 XThC.Tn[3] XThC.Tn[3].n60 0.114505
R24587 XThC.Tn[3] XThC.Tn[3].n64 0.114505
R24588 XThC.Tn[3] XThC.Tn[3].n68 0.114505
R24589 XThC.Tn[3] XThC.Tn[3].n72 0.114505
R24590 XThC.Tn[3].n71 XThC.Tn[3].n70 0.0599512
R24591 XThC.Tn[3].n67 XThC.Tn[3].n66 0.0599512
R24592 XThC.Tn[3].n63 XThC.Tn[3].n62 0.0599512
R24593 XThC.Tn[3].n59 XThC.Tn[3].n58 0.0599512
R24594 XThC.Tn[3].n55 XThC.Tn[3].n54 0.0599512
R24595 XThC.Tn[3].n51 XThC.Tn[3].n50 0.0599512
R24596 XThC.Tn[3].n47 XThC.Tn[3].n46 0.0599512
R24597 XThC.Tn[3].n43 XThC.Tn[3].n42 0.0599512
R24598 XThC.Tn[3].n39 XThC.Tn[3].n38 0.0599512
R24599 XThC.Tn[3].n35 XThC.Tn[3].n34 0.0599512
R24600 XThC.Tn[3].n31 XThC.Tn[3].n30 0.0599512
R24601 XThC.Tn[3].n27 XThC.Tn[3].n26 0.0599512
R24602 XThC.Tn[3].n23 XThC.Tn[3].n22 0.0599512
R24603 XThC.Tn[3].n19 XThC.Tn[3].n18 0.0599512
R24604 XThC.Tn[3].n15 XThC.Tn[3].n14 0.0599512
R24605 XThC.Tn[3].n12 XThC.Tn[3].n11 0.0599512
R24606 XThC.Tn[3].n70 XThC.Tn[3] 0.0469286
R24607 XThC.Tn[3].n66 XThC.Tn[3] 0.0469286
R24608 XThC.Tn[3].n62 XThC.Tn[3] 0.0469286
R24609 XThC.Tn[3].n58 XThC.Tn[3] 0.0469286
R24610 XThC.Tn[3].n54 XThC.Tn[3] 0.0469286
R24611 XThC.Tn[3].n50 XThC.Tn[3] 0.0469286
R24612 XThC.Tn[3].n46 XThC.Tn[3] 0.0469286
R24613 XThC.Tn[3].n42 XThC.Tn[3] 0.0469286
R24614 XThC.Tn[3].n38 XThC.Tn[3] 0.0469286
R24615 XThC.Tn[3].n34 XThC.Tn[3] 0.0469286
R24616 XThC.Tn[3].n30 XThC.Tn[3] 0.0469286
R24617 XThC.Tn[3].n26 XThC.Tn[3] 0.0469286
R24618 XThC.Tn[3].n22 XThC.Tn[3] 0.0469286
R24619 XThC.Tn[3].n18 XThC.Tn[3] 0.0469286
R24620 XThC.Tn[3].n14 XThC.Tn[3] 0.0469286
R24621 XThC.Tn[3].n11 XThC.Tn[3] 0.0469286
R24622 XThC.Tn[3].n70 XThC.Tn[3] 0.0401341
R24623 XThC.Tn[3].n66 XThC.Tn[3] 0.0401341
R24624 XThC.Tn[3].n62 XThC.Tn[3] 0.0401341
R24625 XThC.Tn[3].n58 XThC.Tn[3] 0.0401341
R24626 XThC.Tn[3].n54 XThC.Tn[3] 0.0401341
R24627 XThC.Tn[3].n50 XThC.Tn[3] 0.0401341
R24628 XThC.Tn[3].n46 XThC.Tn[3] 0.0401341
R24629 XThC.Tn[3].n42 XThC.Tn[3] 0.0401341
R24630 XThC.Tn[3].n38 XThC.Tn[3] 0.0401341
R24631 XThC.Tn[3].n34 XThC.Tn[3] 0.0401341
R24632 XThC.Tn[3].n30 XThC.Tn[3] 0.0401341
R24633 XThC.Tn[3].n26 XThC.Tn[3] 0.0401341
R24634 XThC.Tn[3].n22 XThC.Tn[3] 0.0401341
R24635 XThC.Tn[3].n18 XThC.Tn[3] 0.0401341
R24636 XThC.Tn[3].n14 XThC.Tn[3] 0.0401341
R24637 XThC.Tn[3].n11 XThC.Tn[3] 0.0401341
R24638 data[6].n0 data[6].t0 230.576
R24639 data[6].n0 data[6].t1 158.275
R24640 data[6].n1 data[6].n0 152
R24641 data[6].n1 data[6] 11.9995
R24642 data[6] data[6].n1 6.66717
R24643 data[1].n4 data[1].t2 230.576
R24644 data[1].n1 data[1].t0 230.363
R24645 data[1].n0 data[1].t4 229.369
R24646 data[1].n4 data[1].t5 158.275
R24647 data[1].n1 data[1].t3 158.064
R24648 data[1].n0 data[1].t1 157.07
R24649 data[1].n2 data[1].n1 153.28
R24650 data[1].n7 data[1].n0 153.147
R24651 data[1].n5 data[1].n4 152
R24652 data[1].n7 data[1].n6 16.3874
R24653 data[1].n6 data[1].n5 14.9641
R24654 data[1].n3 data[1].n2 9.3005
R24655 data[1].n6 data[1].n3 6.49639
R24656 data[1] data[1].n7 3.24826
R24657 data[1].n2 data[1] 2.92621
R24658 data[1].n3 data[1] 2.15819
R24659 data[1].n5 data[1] 2.13383
R24660 data[2].n0 data[2].t0 230.576
R24661 data[2].n0 data[2].t1 158.275
R24662 data[2].n1 data[2].n0 152
R24663 data[2].n1 data[2] 12.7714
R24664 data[2] data[2].n1 2.13383
R24665 data[5].n4 data[5].t2 230.576
R24666 data[5].n1 data[5].t0 230.363
R24667 data[5].n0 data[5].t1 229.369
R24668 data[5].n4 data[5].t5 158.275
R24669 data[5].n1 data[5].t3 158.064
R24670 data[5].n0 data[5].t4 157.07
R24671 data[5].n2 data[5].n1 152.256
R24672 data[5].n7 data[5].n0 152.238
R24673 data[5].n5 data[5].n4 152
R24674 data[5].n7 data[5].n6 16.3874
R24675 data[5].n6 data[5].n5 14.6005
R24676 data[5].n3 data[5].n2 9.3005
R24677 data[5].n5 data[5] 6.66717
R24678 data[5].n6 data[5].n3 6.49639
R24679 data[5].n2 data[5] 6.1445
R24680 data[5] data[5].n7 5.68939
R24681 data[5].n3 data[5] 2.28319
R24682 data[3].n0 data[3].t1 230.576
R24683 data[3].n0 data[3].t0 158.275
R24684 data[3].n1 data[3].n0 153.553
R24685 data[3].n1 data[3] 11.6078
R24686 data[3] data[3].n1 2.90959
R24687 data[7].n0 data[7].t0 230.576
R24688 data[7].n0 data[7].t1 158.275
R24689 data[7].n1 data[7].n0 152
R24690 data[7].n1 data[7] 11.9995
R24691 data[7] data[7].n1 6.66717
R24692 bias[1] bias[1].t0 23.8076
R24693 bias[2] bias[2].t0 57.7456
R24694 bias[0] bias[0].t0 12.1467
C0 XThR.Tn[9] XA.XIR[10].XIC[12].icell.SM 0.00121f
C1 XThC.Tn[4] XThR.Tn[9] 0.28062f
C2 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02698f
C3 a_5155_9615# Vbias 0.00652f
C4 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.01406f
C5 XA.XIR[10].XIC[9].icell.Ien VPWR 0.19065f
C6 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.03424f
C7 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00212f
C8 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.SM 0.00383f
C9 XThR.Tn[1] XA.XIR[2].XIC[9].icell.Ien 0.00321f
C10 XA.XIR[15].XIC[13].icell.SM Vbias 0.00701f
C11 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.SM 0.00188f
C12 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00212f
C13 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.15089f
C14 XA.XIR[9].XIC[8].icell.SM VPWR 0.00158f
C15 XA.XIR[6].XIC[8].icell.SM Vbias 0.00701f
C16 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.SM 0.00383f
C17 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00529f
C18 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02698f
C19 XA.XIR[5].XIC[11].icell.PUM Vbias 0.00347f
C20 XThR.Tn[3] XA.XIR[4].XIC[6].icell.SM 0.00121f
C21 XA.XIR[9].XIC[5].icell.SM Iout 0.00388f
C22 XA.XIR[13].XIC_dummy_left.icell.Ien Vbias 0.00342f
C23 XA.XIR[7].XIC[0].icell.SM Vbias 0.00675f
C24 XThR.Tn[14] XA.XIR[15].XIC[3].icell.Ien 0.00321f
C25 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.03424f
C26 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.01406f
C27 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04522f
C28 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00212f
C29 XA.XIR[11].XIC_dummy_left.icell.SM VPWR 0.00269f
C30 XA.XIR[3].XIC[11].icell.SM VPWR 0.00158f
C31 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PUM 0.00131f
C32 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PUM 0.00131f
C33 XA.XIR[1].XIC[1].icell.SM Vbias 0.00701f
C34 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02698f
C35 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00529f
C36 XThR.Tn[12] XA.XIR[13].XIC[10].icell.SM 0.00121f
C37 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.15089f
C38 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.15089f
C39 XA.XIR[2].XIC_15.icell.PDM VPWR 0.06959f
C40 XThR.XTB7.B XThR.Tn[5] 0.00705f
C41 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.0353f
C42 XA.XIR[8].XIC[7].icell.SM Vbias 0.00701f
C43 XA.XIR[0].XIC[4].icell.PDM Vbias 0.04061f
C44 XThR.Tn[4] XA.XIR[5].XIC[6].icell.SM 0.00121f
C45 XA.XIR[7].XIC[6].icell.PUM VPWR 0.01036f
C46 XThR.Tn[8] XA.XIR[8].XIC[11].icell.PDM 0.0033f
C47 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PUM 0.00535f
C48 XThR.XTB4.Y a_n997_3979# 0.00497f
C49 XA.XIR[10].XIC[12].icell.PDM VPWR 0.00863f
C50 a_10051_9569# VPWR 0.00319f
C51 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.01406f
C52 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00212f
C53 XThR.Tn[1] XA.XIR[2].XIC[12].icell.SM 0.00121f
C54 XThC.Tn[2] XThR.Tn[11] 0.28062f
C55 XA.XIR[1].XIC[7].icell.PUM VPWR 0.01036f
C56 XA.XIR[13].XIC[1].icell.Ien VPWR 0.19065f
C57 XA.XIR[0].XIC[0].icell.PDM VPWR 0.00806f
C58 XA.XIR[6].XIC[13].icell.PUM Vbias 0.00347f
C59 XA.XIR[9].XIC[13].icell.PUM VPWR 0.01036f
C60 XA.XIR[10].XIC[0].icell.Ien Vbias 0.21102f
C61 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02698f
C62 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PUM 0.00529f
C63 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.SM 0.00383f
C64 XThR.Tn[7] XA.XIR[8].XIC[10].icell.Ien 0.00321f
C65 XThC.XTB6.Y Vbias 0.01416f
C66 XA.XIR[13].XIC[11].icell.PUM VPWR 0.01036f
C67 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.01406f
C68 XA.XIR[0].XIC[7].icell.Ien VPWR 0.19002f
C69 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.15089f
C70 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PUM 0.00131f
C71 XThR.Tn[12] XA.XIR[12].XIC[4].icell.PDM 0.0033f
C72 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PDM 0.00182f
C73 XThR.Tn[3] XA.XIR[3].XIC[14].icell.PDM 0.0033f
C74 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.01406f
C75 XA.XIR[0].XIC[4].icell.Ien Iout 0.06455f
C76 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00529f
C77 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.SM 0.00188f
C78 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PUM 0.00529f
C79 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.SM 0.00383f
C80 XA.XIR[2].XIC[0].icell.PDM Iout 0.00112f
C81 XThR.Tn[5] XA.XIR[5].XIC[11].icell.PDM 0.0033f
C82 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[10].icell.SM 0.00383f
C83 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PUM 0.00131f
C84 XA.XIR[3].XIC_dummy_left.icell.Ien Vbias 0.00342f
C85 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.03592f
C86 XA.XIR[8].XIC[12].icell.PUM Vbias 0.00347f
C87 XThR.Tn[10] Iout 1.16625f
C88 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.SM 0.00383f
C89 XA.XIR[15].XIC[5].icell.PUM Vbias 0.00347f
C90 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01897f
C91 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.15089f
C92 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02698f
C93 XA.XIR[12].XIC[10].icell.SM Vbias 0.00701f
C94 XThC.Tn[8] XThR.Tn[3] 0.28062f
C95 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00212f
C96 XThC.XTB7.A XThC.Tn[6] 0.10589f
C97 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.03982f
C98 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PUM 0.00529f
C99 XThR.Tn[4] XA.XIR[4].XIC[14].icell.PDM 0.0033f
C100 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.03976f
C101 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.03424f
C102 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.38921f
C103 XThR.Tn[7] XA.XIR[8].XIC[13].icell.SM 0.00121f
C104 XThR.XTB7.B a_n1049_6699# 0.0036f
C105 XA.XIR[13].XIC_15.icell.SM VPWR 0.00276f
C106 XThC.Tn[2] XThR.Tn[7] 0.28062f
C107 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.03424f
C108 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PUM 0.00209f
C109 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00529f
C110 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00212f
C111 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PDM 0.00594f
C112 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C113 XThC.Tn[7] XThR.Tn[2] 0.28069f
C114 XThC.Tn[5] XThR.Tn[12] 0.28062f
C115 XA.XIR[3].XIC[1].icell.Ien VPWR 0.19065f
C116 XThR.Tn[6] XA.XIR[7].XIC[0].icell.SM 0.00121f
C117 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.15089f
C118 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.01406f
C119 XA.XIR[9].XIC_dummy_right.icell.Ien Vbias 0.00287f
C120 XA.XIR[8].XIC_15.icell.PDM Iout 0.0013f
C121 XA.XIR[15].XIC[14].icell.PDM Vbias 0.04058f
C122 XA.XIR[2].XIC[3].icell.PUM VPWR 0.01036f
C123 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.03424f
C124 XA.XIR[15].XIC[8].icell.PDM Iout 0.00112f
C125 XA.XIR[0].XIC[13].icell.Ien Vbias 0.21246f
C126 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.15089f
C127 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PUM 0.00529f
C128 XThR.XTBN.A data[4] 0.02581f
C129 XThC.XTB4.Y Vbias 0.01324f
C130 XA.XIR[14].XIC[4].icell.PUM VPWR 0.01036f
C131 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[2].icell.Ien 0.00212f
C132 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.SM 0.00188f
C133 XA.XIR[11].XIC[3].icell.PUM Vbias 0.00347f
C134 XA.XIR[15].XIC[9].icell.PUM Vbias 0.00347f
C135 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PUM 0.00209f
C136 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PUM 0.00131f
C137 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04522f
C138 XA.XIR[13].XIC[5].icell.Ien VPWR 0.19065f
C139 XThR.Tn[1] XA.XIR[2].XIC[2].icell.Ien 0.00321f
C140 XThR.XTB7.A XThR.Tn[2] 0.12549f
C141 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.03424f
C142 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.03528f
C143 XA.XIR[6].XIC[1].icell.SM Vbias 0.00701f
C144 XA.XIR[10].XIC[4].icell.Ien Vbias 0.21238f
C145 XA.XIR[9].XIC[1].icell.SM VPWR 0.00158f
C146 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.SM 0.00188f
C147 XA.XIR[13].XIC[2].icell.Ien Iout 0.06483f
C148 XA.XIR[12].XIC[6].icell.Ien VPWR 0.19065f
C149 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04522f
C150 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.15089f
C151 XA.XIR[5].XIC[4].icell.PUM Vbias 0.00347f
C152 XThC.Tn[4] XThR.Tn[10] 0.28062f
C153 XA.XIR[12].XIC[3].icell.Ien Iout 0.06483f
C154 XA.XIR[11].XIC[9].icell.PDM VPWR 0.00863f
C155 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.15089f
C156 XThC.XTB7.B XThC.Tn[5] 0.00714f
C157 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.03424f
C158 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08027f
C159 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02728f
C160 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PUM 0.00131f
C161 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PUM 0.00529f
C162 XA.XIR[4].XIC[7].icell.PDM Vbias 0.04058f
C163 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.03424f
C164 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PUM 0.00529f
C165 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C166 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PUM 0.00131f
C167 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.03976f
C168 XA.XIR[11].XIC[6].icell.PDM Iout 0.00112f
C169 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06536f
C170 XA.XIR[6].XIC[7].icell.PUM VPWR 0.01036f
C171 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.SM 0.00383f
C172 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.15089f
C173 XThC.XTB6.Y XThC.Tn[13] 0.32552f
C174 XA.XIR[6].XIC[0].icell.PDM Vbias 0.04002f
C175 XThR.XTB5.Y data[7] 0.00931f
C176 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.SM 0.00188f
C177 XA.XIR[3].XIC[7].icell.Ien Vbias 0.21238f
C178 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.SM 0.00383f
C179 XThC.XTB6.A data[0] 0.48493f
C180 XA.XIR[15].XIC[14].icell.PUM Vbias 0.00347f
C181 XA.XIR[10].XIC[5].icell.SM Iout 0.00388f
C182 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00212f
C183 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.03565f
C184 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02698f
C185 XA.XIR[8].XIC[0].icell.SM Vbias 0.00675f
C186 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.03976f
C187 XA.XIR[5].XIC[10].icell.PDM VPWR 0.00863f
C188 XThR.Tn[8] XA.XIR[8].XIC[4].icell.PDM 0.0033f
C189 XA.XIR[2].XIC[9].icell.PUM Vbias 0.00347f
C190 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.15089f
C191 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02698f
C192 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PDM 0.00182f
C193 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.01406f
C194 XA.XIR[13].XIC[9].icell.Ien VPWR 0.19065f
C195 XA.XIR[5].XIC[7].icell.PDM Iout 0.00112f
C196 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.SM 0.00383f
C197 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00529f
C198 XA.XIR[4].XIC[10].icell.Ien VPWR 0.19065f
C199 a_5949_9615# XThC.Tn[6] 0.0018f
C200 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.SM 0.00383f
C201 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PUM 0.00529f
C202 XThR.Tn[12] XA.XIR[13].XIC[1].icell.Ien 0.00321f
C203 XA.XIR[7].XIC[0].icell.PDM Iout 0.00112f
C204 XThR.Tn[7] XA.XIR[8].XIC[3].icell.Ien 0.00321f
C205 XA.XIR[4].XIC[7].icell.Ien Iout 0.06483f
C206 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.02769f
C207 XA.XIR[0].XIC[0].icell.Ien VPWR 0.19003f
C208 XA.XIR[9].XIC[7].icell.SM Vbias 0.00701f
C209 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.SM 0.00188f
C210 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00212f
C211 XA.XIR[8].XIC[6].icell.PUM VPWR 0.01036f
C212 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PUM 0.00131f
C213 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.03976f
C214 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PUM 0.00131f
C215 XA.XIR[3].XIC[8].icell.SM Iout 0.00388f
C216 XThR.XTBN.Y XThR.Tn[5] 0.59911f
C217 XThR.XTB1.Y a_n1335_8331# 0.0097f
C218 XThC.XTBN.Y XThC.Tn[9] 0.49745f
C219 XThR.Tn[5] XA.XIR[5].XIC[4].icell.PDM 0.0033f
C220 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02698f
C221 XA.XIR[14].XIC[0].icell.PUM VPWR 0.01036f
C222 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02801f
C223 XA.XIR[2].XIC[12].icell.PDM Iout 0.00112f
C224 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02698f
C225 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PUM 0.00131f
C226 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Ien 0.00529f
C227 XThR.Tn[9] XA.XIR[10].XIC[13].icell.SM 0.00121f
C228 XA.XIR[10].XIC[10].icell.Ien VPWR 0.19065f
C229 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08194f
C230 XA.XIR[5].XIC[12].icell.Ien VPWR 0.19065f
C231 XA.XIR[2].XIC[14].icell.PDM Vbias 0.04058f
C232 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C233 XA.XIR[15].XIC[14].icell.SM Vbias 0.00701f
C234 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.01406f
C235 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.03547f
C236 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13469f
C237 XThC.XTB7.B a_10051_9569# 0.00209f
C238 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04522f
C239 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PUM 0.00131f
C240 XA.XIR[4].XIC[13].icell.SM VPWR 0.00158f
C241 XA.XIR[13].XIC[12].icell.PDM VPWR 0.00863f
C242 XThR.Tn[14] XA.XIR[15].XIC[6].icell.SM 0.00121f
C243 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.SM 0.00383f
C244 XA.XIR[7].XIC[5].icell.PUM Vbias 0.00347f
C245 XThC.Tn[2] XThR.Tn[14] 0.28062f
C246 XThC.Tn[0] XThR.Tn[0] 0.28136f
C247 a_7875_9569# Vbias 0.00245f
C248 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02698f
C249 XThR.XTB5.Y a_n1049_5317# 0.00907f
C250 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PUM 0.00529f
C251 XA.XIR[13].XIC[0].icell.Ien Vbias 0.21102f
C252 XThC.Tn[8] XThR.Tn[8] 0.28062f
C253 XThR.Tn[11] XA.XIR[11].XIC[13].icell.PDM 0.0033f
C254 XA.XIR[9].XIC[12].icell.PUM Vbias 0.00347f
C255 XA.XIR[1].XIC[6].icell.PUM Vbias 0.00347f
C256 XThC.XTB2.Y Vbias 0.01162f
C257 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.SM 0.00188f
C258 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.SM 0.00383f
C259 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01193f
C260 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.01406f
C261 XThR.Tn[8] XA.XIR[9].XIC[13].icell.Ien 0.00321f
C262 XThC.Tn[9] XThC.Tn[10] 0.08452f
C263 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.02698f
C264 XA.XIR[11].XIC_15.icell.PDM Iout 0.0013f
C265 XA.XIR[12].XIC[1].icell.Ien Vbias 0.21238f
C266 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C267 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.01406f
C268 XA.XIR[0].XIC[6].icell.Ien Vbias 0.21249f
C269 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.03424f
C270 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PUM 0.00131f
C271 XA.XIR[2].XIC[14].icell.Ien Iout 0.06483f
C272 XA.XIR[7].XIC[11].icell.PDM VPWR 0.00863f
C273 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PUM 0.00131f
C274 XA.XIR[3].XIC[14].icell.SM Vbias 0.00701f
C275 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00212f
C276 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PUM 0.00529f
C277 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.SM 0.00188f
C278 XA.XIR[12].XIC[11].icell.PUM Vbias 0.00347f
C279 XThR.XTB7.Y a_n1049_5317# 0.27822f
C280 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6] 0.0033f
C281 XA.XIR[7].XIC[8].icell.PDM Iout 0.00112f
C282 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.PDM 0.00589f
C283 XA.XIR[1].XIC[12].icell.PDM VPWR 0.00863f
C284 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.15089f
C285 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PUM 0.00529f
C286 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PUM 0.00131f
C287 XA.XIR[9].XIC[2].icell.PUM VPWR 0.01036f
C288 XThC.XTB7.Y VPWR 1.07734f
C289 XThR.XTBN.Y a_n1049_6699# 0.07601f
C290 XThR.Tn[13] Iout 1.1663f
C291 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PUM 0.00529f
C292 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01897f
C293 XThR.Tn[12] XA.XIR[13].XIC[5].icell.Ien 0.00321f
C294 XA.XIR[1].XIC[9].icell.PDM Iout 0.00112f
C295 XThC.Tn[9] XThR.Tn[5] 0.28062f
C296 XA.XIR[9].XIC_15.icell.PDM Iout 0.0013f
C297 XA.XIR[0].XIC[10].icell.SM VPWR 0.00158f
C298 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.04037f
C299 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.15089f
C300 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.03981f
C301 XA.XIR[4].XIC[14].icell.SM Iout 0.00388f
C302 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.15089f
C303 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02698f
C304 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00529f
C305 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C306 XA.XIR[0].XIC[7].icell.SM Iout 0.00367f
C307 XA.XIR[15].XIC[12].icell.Ien Vbias 0.17911f
C308 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.SM 0.00383f
C309 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.03424f
C310 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.03976f
C311 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00529f
C312 XA.XIR[10].XIC[1].icell.SM VPWR 0.00158f
C313 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00212f
C314 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PUM 0.00529f
C315 XA.XIR[2].XIC[1].icell.PDM Iout 0.00112f
C316 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PUM 0.00529f
C317 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PUM 0.00131f
C318 XA.XIR[7].XIC[13].icell.Ien VPWR 0.19065f
C319 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PUM 0.00529f
C320 XA.XIR[3].XIC[0].icell.Ien Vbias 0.21102f
C321 XA.XIR[15].XIC[10].icell.PDM Vbias 0.04058f
C322 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.SM 0.00188f
C323 XA.XIR[12].XIC_15.icell.SM Vbias 0.00701f
C324 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.03424f
C325 XA.XIR[5].XIC[3].icell.PDM VPWR 0.00863f
C326 XA.XIR[1].XIC[14].icell.Ien VPWR 0.1907f
C327 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.03983f
C328 XA.XIR[2].XIC[2].icell.PUM Vbias 0.00347f
C329 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.03424f
C330 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00212f
C331 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00212f
C332 XA.XIR[1].XIC[0].icell.Ien Iout 0.06474f
C333 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.SM 0.00383f
C334 XA.XIR[14].XIC[3].icell.PUM Vbias 0.00347f
C335 XA.XIR[4].XIC[3].icell.Ien VPWR 0.19065f
C336 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PUM 0.00131f
C337 XThR.Tn[12] XA.XIR[13].XIC[9].icell.Ien 0.00321f
C338 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PUM 0.00529f
C339 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.SM 0.00383f
C340 XA.XIR[0].XIC[14].icell.SM VPWR 0.00208f
C341 XA.XIR[3].XIC[4].icell.SM VPWR 0.00158f
C342 XA.XIR[13].XIC[4].icell.Ien Vbias 0.21238f
C343 XA.XIR[4].XIC[0].icell.Ien Iout 0.06474f
C344 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PUM 0.00529f
C345 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PUM 0.00131f
C346 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.01406f
C347 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02698f
C348 XThC.Tn[8] data[0] 0.01643f
C349 Vbias Iout 83.1369f
C350 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.SM 0.00383f
C351 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.03976f
C352 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04f
C353 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Ien 0.00529f
C354 XA.XIR[3].XIC[1].icell.SM Iout 0.00388f
C355 XThR.XTB1.Y a_n1049_8581# 0.21263f
C356 XThC.XTB3.Y a_5155_9615# 0.00913f
C357 XA.XIR[12].XIC[5].icell.Ien Vbias 0.21238f
C358 XA.XIR[2].XIC[8].icell.PDM VPWR 0.00863f
C359 XThC.Tn[4] XThR.Tn[13] 0.28062f
C360 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.01406f
C361 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00529f
C362 XA.XIR[14].XIC[9].icell.PDM VPWR 0.00863f
C363 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.01406f
C364 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[3].icell.SM 0.00383f
C365 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00212f
C366 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00529f
C367 XA.XIR[11].XIC[8].icell.PDM Vbias 0.04058f
C368 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PUM 0.00131f
C369 XA.XIR[2].XIC[5].icell.PDM Iout 0.00112f
C370 XThC.Tn[6] XThR.Tn[3] 0.28062f
C371 XA.XIR[14].XIC[6].icell.PDM Iout 0.00112f
C372 XThR.Tn[0] VPWR 6.74637f
C373 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04522f
C374 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PUM 0.00529f
C375 XThR.Tn[1] XA.XIR[2].XIC[5].icell.SM 0.00121f
C376 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C377 XA.XIR[10].XIC[7].icell.SM Vbias 0.00701f
C378 XA.XIR[6].XIC[6].icell.PUM Vbias 0.00347f
C379 XA.XIR[9].XIC[6].icell.PUM VPWR 0.01036f
C380 XThR.Tn[9] XA.XIR[9].XIC[10].icell.PDM 0.0033f
C381 XA.XIR[13].XIC[5].icell.SM Iout 0.00388f
C382 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PUM 0.00131f
C383 XA.XIR[5].XIC[9].icell.PDM Vbias 0.04058f
C384 XA.XIR[1].XIC_15.icell.Ien Iout 0.06485f
C385 XA.XIR[11].XIC[11].icell.SM Iout 0.00388f
C386 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00212f
C387 XA.XIR[0].XIC_dummy_left.icell.SM VPWR 0.00269f
C388 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.SM 0.00188f
C389 XA.XIR[12].XIC[6].icell.SM Iout 0.00388f
C390 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00529f
C391 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.03976f
C392 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.03976f
C393 XThR.Tn[3] XA.XIR[3].XIC[7].icell.PDM 0.0033f
C394 XA.XIR[4].XIC[9].icell.Ien Vbias 0.21238f
C395 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02698f
C396 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.15089f
C397 XA.XIR[11].XIC[8].icell.Ien Iout 0.06483f
C398 XA.XIR[12].XIC[9].icell.Ien Vbias 0.21238f
C399 XA.XIR[6].XIC[12].icell.PDM VPWR 0.00863f
C400 XThR.XTB4.Y XThR.Tn[5] 0.00751f
C401 XThR.XTB5.Y a_n1049_6405# 0.24821f
C402 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PUM 0.00529f
C403 XThR.XTBN.A XThR.Tn[8] 0.1369f
C404 XA.XIR[3].XIC[10].icell.SM Vbias 0.00701f
C405 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PUM 0.00529f
C406 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PUM 0.00131f
C407 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.01406f
C408 XA.XIR[8].XIC[5].icell.PUM Vbias 0.00347f
C409 XA.XIR[6].XIC[9].icell.PDM Iout 0.00112f
C410 XA.XIR[7].XIC[4].icell.PDM VPWR 0.00863f
C411 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.SM 0.00188f
C412 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PUM 0.00131f
C413 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04522f
C414 XThC.Tn[2] XA.XIR[0].XIC[4].icell.PDM 0.00325f
C415 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.15089f
C416 XThR.Tn[3] a_n1049_6405# 0.00542f
C417 XA.XIR[10].XIC[12].icell.SM Vbias 0.00701f
C418 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00529f
C419 XThC.XTB7.Y a_9827_9569# 0.00571f
C420 XThC.Tn[4] Vbias 2.4433f
C421 XA.XIR[1].XIC[5].icell.PDM VPWR 0.00863f
C422 XA.XIR[5].XIC[9].icell.Ien Iout 0.06483f
C423 XThR.Tn[4] XA.XIR[4].XIC[7].icell.PDM 0.0033f
C424 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.15089f
C425 XA.XIR[13].XIC[10].icell.Ien VPWR 0.19065f
C426 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C427 XThR.Tn[7] XA.XIR[8].XIC[6].icell.SM 0.00121f
C428 XA.XIR[4].XIC[10].icell.SM Iout 0.00388f
C429 XA.XIR[15].XIC[10].icell.SM Vbias 0.00701f
C430 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.15089f
C431 XA.XIR[0].XIC[3].icell.SM VPWR 0.00158f
C432 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.SM 0.00383f
C433 XA.XIR[8].XIC[11].icell.PDM VPWR 0.00863f
C434 XThC.XTB5.Y XThC.Tn[7] 0.00912f
C435 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PUM 0.00529f
C436 XA.XIR[11].XIC[1].icell.PUM VPWR 0.01036f
C437 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.03976f
C438 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.0353f
C439 XA.XIR[4].XIC[12].icell.SM Vbias 0.00701f
C440 XA.XIR[11].XIC[13].icell.Ien Iout 0.06483f
C441 XA.XIR[0].XIC[0].icell.SM Iout 0.00367f
C442 XA.XIR[8].XIC[8].icell.PDM Iout 0.00112f
C443 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.15089f
C444 XA.XIR[6].XIC[14].icell.Ien VPWR 0.1907f
C445 XA.XIR[10].XIC[2].icell.PUM VPWR 0.01036f
C446 XThR.Tn[6] Iout 1.16629f
C447 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C448 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00212f
C449 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04522f
C450 XA.XIR[12].XIC[12].icell.PDM Vbias 0.04058f
C451 XA.XIR[14].XIC_15.icell.PDM Iout 0.0013f
C452 XA.XIR[15].XIC[3].icell.PDM Vbias 0.04058f
C453 XThC.Tn[13] Iout 0.84492f
C454 XThR.Tn[9] XA.XIR[10].XIC[14].icell.SM 0.00121f
C455 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00529f
C456 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.03424f
C457 XA.XIR[5].XIC[12].icell.SM Iout 0.00388f
C458 XA.XIR[7].XIC[10].icell.PDM Vbias 0.04058f
C459 XThR.Tn[10] XA.XIR[11].XIC[3].icell.Ien 0.00321f
C460 XThR.XTB4.Y a_n1049_6699# 0.23756f
C461 XThR.XTB5.Y a_n997_2891# 0.00424f
C462 XThC.XTB6.A VPWR 0.68179f
C463 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C464 XA.XIR[5].XIC_15.icell.Ien Vbias 0.21343f
C465 XA.XIR[1].XIC[11].icell.PDM Vbias 0.04058f
C466 XA.XIR[8].XIC[13].icell.Ien VPWR 0.19065f
C467 XA.XIR[9].XIC[1].icell.PUM Vbias 0.00347f
C468 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.SM 0.00383f
C469 XThC.XTBN.A a_7875_9569# 0.01939f
C470 XA.XIR[15].XIC[6].icell.Ien VPWR 0.32782f
C471 XThC.XTBN.Y XThC.Tn[7] 0.91494f
C472 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C473 XA.XIR[6].XIC[1].icell.PDM VPWR 0.00863f
C474 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Iout 0.00347f
C475 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C476 XA.XIR[0].XIC[9].icell.SM Vbias 0.00701f
C477 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C478 XA.XIR[15].XIC[3].icell.Ien Iout 0.06816f
C479 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.03976f
C480 XA.XIR[12].XIC_dummy_right.icell.PUM Vbias 0.00248f
C481 XThR.XTB7.Y a_n997_2891# 0.00474f
C482 XA.XIR[6].XIC_15.icell.Ien Iout 0.06485f
C483 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.SM 0.00383f
C484 XThC.XTB4.Y XThC.Tn[2] 0.0021f
C485 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.03424f
C486 XA.XIR[7].XIC[10].icell.Ien Iout 0.06483f
C487 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.03424f
C488 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.03976f
C489 XA.XIR[13].XIC[1].icell.SM VPWR 0.00158f
C490 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PDM 0.00604f
C491 XThR.XTB1.Y XThR.Tn[1] 0.0099f
C492 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02701f
C493 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.SM 0.00188f
C494 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00212f
C495 XThR.Tn[10] XA.XIR[10].XIC[14].icell.PDM 0.0033f
C496 XA.XIR[1].XIC[11].icell.Ien Iout 0.06483f
C497 XA.XIR[12].XIC[2].icell.SM VPWR 0.00158f
C498 XA.XIR[7].XIC[12].icell.Ien Vbias 0.21238f
C499 XThC.Tn[4] XThR.Tn[6] 0.28062f
C500 XThC.Tn[6] XThR.Tn[8] 0.28062f
C501 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.SM 0.00188f
C502 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PUM 0.00209f
C503 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.03424f
C504 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02698f
C505 XA.XIR[1].XIC[13].icell.Ien Vbias 0.21238f
C506 XThR.Tn[9] XA.XIR[10].XIC[12].icell.Ien 0.00321f
C507 XA.XIR[11].XIC[4].icell.Ien VPWR 0.19065f
C508 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.SM 0.00383f
C509 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PUM 0.00202f
C510 XA.XIR[4].XIC[2].icell.Ien Vbias 0.21238f
C511 XThC.XTB7.A a_8739_10571# 0.00995f
C512 XA.XIR[10].XIC[6].icell.PUM VPWR 0.01036f
C513 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.03976f
C514 XA.XIR[6].XIC[5].icell.PDM VPWR 0.00863f
C515 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00529f
C516 XA.XIR[3].XIC[3].icell.SM Vbias 0.00701f
C517 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02698f
C518 XA.XIR[6].XIC[2].icell.PDM Iout 0.00112f
C519 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C520 XA.XIR[5].XIC[5].icell.Ien VPWR 0.19065f
C521 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04522f
C522 XA.XIR[7].XIC[13].icell.SM Iout 0.00388f
C523 XA.XIR[2].XIC[7].icell.PDM Vbias 0.04058f
C524 XA.XIR[5].XIC[2].icell.Ien Iout 0.06483f
C525 XA.XIR[14].XIC[8].icell.PDM Vbias 0.04058f
C526 XThC.Tn[7] XThR.Tn[5] 0.28062f
C527 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.0353f
C528 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.03976f
C529 XA.XIR[4].XIC[6].icell.SM VPWR 0.00158f
C530 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PUM 0.00135f
C531 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C532 XA.XIR[13].XIC[7].icell.SM Vbias 0.00701f
C533 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.SM 0.00188f
C534 XA.XIR[4].XIC[3].icell.SM Iout 0.00388f
C535 XA.XIR[3].XIC[9].icell.PUM VPWR 0.01036f
C536 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.03976f
C537 XThR.Tn[12] XA.XIR[13].XIC[10].icell.Ien 0.00321f
C538 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04522f
C539 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00529f
C540 XA.XIR[9].XIC[5].icell.PUM Vbias 0.00347f
C541 XA.XIR[8].XIC[4].icell.PDM VPWR 0.00863f
C542 XThC.Tn[5] XThR.Tn[1] 0.28063f
C543 XThR.Tn[8] XA.XIR[9].XIC[6].icell.Ien 0.00321f
C544 XA.XIR[2].XIC[10].icell.Ien VPWR 0.19065f
C545 XThC.XTBN.Y a_3773_9615# 0.08456f
C546 XA.XIR[14].XIC[11].icell.SM Iout 0.00388f
C547 XThR.XTB7.A XThR.Tn[5] 0.02751f
C548 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Iout 0.00347f
C549 a_6243_9615# Vbias 0.00749f
C550 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00529f
C551 XThR.Tn[11] XA.XIR[12].XIC[0].icell.Ien 0.00352f
C552 XA.XIR[2].XIC[7].icell.Ien Iout 0.06483f
C553 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04522f
C554 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02698f
C555 Vbias data[1] 0.00245f
C556 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C557 XA.XIR[10].XIC[13].icell.PUM Vbias 0.00347f
C558 XA.XIR[14].XIC[8].icell.Ien Iout 0.06483f
C559 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PUM 0.00131f
C560 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11] 0.0033f
C561 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00212f
C562 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04522f
C563 XA.XIR[6].XIC[11].icell.PDM Vbias 0.04058f
C564 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04522f
C565 XA.XIR[9].XIC[11].icell.PDM VPWR 0.00863f
C566 XThR.Tn[4] Iout 1.16627f
C567 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02698f
C568 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.SM 0.00188f
C569 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00212f
C570 a_10051_9569# XThC.Tn[12] 0.00623f
C571 XThC.XTB3.Y a_7875_9569# 0.0061f
C572 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.03976f
C573 XA.XIR[15].XIC[11].icell.PUM Vbias 0.00347f
C574 XA.XIR[9].XIC[8].icell.PDM Iout 0.00112f
C575 XA.XIR[7].XIC[3].icell.PDM Vbias 0.04058f
C576 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02742f
C577 XA.XIR[5].XIC[11].icell.Ien Vbias 0.21238f
C578 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PUM 0.00131f
C579 XA.XIR[13].XIC[12].icell.SM Vbias 0.00701f
C580 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.SM 0.00383f
C581 XA.XIR[3].XIC[14].icell.PDM VPWR 0.00873f
C582 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C583 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C584 XThR.Tn[2] XA.XIR[3].XIC[10].icell.Ien 0.00321f
C585 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.15089f
C586 XA.XIR[1].XIC[4].icell.PDM Vbias 0.04058f
C587 XThR.Tn[6] XA.XIR[7].XIC[12].icell.Ien 0.00321f
C588 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04522f
C589 XA.XIR[2].XIC[13].icell.SM VPWR 0.00158f
C590 XThC.XTB2.Y XThC.Tn[2] 0.01113f
C591 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00529f
C592 XA.XIR[1].XIC[0].icell.PDM VPWR 0.00863f
C593 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13469f
C594 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.SM 0.00383f
C595 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.01406f
C596 XA.XIR[14].XIC[2].icell.PDM VPWR 0.00863f
C597 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04522f
C598 XA.XIR[0].XIC[2].icell.SM Vbias 0.00701f
C599 XA.XIR[12].XIC[10].icell.Ien Vbias 0.21238f
C600 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.002f
C601 XA.XIR[6].XIC[11].icell.Ien Iout 0.06483f
C602 XA.XIR[8].XIC[10].icell.PDM Vbias 0.04058f
C603 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.03976f
C604 XA.XIR[7].XIC[6].icell.Ien VPWR 0.19065f
C605 XA.XIR[14].XIC[13].icell.Ien Iout 0.06483f
C606 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.03424f
C607 XThC.Tn[8] VPWR 6.89944f
C608 XA.XIR[13].XIC[2].icell.PUM VPWR 0.01036f
C609 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PDM 0.00182f
C610 XA.XIR[4].XIC[0].icell.PDM VPWR 0.00863f
C611 XThR.Tn[14] XA.XIR[14].XIC[13].icell.PDM 0.0033f
C612 XA.XIR[1].XIC[7].icell.Ien VPWR 0.19065f
C613 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.15089f
C614 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04522f
C615 XA.XIR[7].XIC[3].icell.Ien Iout 0.06483f
C616 XA.XIR[10].XIC[1].icell.PUM Vbias 0.00347f
C617 XA.XIR[9].XIC[13].icell.Ien VPWR 0.19065f
C618 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.01406f
C619 XA.XIR[6].XIC[13].icell.Ien Vbias 0.21238f
C620 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.03981f
C621 XA.XIR[10].XIC[13].icell.SM Vbias 0.00701f
C622 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04522f
C623 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9] 0.15089f
C624 XThR.Tn[9] XA.XIR[10].XIC[10].icell.SM 0.00121f
C625 XA.XIR[15].XIC_15.icell.SM Vbias 0.00701f
C626 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01776f
C627 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PUM 0.00131f
C628 XThR.Tn[12] XA.XIR[13].XIC[1].icell.SM 0.00121f
C629 XThR.XTB7.A a_n1049_6699# 0.02294f
C630 XA.XIR[1].XIC[4].icell.Ien Iout 0.06483f
C631 XA.XIR[0].XIC[8].icell.PUM VPWR 0.00974f
C632 XThR.XTB7.B data[4] 0.01382f
C633 XThR.Tn[5] XA.XIR[6].XIC[8].icell.Ien 0.00321f
C634 XThR.Tn[2] XA.XIR[3].XIC[13].icell.SM 0.00121f
C635 XThR.XTB5.Y a_n997_1579# 0.00133f
C636 XThC.XTB6.A XThC.XTB7.B 1.47641f
C637 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.01406f
C638 XThC.Tn[4] XThR.Tn[4] 0.28062f
C639 XA.XIR[8].XIC[10].icell.Ien Iout 0.06483f
C640 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.39038f
C641 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06536f
C642 XA.XIR[11].XIC[0].icell.SM Iout 0.00388f
C643 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.03424f
C644 XThR.Tn[11] XA.XIR[12].XIC[4].icell.Ien 0.00321f
C645 XA.XIR[11].XIC[14].icell.Ien Iout 0.06483f
C646 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.03424f
C647 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00529f
C648 XA.XIR[8].XIC[12].icell.Ien Vbias 0.21238f
C649 XA.XIR[15].XIC[5].icell.Ien Vbias 0.17911f
C650 XA.XIR[2].XIC[14].icell.SM Iout 0.00388f
C651 XThR.Tn[11] XA.XIR[11].XIC[7].icell.PDM 0.0033f
C652 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00212f
C653 XA.XIR[3].XIC_15.icell.SM Vbias 0.00701f
C654 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.04037f
C655 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Ien 0.00529f
C656 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.15089f
C657 XThR.XTB7.Y a_n997_1579# 0.013f
C658 XThR.Tn[10] XA.XIR[11].XIC[6].icell.SM 0.00121f
C659 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00529f
C660 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PUM 0.00529f
C661 XThR.XTB2.Y a_n1049_7493# 0.02133f
C662 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.SM 0.00383f
C663 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00212f
C664 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.SM 0.00188f
C665 XThR.Tn[6] XA.XIR[6].XIC[11].icell.PDM 0.0033f
C666 XThR.Tn[3] XA.XIR[4].XIC_15.icell.Ien 0.00116f
C667 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04522f
C668 XThR.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.0033f
C669 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PUM 0.00529f
C670 XA.XIR[3].XIC[2].icell.PUM VPWR 0.01036f
C671 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.03976f
C672 XThR.Tn[5] XA.XIR[6].XIC[11].icell.SM 0.00121f
C673 XA.XIR[4].XIC_15.icell.SM Iout 0.0047f
C674 XA.XIR[12].XIC[1].icell.SM Vbias 0.00701f
C675 XA.XIR[8].XIC[13].icell.SM Iout 0.00388f
C676 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7] 0.0033f
C677 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.01406f
C678 XA.XIR[2].XIC[3].icell.Ien VPWR 0.19065f
C679 XA.XIR[15].XIC[6].icell.SM Iout 0.00388f
C680 XA.XIR[0].XIC[14].icell.PUM Vbias 0.00347f
C681 XThC.Tn[2] Iout 0.85247f
C682 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.03424f
C683 XA.XIR[14].XIC[4].icell.Ien VPWR 0.19119f
C684 XThC.Tn[14] XThR.Tn[11] 0.28068f
C685 XA.XIR[11].XIC[3].icell.Ien Vbias 0.21238f
C686 XThR.Tn[4] XA.XIR[5].XIC_15.icell.Ien 0.00116f
C687 XA.XIR[2].XIC[0].icell.Ien Iout 0.06474f
C688 XThR.XTBN.Y a_n997_715# 0.21503f
C689 XA.XIR[15].XIC[9].icell.Ien Vbias 0.17911f
C690 VPWR data[7] 0.212f
C691 XThR.Tn[0] XA.XIR[1].XIC[10].icell.Ien 0.00321f
C692 XA.XIR[13].XIC[6].icell.PUM VPWR 0.01036f
C693 XThR.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.0033f
C694 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PUM 0.00131f
C695 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C696 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Ien 0.00279f
C697 XA.XIR[10].XIC[5].icell.PUM Vbias 0.00347f
C698 XA.XIR[1].XIC[14].icell.SM VPWR 0.00208f
C699 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.SM 0.00188f
C700 XA.XIR[9].XIC[4].icell.PDM VPWR 0.00863f
C701 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C702 XA.XIR[6].XIC[4].icell.PDM Vbias 0.04058f
C703 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.15089f
C704 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02698f
C705 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00529f
C706 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C707 XA.XIR[12].XIC[7].icell.PUM VPWR 0.01036f
C708 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PUM 0.00529f
C709 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C710 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.SM 0.00383f
C711 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.03976f
C712 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.15089f
C713 XA.XIR[5].XIC[4].icell.Ien Vbias 0.21238f
C714 XA.XIR[0].XIC_15.icell.SM VPWR 0.00258f
C715 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04522f
C716 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.01406f
C717 XA.XIR[11].XIC[7].icell.SM VPWR 0.00158f
C718 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.002f
C719 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PUM 0.00529f
C720 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01734f
C721 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PUM 0.00529f
C722 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.03424f
C723 XThR.Tn[2] XA.XIR[3].XIC[3].icell.Ien 0.00321f
C724 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.15089f
C725 XA.XIR[4].XIC[5].icell.SM Vbias 0.00701f
C726 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.03424f
C727 XA.XIR[11].XIC[4].icell.SM Iout 0.00388f
C728 XThR.Tn[5] XA.XIR[5].XIC[1].icell.PDM 0.0033f
C729 XA.XIR[6].XIC[7].icell.Ien VPWR 0.19065f
C730 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C731 XA.XIR[3].XIC[8].icell.PUM Vbias 0.00347f
C732 XA.XIR[10].XIC[14].icell.PDM Vbias 0.04058f
C733 XA.XIR[10].XIC[8].icell.PDM Iout 0.00112f
C734 XA.XIR[5].XIC[8].icell.SM VPWR 0.00158f
C735 XA.XIR[6].XIC[4].icell.Ien Iout 0.06483f
C736 XA.XIR[8].XIC[3].icell.PDM Vbias 0.04058f
C737 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.SM 0.00188f
C738 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00212f
C739 XThC.XTB3.Y XThC.Tn[4] 0.00382f
C740 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02708f
C741 XA.XIR[2].XIC[9].icell.Ien Vbias 0.21238f
C742 XThR.Tn[0] XA.XIR[1].XIC[13].icell.SM 0.00121f
C743 XThR.XTB7.B XThR.Tn[3] 0.00532f
C744 XA.XIR[5].XIC[5].icell.SM Iout 0.00388f
C745 XA.XIR[10].XIC[9].icell.PUM Vbias 0.00347f
C746 XA.XIR[4].XIC[11].icell.PUM VPWR 0.01036f
C747 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.15089f
C748 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01734f
C749 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.03424f
C750 XThC.Tn[2] XThC.Tn[4] 0.02723f
C751 XThC.Tn[10] XThR.Tn[2] 0.28062f
C752 XA.XIR[15].XIC[12].icell.PDM Vbias 0.04058f
C753 XThC.Tn[8] XThR.Tn[12] 0.28062f
C754 XThC.Tn[14] XThR.Tn[7] 0.28068f
C755 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.03424f
C756 XA.XIR[13].XIC[13].icell.PUM Vbias 0.00347f
C757 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.01406f
C758 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PUM 0.00131f
C759 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PUM 0.00529f
C760 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04522f
C761 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PUM 0.00131f
C762 XThR.XTBN.A VPWR 0.90692f
C763 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C764 XA.XIR[11].XIC[12].icell.SM VPWR 0.00158f
C765 XA.XIR[9].XIC[10].icell.PDM Vbias 0.04058f
C766 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02698f
C767 XA.XIR[0].XIC[1].icell.PUM VPWR 0.00971f
C768 XA.XIR[8].XIC[6].icell.Ien VPWR 0.19065f
C769 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04522f
C770 XA.XIR[15].XIC[0].icell.PDM Iout 0.00112f
C771 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02698f
C772 XThR.Tn[5] XA.XIR[6].XIC[1].icell.Ien 0.00321f
C773 XThR.Tn[8] XA.XIR[9].XIC[9].icell.SM 0.00121f
C774 XA.XIR[3].XIC[11].icell.PDM Iout 0.00112f
C775 a_n1049_5317# VPWR 0.72039f
C776 XA.XIR[8].XIC[3].icell.Ien Iout 0.06483f
C777 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08027f
C778 XA.XIR[11].XIC[8].icell.SM Iout 0.00388f
C779 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.002f
C780 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.01406f
C781 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04522f
C782 XThR.Tn[9] XA.XIR[10].XIC[1].icell.Ien 0.00321f
C783 XA.XIR[2].XIC[10].icell.SM Iout 0.00388f
C784 XA.XIR[11].XIC[1].icell.PDM Vbias 0.04058f
C785 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00212f
C786 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.SM 0.00188f
C787 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PUM 0.00529f
C788 a_n1049_8581# XThR.Tn[0] 0.2685f
C789 XA.XIR[5].XIC[13].icell.PUM VPWR 0.01036f
C790 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08027f
C791 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.15089f
C792 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.SM 0.00188f
C793 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.PDM 0.00584f
C794 XA.XIR[2].XIC[12].icell.SM Vbias 0.00701f
C795 XA.XIR[10].XIC[14].icell.PUM Vbias 0.00347f
C796 XThC.XTBN.A data[1] 0.01444f
C797 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PUM 0.00131f
C798 XA.XIR[15].XIC_dummy_right.icell.PUM Vbias 0.00248f
C799 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.SM 0.00383f
C800 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08017f
C801 XA.XIR[9].XIC[10].icell.Ien Iout 0.06483f
C802 XThC.XTB7.B XThC.Tn[8] 0.09736f
C803 XThR.Tn[3] XA.XIR[4].XIC[11].icell.Ien 0.00321f
C804 XA.XIR[7].XIC[5].icell.Ien Vbias 0.21238f
C805 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.03976f
C806 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.01406f
C807 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02698f
C808 a_8963_9569# Vbias 0.00224f
C809 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.01406f
C810 XThC.XTB7.Y XThC.Tn[12] 0.07222f
C811 XThR.Tn[6] XA.XIR[6].XIC[4].icell.PDM 0.0033f
C812 XA.XIR[13].XIC[1].icell.PUM Vbias 0.00347f
C813 XA.XIR[12].XIC[1].icell.PDM Iout 0.00112f
C814 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.03424f
C815 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02698f
C816 XA.XIR[1].XIC[6].icell.Ien Vbias 0.21238f
C817 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00212f
C818 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.SM 0.00188f
C819 XA.XIR[13].XIC[13].icell.SM Vbias 0.00701f
C820 XA.XIR[9].XIC[12].icell.Ien Vbias 0.21238f
C821 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.01406f
C822 XA.XIR[15].XIC[2].icell.SM VPWR 0.00158f
C823 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PUM 0.00131f
C824 XA.XIR[3].XIC[13].icell.Ien Iout 0.06483f
C825 XA.XIR[12].XIC[2].icell.PUM Vbias 0.00347f
C826 XThR.Tn[7] XA.XIR[7].XIC[9].icell.PDM 0.0033f
C827 XA.XIR[0].XIC[7].icell.PUM Vbias 0.00347f
C828 XA.XIR[6].XIC[14].icell.SM VPWR 0.00208f
C829 XThR.Tn[4] XA.XIR[5].XIC[11].icell.Ien 0.00321f
C830 XThR.Tn[13] XA.XIR[14].XIC[3].icell.Ien 0.00321f
C831 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02698f
C832 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00212f
C833 XA.XIR[7].XIC[9].icell.SM VPWR 0.00158f
C834 XA.XIR[3].XIC_dummy_right.icell.PUM Vbias 0.00248f
C835 XA.XIR[1].XIC[0].icell.PUM VPWR 0.01036f
C836 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C837 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.03424f
C838 XA.XIR[14].XIC[0].icell.SM Iout 0.00388f
C839 XA.XIR[14].XIC[14].icell.Ien Iout 0.06483f
C840 XA.XIR[7].XIC[6].icell.SM Iout 0.00388f
C841 XA.XIR[1].XIC[10].icell.SM VPWR 0.00158f
C842 XThR.Tn[0] XA.XIR[1].XIC[3].icell.Ien 0.00321f
C843 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.03424f
C844 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.03424f
C845 XA.XIR[4].XIC[0].icell.PUM VPWR 0.01036f
C846 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.03424f
C847 XA.XIR[9].XIC[13].icell.SM Iout 0.00388f
C848 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PUM 0.00131f
C849 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PUM 0.00131f
C850 XA.XIR[1].XIC[7].icell.SM Iout 0.00388f
C851 XA.XIR[10].XIC[14].icell.SM Vbias 0.00701f
C852 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04522f
C853 XA.XIR[0].XIC[13].icell.PDM VPWR 0.00806f
C854 XThR.Tn[1] XA.XIR[1].XIC[12].icell.PDM 0.0033f
C855 XA.XIR[5].XIC_dummy_right.icell.Ien Vbias 0.00287f
C856 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00529f
C857 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.01406f
C858 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02698f
C859 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PUM 0.00529f
C860 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.01406f
C861 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.SM 0.00188f
C862 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02698f
C863 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[13].icell.Ien 0.00212f
C864 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PUM 0.00529f
C865 XThR.Tn[11] XA.XIR[12].XIC[7].icell.SM 0.00121f
C866 XA.XIR[10].XIC[4].icell.PDM VPWR 0.00863f
C867 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.03424f
C868 XA.XIR[6].XIC[0].icell.Ien VPWR 0.19066f
C869 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04522f
C870 XThR.Tn[13] XA.XIR[13].XIC[14].icell.PDM 0.0033f
C871 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04522f
C872 XThR.Tn[9] XA.XIR[10].XIC[5].icell.Ien 0.00321f
C873 XThC.Tn[6] VPWR 5.96212f
C874 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.03424f
C875 XA.XIR[11].XIC_15.icell.Ien Iout 0.06485f
C876 XA.XIR[3].XIC[1].icell.PUM Vbias 0.00347f
C877 XA.XIR[7].XIC[14].icell.PUM VPWR 0.01036f
C878 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.03424f
C879 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04522f
C880 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PUM 0.00302f
C881 XA.XIR[5].XIC[1].icell.SM VPWR 0.00158f
C882 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04522f
C883 XA.XIR[2].XIC[2].icell.Ien Vbias 0.21238f
C884 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02698f
C885 XA.XIR[11].XIC[13].icell.PDM Iout 0.00112f
C886 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C887 XThC.Tn[14] XThR.Tn[14] 0.28068f
C888 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04522f
C889 XA.XIR[14].XIC[3].icell.Ien Vbias 0.21238f
C890 XA.XIR[4].XIC[4].icell.PUM VPWR 0.01036f
C891 XThC.Tn[12] XThR.Tn[0] 0.28122f
C892 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.03424f
C893 XThC.Tn[5] XThR.Tn[9] 0.28062f
C894 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.03424f
C895 XA.XIR[13].XIC[5].icell.PUM Vbias 0.00347f
C896 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01681f
C897 XA.XIR[3].XIC[7].icell.PDM VPWR 0.00863f
C898 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00212f
C899 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.SM 0.00188f
C900 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.15089f
C901 XThR.Tn[6] XA.XIR[7].XIC[5].icell.Ien 0.00321f
C902 XThR.XTB7.B XThR.Tn[8] 0.05091f
C903 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C904 XThR.XTBN.A XThR.Tn[12] 0.22096f
C905 XThR.XTB6.Y a_n1049_5611# 0.26831f
C906 XA.XIR[12].XIC[6].icell.PUM Vbias 0.00347f
C907 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C908 XThR.Tn[8] XA.XIR[9].XIC[2].icell.SM 0.00121f
C909 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.0169f
C910 XThR.Tn[11] XA.XIR[12].XIC[12].icell.SM 0.00121f
C911 XA.XIR[3].XIC[4].icell.PDM Iout 0.00112f
C912 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00529f
C913 XThC.XTB3.Y a_6243_9615# 0.00899f
C914 XA.XIR[2].XIC[6].icell.SM VPWR 0.00158f
C915 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.01406f
C916 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC_15.icell.Ien 0.00212f
C917 XA.XIR[14].XIC[7].icell.SM VPWR 0.00158f
C918 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13469f
C919 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02698f
C920 XA.XIR[10].XIC[12].icell.Ien Vbias 0.21238f
C921 XThR.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.00321f
C922 XA.XIR[11].XIC[6].icell.SM Vbias 0.00701f
C923 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04522f
C924 XA.XIR[2].XIC[3].icell.SM Iout 0.00388f
C925 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02698f
C926 XThR.XTBN.Y XThR.Tn[3] 0.62502f
C927 a_n1049_6405# VPWR 0.72117f
C928 XA.XIR[14].XIC[4].icell.SM Iout 0.00388f
C929 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.03976f
C930 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04522f
C931 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04522f
C932 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.03424f
C933 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.0353f
C934 XA.XIR[10].XIC[10].icell.PDM Vbias 0.04058f
C935 XA.XIR[6].XIC[6].icell.Ien Vbias 0.21238f
C936 XA.XIR[9].XIC[6].icell.Ien VPWR 0.19065f
C937 XA.XIR[15].XIC[10].icell.Ien Vbias 0.17911f
C938 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00212f
C939 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.SM 0.00188f
C940 XA.XIR[13].XIC[14].icell.PDM Vbias 0.04058f
C941 XThR.Tn[10] XA.XIR[11].XIC[0].icell.Ien 0.00321f
C942 XA.XIR[13].XIC[8].icell.PDM Iout 0.00112f
C943 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C944 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.38945f
C945 XA.XIR[9].XIC[3].icell.Ien Iout 0.06483f
C946 XThR.Tn[3] XA.XIR[4].XIC[4].icell.Ien 0.00321f
C947 XThR.Tn[0] XThR.Tn[1] 0.238f
C948 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.SM 0.00188f
C949 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.03976f
C950 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00529f
C951 XA.XIR[11].XIC[13].icell.PUM VPWR 0.01036f
C952 XA.XIR[5].XIC[7].icell.SM Vbias 0.00701f
C953 XA.XIR[12].XIC[9].icell.PDM Iout 0.00112f
C954 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.15089f
C955 XA.XIR[13].XIC[9].icell.PUM Vbias 0.00347f
C956 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04522f
C957 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02698f
C958 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C959 XThR.Tn[2] XA.XIR[3].XIC[6].icell.SM 0.00121f
C960 XA.XIR[4].XIC[10].icell.PUM Vbias 0.00347f
C961 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14] 0.0033f
C962 XThC.Tn[3] XThR.Tn[11] 0.28062f
C963 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00212f
C964 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02698f
C965 XA.XIR[6].XIC[10].icell.SM VPWR 0.00158f
C966 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.03424f
C967 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.SM 0.00188f
C968 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00212f
C969 XA.XIR[14].XIC[12].icell.SM VPWR 0.00158f
C970 XA.XIR[11].XIC_dummy_left.icell.Ien Vbias 0.00342f
C971 XThR.Tn[2] XA.XIR[2].XIC[10].icell.PDM 0.0033f
C972 XA.XIR[3].XIC[13].icell.PDM Vbias 0.04058f
C973 XThR.Tn[7] XA.XIR[7].XIC[2].icell.PDM 0.0033f
C974 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00212f
C975 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.SM 0.00188f
C976 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.03424f
C977 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.01406f
C978 XA.XIR[6].XIC[7].icell.SM Iout 0.00388f
C979 XThR.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.00321f
C980 XA.XIR[8].XIC[5].icell.Ien Vbias 0.21238f
C981 XA.XIR[7].XIC[2].icell.SM VPWR 0.00158f
C982 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.SM 0.00383f
C983 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00212f
C984 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04674f
C985 XA.XIR[14].XIC[8].icell.SM Iout 0.00388f
C986 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.03976f
C987 XThC.XTB7.Y a_10915_9569# 0.06874f
C988 XA.XIR[1].XIC[3].icell.SM VPWR 0.00158f
C989 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02698f
C990 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.SM 0.00188f
C991 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00212f
C992 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00529f
C993 XA.XIR[1].XIC[0].icell.SM Iout 0.00388f
C994 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.03976f
C995 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02698f
C996 XA.XIR[4].XIC[13].icell.PDM Iout 0.00112f
C997 XA.XIR[5].XIC[12].icell.PUM Vbias 0.00347f
C998 XA.XIR[13].XIC[14].icell.PUM Vbias 0.00347f
C999 XA.XIR[0].XIC[6].icell.PDM VPWR 0.00812f
C1000 XA.XIR[8].XIC[9].icell.SM VPWR 0.00158f
C1001 XThR.Tn[1] XA.XIR[1].XIC[5].icell.PDM 0.0033f
C1002 XThR.Tn[5] XA.XIR[6].XIC[4].icell.SM 0.00121f
C1003 a_n997_2891# VPWR 0.01372f
C1004 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.03424f
C1005 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01799f
C1006 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04522f
C1007 XA.XIR[11].XIC[13].icell.SM VPWR 0.00158f
C1008 XA.XIR[4].XIC_15.icell.PDM Vbias 0.04206f
C1009 XA.XIR[8].XIC[6].icell.SM Iout 0.00388f
C1010 XThC.Tn[9] XThR.Tn[3] 0.28062f
C1011 XThC.XTB7.A XThC.Tn[7] 0.00184f
C1012 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01776f
C1013 XThR.XTBN.A a_n997_1803# 0.09118f
C1014 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.SM 0.00383f
C1015 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.15089f
C1016 XA.XIR[11].XIC[9].icell.SM Iout 0.00388f
C1017 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.SM 0.00383f
C1018 XThC.Tn[3] XThR.Tn[7] 0.28062f
C1019 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02698f
C1020 XA.XIR[15].XIC[1].icell.SM Vbias 0.00701f
C1021 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.15089f
C1022 XThC.Tn[6] XThR.Tn[12] 0.28062f
C1023 XA.XIR[5].XIC_15.icell.PDM Iout 0.0013f
C1024 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PUM 0.00131f
C1025 XA.XIR[7].XIC[8].icell.SM Vbias 0.00701f
C1026 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.SM 0.00188f
C1027 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04522f
C1028 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.15089f
C1029 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00529f
C1030 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.PUM 0.00112f
C1031 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.SM 0.00188f
C1032 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C1033 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.01406f
C1034 XA.XIR[1].XIC[9].icell.SM Vbias 0.00701f
C1035 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.15089f
C1036 XA.XIR[10].XIC[10].icell.SM Vbias 0.00701f
C1037 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00529f
C1038 XA.XIR[15].XIC[7].icell.PUM VPWR 0.01036f
C1039 XA.XIR[8].XIC[14].icell.PUM VPWR 0.01036f
C1040 XA.XIR[9].XIC[1].icell.Ien Vbias 0.21238f
C1041 XThC.XTBN.A a_8963_9569# 0.01679f
C1042 XThR.Tn[14] XA.XIR[14].XIC[7].icell.PDM 0.0033f
C1043 XA.XIR[13].XIC[14].icell.SM Vbias 0.00701f
C1044 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PUM 0.00209f
C1045 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.01406f
C1046 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.15089f
C1047 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.01406f
C1048 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.002f
C1049 XA.XIR[6].XIC_dummy_left.icell.SM VPWR 0.00269f
C1050 XA.XIR[0].XIC[12].icell.PDM Vbias 0.04065f
C1051 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.15089f
C1052 XThR.Tn[13] XA.XIR[14].XIC[6].icell.SM 0.00121f
C1053 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.SM 0.00188f
C1054 XThC.Tn[5] XThR.Tn[10] 0.28062f
C1055 XThR.Tn[13] XA.XIR[13].XIC[10].icell.PDM 0.0033f
C1056 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.01406f
C1057 XA.XIR[2].XIC_15.icell.SM Iout 0.0047f
C1058 XThR.Tn[0] XA.XIR[1].XIC[6].icell.SM 0.00121f
C1059 XA.XIR[13].XIC[4].icell.PDM VPWR 0.00863f
C1060 XA.XIR[11].XIC[11].icell.Ien Iout 0.06483f
C1061 XThC.XTB7.B XThC.Tn[6] 0.05039f
C1062 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.01406f
C1063 VPWR data[3] 0.20846f
C1064 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C1065 XA.XIR[14].XIC_15.icell.Ien Iout 0.06485f
C1066 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02698f
C1067 XThC.XTB5.Y XThC.Tn[10] 0.01742f
C1068 XA.XIR[12].XIC[5].icell.PDM VPWR 0.00863f
C1069 XA.XIR[7].XIC[13].icell.PUM Vbias 0.00347f
C1070 XThR.XTBN.Y XThR.Tn[8] 0.47815f
C1071 XThR.Tn[0] XA.XIR[0].XIC[9].icell.PDM 0.0033f
C1072 XThC.XTB6.Y XThC.Tn[14] 0.00128f
C1073 XThR.Tn[7] XA.XIR[8].XIC_15.icell.Ien 0.00116f
C1074 XA.XIR[5].XIC[0].icell.SM Vbias 0.00675f
C1075 XA.XIR[1].XIC[14].icell.PUM Vbias 0.00347f
C1076 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.15089f
C1077 XA.XIR[14].XIC[13].icell.PDM Iout 0.00112f
C1078 XThC.XTB5.Y a_4861_9615# 0.0021f
C1079 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.01406f
C1080 XA.XIR[11].XIC[5].icell.PUM VPWR 0.01036f
C1081 XA.XIR[0].XIC[12].icell.Ien Iout 0.06455f
C1082 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00529f
C1083 XThR.XTB6.Y VPWR 1.05511f
C1084 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04522f
C1085 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PUM 0.00131f
C1086 XThR.Tn[14] XA.XIR[14].XIC[11].icell.PDM 0.0033f
C1087 XA.XIR[4].XIC[3].icell.PUM Vbias 0.00347f
C1088 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.01406f
C1089 XA.XIR[10].XIC[6].icell.Ien VPWR 0.19065f
C1090 XA.XIR[6].XIC[3].icell.SM VPWR 0.00158f
C1091 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C1092 XThR.Tn[2] XA.XIR[2].XIC[3].icell.PDM 0.0033f
C1093 XA.XIR[3].XIC[6].icell.PDM Vbias 0.04058f
C1094 XA.XIR[10].XIC[3].icell.Ien Iout 0.06483f
C1095 XA.XIR[5].XIC[6].icell.PUM VPWR 0.01036f
C1096 XA.XIR[6].XIC[0].icell.SM Iout 0.00388f
C1097 XThR.XTB7.B a_n1049_5611# 0.00927f
C1098 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PUM 0.00529f
C1099 XA.XIR[2].XIC[5].icell.SM Vbias 0.00701f
C1100 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C1101 XA.XIR[13].XIC[12].icell.Ien Vbias 0.21238f
C1102 XA.XIR[14].XIC[6].icell.SM Vbias 0.00701f
C1103 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00529f
C1104 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01799f
C1105 XA.XIR[4].XIC[9].icell.PDM VPWR 0.00863f
C1106 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PUM 0.00529f
C1107 XA.XIR[1].XIC_15.icell.SM VPWR 0.00276f
C1108 XA.XIR[11].XIC[14].icell.PDM VPWR 0.00873f
C1109 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00529f
C1110 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C1111 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00212f
C1112 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.SM 0.00188f
C1113 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06536f
C1114 XA.XIR[13].XIC[10].icell.PDM Vbias 0.04058f
C1115 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.01406f
C1116 XThC.XTBN.Y XThC.Tn[10] 0.51405f
C1117 XA.XIR[3].XIC[9].icell.Ien VPWR 0.19065f
C1118 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.SM 0.00383f
C1119 XA.XIR[4].XIC[6].icell.PDM Iout 0.00112f
C1120 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.0353f
C1121 XThR.Tn[6] XA.XIR[7].XIC[8].icell.SM 0.00121f
C1122 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04522f
C1123 XA.XIR[9].XIC[5].icell.Ien Vbias 0.21238f
C1124 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.SM 0.00188f
C1125 XA.XIR[11].XIC[9].icell.PUM VPWR 0.01036f
C1126 XA.XIR[8].XIC[2].icell.SM VPWR 0.00158f
C1127 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00212f
C1128 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00212f
C1129 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PUM 0.00131f
C1130 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01734f
C1131 XA.XIR[2].XIC[11].icell.PUM VPWR 0.01036f
C1132 XA.XIR[3].XIC[6].icell.Ien Iout 0.06483f
C1133 XThC.XTBN.Y a_4861_9615# 0.07601f
C1134 XA.XIR[14].XIC[13].icell.PUM VPWR 0.01036f
C1135 XThR.Tn[10] XA.XIR[10].XIC[12].icell.PDM 0.0033f
C1136 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00529f
C1137 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02698f
C1138 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PUM 0.00131f
C1139 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.15107f
C1140 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[6].icell.Ien 0.00212f
C1141 XA.XIR[0].XIC[1].icell.PDM Vbias 0.04065f
C1142 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.SM 0.00188f
C1143 XThC.Tn[0] XA.XIR[4].XIC_dummy_left.icell.Iout 0.00111f
C1144 XThR.Tn[11] XA.XIR[12].XIC[13].icell.SM 0.00121f
C1145 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06536f
C1146 XThC.Tn[3] XThR.Tn[14] 0.28062f
C1147 XThC.Tn[1] XThR.Tn[0] 0.28118f
C1148 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04522f
C1149 XThR.Tn[1] XA.XIR[2].XIC[10].icell.Ien 0.00321f
C1150 XThR.Tn[9] XA.XIR[10].XIC[10].icell.Ien 0.00321f
C1151 XThC.Tn[9] XThR.Tn[8] 0.28062f
C1152 XA.XIR[9].XIC[9].icell.SM VPWR 0.00158f
C1153 XA.XIR[6].XIC[9].icell.SM Vbias 0.00701f
C1154 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.SM 0.00383f
C1155 XThC.XTB5.Y a_5155_10571# 0.01188f
C1156 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PUM 0.00209f
C1157 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C1158 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.002f
C1159 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.01406f
C1160 XThC.Tn[9] XThC.Tn[11] 0.00252f
C1161 XA.XIR[9].XIC[6].icell.SM Iout 0.00388f
C1162 XThC.XTB3.Y a_8963_9569# 0.002f
C1163 XThR.Tn[3] XA.XIR[4].XIC[7].icell.SM 0.00121f
C1164 XThR.Tn[14] XA.XIR[15].XIC[4].icell.Ien 0.00321f
C1165 XA.XIR[7].XIC[1].icell.SM Vbias 0.00701f
C1166 XThR.XTB7.A data[4] 0.8689f
C1167 XA.XIR[3].XIC[12].icell.SM VPWR 0.00158f
C1168 XA.XIR[1].XIC[2].icell.SM Vbias 0.00701f
C1169 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.SM 0.00188f
C1170 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PUM 0.00131f
C1171 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PUM 0.00131f
C1172 XA.XIR[11].XIC[14].icell.PUM VPWR 0.01036f
C1173 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.SM 0.00188f
C1174 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.SM 0.00188f
C1175 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08017f
C1176 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.SM 0.00383f
C1177 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PUM 0.00529f
C1178 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.15089f
C1179 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PUM 0.00529f
C1180 XA.XIR[0].XIC[5].icell.PDM Vbias 0.04061f
C1181 a_n997_1579# VPWR 0.02422f
C1182 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.SM 0.00383f
C1183 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00529f
C1184 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C1185 XThR.Tn[4] XA.XIR[5].XIC[7].icell.SM 0.00121f
C1186 XA.XIR[14].XIC[13].icell.SM VPWR 0.00158f
C1187 XA.XIR[7].XIC[7].icell.PUM VPWR 0.01036f
C1188 XA.XIR[8].XIC[8].icell.SM Vbias 0.00701f
C1189 XA.XIR[11].XIC[0].icell.Ien Vbias 0.21102f
C1190 XThC.Tn[10] XThR.Tn[5] 0.28062f
C1191 XThR.Tn[8] XA.XIR[8].XIC[12].icell.PDM 0.0033f
C1192 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PUM 0.00529f
C1193 XThR.Tn[1] XA.XIR[2].XIC[13].icell.SM 0.00121f
C1194 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.01406f
C1195 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04522f
C1196 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00212f
C1197 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Ien 0.00529f
C1198 XA.XIR[1].XIC[8].icell.PUM VPWR 0.01036f
C1199 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.SM 0.00383f
C1200 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.SM 0.00188f
C1201 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.SM 0.00383f
C1202 XThR.Tn[1] XA.XIR[1].XIC[0].icell.PDM 0.00336f
C1203 XA.XIR[9].XIC[14].icell.PUM VPWR 0.01036f
C1204 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.SM 0.00383f
C1205 XA.XIR[10].XIC[1].icell.Ien Vbias 0.21238f
C1206 XA.XIR[6].XIC[14].icell.PUM Vbias 0.00347f
C1207 XA.XIR[14].XIC[9].icell.SM Iout 0.00388f
C1208 XA.XIR[4].XIC_15.icell.Ien VPWR 0.25675f
C1209 XThR.Tn[7] XA.XIR[8].XIC[11].icell.Ien 0.00321f
C1210 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PUM 0.00131f
C1211 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.03976f
C1212 XThC.Tn[8] XThR.Tn[1] 0.28062f
C1213 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04522f
C1214 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.SM 0.00188f
C1215 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00212f
C1216 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06536f
C1217 XThR.Tn[0] XA.XIR[0].XIC[2].icell.PDM 0.0033f
C1218 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.15089f
C1219 XA.XIR[0].XIC[8].icell.Ien VPWR 0.19189f
C1220 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PUM 0.00529f
C1221 XA.XIR[10].XIC[11].icell.PUM Vbias 0.00347f
C1222 XA.XIR[12].XIC[0].icell.Ien Iout 0.06474f
C1223 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PUM 0.00131f
C1224 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PUM 0.00529f
C1225 XA.XIR[8].XIC[0].icell.PDM Iout 0.00112f
C1226 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.SM 0.00188f
C1227 XThR.Tn[12] XA.XIR[12].XIC[5].icell.PDM 0.0033f
C1228 XThR.Tn[3] XA.XIR[3].XIC_15.icell.PDM 0.0033f
C1229 XA.XIR[0].XIC[5].icell.Ien Iout 0.06455f
C1230 XA.XIR[2].XIC[0].icell.PUM VPWR 0.01036f
C1231 XA.XIR[11].XIC[3].icell.PDM Iout 0.00112f
C1232 XThR.Tn[5] XA.XIR[5].XIC[12].icell.PDM 0.0033f
C1233 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PUM 0.00131f
C1234 XA.XIR[11].XIC[14].icell.SM VPWR 0.00208f
C1235 XA.XIR[13].XIC[10].icell.SM Vbias 0.00701f
C1236 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C1237 XThR.Tn[9] XA.XIR[10].XIC[1].icell.SM 0.00121f
C1238 XA.XIR[6].XIC_15.icell.SM VPWR 0.00276f
C1239 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00212f
C1240 XA.XIR[15].XIC[6].icell.PUM Vbias 0.00347f
C1241 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PUM 0.00131f
C1242 XA.XIR[8].XIC[13].icell.PUM Vbias 0.00347f
C1243 XA.XIR[1].XIC[2].icell.PDM VPWR 0.00863f
C1244 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.15089f
C1245 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02698f
C1246 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04522f
C1247 XThR.Tn[4] XA.XIR[4].XIC_15.icell.PDM 0.0033f
C1248 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.03976f
C1249 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.03424f
C1250 XThC.Tn[5] XThR.Tn[13] 0.28062f
C1251 XThC.XTB6.A XThC.Tn[1] 0.00411f
C1252 XA.XIR[4].XIC[2].icell.PDM VPWR 0.00863f
C1253 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00212f
C1254 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.03976f
C1255 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00529f
C1256 XA.XIR[10].XIC_15.icell.SM Vbias 0.00701f
C1257 XA.XIR[14].XIC[11].icell.Ien Iout 0.06483f
C1258 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C1259 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04f
C1260 XThC.Tn[7] XThR.Tn[3] 0.28062f
C1261 XA.XIR[3].XIC[2].icell.Ien VPWR 0.19065f
C1262 a_5155_9615# XThC.Tn[3] 0.00508f
C1263 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.11124f
C1264 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04f
C1265 XThR.Tn[6] XA.XIR[7].XIC[1].icell.SM 0.00121f
C1266 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PUM 0.00131f
C1267 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PUM 0.00529f
C1268 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Ien 0.00529f
C1269 XThR.XTB2.Y a_n997_3755# 0.06476f
C1270 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.03982f
C1271 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02698f
C1272 XA.XIR[12].XIC[4].icell.PDM Vbias 0.04058f
C1273 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.15089f
C1274 XA.XIR[2].XIC[4].icell.PUM VPWR 0.01036f
C1275 XA.XIR[15].XIC[9].icell.PDM Iout 0.00112f
C1276 XA.XIR[0].XIC[14].icell.Ien Vbias 0.21246f
C1277 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PUM 0.00131f
C1278 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04522f
C1279 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C1280 XA.XIR[14].XIC[5].icell.PUM VPWR 0.01036f
C1281 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04522f
C1282 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.03976f
C1283 XThR.XTBN.Y a_n1049_5611# 0.0768f
C1284 XA.XIR[11].XIC[4].icell.PUM Vbias 0.00347f
C1285 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.SM 0.00188f
C1286 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.SM 0.00188f
C1287 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00212f
C1288 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.SM 0.00383f
C1289 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PUM 0.00131f
C1290 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04522f
C1291 XA.XIR[13].XIC[6].icell.Ien VPWR 0.19065f
C1292 XA.XIR[7].XIC[1].icell.PDM Iout 0.00112f
C1293 XThR.Tn[1] XA.XIR[2].XIC[3].icell.Ien 0.00321f
C1294 XThR.XTB7.B VPWR 1.67384f
C1295 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00212f
C1296 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.SM 0.00188f
C1297 XThR.XTB7.A XThR.Tn[3] 0.0306f
C1298 XA.XIR[10].XIC[5].icell.Ien Vbias 0.21238f
C1299 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01897f
C1300 XA.XIR[9].XIC[2].icell.SM VPWR 0.00158f
C1301 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00212f
C1302 XA.XIR[6].XIC[2].icell.SM Vbias 0.00701f
C1303 XA.XIR[11].XIC[12].icell.Ien VPWR 0.19065f
C1304 XA.XIR[13].XIC[3].icell.Ien Iout 0.06483f
C1305 XA.XIR[12].XIC[7].icell.Ien VPWR 0.19065f
C1306 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.15089f
C1307 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00529f
C1308 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C1309 XA.XIR[5].XIC[5].icell.PUM Vbias 0.00347f
C1310 XThR.Tn[3] XA.XIR[4].XIC[0].icell.SM 0.00121f
C1311 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PUM 0.00529f
C1312 XThR.XTB6.A XThR.XTBN.A 0.0512f
C1313 XA.XIR[12].XIC[4].icell.Ien Iout 0.06483f
C1314 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04522f
C1315 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00529f
C1316 XA.XIR[11].XIC[10].icell.PDM VPWR 0.00863f
C1317 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.03424f
C1318 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.SM 0.00188f
C1319 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00212f
C1320 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PUM 0.00131f
C1321 XA.XIR[4].XIC[8].icell.PDM Vbias 0.04058f
C1322 XA.XIR[14].XIC[14].icell.PDM VPWR 0.00873f
C1323 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.15089f
C1324 XA.XIR[11].XIC[7].icell.PDM Iout 0.00112f
C1325 XThC.Tn[5] Vbias 2.30671f
C1326 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.01406f
C1327 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00529f
C1328 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PUM 0.00131f
C1329 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.01406f
C1330 XA.XIR[6].XIC[8].icell.PUM VPWR 0.01036f
C1331 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.15089f
C1332 XA.XIR[3].XIC[8].icell.Ien Vbias 0.21238f
C1333 XA.XIR[14].XIC[9].icell.PUM VPWR 0.01036f
C1334 XA.XIR[10].XIC[6].icell.SM Iout 0.00388f
C1335 XA.XIR[8].XIC[1].icell.SM Vbias 0.00701f
C1336 XA.XIR[5].XIC[11].icell.PDM VPWR 0.00863f
C1337 XThR.Tn[4] XA.XIR[5].XIC[0].icell.SM 0.00121f
C1338 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02698f
C1339 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04522f
C1340 XA.XIR[14].XIC[0].icell.PDM Vbias 0.04002f
C1341 XA.XIR[2].XIC[10].icell.PUM Vbias 0.00347f
C1342 XThR.Tn[8] XA.XIR[8].XIC[5].icell.PDM 0.0033f
C1343 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.15089f
C1344 XThR.XTB6.Y a_n997_1803# 0.00871f
C1345 XThC.XTB5.Y a_7651_9569# 0.00418f
C1346 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00212f
C1347 XA.XIR[4].XIC[11].icell.Ien VPWR 0.19065f
C1348 XA.XIR[5].XIC[8].icell.PDM Iout 0.00112f
C1349 XA.XIR[10].XIC[9].icell.Ien Vbias 0.21238f
C1350 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C1351 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.03424f
C1352 XThR.Tn[7] XA.XIR[8].XIC[4].icell.Ien 0.00321f
C1353 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13469f
C1354 a_8963_9569# XA.XIR[0].XIC[10].icell.PDM 0.00281f
C1355 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PUM 0.00529f
C1356 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.SM 0.00383f
C1357 XA.XIR[4].XIC[8].icell.Ien Iout 0.06483f
C1358 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.01406f
C1359 XA.XIR[9].XIC[8].icell.SM Vbias 0.00701f
C1360 XA.XIR[0].XIC[1].icell.Ien VPWR 0.19003f
C1361 XA.XIR[8].XIC[7].icell.PUM VPWR 0.01036f
C1362 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.SM 0.00383f
C1363 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PUM 0.00131f
C1364 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.SM 0.00188f
C1365 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01193f
C1366 XA.XIR[3].XIC[9].icell.SM Iout 0.00388f
C1367 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.03976f
C1368 XThR.XTB3.Y a_n1049_5317# 0.00899f
C1369 XThC.Tn[14] Iout 0.84551f
C1370 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00529f
C1371 XA.XIR[11].XIC[11].icell.PDM Iout 0.00112f
C1372 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02698f
C1373 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[7].icell.SM 0.00383f
C1374 XThR.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.0033f
C1375 XA.XIR[14].XIC[14].icell.PUM VPWR 0.01036f
C1376 XA.XIR[2].XIC[13].icell.PDM Iout 0.00112f
C1377 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PUM 0.00131f
C1378 XA.XIR[3].XIC[11].icell.SM Vbias 0.00701f
C1379 XThR.Tn[11] XA.XIR[12].XIC[14].icell.SM 0.00121f
C1380 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.03424f
C1381 XA.XIR[5].XIC[13].icell.Ien VPWR 0.19065f
C1382 XA.XIR[2].XIC_15.icell.PDM Vbias 0.04206f
C1383 XA.XIR[9].XIC[0].icell.PDM Iout 0.00112f
C1384 XThC.XTBN.Y a_7651_9569# 0.23021f
C1385 XA.XIR[7].XIC[6].icell.PUM Vbias 0.00347f
C1386 XThR.Tn[14] XA.XIR[15].XIC[7].icell.SM 0.00121f
C1387 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.SM 0.00188f
C1388 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00212f
C1389 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.01406f
C1390 a_10051_9569# Vbias 0.00636f
C1391 XA.XIR[10].XIC[12].icell.PDM Vbias 0.04058f
C1392 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02698f
C1393 XA.XIR[13].XIC[1].icell.Ien Vbias 0.21238f
C1394 XA.XIR[4].XIC[11].icell.SM Iout 0.00388f
C1395 XA.XIR[0].XIC[0].icell.PDM Vbias 0.04009f
C1396 XA.XIR[1].XIC[7].icell.PUM Vbias 0.00347f
C1397 XA.XIR[9].XIC[13].icell.PUM Vbias 0.00347f
C1398 XThR.XTB3.Y a_n1335_7243# 0.00941f
C1399 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.0449f
C1400 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01193f
C1401 XThC.XTB4.Y XThC.Tn[3] 0.18952f
C1402 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PUM 0.00529f
C1403 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.15089f
C1404 XThR.Tn[8] XA.XIR[9].XIC[14].icell.Ien 0.00321f
C1405 XA.XIR[13].XIC[11].icell.PUM Vbias 0.00347f
C1406 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.01406f
C1407 XA.XIR[15].XIC[2].icell.PDM Iout 0.00112f
C1408 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01897f
C1409 XA.XIR[0].XIC[7].icell.Ien Vbias 0.21249f
C1410 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PUM 0.00529f
C1411 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.01406f
C1412 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PUM 0.00131f
C1413 XA.XIR[7].XIC[12].icell.PDM VPWR 0.00863f
C1414 XThC.Tn[5] XThR.Tn[6] 0.28062f
C1415 XA.XIR[11].XIC[10].icell.SM VPWR 0.00158f
C1416 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00529f
C1417 XThC.Tn[7] XThR.Tn[8] 0.28062f
C1418 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Iout 0.00347f
C1419 XA.XIR[14].XIC[3].icell.PDM Iout 0.00112f
C1420 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8] 0.0033f
C1421 XA.XIR[5].XIC[0].icell.PDM Iout 0.00112f
C1422 XA.XIR[14].XIC[14].icell.SM VPWR 0.00208f
C1423 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00529f
C1424 XA.XIR[1].XIC[13].icell.PDM VPWR 0.00863f
C1425 XA.XIR[7].XIC[9].icell.PDM Iout 0.00112f
C1426 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.15089f
C1427 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PUM 0.00131f
C1428 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.01406f
C1429 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02698f
C1430 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PUM 0.00529f
C1431 XA.XIR[1].XIC[10].icell.PDM Iout 0.00112f
C1432 XThR.XTB7.B XThR.Tn[12] 0.00772f
C1433 XThR.Tn[14] XA.XIR[15].XIC[12].icell.SM 0.00121f
C1434 XThR.Tn[12] XA.XIR[13].XIC[6].icell.Ien 0.00321f
C1435 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.SM 0.00383f
C1436 XA.XIR[10].XIC_dummy_right.icell.PUM Vbias 0.00248f
C1437 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.01406f
C1438 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.15089f
C1439 XA.XIR[0].XIC[11].icell.SM VPWR 0.00158f
C1440 XA.XIR[4].XIC_dummy_right.icell.SM VPWR 0.00123f
C1441 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PUM 0.00529f
C1442 XThR.Tn[11] XA.XIR[12].XIC[12].icell.Ien 0.00321f
C1443 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.15089f
C1444 XA.XIR[0].XIC[8].icell.SM Iout 0.00367f
C1445 XThC.XTB2.Y a_4067_9615# 0.02133f
C1446 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PDM 0.00594f
C1447 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02698f
C1448 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.01406f
C1449 XA.XIR[0].XIC_dummy_left.icell.Ien Vbias 0.00354f
C1450 XA.XIR[13].XIC_15.icell.SM Vbias 0.00701f
C1451 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.03976f
C1452 XA.XIR[10].XIC[2].icell.SM VPWR 0.00158f
C1453 XA.XIR[6].XIC[1].icell.PUM VPWR 0.01036f
C1454 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Ien 0.00217f
C1455 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04522f
C1456 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PUM 0.00131f
C1457 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.SM 0.00383f
C1458 XA.XIR[3].XIC[1].icell.Ien Vbias 0.21238f
C1459 XA.XIR[7].XIC[14].icell.Ien VPWR 0.1907f
C1460 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PUM 0.00529f
C1461 XThR.XTBN.Y VPWR 4.542f
C1462 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.SM 0.00383f
C1463 XThR.XTB4.Y a_n1049_5611# 0.00465f
C1464 XA.XIR[5].XIC[4].icell.PDM VPWR 0.00863f
C1465 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PUM 0.00529f
C1466 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.15089f
C1467 XA.XIR[2].XIC[3].icell.PUM Vbias 0.00347f
C1468 XA.XIR[14].XIC[4].icell.PUM Vbias 0.00347f
C1469 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.01406f
C1470 XThC.Tn[6] XThR.Tn[1] 0.28063f
C1471 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.SM 0.00383f
C1472 XA.XIR[4].XIC[4].icell.Ien VPWR 0.19065f
C1473 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00529f
C1474 XA.XIR[1].XIC[12].icell.Ien Iout 0.06483f
C1475 XA.XIR[4].XIC[1].icell.Ien Iout 0.06483f
C1476 XA.XIR[13].XIC[5].icell.Ien Vbias 0.21238f
C1477 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PUM 0.00131f
C1478 XA.XIR[3].XIC[5].icell.SM VPWR 0.00158f
C1479 XA.XIR[14].XIC[12].icell.Ien VPWR 0.19119f
C1480 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00212f
C1481 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00212f
C1482 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.SM 0.00188f
C1483 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.SM 0.00188f
C1484 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.SM 0.00188f
C1485 XA.XIR[9].XIC[1].icell.SM Vbias 0.00701f
C1486 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.03976f
C1487 XA.XIR[3].XIC[2].icell.SM Iout 0.00388f
C1488 XA.XIR[12].XIC[6].icell.Ien Vbias 0.21238f
C1489 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.01406f
C1490 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.SM 0.00188f
C1491 XA.XIR[2].XIC[9].icell.PDM VPWR 0.00863f
C1492 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PUM 0.00134f
C1493 XA.XIR[14].XIC[10].icell.PDM VPWR 0.00863f
C1494 a_10051_9569# XThC.Tn[13] 0.19413f
C1495 XA.XIR[11].XIC[9].icell.PDM Vbias 0.04058f
C1496 XA.XIR[2].XIC[6].icell.PDM Iout 0.00112f
C1497 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.SM 0.00383f
C1498 XThR.XTB3.Y a_n1049_6405# 0.00913f
C1499 XA.XIR[14].XIC[7].icell.PDM Iout 0.00112f
C1500 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PUM 0.00529f
C1501 XThR.Tn[1] XA.XIR[2].XIC[6].icell.SM 0.00121f
C1502 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.SM 0.00383f
C1503 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.SM 0.00383f
C1504 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.SM 0.00383f
C1505 XA.XIR[9].XIC[7].icell.PUM VPWR 0.01036f
C1506 XA.XIR[6].XIC[7].icell.PUM Vbias 0.00347f
C1507 XA.XIR[12].XIC[0].icell.PDM VPWR 0.00863f
C1508 XA.XIR[7].XIC_15.icell.Ien Iout 0.06485f
C1509 XThR.Tn[9] XA.XIR[9].XIC[11].icell.PDM 0.0033f
C1510 XThR.Tn[2] XThR.Tn[3] 0.12f
C1511 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.01406f
C1512 XA.XIR[13].XIC[6].icell.SM Iout 0.00388f
C1513 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PUM 0.00131f
C1514 XA.XIR[5].XIC[10].icell.PDM Vbias 0.04058f
C1515 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PUM 0.00131f
C1516 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.SM 0.00383f
C1517 XThR.Tn[13] XA.XIR[13].XIC[12].icell.PDM 0.0033f
C1518 XThR.Tn[14] XA.XIR[15].XIC[0].icell.SM 0.00128f
C1519 XA.XIR[12].XIC[7].icell.SM Iout 0.00388f
C1520 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00529f
C1521 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Iout 0.00347f
C1522 XA.XIR[13].XIC[9].icell.Ien Vbias 0.21238f
C1523 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38579f
C1524 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.SM 0.00383f
C1525 XThR.XTB7.B a_n997_1803# 0.00228f
C1526 XA.XIR[4].XIC[10].icell.Ien Vbias 0.21238f
C1527 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.03976f
C1528 XThC.Tn[9] VPWR 6.88847f
C1529 XThR.Tn[3] XA.XIR[3].XIC[8].icell.PDM 0.0033f
C1530 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00529f
C1531 XA.XIR[6].XIC[13].icell.PDM VPWR 0.00863f
C1532 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00529f
C1533 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04522f
C1534 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.01406f
C1535 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Iout 0.00347f
C1536 XA.XIR[0].XIC[0].icell.Ien Vbias 0.2111f
C1537 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PUM 0.00131f
C1538 XA.XIR[7].XIC[5].icell.PDM VPWR 0.00863f
C1539 XA.XIR[6].XIC[10].icell.PDM Iout 0.00112f
C1540 XA.XIR[8].XIC[6].icell.PUM Vbias 0.00347f
C1541 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.15089f
C1542 XA.XIR[14].XIC[11].icell.PDM Iout 0.00112f
C1543 XThC.Tn[8] XThR.Tn[9] 0.28062f
C1544 XA.XIR[1].XIC[6].icell.PDM VPWR 0.00863f
C1545 XThR.Tn[4] XA.XIR[4].XIC[8].icell.PDM 0.0033f
C1546 XA.XIR[7].XIC[2].icell.PDM Iout 0.00112f
C1547 XA.XIR[5].XIC[10].icell.Ien Iout 0.06483f
C1548 XThR.Tn[11] XA.XIR[12].XIC[10].icell.SM 0.00121f
C1549 XThC.Tn[5] XThR.Tn[4] 0.28062f
C1550 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.15089f
C1551 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06536f
C1552 XThR.Tn[7] XA.XIR[8].XIC[7].icell.SM 0.00121f
C1553 XA.XIR[10].XIC[10].icell.Ien Vbias 0.21238f
C1554 XA.XIR[1].XIC[3].icell.PDM Iout 0.00112f
C1555 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.0353f
C1556 XA.XIR[12].XIC[12].icell.SM Iout 0.00388f
C1557 XA.XIR[5].XIC[12].icell.Ien Vbias 0.21238f
C1558 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00529f
C1559 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PUM 0.00487f
C1560 data[5] data[6] 0.01513f
C1561 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C1562 XA.XIR[0].XIC[4].icell.SM VPWR 0.00158f
C1563 XThR.XTB3.Y a_n997_2891# 0.07285f
C1564 XA.XIR[8].XIC[12].icell.PDM VPWR 0.00863f
C1565 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.SM 0.00383f
C1566 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.03976f
C1567 XA.XIR[11].XIC[1].icell.Ien VPWR 0.19065f
C1568 XA.XIR[4].XIC[13].icell.SM Vbias 0.00701f
C1569 XA.XIR[0].XIC[1].icell.SM Iout 0.00367f
C1570 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00529f
C1571 XA.XIR[8].XIC[9].icell.PDM Iout 0.00112f
C1572 XA.XIR[13].XIC[12].icell.PDM Vbias 0.04058f
C1573 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.15089f
C1574 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00529f
C1575 XThR.XTB5.Y a_n997_3979# 0.00418f
C1576 XA.XIR[2].XIC_15.icell.Ien VPWR 0.25675f
C1577 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PUM 0.00529f
C1578 XA.XIR[11].XIC[11].icell.PUM VPWR 0.01036f
C1579 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.PUM 0.00112f
C1580 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PUM 0.00529f
C1581 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.01405f
C1582 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00529f
C1583 XA.XIR[15].XIC[4].icell.PDM Vbias 0.04058f
C1584 XA.XIR[6].XIC[12].icell.Ien Iout 0.06483f
C1585 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04522f
C1586 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04522f
C1587 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04522f
C1588 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C1589 a_4067_9615# XThC.Tn[4] 0.00141f
C1590 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PUM 0.00209f
C1591 XA.XIR[5].XIC[13].icell.SM Iout 0.00388f
C1592 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.SM 0.00188f
C1593 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PUM 0.00131f
C1594 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00212f
C1595 XA.XIR[14].XIC[10].icell.SM VPWR 0.00158f
C1596 XThR.Tn[10] XA.XIR[11].XIC[4].icell.Ien 0.00321f
C1597 XA.XIR[7].XIC[11].icell.PDM Vbias 0.04058f
C1598 XA.XIR[9].XIC[1].icell.PDM Iout 0.00112f
C1599 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.SM 0.00383f
C1600 XThC.Tn[3] Iout 0.83945f
C1601 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35783f
C1602 XThR.XTB7.Y a_n997_3979# 0.00477f
C1603 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PUM 0.00131f
C1604 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00212f
C1605 XThC.Tn[12] data[3] 0.00161f
C1606 XA.XIR[1].XIC[12].icell.PDM Vbias 0.04058f
C1607 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Iout 0.00347f
C1608 XA.XIR[8].XIC[14].icell.Ien VPWR 0.1907f
C1609 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Ien 0.00529f
C1610 XA.XIR[9].XIC[2].icell.PUM Vbias 0.00347f
C1611 XThC.XTB7.Y Vbias 0.01557f
C1612 XA.XIR[15].XIC[7].icell.Ien VPWR 0.32782f
C1613 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C1614 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PUM 0.00529f
C1615 XThC.XTBN.A a_10051_9569# 0.00199f
C1616 XA.XIR[13].XIC_dummy_right.icell.PUM Vbias 0.00248f
C1617 XThR.Tn[2] XA.XIR[3].XIC_15.icell.Ien 0.00116f
C1618 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PUM 0.00529f
C1619 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PUM 0.00487f
C1620 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PUM 0.00529f
C1621 XA.XIR[15].XIC[4].icell.Ien Iout 0.06816f
C1622 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C1623 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.PUM 0.00112f
C1624 XA.XIR[2].XIC[2].icell.PDM VPWR 0.00863f
C1625 XA.XIR[0].XIC[10].icell.SM Vbias 0.00701f
C1626 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.03976f
C1627 XA.XIR[11].XIC_15.icell.SM VPWR 0.00276f
C1628 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[0].icell.SM 0.00383f
C1629 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.SM 0.00188f
C1630 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.03011f
C1631 XThR.XTB4.Y VPWR 0.92824f
C1632 XThR.XTB7.A a_n1049_5611# 0.01824f
C1633 XA.XIR[7].XIC[11].icell.Ien Iout 0.06483f
C1634 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.03976f
C1635 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04522f
C1636 XA.XIR[13].XIC[2].icell.SM VPWR 0.00158f
C1637 XA.XIR[10].XIC[1].icell.SM Vbias 0.00701f
C1638 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00212f
C1639 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PUM 0.00529f
C1640 XThR.Tn[9] XA.XIR[9].XIC[4].icell.PDM 0.0033f
C1641 XA.XIR[12].XIC[3].icell.SM VPWR 0.00158f
C1642 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12] 0.0033f
C1643 XA.XIR[7].XIC[13].icell.Ien Vbias 0.21238f
C1644 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00212f
C1645 XA.XIR[5].XIC[3].icell.PDM Vbias 0.04058f
C1646 XThR.Tn[14] XA.XIR[15].XIC[13].icell.SM 0.00121f
C1647 XThC.XTB7.A XThC.Tn[10] 0.00406f
C1648 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00212f
C1649 XA.XIR[1].XIC[14].icell.Ien Vbias 0.21238f
C1650 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PUM 0.005f
C1651 XThC.XTB5.Y a_5949_9615# 0.0093f
C1652 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.SM 0.00188f
C1653 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Iout 0.00347f
C1654 XA.XIR[11].XIC[5].icell.Ien VPWR 0.19065f
C1655 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C1656 XThC.XTB3.Y XThC.Tn[5] 0.00384f
C1657 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.03976f
C1658 XA.XIR[4].XIC[3].icell.Ien Vbias 0.21238f
C1659 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.SM 0.00188f
C1660 XThC.XTB7.A a_4861_9615# 0.02294f
C1661 XA.XIR[10].XIC[7].icell.PUM VPWR 0.01036f
C1662 XA.XIR[11].XIC[2].icell.Ien Iout 0.06483f
C1663 XA.XIR[6].XIC[6].icell.PDM VPWR 0.00863f
C1664 XA.XIR[8].XIC_15.icell.Ien Iout 0.06485f
C1665 XThC.Tn[11] XThR.Tn[2] 0.28062f
C1666 XA.XIR[0].XIC[14].icell.SM Vbias 0.00701f
C1667 XThC.Tn[3] XThC.Tn[4] 0.50242f
C1668 XThC.Tn[9] XThR.Tn[12] 0.28062f
C1669 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.SM 0.00188f
C1670 XA.XIR[3].XIC[4].icell.SM Vbias 0.00701f
C1671 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01734f
C1672 XThR.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.00321f
C1673 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.SM 0.00383f
C1674 XA.XIR[5].XIC[6].icell.Ien VPWR 0.19065f
C1675 XA.XIR[6].XIC[3].icell.PDM Iout 0.00112f
C1676 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04522f
C1677 XThR.XTBN.Y XA.XIR[10].XIC_dummy_left.icell.Iout 0.00376f
C1678 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00212f
C1679 XA.XIR[2].XIC[8].icell.PDM Vbias 0.04058f
C1680 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C1681 XA.XIR[14].XIC[9].icell.PDM Vbias 0.04058f
C1682 XA.XIR[5].XIC[3].icell.Ien Iout 0.06483f
C1683 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00529f
C1684 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00212f
C1685 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.03011f
C1686 XA.XIR[4].XIC[7].icell.SM VPWR 0.00158f
C1687 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.15089f
C1688 XThR.Tn[7] XA.XIR[8].XIC[0].icell.SM 0.00121f
C1689 XThR.XTBN.Y a_n997_1803# 0.22873f
C1690 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01799f
C1691 XThR.Tn[0] Vbias 3.72674f
C1692 XA.XIR[4].XIC[4].icell.SM Iout 0.00388f
C1693 XThR.XTBN.A XThR.Tn[9] 0.12398f
C1694 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.03976f
C1695 XA.XIR[3].XIC[10].icell.PUM VPWR 0.01036f
C1696 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.SM 0.00383f
C1697 XA.XIR[8].XIC[5].icell.PDM VPWR 0.00863f
C1698 XA.XIR[9].XIC[6].icell.PUM Vbias 0.00347f
C1699 XA.XIR[11].XIC[9].icell.Ien VPWR 0.19065f
C1700 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04522f
C1701 XThC.XTBN.Y a_5949_9615# 0.0768f
C1702 XThR.Tn[8] XA.XIR[9].XIC[7].icell.Ien 0.00321f
C1703 XA.XIR[2].XIC[11].icell.Ien VPWR 0.19065f
C1704 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02698f
C1705 XThC.Tn[8] XThR.Tn[10] 0.28062f
C1706 XThR.Tn[11] XA.XIR[12].XIC[1].icell.Ien 0.00321f
C1707 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06536f
C1708 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PUM 0.00502f
C1709 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Iout 0.00347f
C1710 XThC.XTB7.B XThC.Tn[9] 0.09572f
C1711 XA.XIR[2].XIC[8].icell.Ien Iout 0.06483f
C1712 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_15.icell.SM 0.00383f
C1713 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00529f
C1714 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00529f
C1715 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04522f
C1716 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04522f
C1717 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PUM 0.00131f
C1718 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.SM 0.00383f
C1719 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.0353f
C1720 XThC.XTB7.Y XThC.Tn[13] 0.11626f
C1721 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PUM 0.00131f
C1722 XA.XIR[9].XIC[12].icell.PDM VPWR 0.00863f
C1723 XA.XIR[6].XIC[12].icell.PDM Vbias 0.04058f
C1724 XThR.Tn[0] XA.XIR[1].XIC_15.icell.Ien 0.00116f
C1725 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00529f
C1726 XA.XIR[12].XIC[0].icell.PUM VPWR 0.01036f
C1727 XThC.XTB5.A XThC.XTBN.Y 0.00282f
C1728 XA.XIR[4].XIC[12].icell.PUM VPWR 0.01036f
C1729 XA.XIR[9].XIC[9].icell.PDM Iout 0.00112f
C1730 XA.XIR[7].XIC[4].icell.PDM Vbias 0.04058f
C1731 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.03976f
C1732 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PUM 0.00131f
C1733 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PUM 0.00529f
C1734 XA.XIR[3].XIC_15.icell.PDM VPWR 0.06959f
C1735 XThR.Tn[2] XA.XIR[3].XIC[11].icell.Ien 0.00321f
C1736 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02698f
C1737 XThR.Tn[6] XA.XIR[7].XIC[13].icell.Ien 0.00321f
C1738 XThR.Tn[8] a_n997_3979# 0.1927f
C1739 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.15089f
C1740 XA.XIR[1].XIC[5].icell.PDM Vbias 0.04058f
C1741 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00529f
C1742 XA.XIR[13].XIC[10].icell.Ien Vbias 0.21238f
C1743 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.01406f
C1744 XA.XIR[15].XIC[0].icell.Ien VPWR 0.32783f
C1745 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.03424f
C1746 XA.XIR[11].XIC[12].icell.PDM VPWR 0.00863f
C1747 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04522f
C1748 XA.XIR[0].XIC[3].icell.SM Vbias 0.00701f
C1749 XA.XIR[14].XIC[1].icell.Ien VPWR 0.19119f
C1750 XA.XIR[10].XIC[1].icell.PDM Iout 0.00112f
C1751 XA.XIR[8].XIC[11].icell.PDM Vbias 0.04058f
C1752 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.03976f
C1753 XA.XIR[2].XIC[11].icell.SM Iout 0.00388f
C1754 XA.XIR[7].XIC[7].icell.Ien VPWR 0.19065f
C1755 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.01406f
C1756 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02698f
C1757 XA.XIR[11].XIC[1].icell.PUM Vbias 0.00347f
C1758 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02698f
C1759 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.SM 0.00383f
C1760 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04f
C1761 XA.XIR[9].XIC[14].icell.Ien VPWR 0.1907f
C1762 XA.XIR[1].XIC[8].icell.Ien VPWR 0.19065f
C1763 XA.XIR[7].XIC[4].icell.Ien Iout 0.06483f
C1764 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.15089f
C1765 XA.XIR[6].XIC[14].icell.Ien Vbias 0.21238f
C1766 XA.XIR[14].XIC[11].icell.PUM VPWR 0.01036f
C1767 XA.XIR[10].XIC[2].icell.PUM Vbias 0.00347f
C1768 XThR.XTB4.Y XThR.Tn[12] 0.00209f
C1769 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04522f
C1770 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.03424f
C1771 XThR.Tn[12] XA.XIR[13].XIC[2].icell.SM 0.00121f
C1772 XA.XIR[1].XIC[5].icell.Ien Iout 0.06483f
C1773 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01734f
C1774 XThR.Tn[3] XA.XIR[4].XIC[12].icell.Ien 0.00321f
C1775 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PUM 0.00131f
C1776 XA.XIR[0].XIC[9].icell.PUM VPWR 0.00971f
C1777 XThC.Tn[7] VPWR 6.34857f
C1778 XA.XIR[8].XIC[1].icell.PDM VPWR 0.00863f
C1779 XA.XIR[3].XIC[0].icell.PDM Iout 0.00112f
C1780 XThR.Tn[5] XA.XIR[6].XIC[9].icell.Ien 0.00321f
C1781 XA.XIR[12].XIC[13].icell.SM Iout 0.00388f
C1782 XA.XIR[8].XIC[11].icell.Ien Iout 0.06483f
C1783 XThR.Tn[11] Iout 1.16629f
C1784 XThC.XTB6.A Vbias 0.00608f
C1785 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00212f
C1786 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.SM 0.00188f
C1787 XThR.Tn[8] XA.XIR[9].XIC[14].icell.SM 0.00121f
C1788 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04522f
C1789 XThR.Tn[11] XA.XIR[12].XIC[5].icell.Ien 0.00321f
C1790 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01897f
C1791 XThC.Tn[13] XThR.Tn[0] 0.28124f
C1792 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00212f
C1793 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.03976f
C1794 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.SM 0.00188f
C1795 XA.XIR[8].XIC[13].icell.Ien Vbias 0.21238f
C1796 XA.XIR[2].XIC_dummy_right.icell.SM VPWR 0.00123f
C1797 XA.XIR[15].XIC[6].icell.Ien Vbias 0.17911f
C1798 XThR.Tn[4] XA.XIR[5].XIC[12].icell.Ien 0.00321f
C1799 XThR.Tn[11] XA.XIR[11].XIC[8].icell.PDM 0.0033f
C1800 XThC.Tn[6] XThR.Tn[9] 0.28062f
C1801 XThR.XTB7.A VPWR 0.88601f
C1802 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PUM 0.00131f
C1803 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.15089f
C1804 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.SM 0.00188f
C1805 XA.XIR[14].XIC_15.icell.SM VPWR 0.00276f
C1806 XA.XIR[6].XIC[1].icell.PDM Vbias 0.04058f
C1807 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C1808 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.SM 0.00383f
C1809 XThR.XTB7.B XThR.XTB6.A 1.47641f
C1810 XA.XIR[1].XIC[11].icell.SM VPWR 0.00158f
C1811 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PUM 0.00529f
C1812 XThR.Tn[10] XA.XIR[11].XIC[7].icell.SM 0.00121f
C1813 XA.XIR[4].XIC[0].icell.SM VPWR 0.00158f
C1814 a_5949_10571# VPWR 0.00653f
C1815 XThR.Tn[6] XA.XIR[6].XIC[12].icell.PDM 0.0033f
C1816 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.SM 0.00383f
C1817 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.01406f
C1818 XThR.Tn[1] XA.XIR[1].XIC[2].icell.PDM 0.0033f
C1819 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PUM 0.00131f
C1820 XA.XIR[9].XIC_15.icell.Ien Iout 0.06485f
C1821 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.SM 0.00188f
C1822 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06536f
C1823 XA.XIR[13].XIC[1].icell.SM Vbias 0.00701f
C1824 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.03424f
C1825 XA.XIR[3].XIC[3].icell.PUM VPWR 0.01036f
C1826 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.03976f
C1827 XThR.Tn[5] XA.XIR[6].XIC[12].icell.SM 0.00121f
C1828 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.03424f
C1829 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00529f
C1830 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.SM 0.00383f
C1831 XThC.XTB4.Y data[2] 0.0086f
C1832 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.SM 0.00383f
C1833 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C1834 XA.XIR[12].XIC[2].icell.SM Vbias 0.00701f
C1835 XThC.XTB6.A a_7331_10587# 0.00304f
C1836 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.SM 0.00383f
C1837 XA.XIR[15].XIC[7].icell.SM Iout 0.00388f
C1838 XA.XIR[2].XIC[4].icell.Ien VPWR 0.19065f
C1839 XA.XIR[8].XIC[2].icell.PDM Iout 0.00112f
C1840 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.SM 0.00383f
C1841 XThR.Tn[11] XA.XIR[12].XIC[9].icell.Ien 0.00321f
C1842 XA.XIR[14].XIC[5].icell.Ien VPWR 0.19119f
C1843 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.SM 0.00188f
C1844 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00529f
C1845 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00529f
C1846 XA.XIR[2].XIC[1].icell.Ien Iout 0.06483f
C1847 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.SM 0.00383f
C1848 XA.XIR[11].XIC[4].icell.Ien Vbias 0.21238f
C1849 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C1850 XA.XIR[7].XIC[14].icell.SM VPWR 0.00208f
C1851 XA.XIR[14].XIC[2].icell.Ien Iout 0.06483f
C1852 XThR.Tn[0] XA.XIR[1].XIC[11].icell.Ien 0.00321f
C1853 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02698f
C1854 XThR.Tn[7] Iout 1.16628f
C1855 XThR.XTBN.A XThR.Tn[10] 0.12147f
C1856 XA.XIR[13].XIC[7].icell.PUM VPWR 0.01036f
C1857 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PUM 0.00131f
C1858 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.01406f
C1859 XA.XIR[6].XIC[5].icell.PDM Vbias 0.04058f
C1860 XThR.Tn[10] XA.XIR[11].XIC[12].icell.SM 0.00121f
C1861 XA.XIR[9].XIC[5].icell.PDM VPWR 0.00863f
C1862 XA.XIR[10].XIC[6].icell.PUM Vbias 0.00347f
C1863 XThC.Tn[4] XThR.Tn[11] 0.28062f
C1864 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.15089f
C1865 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.01406f
C1866 XA.XIR[12].XIC[8].icell.PUM VPWR 0.01036f
C1867 XThR.XTBN.Y XA.XIR[13].XIC_dummy_left.icell.Iout 0.0045f
C1868 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.15089f
C1869 XA.XIR[5].XIC[5].icell.Ien Vbias 0.21238f
C1870 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.03976f
C1871 a_3773_9615# VPWR 0.70508f
C1872 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.03424f
C1873 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00212f
C1874 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.SM 0.00383f
C1875 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.01406f
C1876 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04522f
C1877 XThR.Tn[2] XA.XIR[3].XIC[4].icell.Ien 0.00321f
C1878 XThR.Tn[14] XA.XIR[15].XIC[14].icell.SM 0.00121f
C1879 XThR.XTB2.Y data[5] 0.017f
C1880 XA.XIR[4].XIC[6].icell.SM Vbias 0.00701f
C1881 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.15089f
C1882 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.0353f
C1883 XA.XIR[15].XIC[12].icell.SM Iout 0.00388f
C1884 XA.XIR[11].XIC[5].icell.SM Iout 0.00388f
C1885 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06536f
C1886 XA.XIR[6].XIC[8].icell.Ien VPWR 0.19065f
C1887 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04522f
C1888 XThC.XTB4.Y a_5155_9615# 0.01546f
C1889 XThR.XTBN.Y a_n1049_8581# 0.0607f
C1890 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.03976f
C1891 XA.XIR[3].XIC[9].icell.PUM Vbias 0.00347f
C1892 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02698f
C1893 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00529f
C1894 XA.XIR[14].XIC[9].icell.Ien VPWR 0.19119f
C1895 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04522f
C1896 XA.XIR[10].XIC[9].icell.PDM Iout 0.00112f
C1897 XA.XIR[8].XIC[4].icell.PDM Vbias 0.04058f
C1898 XA.XIR[6].XIC[5].icell.Ien Iout 0.06483f
C1899 XA.XIR[7].XIC[0].icell.Ien VPWR 0.19066f
C1900 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.03976f
C1901 XA.XIR[5].XIC[9].icell.SM VPWR 0.00158f
C1902 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.SM 0.00383f
C1903 XThC.Tn[8] XThR.Tn[13] 0.28062f
C1904 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.03976f
C1905 XA.XIR[2].XIC[10].icell.Ien Vbias 0.21238f
C1906 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04522f
C1907 XThC.XTB5.Y a_8739_9569# 0.00424f
C1908 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04522f
C1909 XA.XIR[5].XIC[6].icell.SM Iout 0.00388f
C1910 XA.XIR[1].XIC[1].icell.Ien VPWR 0.19065f
C1911 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.15089f
C1912 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11595f
C1913 XA.XIR[12].XIC[14].icell.PDM Iout 0.00112f
C1914 XThC.Tn[10] XThR.Tn[3] 0.28062f
C1915 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04522f
C1916 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02698f
C1917 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PUM 0.00131f
C1918 XThR.Tn[6] XA.XIR[6].XIC[1].icell.PDM 0.0033f
C1919 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.03424f
C1920 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00212f
C1921 XA.XIR[0].XIC[2].icell.PUM VPWR 0.00971f
C1922 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.PUM 0.00112f
C1923 XA.XIR[8].XIC[7].icell.Ien VPWR 0.19065f
C1924 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00212f
C1925 XA.XIR[9].XIC[11].icell.PDM Vbias 0.04058f
C1926 XThC.Tn[0] XThR.Tn[2] 0.28071f
C1927 XThC.Tn[4] XThR.Tn[7] 0.28062f
C1928 XThR.Tn[5] XA.XIR[6].XIC[2].icell.Ien 0.00321f
C1929 XA.XIR[15].XIC_dummy_left.icell.SM VPWR 0.00269f
C1930 XThR.Tn[8] XA.XIR[9].XIC[10].icell.SM 0.00121f
C1931 XA.XIR[3].XIC[12].icell.PDM Iout 0.00112f
C1932 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C1933 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.01406f
C1934 XA.XIR[11].XIC[10].icell.Ien VPWR 0.19065f
C1935 XThC.Tn[7] XThR.Tn[12] 0.28062f
C1936 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PUM 0.00529f
C1937 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04522f
C1938 XA.XIR[8].XIC[4].icell.Ien Iout 0.06483f
C1939 XA.XIR[6].XIC[11].icell.SM VPWR 0.00158f
C1940 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00212f
C1941 XA.XIR[3].XIC[14].icell.PDM Vbias 0.04058f
C1942 XA.XIR[5].XIC[14].icell.PUM VPWR 0.01036f
C1943 XThR.Tn[14] XA.XIR[15].XIC[12].icell.Ien 0.00321f
C1944 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00212f
C1945 XA.XIR[2].XIC[13].icell.SM Vbias 0.00701f
C1946 XA.XIR[14].XIC[12].icell.PDM VPWR 0.00863f
C1947 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.SM 0.00188f
C1948 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02698f
C1949 XA.XIR[1].XIC[0].icell.PDM Vbias 0.04002f
C1950 XA.XIR[13].XIC[1].icell.PDM Iout 0.00112f
C1951 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02698f
C1952 XThC.XTBN.Y a_8739_9569# 0.22804f
C1953 XA.XIR[14].XIC[2].icell.PDM Vbias 0.04058f
C1954 XA.XIR[7].XIC[6].icell.Ien Vbias 0.21238f
C1955 XA.XIR[9].XIC[11].icell.Ien Iout 0.06483f
C1956 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.03976f
C1957 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04522f
C1958 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Iout 0.00347f
C1959 XThR.Tn[6] XA.XIR[6].XIC[5].icell.PDM 0.0033f
C1960 XThC.Tn[8] Vbias 2.30737f
C1961 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.39054f
C1962 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C1963 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C1964 XA.XIR[4].XIC[14].icell.PDM Iout 0.00112f
C1965 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00529f
C1966 XA.XIR[4].XIC[0].icell.PDM Vbias 0.04002f
C1967 XA.XIR[13].XIC[2].icell.PUM Vbias 0.00347f
C1968 XThR.Tn[10] XA.XIR[10].XIC[4].icell.PDM 0.0033f
C1969 XA.XIR[1].XIC[7].icell.Ien Vbias 0.21238f
C1970 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PUM 0.00529f
C1971 XA.XIR[9].XIC[13].icell.Ien Vbias 0.21238f
C1972 XA.XIR[15].XIC[3].icell.SM VPWR 0.00158f
C1973 XThC.Tn[6] XThR.Tn[10] 0.28062f
C1974 XA.XIR[3].XIC[14].icell.Ien Iout 0.06483f
C1975 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.03424f
C1976 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PUM 0.00529f
C1977 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04522f
C1978 XThC.XTB7.B XThC.Tn[7] 0.0847f
C1979 XThR.Tn[7] XA.XIR[7].XIC[10].icell.PDM 0.0033f
C1980 XA.XIR[4].XIC_15.icell.PUM Vbias 0.00347f
C1981 XA.XIR[15].XIC[0].icell.SM Iout 0.00388f
C1982 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Iout 0.00347f
C1983 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.01406f
C1984 XThR.XTB1.Y bias[2] 0.00266f
C1985 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00212f
C1986 XThC.XTB5.Y XThC.Tn[11] 0.02206f
C1987 XA.XIR[0].XIC[8].icell.PUM Vbias 0.00347f
C1988 XThR.Tn[13] XA.XIR[14].XIC[4].icell.Ien 0.00321f
C1989 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35783f
C1990 XA.XIR[7].XIC[10].icell.SM VPWR 0.00158f
C1991 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.SM 0.00188f
C1992 XA.XIR[5].XIC[1].icell.PDM VPWR 0.00863f
C1993 XThR.Tn[14] Iout 1.16628f
C1994 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C1995 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01897f
C1996 XA.XIR[6].XIC_dummy_left.icell.Ien Vbias 0.00342f
C1997 XThR.Tn[0] XA.XIR[1].XIC[4].icell.Ien 0.00321f
C1998 XA.XIR[7].XIC[7].icell.SM Iout 0.00388f
C1999 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.SM 0.00188f
C2000 a_8739_9569# XThC.Tn[10] 0.19671f
C2001 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Ien 0.00529f
C2002 a_n1049_6699# XThR.XTB5.Y 0.0021f
C2003 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.03424f
C2004 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PUM 0.00131f
C2005 XA.XIR[1].XIC[8].icell.SM Iout 0.00388f
C2006 XA.XIR[0].XIC[14].icell.PDM VPWR 0.00816f
C2007 XA.XIR[9].XIC[0].icell.Ien Iout 0.06474f
C2008 XThR.Tn[1] XA.XIR[1].XIC[13].icell.PDM 0.0033f
C2009 XThR.Tn[3] a_n1049_6699# 0.27008f
C2010 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PUM 0.00529f
C2011 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.03424f
C2012 XA.XIR[11].XIC[1].icell.SM VPWR 0.00158f
C2013 XThC.XTB2.Y a_5155_9615# 0.00847f
C2014 XA.XIR[8].XIC[14].icell.SM VPWR 0.00208f
C2015 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C2016 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02698f
C2017 XA.XIR[3].XIC[1].icell.PDM Iout 0.00112f
C2018 XA.XIR[12].XIC[14].icell.SM Iout 0.00388f
C2019 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C2020 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.01406f
C2021 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.15089f
C2022 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.03424f
C2023 XA.XIR[10].XIC[5].icell.PDM VPWR 0.00863f
C2024 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C2025 XA.XIR[6].XIC[1].icell.Ien VPWR 0.19065f
C2026 XThR.Tn[9] XA.XIR[10].XIC[6].icell.Ien 0.00321f
C2027 XA.XIR[3].XIC[2].icell.PUM Vbias 0.00347f
C2028 XThC.XTB6.A XThC.XTBN.A 0.0513f
C2029 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.03424f
C2030 XThC.XTBN.Y XThC.Tn[11] 0.53369f
C2031 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00212f
C2032 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00529f
C2033 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00212f
C2034 XA.XIR[5].XIC[2].icell.SM VPWR 0.00158f
C2035 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.03424f
C2036 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PUM 0.00131f
C2037 XA.XIR[2].XIC[3].icell.Ien Vbias 0.21238f
C2038 XThR.Tn[2] VPWR 6.70644f
C2039 XThR.XTBN.Y XThR.Tn[1] 0.61095f
C2040 XA.XIR[5].XIC[2].icell.PDM Iout 0.00112f
C2041 XA.XIR[14].XIC[4].icell.Ien Vbias 0.21238f
C2042 XA.XIR[4].XIC[5].icell.PUM VPWR 0.01036f
C2043 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00529f
C2044 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.01406f
C2045 XThR.XTBN.A XThR.Tn[13] 0.00106f
C2046 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02698f
C2047 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04522f
C2048 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.SM 0.00188f
C2049 XA.XIR[13].XIC[6].icell.PUM Vbias 0.00347f
C2050 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00212f
C2051 XThR.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.00321f
C2052 XThC.Tn[4] XThR.Tn[14] 0.28062f
C2053 XA.XIR[3].XIC[8].icell.PDM VPWR 0.00863f
C2054 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02698f
C2055 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04522f
C2056 XA.XIR[9].XIC[4].icell.PDM Vbias 0.04058f
C2057 XThC.Tn[2] XThR.Tn[0] 0.28238f
C2058 XThC.Tn[8] XThR.Tn[6] 0.28062f
C2059 XA.XIR[1].XIC[14].icell.SM Vbias 0.00701f
C2060 XThC.Tn[10] XThR.Tn[8] 0.28062f
C2061 XThR.Tn[8] XA.XIR[9].XIC[3].icell.SM 0.00121f
C2062 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04522f
C2063 XA.XIR[3].XIC[5].icell.PDM Iout 0.00112f
C2064 XA.XIR[12].XIC[7].icell.PUM Vbias 0.00347f
C2065 XA.XIR[2].XIC[7].icell.SM VPWR 0.00158f
C2066 XThR.Tn[14] XA.XIR[15].XIC[10].icell.SM 0.00121f
C2067 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00529f
C2068 XThC.Tn[10] XThC.Tn[11] 0.10442f
C2069 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04522f
C2070 XA.XIR[2].XIC[4].icell.SM Iout 0.00388f
C2071 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.03424f
C2072 XA.XIR[0].XIC_15.icell.SM Vbias 0.00701f
C2073 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02698f
C2074 XA.XIR[11].XIC[7].icell.SM Vbias 0.00701f
C2075 XA.XIR[7].XIC_dummy_left.icell.SM VPWR 0.00269f
C2076 XThC.XTB6.Y a_7875_9569# 0.0046f
C2077 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.01406f
C2078 XThR.Tn[11] XA.XIR[12].XIC[10].icell.Ien 0.00321f
C2079 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00212f
C2080 XA.XIR[14].XIC[5].icell.SM Iout 0.00388f
C2081 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.SM 0.00188f
C2082 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.03424f
C2083 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.03976f
C2084 XA.XIR[9].XIC[7].icell.Ien VPWR 0.19065f
C2085 XA.XIR[6].XIC[7].icell.Ien Vbias 0.21238f
C2086 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C2087 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C2088 XA.XIR[12].XIC[12].icell.Ien Iout 0.06483f
C2089 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PUM 0.00529f
C2090 XA.XIR[13].XIC[9].icell.PDM Iout 0.00112f
C2091 XThR.Tn[10] a_n997_2891# 0.1927f
C2092 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01421f
C2093 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Iout 0.00347f
C2094 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.01406f
C2095 XThR.Tn[10] XA.XIR[11].XIC[13].icell.SM 0.00121f
C2096 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.SM 0.00383f
C2097 XA.XIR[9].XIC[4].icell.Ien Iout 0.06483f
C2098 XThR.Tn[3] XA.XIR[4].XIC[5].icell.Ien 0.00321f
C2099 XA.XIR[5].XIC[8].icell.SM Vbias 0.00701f
C2100 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.03976f
C2101 XA.XIR[12].XIC[10].icell.PDM Iout 0.00112f
C2102 XThC.Tn[11] XThR.Tn[5] 0.28062f
C2103 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00212f
C2104 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.SM 0.00188f
C2105 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PUM 0.00535f
C2106 XThR.Tn[2] XA.XIR[3].XIC[7].icell.SM 0.00121f
C2107 XA.XIR[4].XIC[11].icell.PUM Vbias 0.00347f
C2108 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.SM 0.00188f
C2109 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.01406f
C2110 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.SM 0.00188f
C2111 XThR.Tn[7] XA.XIR[7].XIC[3].icell.PDM 0.0033f
C2112 XA.XIR[2].XIC[12].icell.PUM VPWR 0.01036f
C2113 XThR.Tn[2] XA.XIR[2].XIC[11].icell.PDM 0.0033f
C2114 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02698f
C2115 XA.XIR[15].XIC[13].icell.SM Iout 0.00388f
C2116 XA.XIR[11].XIC[12].icell.SM Vbias 0.00701f
C2117 XA.XIR[8].XIC[6].icell.Ien Vbias 0.21238f
C2118 XA.XIR[0].XIC[1].icell.PUM Vbias 0.00347f
C2119 XA.XIR[6].XIC[8].icell.SM Iout 0.00388f
C2120 XA.XIR[7].XIC[3].icell.SM VPWR 0.00158f
C2121 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00212f
C2122 XThR.Tn[4] XA.XIR[5].XIC[5].icell.Ien 0.00321f
C2123 XThC.Tn[9] XThR.Tn[1] 0.28062f
C2124 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.SM 0.00188f
C2125 XA.XIR[14].XIC[10].icell.Ien VPWR 0.19119f
C2126 a_n997_3979# VPWR 0.01671f
C2127 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.SM 0.00188f
C2128 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00212f
C2129 XA.XIR[7].XIC[0].icell.SM Iout 0.00388f
C2130 XA.XIR[1].XIC[4].icell.SM VPWR 0.00158f
C2131 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C2132 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.SM 0.00188f
C2133 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.SM 0.00188f
C2134 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.03976f
C2135 XA.XIR[12].XIC[2].icell.PDM VPWR 0.00863f
C2136 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PUM 0.00529f
C2137 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.01406f
C2138 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00212f
C2139 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.0353f
C2140 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01799f
C2141 XA.XIR[1].XIC[1].icell.SM Iout 0.00388f
C2142 XA.XIR[5].XIC[13].icell.PUM Vbias 0.00347f
C2143 XA.XIR[0].XIC[7].icell.PDM VPWR 0.00806f
C2144 XThR.XTB5.A data[5] 0.11096f
C2145 XThC.XTB4.Y a_7875_9569# 0.00497f
C2146 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.03594f
C2147 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04522f
C2148 XThR.Tn[1] XA.XIR[1].XIC[6].icell.PDM 0.0033f
C2149 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02698f
C2150 XA.XIR[8].XIC[10].icell.SM VPWR 0.00158f
C2151 XThR.Tn[5] XA.XIR[6].XIC[5].icell.SM 0.00121f
C2152 XA.XIR[11].XIC[2].icell.PUM VPWR 0.01036f
C2153 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PUM 0.00131f
C2154 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PUM 0.00131f
C2155 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04522f
C2156 XThR.XTB7.B a_n1319_5317# 0.00108f
C2157 XThC.XTB1.Y a_3299_10575# 0.0097f
C2158 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C2159 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C2160 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00529f
C2161 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.01406f
C2162 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06536f
C2163 XA.XIR[8].XIC[7].icell.SM Iout 0.00388f
C2164 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[10].icell.Ien 0.00212f
C2165 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.SM 0.00188f
C2166 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.15089f
C2167 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.03424f
C2168 XThR.Tn[11] XA.XIR[12].XIC[1].icell.SM 0.00121f
C2169 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00212f
C2170 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.SM 0.00188f
C2171 XThC.XTB6.A XThC.Tn[2] 0.00108f
C2172 XThC.Tn[6] XThR.Tn[13] 0.28062f
C2173 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.03424f
C2174 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38979f
C2175 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04522f
C2176 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.SM 0.00383f
C2177 XA.XIR[15].XIC[2].icell.SM Vbias 0.00701f
C2178 XA.XIR[10].XIC[0].icell.Ien Iout 0.06474f
C2179 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.15089f
C2180 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.SM 0.00383f
C2181 a_5155_9615# XThC.Tn[4] 0.26653f
C2182 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C2183 XThR.Tn[1] XA.XIR[2].XIC_15.icell.Ien 0.00116f
C2184 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.SM 0.00188f
C2185 XA.XIR[9].XIC[14].icell.SM VPWR 0.00208f
C2186 XA.XIR[6].XIC[14].icell.SM Vbias 0.00701f
C2187 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PUM 0.00131f
C2188 XA.XIR[7].XIC[9].icell.SM Vbias 0.00701f
C2189 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04522f
C2190 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C2191 XThR.Tn[7] XA.XIR[8].XIC[12].icell.Ien 0.00321f
C2192 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.15089f
C2193 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.PUM 0.00137f
C2194 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PUM 0.00529f
C2195 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04522f
C2196 XA.XIR[1].XIC[10].icell.SM Vbias 0.00701f
C2197 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.15089f
C2198 XThC.XTBN.A XThC.Tn[8] 0.1369f
C2199 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C2200 XA.XIR[8].XIC[0].icell.Ien VPWR 0.19066f
C2201 XThR.Tn[14] XA.XIR[14].XIC[8].icell.PDM 0.0033f
C2202 XA.XIR[15].XIC[8].icell.PUM VPWR 0.01036f
C2203 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06536f
C2204 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.03424f
C2205 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.0352f
C2206 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00529f
C2207 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.03424f
C2208 XA.XIR[2].XIC[0].icell.SM VPWR 0.00158f
C2209 XThR.Tn[13] XA.XIR[14].XIC[7].icell.SM 0.00121f
C2210 XA.XIR[0].XIC[13].icell.PDM Vbias 0.04065f
C2211 XA.XIR[7].XIC[0].icell.PUM VPWR 0.01036f
C2212 XA.XIR[14].XIC[1].icell.SM VPWR 0.00158f
C2213 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.SM 0.00383f
C2214 XA.XIR[12].XIC[10].icell.SM Iout 0.00388f
C2215 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C2216 XThC.Tn[8] XThR.Tn[4] 0.28062f
C2217 XThR.Tn[6] XThR.XTBN.A 0.00131f
C2218 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04522f
C2219 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04f
C2220 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C2221 XThR.Tn[4] XA.XIR[4].XIC[0].icell.PDM 0.00335f
C2222 XA.XIR[13].XIC[5].icell.PDM VPWR 0.00863f
C2223 XThR.Tn[0] XA.XIR[1].XIC[7].icell.SM 0.00121f
C2224 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.03976f
C2225 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.SM 0.00383f
C2226 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02698f
C2227 XThR.XTB7.B XThR.Tn[9] 0.0565f
C2228 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02736f
C2229 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PUM 0.00529f
C2230 XA.XIR[10].XIC[4].icell.PDM Vbias 0.04058f
C2231 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.03424f
C2232 XA.XIR[6].XIC[0].icell.Ien Vbias 0.21102f
C2233 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PUM 0.00534f
C2234 a_n1049_5317# XThR.Tn[6] 0.26047f
C2235 XThC.Tn[6] Vbias 2.24855f
C2236 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PUM 0.00131f
C2237 XA.XIR[12].XIC[6].icell.PDM VPWR 0.00863f
C2238 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.01406f
C2239 XA.XIR[7].XIC[14].icell.PUM Vbias 0.00347f
C2240 XThR.Tn[0] XA.XIR[0].XIC[10].icell.PDM 0.0033f
C2241 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.SM 0.00188f
C2242 XA.XIR[5].XIC[1].icell.SM Vbias 0.00701f
C2243 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02698f
C2244 XA.XIR[11].XIC[6].icell.PUM VPWR 0.01036f
C2245 XA.XIR[15].XIC[14].icell.PDM Iout 0.00112f
C2246 XThR.XTB5.A a_n1335_4229# 0.01243f
C2247 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.03552f
C2248 XA.XIR[0].XIC[13].icell.Ien Iout 0.06455f
C2249 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04522f
C2250 XThR.Tn[2] XA.XIR[3].XIC[0].icell.SM 0.00121f
C2251 XA.XIR[4].XIC[4].icell.PUM Vbias 0.00347f
C2252 XThC.XTB6.Y XThC.Tn[4] 0.00264f
C2253 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02698f
C2254 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PUM 0.00131f
C2255 XThC.XTB7.A a_5949_9615# 0.01824f
C2256 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PUM 0.00529f
C2257 XA.XIR[10].XIC[7].icell.Ien VPWR 0.19065f
C2258 XThR.Tn[13] XA.XIR[14].XIC[12].icell.SM 0.00121f
C2259 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00212f
C2260 XA.XIR[6].XIC[4].icell.SM VPWR 0.00158f
C2261 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.SM 0.00188f
C2262 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PUM 0.00529f
C2263 XA.XIR[0].XIC_dummy_right.icell.PUM Vbias 0.00248f
C2264 XThR.Tn[2] XA.XIR[2].XIC[4].icell.PDM 0.0033f
C2265 XA.XIR[3].XIC[7].icell.PDM Vbias 0.04058f
C2266 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00212f
C2267 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.SM 0.00188f
C2268 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02761f
C2269 XA.XIR[10].XIC[4].icell.Ien Iout 0.06483f
C2270 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PUM 0.00131f
C2271 XA.XIR[6].XIC[1].icell.SM Iout 0.00388f
C2272 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11] 0.0033f
C2273 XA.XIR[5].XIC[7].icell.PUM VPWR 0.01036f
C2274 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.SM 0.00383f
C2275 XA.XIR[7].XIC_15.icell.SM VPWR 0.00276f
C2276 XA.XIR[2].XIC[6].icell.SM Vbias 0.00701f
C2277 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PUM 0.00131f
C2278 XThC.XTB2.Y a_7875_9569# 0.06476f
C2279 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06536f
C2280 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.SM 0.00188f
C2281 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00212f
C2282 XA.XIR[14].XIC[7].icell.SM Vbias 0.00701f
C2283 XA.XIR[4].XIC[10].icell.PDM VPWR 0.00863f
C2284 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PUM 0.00131f
C2285 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.01406f
C2286 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00529f
C2287 XThC.XTB5.A XThC.XTB7.A 0.07824f
C2288 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C2289 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.03976f
C2290 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.01406f
C2291 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02698f
C2292 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.03424f
C2293 XA.XIR[4].XIC[7].icell.PDM Iout 0.00112f
C2294 XThR.Tn[6] XA.XIR[7].XIC[9].icell.SM 0.00121f
C2295 XA.XIR[3].XIC[10].icell.Ien VPWR 0.19065f
C2296 XA.XIR[9].XIC[6].icell.Ien Vbias 0.21238f
C2297 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PUM 0.00529f
C2298 XA.XIR[8].XIC[3].icell.SM VPWR 0.00158f
C2299 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12] 0.0033f
C2300 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.SM 0.00188f
C2301 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PUM 0.00131f
C2302 XA.XIR[6].XIC[0].icell.PDM Iout 0.00112f
C2303 XA.XIR[3].XIC[7].icell.Ien Iout 0.06483f
C2304 XA.XIR[7].XIC_dummy_left.icell.Ien Vbias 0.00342f
C2305 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11595f
C2306 XThC.XTBN.Y XThC.Tn[0] 0.53577f
C2307 data[1] data[2] 0.01393f
C2308 XA.XIR[8].XIC[0].icell.SM Iout 0.00388f
C2309 XA.XIR[11].XIC[13].icell.PUM Vbias 0.00347f
C2310 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.03548f
C2311 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PUM 0.00131f
C2312 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PUM 0.00529f
C2313 XThR.Tn[5] a_n1049_5611# 0.27042f
C2314 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.SM 0.00383f
C2315 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01799f
C2316 XThR.Tn[1] XA.XIR[2].XIC[11].icell.Ien 0.00321f
C2317 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PUM 0.00529f
C2318 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00212f
C2319 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02698f
C2320 XA.XIR[9].XIC[10].icell.SM VPWR 0.00158f
C2321 XA.XIR[6].XIC[10].icell.SM Vbias 0.00701f
C2322 XThC.XTB4.Y XThC.Tn[4] 0.00758f
C2323 XA.XIR[14].XIC[12].icell.SM Vbias 0.00701f
C2324 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04522f
C2325 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.SM 0.00188f
C2326 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00529f
C2327 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.02698f
C2328 XA.XIR[4].XIC[12].icell.Ien VPWR 0.19065f
C2329 XThR.Tn[3] XA.XIR[4].XIC[8].icell.SM 0.00121f
C2330 XThC.XTB3.Y XThC.Tn[8] 0.00178f
C2331 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.SM 0.00188f
C2332 XA.XIR[12].XIC_15.icell.PDM VPWR 0.06959f
C2333 XA.XIR[9].XIC[7].icell.SM Iout 0.00388f
C2334 XA.XIR[7].XIC[2].icell.SM Vbias 0.00701f
C2335 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.SM 0.00188f
C2336 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04522f
C2337 XThR.Tn[14] XA.XIR[15].XIC[5].icell.Ien 0.00321f
C2338 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02698f
C2339 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.15089f
C2340 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04522f
C2341 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.03424f
C2342 XThR.Tn[10] XA.XIR[11].XIC[14].icell.SM 0.00121f
C2343 XThC.Tn[6] XThR.Tn[6] 0.28062f
C2344 XA.XIR[3].XIC[13].icell.SM VPWR 0.00158f
C2345 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PUM 0.00131f
C2346 XA.XIR[1].XIC[3].icell.SM Vbias 0.00701f
C2347 XThR.XTBN.Y a_n1049_7787# 0.08456f
C2348 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PUM 0.00529f
C2349 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00529f
C2350 XA.XIR[15].XIC[1].icell.PUM VPWR 0.01036f
C2351 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PUM 0.00529f
C2352 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.15089f
C2353 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.SM 0.00383f
C2354 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PUM 0.00529f
C2355 XA.XIR[0].XIC[6].icell.PDM Vbias 0.04065f
C2356 XA.XIR[8].XIC[9].icell.SM Vbias 0.00701f
C2357 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01799f
C2358 XA.XIR[14].XIC[2].icell.PUM VPWR 0.01036f
C2359 XThR.Tn[4] XA.XIR[5].XIC[8].icell.SM 0.00121f
C2360 XA.XIR[7].XIC[8].icell.PUM VPWR 0.01036f
C2361 XA.XIR[2].XIC[14].icell.PDM Iout 0.00112f
C2362 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02698f
C2363 XA.XIR[15].XIC[14].icell.SM Iout 0.00388f
C2364 XThR.Tn[8] XA.XIR[8].XIC[13].icell.PDM 0.0033f
C2365 XA.XIR[11].XIC[13].icell.SM Vbias 0.00701f
C2366 XThR.Tn[13] XA.XIR[13].XIC[4].icell.PDM 0.0033f
C2367 XA.XIR[1].XIC[9].icell.PUM VPWR 0.01036f
C2368 XThR.Tn[0] XA.XIR[1].XIC[0].icell.SM 0.00121f
C2369 XThR.XTB6.A XThR.XTB7.A 0.44014f
C2370 XThC.Tn[0] XThR.Tn[5] 0.28067f
C2371 XA.XIR[2].XIC_15.icell.PUM Vbias 0.00347f
C2372 XThC.XTB5.Y VPWR 1.0121f
C2373 XA.XIR[13].XIC[0].icell.Ien Iout 0.06474f
C2374 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.SM 0.00383f
C2375 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PUM 0.00131f
C2376 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.03976f
C2377 XThR.Tn[14] XA.XIR[15].XIC[9].icell.Ien 0.00321f
C2378 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PUM 0.00529f
C2379 XThR.XTBN.A a_n997_2667# 0.01679f
C2380 XA.XIR[0].XIC[9].icell.Ien VPWR 0.19155f
C2381 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.01406f
C2382 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.15089f
C2383 XThR.Tn[0] XA.XIR[0].XIC[3].icell.PDM 0.0033f
C2384 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.03424f
C2385 XA.XIR[12].XIC[1].icell.Ien Iout 0.06483f
C2386 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PUM 0.00529f
C2387 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PUM 0.00131f
C2388 XA.XIR[8].XIC_dummy_left.icell.SM VPWR 0.00269f
C2389 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01776f
C2390 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04522f
C2391 XThR.Tn[12] XA.XIR[12].XIC[6].icell.PDM 0.0033f
C2392 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C2393 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.01406f
C2394 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06536f
C2395 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C2396 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00529f
C2397 XA.XIR[0].XIC[6].icell.Ien Iout 0.06455f
C2398 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04522f
C2399 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[11].icell.SM 0.00383f
C2400 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02698f
C2401 XA.XIR[3].XIC[14].icell.SM Iout 0.00388f
C2402 XThR.Tn[5] XA.XIR[5].XIC[13].icell.PDM 0.0033f
C2403 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PUM 0.00131f
C2404 XThR.XTB7.B XThR.Tn[10] 0.06102f
C2405 XThC.Tn[7] XThR.Tn[1] 0.28093f
C2406 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.SM 0.00188f
C2407 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Ien 0.00217f
C2408 XThR.Tn[9] XA.XIR[10].XIC[2].icell.SM 0.00121f
C2409 XA.XIR[8].XIC[14].icell.PUM Vbias 0.00347f
C2410 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PUM 0.00131f
C2411 XA.XIR[15].XIC[7].icell.PUM Vbias 0.00347f
C2412 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C2413 XThR.Tn[10] XA.XIR[11].XIC[12].icell.Ien 0.00321f
C2414 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04522f
C2415 XThR.XTBN.Y XThR.Tn[9] 0.48051f
C2416 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PUM 0.00529f
C2417 XA.XIR[5].XIC[0].icell.Ien VPWR 0.19066f
C2418 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00529f
C2419 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02698f
C2420 XA.XIR[1].XIC[14].icell.PDM VPWR 0.00873f
C2421 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PUM 0.00529f
C2422 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.03976f
C2423 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PUM 0.00529f
C2424 XA.XIR[4].XIC[3].icell.PDM VPWR 0.00863f
C2425 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.SM 0.00188f
C2426 XThC.XTBN.Y VPWR 4.08965f
C2427 XThC.XTB6.Y a_6243_9615# 0.01199f
C2428 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00212f
C2429 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PUM 0.00529f
C2430 XA.XIR[15].XIC[12].icell.Ien Iout 0.06816f
C2431 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.SM 0.00188f
C2432 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00529f
C2433 XA.XIR[13].XIC[4].icell.PDM Vbias 0.04058f
C2434 XA.XIR[3].XIC[3].icell.Ien VPWR 0.19065f
C2435 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PDM 0.00182f
C2436 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.SM 0.00383f
C2437 XThR.Tn[6] XA.XIR[7].XIC[2].icell.SM 0.00121f
C2438 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.03976f
C2439 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PUM 0.00529f
C2440 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00212f
C2441 XA.XIR[8].XIC_15.icell.SM VPWR 0.00276f
C2442 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PUM 0.00131f
C2443 XA.XIR[3].XIC[0].icell.Ien Iout 0.06474f
C2444 XA.XIR[2].XIC[5].icell.PUM VPWR 0.01036f
C2445 XA.XIR[15].XIC[10].icell.PDM Iout 0.00112f
C2446 XA.XIR[12].XIC[5].icell.PDM Vbias 0.04058f
C2447 XA.XIR[12].XIC_15.icell.SM Iout 0.0047f
C2448 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00529f
C2449 XA.XIR[14].XIC[6].icell.PUM VPWR 0.01036f
C2450 XA.XIR[11].XIC[5].icell.PUM Vbias 0.00347f
C2451 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[3].icell.Ien 0.00212f
C2452 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01402f
C2453 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.SM 0.00188f
C2454 XThC.XTB1.Y XThC.Tn[8] 0.29191f
C2455 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.SM 0.00383f
C2456 XA.XIR[12].XIC[11].icell.SM VPWR 0.00158f
C2457 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01897f
C2458 XA.XIR[13].XIC[7].icell.Ien VPWR 0.19065f
C2459 XThR.Tn[1] XA.XIR[2].XIC[4].icell.Ien 0.00321f
C2460 XA.XIR[10].XIC[6].icell.Ien Vbias 0.21238f
C2461 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00212f
C2462 XA.XIR[9].XIC[3].icell.SM VPWR 0.00158f
C2463 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.SM 0.00188f
C2464 XA.XIR[6].XIC[3].icell.SM Vbias 0.00701f
C2465 XThC.Tn[10] VPWR 6.89727f
C2466 XA.XIR[13].XIC[4].icell.Ien Iout 0.06483f
C2467 XA.XIR[12].XIC[8].icell.Ien VPWR 0.19065f
C2468 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PUM 0.00529f
C2469 XThR.Tn[3] XA.XIR[4].XIC[1].icell.SM 0.00121f
C2470 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.15089f
C2471 XA.XIR[5].XIC[6].icell.PUM Vbias 0.00347f
C2472 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00529f
C2473 a_4861_9615# VPWR 0.70525f
C2474 XThC.XTBN.A XThC.Tn[6] 0.00131f
C2475 XA.XIR[12].XIC[5].icell.Ien Iout 0.06483f
C2476 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C2477 XThR.XTB7.Y a_n997_715# 0.06874f
C2478 XThR.Tn[12] XA.XIR[12].XIC_15.icell.PDM 0.0033f
C2479 XA.XIR[10].XIC[0].icell.PDM VPWR 0.00863f
C2480 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PUM 0.00131f
C2481 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00212f
C2482 XA.XIR[4].XIC[9].icell.PDM Vbias 0.04058f
C2483 XA.XIR[1].XIC_15.icell.SM Vbias 0.00701f
C2484 XThC.Tn[9] XThR.Tn[9] 0.28062f
C2485 XA.XIR[11].XIC[8].icell.PDM Iout 0.00112f
C2486 XA.XIR[11].XIC[14].icell.PDM Vbias 0.04058f
C2487 XA.XIR[6].XIC[9].icell.PUM VPWR 0.01036f
C2488 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.SM 0.00383f
C2489 XThC.Tn[6] XThR.Tn[4] 0.28062f
C2490 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.15089f
C2491 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.01406f
C2492 XThR.Tn[13] a_n997_1579# 0.19413f
C2493 XThR.Tn[5] VPWR 6.69157f
C2494 XA.XIR[3].XIC[9].icell.Ien Vbias 0.21238f
C2495 XThC.XTB4.Y a_6243_9615# 0.00463f
C2496 XThR.Tn[13] XA.XIR[14].XIC[13].icell.SM 0.00121f
C2497 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.SM 0.00383f
C2498 XA.XIR[11].XIC[9].icell.PUM Vbias 0.00347f
C2499 XA.XIR[8].XIC[2].icell.SM Vbias 0.00701f
C2500 XA.XIR[10].XIC[7].icell.SM Iout 0.00388f
C2501 XA.XIR[7].XIC[1].icell.PUM VPWR 0.01036f
C2502 XA.XIR[5].XIC[12].icell.PDM VPWR 0.00863f
C2503 XThR.Tn[4] XA.XIR[5].XIC[1].icell.SM 0.00121f
C2504 XThR.Tn[8] XA.XIR[8].XIC[6].icell.PDM 0.0033f
C2505 XA.XIR[14].XIC[13].icell.PUM Vbias 0.00347f
C2506 XA.XIR[2].XIC[11].icell.PUM Vbias 0.00347f
C2507 XThC.XTB5.Y a_9827_9569# 0.06458f
C2508 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.01406f
C2509 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PUM 0.00529f
C2510 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.SM 0.00383f
C2511 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.SM 0.00383f
C2512 XA.XIR[1].XIC[2].icell.PUM VPWR 0.01036f
C2513 XA.XIR[5].XIC[9].icell.PDM Iout 0.00112f
C2514 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.SM 0.00383f
C2515 XA.XIR[12].XIC[13].icell.Ien VPWR 0.19065f
C2516 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00529f
C2517 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.SM 0.00383f
C2518 XThC.XTB7.A a_8739_9569# 0.00342f
C2519 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02698f
C2520 XThR.Tn[7] XA.XIR[8].XIC[5].icell.Ien 0.00321f
C2521 XA.XIR[4].XIC[9].icell.Ien Iout 0.06483f
C2522 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.SM 0.00383f
C2523 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.SM 0.00188f
C2524 XThR.XTBN.Y XA.XIR[0].XIC_dummy_left.icell.Iout 0.00136f
C2525 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00212f
C2526 XA.XIR[0].XIC[2].icell.Ien VPWR 0.19003f
C2527 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.SM 0.00188f
C2528 XA.XIR[9].XIC[9].icell.SM Vbias 0.00701f
C2529 XA.XIR[8].XIC[8].icell.PUM VPWR 0.01036f
C2530 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.15089f
C2531 XA.XIR[12].XIC[9].icell.Ien Iout 0.06483f
C2532 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PUM 0.00131f
C2533 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.03981f
C2534 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.SM 0.00188f
C2535 XA.XIR[3].XIC[10].icell.SM Iout 0.00388f
C2536 XThR.Tn[10] XA.XIR[11].XIC[10].icell.SM 0.00121f
C2537 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.03424f
C2538 XThR.Tn[5] XA.XIR[5].XIC[6].icell.PDM 0.0033f
C2539 XA.XIR[6].XIC[14].icell.PDM VPWR 0.00873f
C2540 XA.XIR[3].XIC[12].icell.SM Vbias 0.00701f
C2541 XA.XIR[11].XIC[14].icell.PUM Vbias 0.00347f
C2542 XA.XIR[10].XIC[12].icell.SM Iout 0.00388f
C2543 XThC.Tn[4] Iout 0.84024f
C2544 a_n1049_6405# XThR.Tn[4] 0.26564f
C2545 XA.XIR[5].XIC[14].icell.Ien VPWR 0.1907f
C2546 a_5155_10571# VPWR 0.00653f
C2547 XA.XIR[9].XIC[0].icell.PUM VPWR 0.01036f
C2548 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.SM 0.00188f
C2549 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.01406f
C2550 XA.XIR[15].XIC[10].icell.SM Iout 0.00388f
C2551 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C2552 XThR.XTB6.Y XThR.Tn[6] 0.00639f
C2553 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04522f
C2554 XThC.XTBN.Y a_9827_9569# 0.22873f
C2555 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02698f
C2556 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C2557 XA.XIR[14].XIC[13].icell.SM Vbias 0.00701f
C2558 XA.XIR[7].XIC[7].icell.PUM Vbias 0.00347f
C2559 a_n1049_6699# VPWR 0.72168f
C2560 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C2561 XA.XIR[4].XIC[12].icell.SM Iout 0.00388f
C2562 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08017f
C2563 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00529f
C2564 XA.XIR[1].XIC[8].icell.PUM Vbias 0.00347f
C2565 XA.XIR[9].XIC[14].icell.PUM Vbias 0.00347f
C2566 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01193f
C2567 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C2568 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.15089f
C2569 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.03976f
C2570 XA.XIR[4].XIC_15.icell.Ien Vbias 0.21343f
C2571 XA.XIR[12].XIC[12].icell.PDM Iout 0.00112f
C2572 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.SM 0.00188f
C2573 XA.XIR[0].XIC[8].icell.Ien Vbias 0.21246f
C2574 XA.XIR[15].XIC[3].icell.PDM Iout 0.00112f
C2575 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.PUM 0.00112f
C2576 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.03424f
C2577 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PUM 0.00131f
C2578 XA.XIR[7].XIC[13].icell.PDM VPWR 0.00863f
C2579 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.SM 0.00188f
C2580 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02698f
C2581 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C2582 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Ien 0.00529f
C2583 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00212f
C2584 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00212f
C2585 XA.XIR[5].XIC_dummy_left.icell.SM VPWR 0.00269f
C2586 XA.XIR[7].XIC[10].icell.PDM Iout 0.00112f
C2587 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.15089f
C2588 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PUM 0.00529f
C2589 XThR.XTB7.B XThR.Tn[13] 0.00276f
C2590 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C2591 XA.XIR[11].XIC[14].icell.SM Vbias 0.00701f
C2592 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PUM 0.00131f
C2593 XThC.XTB3.Y XThC.Tn[6] 0.00301f
C2594 XA.XIR[5].XIC_15.icell.Ien Iout 0.06485f
C2595 XThR.Tn[12] XA.XIR[13].XIC[7].icell.Ien 0.00321f
C2596 XA.XIR[9].XIC_15.icell.SM VPWR 0.00276f
C2597 XA.XIR[6].XIC_15.icell.SM Vbias 0.00701f
C2598 XA.XIR[1].XIC[11].icell.PDM Iout 0.00112f
C2599 XThC.Tn[3] XThC.Tn[5] 0.00492f
C2600 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00212f
C2601 XA.XIR[1].XIC[2].icell.PDM Vbias 0.04058f
C2602 XA.XIR[0].XIC[12].icell.SM VPWR 0.00158f
C2603 XThC.Tn[10] XThR.Tn[12] 0.28062f
C2604 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02698f
C2605 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.15089f
C2606 XThC.Tn[12] XThR.Tn[2] 0.28062f
C2607 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02698f
C2608 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PUM 0.00529f
C2609 XThR.Tn[14] XA.XIR[15].XIC[10].icell.Ien 0.00321f
C2610 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.15089f
C2611 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00529f
C2612 XThC.XTB2.Y a_6243_9615# 0.00844f
C2613 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C2614 XA.XIR[11].XIC[4].icell.PDM VPWR 0.00863f
C2615 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01897f
C2616 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04f
C2617 XA.XIR[0].XIC[9].icell.SM Iout 0.00367f
C2618 XThC.XTB2.Y data[1] 0.017f
C2619 XA.XIR[4].XIC[2].icell.PDM Vbias 0.04058f
C2620 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00529f
C2621 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Iout 0.00347f
C2622 XA.XIR[10].XIC[3].icell.SM VPWR 0.00158f
C2623 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PUM 0.00131f
C2624 XA.XIR[6].XIC[2].icell.PUM VPWR 0.01036f
C2625 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PUM 0.00131f
C2626 XA.XIR[12].XIC[12].icell.PUM VPWR 0.01036f
C2627 XThC.XTB3.Y a_4387_10575# 0.00941f
C2628 XA.XIR[3].XIC[2].icell.Ien Vbias 0.21238f
C2629 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.SM 0.00188f
C2630 XA.XIR[5].XIC[5].icell.PDM VPWR 0.00863f
C2631 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C2632 XA.XIR[7].XIC[12].icell.Ien Iout 0.06483f
C2633 XA.XIR[2].XIC[4].icell.PUM Vbias 0.00347f
C2634 XA.XIR[14].XIC[5].icell.PUM Vbias 0.00347f
C2635 XA.XIR[4].XIC[5].icell.Ien VPWR 0.19065f
C2636 XThC.Tn[9] XThR.Tn[10] 0.28062f
C2637 XA.XIR[1].XIC[13].icell.Ien Iout 0.06483f
C2638 XThC.XTB7.B XThC.Tn[10] 0.14845f
C2639 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.SM 0.00383f
C2640 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04522f
C2641 XA.XIR[13].XIC[6].icell.Ien Vbias 0.21238f
C2642 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.15089f
C2643 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.0353f
C2644 XA.XIR[3].XIC[6].icell.SM VPWR 0.00158f
C2645 XA.XIR[4].XIC[2].icell.Ien Iout 0.06483f
C2646 XThR.Tn[1] XThR.Tn[2] 0.11944f
C2647 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PUM 0.00131f
C2648 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08027f
C2649 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.SM 0.00188f
C2650 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07289f
C2651 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C2652 XA.XIR[9].XIC[2].icell.SM Vbias 0.00701f
C2653 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.01406f
C2654 XA.XIR[11].XIC[12].icell.Ien Vbias 0.21238f
C2655 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.SM 0.00383f
C2656 XA.XIR[1].XIC_dummy_right.icell.PUM Vbias 0.00248f
C2657 XA.XIR[12].XIC[7].icell.Ien Vbias 0.21238f
C2658 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.03976f
C2659 XThC.XTB7.B a_4861_9615# 0.0036f
C2660 XA.XIR[3].XIC[3].icell.SM Iout 0.00388f
C2661 XA.XIR[2].XIC[10].icell.PDM VPWR 0.00863f
C2662 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08027f
C2663 XThC.XTBN.A data[3] 0.07741f
C2664 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.01406f
C2665 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PUM 0.00131f
C2666 XA.XIR[13].XIC[0].icell.PDM VPWR 0.00863f
C2667 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[4].icell.SM 0.00383f
C2668 XA.XIR[11].XIC[10].icell.PDM Vbias 0.04058f
C2669 XA.XIR[2].XIC[7].icell.PDM Iout 0.00112f
C2670 XThC.XTB7.A data[0] 0.86893f
C2671 XThC.XTB6.Y a_8963_9569# 0.00468f
C2672 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PUM 0.00529f
C2673 XA.XIR[14].XIC[14].icell.PDM Vbias 0.04058f
C2674 XA.XIR[14].XIC[8].icell.PDM Iout 0.00112f
C2675 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.15089f
C2676 XThR.Tn[1] XA.XIR[2].XIC[7].icell.SM 0.00121f
C2677 XA.XIR[6].XIC[8].icell.PUM Vbias 0.00347f
C2678 XA.XIR[9].XIC[8].icell.PUM VPWR 0.01036f
C2679 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C2680 XThR.Tn[9] XA.XIR[9].XIC[12].icell.PDM 0.0033f
C2681 XA.XIR[13].XIC[7].icell.SM Iout 0.00388f
C2682 XThR.Tn[10] XA.XIR[11].XIC[1].icell.Ien 0.00321f
C2683 XA.XIR[14].XIC[9].icell.PUM Vbias 0.00347f
C2684 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PUM 0.00131f
C2685 a_3773_9615# XThC.Tn[1] 0.27139f
C2686 XThR.Tn[14] XA.XIR[15].XIC[1].icell.SM 0.00121f
C2687 XA.XIR[5].XIC[11].icell.PDM Vbias 0.04058f
C2688 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.SM 0.00188f
C2689 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00212f
C2690 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.01406f
C2691 XThR.Tn[4] XThR.XTB6.Y 0.00264f
C2692 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.03976f
C2693 XThR.Tn[3] XA.XIR[3].XIC[9].icell.PDM 0.0033f
C2694 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.03428f
C2695 XThR.XTB7.A a_n1319_5317# 0.0017f
C2696 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PUM 0.00131f
C2697 XA.XIR[4].XIC[11].icell.Ien Vbias 0.21238f
C2698 XThR.XTB6.Y a_n997_2667# 0.00468f
C2699 XA.XIR[2].XIC[12].icell.Ien VPWR 0.19065f
C2700 XA.XIR[10].XIC[0].icell.PUM VPWR 0.01036f
C2701 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01776f
C2702 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.01406f
C2703 XA.XIR[0].XIC[1].icell.Ien Vbias 0.21246f
C2704 XA.XIR[6].XIC[11].icell.PDM Iout 0.00112f
C2705 XA.XIR[8].XIC[7].icell.PUM Vbias 0.00347f
C2706 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PUM 0.00131f
C2707 XThR.XTB3.Y a_n997_3979# 0.00604f
C2708 XA.XIR[15].XIC[1].icell.PDM Vbias 0.04058f
C2709 XA.XIR[7].XIC[6].icell.PDM VPWR 0.00863f
C2710 XThR.Tn[8] data[4] 0.01643f
C2711 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.15089f
C2712 a_7651_9569# VPWR 0.00385f
C2713 XThR.Tn[13] XA.XIR[14].XIC[14].icell.SM 0.00121f
C2714 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.03424f
C2715 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00529f
C2716 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04522f
C2717 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PUM 0.00131f
C2718 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.SM 0.00188f
C2719 XThR.Tn[4] XA.XIR[4].XIC[9].icell.PDM 0.0033f
C2720 XA.XIR[1].XIC[7].icell.PDM VPWR 0.00863f
C2721 XA.XIR[5].XIC[11].icell.Ien Iout 0.06483f
C2722 XA.XIR[7].XIC[3].icell.PDM Iout 0.00112f
C2723 XA.XIR[13].XIC[12].icell.SM Iout 0.00388f
C2724 XA.XIR[14].XIC[14].icell.PUM Vbias 0.00347f
C2725 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.15089f
C2726 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00212f
C2727 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01799f
C2728 XA.XIR[12].XIC[0].icell.SM VPWR 0.00158f
C2729 XThR.Tn[7] XA.XIR[8].XIC[8].icell.SM 0.00121f
C2730 XA.XIR[1].XIC[4].icell.PDM Iout 0.00112f
C2731 XA.XIR[12].XIC[14].icell.Ien VPWR 0.1907f
C2732 XThC.Tn[14] XThR.Tn[0] 0.281f
C2733 XA.XIR[5].XIC[13].icell.Ien Vbias 0.21238f
C2734 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.SM 0.00383f
C2735 XA.XIR[0].XIC[5].icell.SM VPWR 0.00158f
C2736 XThC.XTB4.Y a_8963_9569# 0.07199f
C2737 XA.XIR[8].XIC[13].icell.PDM VPWR 0.00863f
C2738 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01776f
C2739 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.03976f
C2740 XThC.Tn[7] XThR.Tn[9] 0.28062f
C2741 XThR.Tn[2] XA.XIR[3].XIC[12].icell.Ien 0.00321f
C2742 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.SM 0.00383f
C2743 XA.XIR[0].XIC[2].icell.SM Iout 0.00367f
C2744 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00212f
C2745 XThR.XTB7.B XThR.Tn[6] 0.04822f
C2746 XA.XIR[12].XIC[10].icell.Ien Iout 0.06483f
C2747 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.SM 0.00383f
C2748 XA.XIR[8].XIC[10].icell.PDM Iout 0.00112f
C2749 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C2750 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.15089f
C2751 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PUM 0.00529f
C2752 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.03976f
C2753 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C2754 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04522f
C2755 XA.XIR[6].XIC[13].icell.Ien Iout 0.06483f
C2756 XA.XIR[10].XIC[13].icell.SM Iout 0.00388f
C2757 XA.XIR[15].XIC[5].icell.PDM Vbias 0.04058f
C2758 XA.XIR[15].XIC_15.icell.SM Iout 0.0047f
C2759 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00529f
C2760 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04522f
C2761 XA.XIR[6].XIC_dummy_right.icell.PUM Vbias 0.00248f
C2762 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01897f
C2763 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.SM 0.00188f
C2764 XThR.Tn[10] XA.XIR[11].XIC[5].icell.Ien 0.00321f
C2765 XA.XIR[7].XIC[12].icell.PDM Vbias 0.04058f
C2766 XA.XIR[15].XIC[11].icell.SM VPWR 0.00158f
C2767 XA.XIR[11].XIC[10].icell.SM Vbias 0.00701f
C2768 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PUM 0.00529f
C2769 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.03424f
C2770 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PUM 0.00131f
C2771 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.03424f
C2772 XThC.XTB7.Y a_6243_10571# 0.01283f
C2773 XA.XIR[14].XIC[14].icell.SM Vbias 0.00701f
C2774 XA.XIR[1].XIC[13].icell.PDM Vbias 0.04058f
C2775 XThR.XTB1.Y XThR.Tn[7] 0.00426f
C2776 XA.XIR[15].XIC[8].icell.Ien VPWR 0.32782f
C2777 XThR.Tn[13] XA.XIR[14].XIC[12].icell.Ien 0.00321f
C2778 XA.XIR[8].XIC[1].icell.PUM VPWR 0.01036f
C2779 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13469f
C2780 XThC.XTB5.A data[0] 0.14415f
C2781 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Iout 0.00347f
C2782 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PUM 0.00529f
C2783 XA.XIR[8].XIC[12].icell.Ien Iout 0.06483f
C2784 XThC.Tn[5] XThR.Tn[11] 0.28062f
C2785 XA.XIR[0].XIC[11].icell.SM Vbias 0.00701f
C2786 XA.XIR[2].XIC[3].icell.PDM VPWR 0.00863f
C2787 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00212f
C2788 XA.XIR[15].XIC[5].icell.Ien Iout 0.06816f
C2789 XA.XIR[3].XIC_15.icell.SM Iout 0.0047f
C2790 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.03976f
C2791 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.SM 0.00188f
C2792 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02698f
C2793 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11595f
C2794 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04522f
C2795 XA.XIR[14].XIC[4].icell.PDM VPWR 0.00863f
C2796 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.SM 0.00188f
C2797 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02698f
C2798 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.SM 0.00383f
C2799 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00212f
C2800 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.03976f
C2801 XA.XIR[13].XIC[3].icell.SM VPWR 0.00158f
C2802 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PUM 0.00529f
C2803 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.SM 0.00383f
C2804 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.03982f
C2805 XThR.Tn[1] XA.XIR[2].XIC[0].icell.SM 0.00121f
C2806 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.SM 0.00383f
C2807 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.03424f
C2808 XA.XIR[10].XIC[2].icell.SM Vbias 0.00701f
C2809 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.03424f
C2810 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13469f
C2811 XA.XIR[6].XIC[1].icell.PUM Vbias 0.00347f
C2812 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.SM 0.00188f
C2813 XThR.XTBN.Y Vbias 0.00722f
C2814 XThR.Tn[9] XA.XIR[9].XIC[5].icell.PDM 0.0033f
C2815 XThR.Tn[10] XA.XIR[11].XIC[9].icell.Ien 0.00321f
C2816 XA.XIR[7].XIC[14].icell.Ien Vbias 0.21238f
C2817 XA.XIR[12].XIC[4].icell.SM VPWR 0.00158f
C2818 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C2819 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00212f
C2820 XA.XIR[5].XIC[4].icell.PDM Vbias 0.04058f
C2821 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04522f
C2822 XA.XIR[15].XIC[13].icell.Ien VPWR 0.32782f
C2823 XA.XIR[11].XIC[6].icell.Ien VPWR 0.19065f
C2824 XA.XIR[12].XIC[1].icell.SM Iout 0.00388f
C2825 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.SM 0.00383f
C2826 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.SM 0.00383f
C2827 XThR.Tn[3] XA.XIR[3].XIC[2].icell.PDM 0.0033f
C2828 XThC.Tn[9] XThR.Tn[13] 0.28062f
C2829 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.03976f
C2830 XA.XIR[4].XIC[4].icell.Ien Vbias 0.21238f
C2831 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02709f
C2832 XA.XIR[11].XIC[3].icell.Ien Iout 0.06483f
C2833 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.03424f
C2834 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00529f
C2835 XA.XIR[10].XIC[8].icell.PUM VPWR 0.01036f
C2836 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08027f
C2837 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00529f
C2838 XA.XIR[15].XIC[9].icell.Ien Iout 0.06816f
C2839 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PUM 0.00529f
C2840 XA.XIR[6].XIC[7].icell.PDM VPWR 0.00863f
C2841 XThC.Tn[11] XThR.Tn[3] 0.28062f
C2842 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.03424f
C2843 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.04495f
C2844 XA.XIR[3].XIC[5].icell.SM Vbias 0.00701f
C2845 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C2846 XA.XIR[14].XIC[12].icell.Ien Vbias 0.21238f
C2847 XA.XIR[5].XIC[7].icell.Ien VPWR 0.19065f
C2848 XA.XIR[6].XIC[4].icell.PDM Iout 0.00112f
C2849 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04522f
C2850 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04522f
C2851 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.15089f
C2852 XThC.Tn[1] XThR.Tn[2] 0.28062f
C2853 XA.XIR[2].XIC[9].icell.PDM Vbias 0.04058f
C2854 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04522f
C2855 XThC.Tn[5] XThR.Tn[7] 0.28062f
C2856 XThR.Tn[0] XA.XIR[1].XIC[12].icell.Ien 0.00321f
C2857 XA.XIR[14].XIC[10].icell.PDM Vbias 0.04058f
C2858 XA.XIR[4].XIC[8].icell.SM VPWR 0.00158f
C2859 XA.XIR[5].XIC[4].icell.Ien Iout 0.06483f
C2860 XThR.Tn[4] XA.XIR[4].XIC[2].icell.PDM 0.0033f
C2861 XA.XIR[12].XIC[8].icell.SM VPWR 0.00158f
C2862 XThR.Tn[7] XA.XIR[8].XIC[1].icell.SM 0.00121f
C2863 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00529f
C2864 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.04559f
C2865 XA.XIR[3].XIC[11].icell.PUM VPWR 0.01036f
C2866 XA.XIR[4].XIC[5].icell.SM Iout 0.00388f
C2867 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00212f
C2868 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04522f
C2869 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.03976f
C2870 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.03976f
C2871 XA.XIR[12].XIC[0].icell.PDM Vbias 0.04002f
C2872 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PUM 0.00529f
C2873 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.03424f
C2874 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00529f
C2875 XA.XIR[9].XIC[7].icell.PUM Vbias 0.00347f
C2876 XA.XIR[8].XIC[6].icell.PDM VPWR 0.00863f
C2877 XThR.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.00321f
C2878 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.15089f
C2879 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.01406f
C2880 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.08055f
C2881 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00529f
C2882 XA.XIR[10].XIC[14].icell.PDM Iout 0.00112f
C2883 XA.XIR[8].XIC[3].icell.PDM Iout 0.00112f
C2884 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00529f
C2885 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.15089f
C2886 XA.XIR[15].XIC_dummy_left.icell.Ien Vbias 0.00342f
C2887 XA.XIR[2].XIC[9].icell.Ien Iout 0.06483f
C2888 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02698f
C2889 XThR.XTB7.B XThR.Tn[4] 0.00356f
C2890 XThC.Tn[9] Vbias 2.30815f
C2891 XA.XIR[13].XIC[0].icell.PUM VPWR 0.01036f
C2892 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.03424f
C2893 XA.XIR[15].XIC[12].icell.PDM Iout 0.00112f
C2894 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04522f
C2895 XThC.Tn[0] XA.XIR[12].XIC_dummy_left.icell.Iout 0.00111f
C2896 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04522f
C2897 XA.XIR[6].XIC[13].icell.PDM Vbias 0.04058f
C2898 XA.XIR[9].XIC[13].icell.PDM VPWR 0.00863f
C2899 XThR.XTB7.B a_n997_2667# 0.02071f
C2900 XThC.Tn[7] XThR.Tn[10] 0.28062f
C2901 XThR.Tn[13] XA.XIR[14].XIC[10].icell.SM 0.00121f
C2902 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00212f
C2903 XA.XIR[4].XIC[13].icell.PUM VPWR 0.01036f
C2904 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.SM 0.00188f
C2905 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.SM 0.00188f
C2906 XA.XIR[9].XIC[10].icell.PDM Iout 0.00112f
C2907 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.03976f
C2908 XThC.XTB7.B a_7651_9569# 0.01152f
C2909 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.SM 0.00383f
C2910 XA.XIR[7].XIC[5].icell.PDM Vbias 0.04058f
C2911 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PUM 0.00131f
C2912 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.SM 0.00383f
C2913 XThC.XTB5.Y XThC.Tn[12] 0.32495f
C2914 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02698f
C2915 XThR.XTBN.Y XThR.Tn[6] 0.59885f
C2916 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08017f
C2917 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04522f
C2918 XThR.Tn[6] XA.XIR[7].XIC[14].icell.Ien 0.00321f
C2919 XThR.XTB7.A a_n1331_2891# 0.00995f
C2920 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.15089f
C2921 XA.XIR[1].XIC[6].icell.PDM Vbias 0.04058f
C2922 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.SM 0.00188f
C2923 XA.XIR[15].XIC[1].icell.Ien VPWR 0.32782f
C2924 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.SM 0.00383f
C2925 XThR.Tn[8] XA.XIR[9].XIC[11].icell.SM 0.00121f
C2926 XA.XIR[11].XIC[1].icell.PDM Iout 0.00112f
C2927 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04522f
C2928 XThR.XTB7.A XThR.Tn[10] 0.00404f
C2929 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.03424f
C2930 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00529f
C2931 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C2932 XA.XIR[0].XIC[4].icell.SM Vbias 0.00701f
C2933 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.03424f
C2934 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04522f
C2935 a_n1049_7787# XThR.Tn[2] 0.00158f
C2936 XA.XIR[8].XIC[12].icell.PDM Vbias 0.04058f
C2937 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.03976f
C2938 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Iout 0.00347f
C2939 XA.XIR[11].XIC[1].icell.Ien Vbias 0.21238f
C2940 XA.XIR[2].XIC[12].icell.SM Iout 0.00388f
C2941 XA.XIR[7].XIC[8].icell.Ien VPWR 0.19065f
C2942 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PUM 0.00529f
C2943 XA.XIR[5].XIC[14].icell.SM VPWR 0.00208f
C2944 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.15089f
C2945 XA.XIR[1].XIC[9].icell.Ien VPWR 0.19065f
C2946 XA.XIR[7].XIC[5].icell.Ien Iout 0.06483f
C2947 XA.XIR[2].XIC_15.icell.Ien Vbias 0.21343f
C2948 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.03976f
C2949 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02698f
C2950 XA.XIR[15].XIC[12].icell.PUM VPWR 0.01036f
C2951 XA.XIR[9].XIC[2].icell.PDM VPWR 0.00863f
C2952 XA.XIR[11].XIC[11].icell.PUM Vbias 0.00347f
C2953 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02698f
C2954 XA.XIR[1].XIC[6].icell.Ien Iout 0.06483f
C2955 XThR.Tn[3] XA.XIR[4].XIC[13].icell.Ien 0.00321f
C2956 XA.XIR[9].XIC[12].icell.Ien Iout 0.06483f
C2957 XThR.Tn[12] XA.XIR[13].XIC[3].icell.SM 0.00121f
C2958 XA.XIR[13].XIC[13].icell.SM Iout 0.00388f
C2959 XThC.XTB7.A VPWR 0.87306f
C2960 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.03424f
C2961 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00529f
C2962 XA.XIR[0].XIC[10].icell.PUM VPWR 0.00971f
C2963 XA.XIR[3].XIC[0].icell.PUM VPWR 0.01036f
C2964 XThR.Tn[5] XA.XIR[6].XIC[10].icell.Ien 0.00321f
C2965 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02723f
C2966 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.03424f
C2967 XThR.XTB2.Y a_n1335_8107# 0.01006f
C2968 XA.XIR[12].XIC_15.icell.Ien VPWR 0.25675f
C2969 XThC.XTBN.Y XThC.Tn[12] 0.56523f
C2970 XThC.XTB6.A a_6243_10571# 0.00295f
C2971 XA.XIR[14].XIC[10].icell.SM Vbias 0.00701f
C2972 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.01406f
C2973 XA.XIR[4].XIC_dummy_right.icell.Ien Vbias 0.00287f
C2974 XA.XIR[12].XIC[13].icell.PDM VPWR 0.00863f
C2975 XThR.Tn[11] XA.XIR[12].XIC[6].icell.Ien 0.00321f
C2976 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02698f
C2977 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.03976f
C2978 XA.XIR[8].XIC[14].icell.Ien Vbias 0.21238f
C2979 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.01406f
C2980 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.002f
C2981 XThR.Tn[4] XA.XIR[5].XIC[13].icell.Ien 0.00321f
C2982 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02698f
C2983 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02698f
C2984 XA.XIR[15].XIC[7].icell.Ien Vbias 0.17911f
C2985 XA.XIR[7].XIC[11].icell.SM VPWR 0.00158f
C2986 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.03424f
C2987 XThR.Tn[11] XA.XIR[11].XIC[9].icell.PDM 0.0033f
C2988 XA.XIR[5].XIC[1].icell.PUM VPWR 0.01036f
C2989 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PDM 0.00591f
C2990 XThC.Tn[5] XThR.Tn[14] 0.28062f
C2991 XThC.Tn[3] XThR.Tn[0] 0.28066f
C2992 a_n997_715# VPWR 0.02818f
C2993 XA.XIR[1].XIC[12].icell.SM VPWR 0.00158f
C2994 XA.XIR[2].XIC[2].icell.PDM Vbias 0.04058f
C2995 XA.XIR[10].XIC[14].icell.SM Iout 0.00388f
C2996 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.03424f
C2997 XThC.Tn[9] XThR.Tn[6] 0.28062f
C2998 XA.XIR[11].XIC_15.icell.SM Vbias 0.00701f
C2999 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00529f
C3000 XThC.Tn[11] XThR.Tn[8] 0.28062f
C3001 XA.XIR[4].XIC[1].icell.SM VPWR 0.00158f
C3002 XThR.Tn[6] XA.XIR[6].XIC[13].icell.PDM 0.0033f
C3003 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.SM 0.00188f
C3004 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02698f
C3005 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C3006 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14] 0.0033f
C3007 XThR.Tn[13] XA.XIR[15].XIC_dummy_left.icell.PUM 0.0012f
C3008 XThC.Tn[10] XThC.Tn[12] 0.00453f
C3009 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04522f
C3010 XA.XIR[13].XIC[2].icell.SM Vbias 0.00701f
C3011 XThR.Tn[5] XA.XIR[6].XIC[13].icell.SM 0.00121f
C3012 XThR.Tn[1] XA.XIR[1].XIC[14].icell.PDM 0.0033f
C3013 XA.XIR[3].XIC[4].icell.PUM VPWR 0.01036f
C3014 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.03976f
C3015 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02698f
C3016 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.SM 0.00383f
C3017 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.03424f
C3018 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00529f
C3019 XA.XIR[12].XIC[3].icell.SM Vbias 0.00701f
C3020 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.11171f
C3021 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.01406f
C3022 XA.XIR[2].XIC[5].icell.Ien VPWR 0.19065f
C3023 XThR.XTB5.Y a_n1049_5611# 0.0093f
C3024 XA.XIR[14].XIC[6].icell.Ien VPWR 0.19119f
C3025 XA.XIR[11].XIC[5].icell.Ien Vbias 0.21238f
C3026 XThR.XTB6.A XThR.Tn[5] 0.00361f
C3027 XA.XIR[2].XIC[2].icell.Ien Iout 0.06483f
C3028 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04522f
C3029 XA.XIR[14].XIC[3].icell.Ien Iout 0.06483f
C3030 XA.XIR[13].XIC[8].icell.PUM VPWR 0.01036f
C3031 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04522f
C3032 XThC.Tn[12] XThR.Tn[5] 0.28062f
C3033 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02698f
C3034 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PUM 0.00131f
C3035 XA.XIR[10].XIC[7].icell.PUM Vbias 0.00347f
C3036 XA.XIR[6].XIC[6].icell.PDM Vbias 0.04058f
C3037 XA.XIR[9].XIC[6].icell.PDM VPWR 0.00863f
C3038 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.15089f
C3039 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00529f
C3040 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02698f
C3041 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04522f
C3042 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PUM 0.00134f
C3043 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00529f
C3044 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.03424f
C3045 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.03976f
C3046 XThR.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.00321f
C3047 a_n1049_5611# XThR.XTB7.Y 0.00153f
C3048 XA.XIR[5].XIC[6].icell.Ien Vbias 0.21238f
C3049 a_5949_9615# VPWR 0.7053f
C3050 XThC.Tn[10] XThR.Tn[1] 0.28062f
C3051 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00212f
C3052 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.15089f
C3053 XThR.Tn[2] XA.XIR[3].XIC[5].icell.Ien 0.00321f
C3054 XA.XIR[10].XIC[12].icell.Ien Iout 0.06483f
C3055 XA.XIR[4].XIC[7].icell.SM Vbias 0.00701f
C3056 XA.XIR[15].XIC[14].icell.Ien VPWR 0.32787f
C3057 XA.XIR[11].XIC[6].icell.SM Iout 0.00388f
C3058 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02698f
C3059 XA.XIR[6].XIC[9].icell.Ien VPWR 0.19065f
C3060 XThR.XTB3.Y XThR.Tn[5] 0.00381f
C3061 XA.XIR[3].XIC[10].icell.PUM Vbias 0.00347f
C3062 XThR.XTBN.Y XThR.Tn[4] 0.60351f
C3063 XThR.Tn[13] XA.XIR[14].XIC[1].icell.Ien 0.00321f
C3064 XA.XIR[10].XIC[10].icell.PDM Iout 0.00112f
C3065 XThR.XTBN.Y a_n997_2667# 0.22784f
C3066 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02698f
C3067 XA.XIR[6].XIC[6].icell.Ien Iout 0.06483f
C3068 XA.XIR[15].XIC[10].icell.Ien Iout 0.06816f
C3069 XA.XIR[11].XIC[9].icell.Ien Vbias 0.21238f
C3070 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.03976f
C3071 XA.XIR[5].XIC[10].icell.SM VPWR 0.00158f
C3072 XA.XIR[8].XIC[5].icell.PDM Vbias 0.04058f
C3073 XA.XIR[7].XIC[1].icell.Ien VPWR 0.19065f
C3074 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.SM 0.00188f
C3075 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02698f
C3076 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00212f
C3077 XA.XIR[13].XIC[14].icell.PDM Iout 0.00112f
C3078 XA.XIR[2].XIC[11].icell.Ien Vbias 0.21238f
C3079 XThC.XTB5.A VPWR 0.82807f
C3080 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.03424f
C3081 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PUM 0.00131f
C3082 XA.XIR[1].XIC[2].icell.Ien VPWR 0.19065f
C3083 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.15089f
C3084 XA.XIR[5].XIC[7].icell.SM Iout 0.00388f
C3085 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.01406f
C3086 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04522f
C3087 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PUM 0.00131f
C3088 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.SM 0.00188f
C3089 XThC.Tn[7] XThR.Tn[13] 0.28062f
C3090 XA.XIR[9].XIC[12].icell.PDM Vbias 0.04058f
C3091 XA.XIR[0].XIC[3].icell.PUM VPWR 0.00971f
C3092 XThC.Tn[0] XThR.Tn[3] 0.2807f
C3093 XA.XIR[12].XIC[9].icell.SM VPWR 0.00158f
C3094 XA.XIR[8].XIC[8].icell.Ien VPWR 0.19065f
C3095 VPWR data[4] 0.5303f
C3096 XThR.Tn[5] XA.XIR[6].XIC[3].icell.Ien 0.00321f
C3097 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02698f
C3098 XThR.XTB4.Y XThR.Tn[6] 0.00605f
C3099 XA.XIR[3].XIC[13].icell.PDM Iout 0.00112f
C3100 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.03011f
C3101 XA.XIR[4].XIC[12].icell.PUM Vbias 0.00347f
C3102 XA.XIR[8].XIC[5].icell.Ien Iout 0.06483f
C3103 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13469f
C3104 XA.XIR[6].XIC[12].icell.SM VPWR 0.00158f
C3105 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04522f
C3106 XA.XIR[10].XIC[2].icell.PDM VPWR 0.00863f
C3107 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06536f
C3108 XA.XIR[3].XIC_15.icell.PDM Vbias 0.04206f
C3109 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00212f
C3110 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.SM 0.00188f
C3111 XA.XIR[15].XIC[0].icell.Ien Vbias 0.17775f
C3112 XThR.Tn[12] XA.XIR[12].XIC[13].icell.PDM 0.0033f
C3113 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00212f
C3114 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.SM 0.00383f
C3115 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00212f
C3116 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04522f
C3117 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11595f
C3118 XThC.XTBN.A XThC.Tn[9] 0.12399f
C3119 XA.XIR[11].XIC[12].icell.PDM Vbias 0.04058f
C3120 XA.XIR[14].XIC[1].icell.Ien Vbias 0.21238f
C3121 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00212f
C3122 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.SM 0.00383f
C3123 XThC.XTBN.Y a_10915_9569# 0.21503f
C3124 XThR.Tn[10] XA.XIR[11].XIC[1].icell.SM 0.00121f
C3125 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PUM 0.00529f
C3126 XA.XIR[7].XIC[7].icell.Ien Vbias 0.21238f
C3127 XThR.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.0033f
C3128 XThR.XTB3.Y a_n1049_6699# 0.0093f
C3129 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.01406f
C3130 XA.XIR[4].XIC_15.icell.PDM Iout 0.0013f
C3131 XA.XIR[1].XIC[8].icell.Ien Vbias 0.21238f
C3132 XThR.Tn[10] XA.XIR[10].XIC[5].icell.PDM 0.0033f
C3133 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.SM 0.00188f
C3134 XA.XIR[9].XIC[14].icell.Ien Vbias 0.21238f
C3135 XA.XIR[14].XIC[11].icell.PUM Vbias 0.00347f
C3136 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PUM 0.00529f
C3137 XThC.Tn[9] XThR.Tn[4] 0.28062f
C3138 XA.XIR[15].XIC[4].icell.SM VPWR 0.00158f
C3139 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.01406f
C3140 XA.XIR[8].XIC[11].icell.SM VPWR 0.00158f
C3141 XThC.XTB7.A XThC.XTB7.B 0.35844f
C3142 XThR.Tn[2] XA.XIR[2].XIC[0].icell.PDM 0.00336f
C3143 XThR.Tn[8] XA.XIR[9].XIC[0].icell.SM 0.00121f
C3144 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.SM 0.00383f
C3145 XA.XIR[12].XIC[11].icell.Ien VPWR 0.19065f
C3146 XThR.Tn[7] XA.XIR[7].XIC[11].icell.PDM 0.0033f
C3147 XA.XIR[0].XIC[9].icell.PUM Vbias 0.00347f
C3148 XA.XIR[15].XIC[1].icell.SM Iout 0.00388f
C3149 XThC.Tn[7] Vbias 2.28504f
C3150 XThR.Tn[13] XA.XIR[14].XIC[5].icell.Ien 0.00321f
C3151 XA.XIR[8].XIC[1].icell.PDM Vbias 0.04058f
C3152 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04522f
C3153 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.04037f
C3154 XThR.Tn[0] XA.XIR[1].XIC[5].icell.Ien 0.00321f
C3155 XA.XIR[7].XIC[8].icell.SM Iout 0.00388f
C3156 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21491f
C3157 XA.XIR[11].XIC_dummy_right.icell.PUM Vbias 0.00248f
C3158 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PUM 0.00529f
C3159 XThC.XTB6.Y XThC.Tn[5] 0.20189f
C3160 XA.XIR[1].XIC[9].icell.SM Iout 0.00388f
C3161 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PUM 0.00131f
C3162 XA.XIR[9].XIC[1].icell.Ien Iout 0.06483f
C3163 XA.XIR[10].XIC[10].icell.SM Iout 0.00388f
C3164 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04522f
C3165 XA.XIR[0].XIC_15.icell.PDM VPWR 0.06796f
C3166 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04522f
C3167 XA.XIR[14].XIC_15.icell.SM Vbias 0.00701f
C3168 XA.XIR[13].XIC[14].icell.SM Iout 0.00388f
C3169 XA.XIR[1].XIC[11].icell.SM Vbias 0.00701f
C3170 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.SM 0.00383f
C3171 XA.XIR[11].XIC[2].icell.SM VPWR 0.00158f
C3172 XA.XIR[15].XIC[8].icell.SM VPWR 0.00158f
C3173 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.01406f
C3174 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[14].icell.Ien 0.00212f
C3175 XA.XIR[12].XIC_dummy_right.icell.SM VPWR 0.00123f
C3176 XA.XIR[4].XIC[0].icell.SM Vbias 0.00675f
C3177 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C3178 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.15089f
C3179 XA.XIR[6].XIC[2].icell.Ien VPWR 0.19065f
C3180 XA.XIR[10].XIC[6].icell.PDM VPWR 0.00863f
C3181 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04522f
C3182 XThR.Tn[9] XA.XIR[10].XIC[7].icell.Ien 0.00321f
C3183 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PUM 0.00529f
C3184 XThR.XTB5.Y VPWR 1.0269f
C3185 XThR.Tn[13] XA.XIR[14].XIC[9].icell.Ien 0.00321f
C3186 XA.XIR[3].XIC[3].icell.PUM Vbias 0.00347f
C3187 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04522f
C3188 XA.XIR[5].XIC[3].icell.SM VPWR 0.00158f
C3189 XA.XIR[2].XIC[4].icell.Ien Vbias 0.21238f
C3190 XThR.Tn[3] VPWR 6.72245f
C3191 XA.XIR[14].XIC[5].icell.Ien Vbias 0.21238f
C3192 XA.XIR[5].XIC[0].icell.SM Iout 0.00388f
C3193 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04522f
C3194 XA.XIR[4].XIC[6].icell.PUM VPWR 0.01036f
C3195 XThC.XTBN.Y XThC.Tn[1] 0.7252f
C3196 XThC.Tn[0] XA.XIR[15].XIC_dummy_left.icell.Iout 0.00111f
C3197 XA.XIR[7].XIC[14].icell.SM Vbias 0.00701f
C3198 XA.XIR[13].XIC[7].icell.PUM Vbias 0.00347f
C3199 XThR.XTB7.Y VPWR 1.14767f
C3200 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.SM 0.00188f
C3201 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00212f
C3202 XA.XIR[3].XIC[9].icell.PDM VPWR 0.00863f
C3203 XThR.Tn[6] XA.XIR[7].XIC[7].icell.Ien 0.00321f
C3204 XA.XIR[9].XIC[5].icell.PDM Vbias 0.04058f
C3205 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00212f
C3206 XA.XIR[8].XIC[1].icell.Ien VPWR 0.19065f
C3207 XThR.Tn[8] XA.XIR[9].XIC[4].icell.SM 0.00121f
C3208 XA.XIR[12].XIC[8].icell.PUM Vbias 0.00347f
C3209 XA.XIR[3].XIC[6].icell.PDM Iout 0.00112f
C3210 XThC.XTB7.B a_5949_9615# 0.00927f
C3211 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00529f
C3212 XA.XIR[2].XIC[8].icell.SM VPWR 0.00158f
C3213 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.01406f
C3214 XThC.XTB4.Y XThC.Tn[5] 0.00814f
C3215 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.01406f
C3216 a_3773_9615# Vbias 0.00826f
C3217 XA.XIR[2].XIC[5].icell.SM Iout 0.00388f
C3218 XThC.XTB3.Y XThC.Tn[9] 0.00285f
C3219 XThR.XTB4.Y XThR.Tn[4] 0.00757f
C3220 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.SM 0.00188f
C3221 XA.XIR[13].XIC[12].icell.Ien Iout 0.06483f
C3222 XThC.Tn[0] XThR.Tn[8] 0.28063f
C3223 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04522f
C3224 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.03424f
C3225 XThC.XTB6.Y a_10051_9569# 0.07626f
C3226 XA.XIR[14].XIC[6].icell.SM Iout 0.00388f
C3227 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.03976f
C3228 XThC.Tn[7] XThR.Tn[6] 0.28062f
C3229 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04522f
C3230 XThR.XTB4.Y a_n997_2667# 0.07199f
C3231 XThC.Tn[0] XA.XIR[3].XIC_dummy_left.icell.Iout 0.00111f
C3232 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.03976f
C3233 XA.XIR[6].XIC[8].icell.Ien Vbias 0.21238f
C3234 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00212f
C3235 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.SM 0.00188f
C3236 XA.XIR[9].XIC[8].icell.Ien VPWR 0.19065f
C3237 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00212f
C3238 XA.XIR[13].XIC[10].icell.PDM Iout 0.00112f
C3239 XA.XIR[14].XIC[9].icell.Ien Vbias 0.21238f
C3240 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PUM 0.00131f
C3241 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.01406f
C3242 XThC.XTB5.A XThC.XTB7.B 0.30355f
C3243 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PUM 0.00529f
C3244 XThR.Tn[3] XA.XIR[4].XIC[6].icell.Ien 0.00321f
C3245 XA.XIR[9].XIC[5].icell.Ien Iout 0.06483f
C3246 XA.XIR[5].XIC[9].icell.SM Vbias 0.00701f
C3247 XA.XIR[7].XIC[0].icell.Ien Vbias 0.21102f
C3248 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.03976f
C3249 XA.XIR[12].XIC[10].icell.PUM VPWR 0.01036f
C3250 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04522f
C3251 XThR.Tn[2] XA.XIR[3].XIC[8].icell.SM 0.00121f
C3252 XA.XIR[1].XIC[1].icell.Ien Vbias 0.21238f
C3253 XThR.XTB7.A XThR.Tn[6] 0.1056f
C3254 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00529f
C3255 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00212f
C3256 XThC.Tn[1] XThR.Tn[5] 0.28062f
C3257 XA.XIR[2].XIC[13].icell.PUM VPWR 0.01036f
C3258 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.SM 0.00188f
C3259 XA.XIR[10].XIC_15.icell.PDM VPWR 0.06959f
C3260 XA.XIR[15].XIC_15.icell.Ien VPWR 0.36693f
C3261 XThR.Tn[7] XA.XIR[7].XIC[4].icell.PDM 0.0033f
C3262 XThR.Tn[2] XA.XIR[2].XIC[12].icell.PDM 0.0033f
C3263 XA.XIR[0].XIC[2].icell.PUM Vbias 0.00347f
C3264 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.SM 0.00188f
C3265 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.SM 0.00188f
C3266 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.SM 0.00383f
C3267 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.01406f
C3268 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00212f
C3269 XA.XIR[8].XIC[7].icell.Ien Vbias 0.21238f
C3270 XA.XIR[6].XIC[9].icell.SM Iout 0.00388f
C3271 XThR.Tn[4] XA.XIR[5].XIC[6].icell.Ien 0.00321f
C3272 XA.XIR[7].XIC[4].icell.SM VPWR 0.00158f
C3273 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PUM 0.00529f
C3274 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.15089f
C3275 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Ien 0.00529f
C3276 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01193f
C3277 a_8739_9569# VPWR 0.00582f
C3278 XA.XIR[13].XIC[2].icell.PDM VPWR 0.00863f
C3279 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00212f
C3280 XThR.Tn[1] XA.XIR[2].XIC[12].icell.Ien 0.00321f
C3281 XA.XIR[11].XIC[10].icell.Ien Vbias 0.21238f
C3282 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04522f
C3283 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00212f
C3284 XA.XIR[7].XIC[1].icell.SM Iout 0.00388f
C3285 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.SM 0.00188f
C3286 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C3287 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.SM 0.00188f
C3288 XA.XIR[1].XIC[5].icell.SM VPWR 0.00158f
C3289 XA.XIR[6].XIC[11].icell.SM Vbias 0.00701f
C3290 XA.XIR[9].XIC[11].icell.SM VPWR 0.00158f
C3291 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.SM 0.00188f
C3292 XA.XIR[12].XIC[3].icell.PDM VPWR 0.00863f
C3293 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.03976f
C3294 XA.XIR[1].XIC[2].icell.SM Iout 0.00388f
C3295 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.01406f
C3296 XA.XIR[5].XIC[14].icell.PUM Vbias 0.00347f
C3297 XA.XIR[14].XIC[12].icell.PDM Vbias 0.04058f
C3298 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01096f
C3299 XThR.Tn[1] XA.XIR[1].XIC[7].icell.PDM 0.0033f
C3300 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.01406f
C3301 XThR.Tn[5] XA.XIR[6].XIC[6].icell.SM 0.00121f
C3302 XA.XIR[3].XIC_15.icell.Ien VPWR 0.25675f
C3303 XThR.Tn[6] XA.XIR[7].XIC[14].icell.SM 0.00121f
C3304 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PUM 0.00131f
C3305 XA.XIR[8].XIC[8].icell.SM Iout 0.00388f
C3306 XA.XIR[11].XIC[0].icell.Ien Iout 0.06474f
C3307 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.002f
C3308 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.01406f
C3309 XThR.Tn[11] XA.XIR[12].XIC[2].icell.SM 0.00121f
C3310 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.15089f
C3311 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.03424f
C3312 XA.XIR[8].XIC_dummy_left.icell.Ien Vbias 0.00342f
C3313 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.SM 0.00383f
C3314 XA.XIR[10].XIC[1].icell.Ien Iout 0.06483f
C3315 XA.XIR[15].XIC[3].icell.SM Vbias 0.00701f
C3316 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.15089f
C3317 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.25822f
C3318 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01776f
C3319 XThR.Tn[8] XA.XIR[8].XIC[14].icell.PDM 0.0033f
C3320 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C3321 XA.XIR[5].XIC_15.icell.SM VPWR 0.00276f
C3322 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PUM 0.00529f
C3323 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.SM 0.00383f
C3324 XA.XIR[2].XIC_dummy_right.icell.Ien Vbias 0.00287f
C3325 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PUM 0.00131f
C3326 XA.XIR[7].XIC[10].icell.SM Vbias 0.00701f
C3327 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.SM 0.00383f
C3328 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.01406f
C3329 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02698f
C3330 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.15089f
C3331 XThR.Tn[7] XA.XIR[8].XIC[13].icell.Ien 0.00321f
C3332 XA.XIR[5].XIC[1].icell.PDM Vbias 0.04058f
C3333 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00529f
C3334 XA.XIR[14].XIC_dummy_right.icell.PUM Vbias 0.00248f
C3335 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.01406f
C3336 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.15089f
C3337 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.01406f
C3338 XA.XIR[3].XIC[2].icell.PDM VPWR 0.00863f
C3339 XThR.Tn[8] VPWR 7.59166f
C3340 XThR.Tn[6] XA.XIR[7].XIC[0].icell.Ien 0.00321f
C3341 XThR.Tn[14] XA.XIR[14].XIC[9].icell.PDM 0.0033f
C3342 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35783f
C3343 XA.XIR[13].XIC[10].icell.SM Iout 0.00388f
C3344 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.03424f
C3345 XThC.Tn[5] XA.XIR[0].XIC[6].icell.Ien 0.00164f
C3346 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C3347 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.01406f
C3348 XA.XIR[2].XIC[1].icell.SM VPWR 0.00158f
C3349 XA.XIR[0].XIC[14].icell.PDM Vbias 0.04065f
C3350 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11403f
C3351 XThC.Tn[11] VPWR 6.92826f
C3352 XThR.Tn[5] XA.XIR[5].XIC[14].icell.PDM 0.0033f
C3353 XThR.Tn[2] XA.XIR[2].XIC[1].icell.PDM 0.0033f
C3354 XA.XIR[14].XIC[2].icell.SM VPWR 0.00158f
C3355 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04522f
C3356 XA.XIR[11].XIC[1].icell.SM Vbias 0.00701f
C3357 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PUM 0.00529f
C3358 XA.XIR[8].XIC[14].icell.SM Vbias 0.00701f
C3359 XThC.XTBN.A XThC.Tn[7] 0.01439f
C3360 XThR.Tn[0] XA.XIR[1].XIC[8].icell.SM 0.00121f
C3361 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.03424f
C3362 XA.XIR[13].XIC[6].icell.PDM VPWR 0.00863f
C3363 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00212f
C3364 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.03976f
C3365 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.01406f
C3366 XThR.Tn[0] XThR.XTB2.Y 0.00125f
C3367 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00529f
C3368 XA.XIR[10].XIC[5].icell.PDM Vbias 0.04058f
C3369 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Iout 0.00347f
C3370 XA.XIR[10].XIC_15.icell.SM Iout 0.0047f
C3371 XA.XIR[6].XIC[1].icell.Ien Vbias 0.21238f
C3372 XThC.Tn[10] XThR.Tn[9] 0.28062f
C3373 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02698f
C3374 XA.XIR[12].XIC[7].icell.PDM VPWR 0.00863f
C3375 XThC.Tn[7] XThR.Tn[4] 0.28062f
C3376 XThR.Tn[0] XA.XIR[0].XIC[11].icell.PDM 0.0033f
C3377 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.01406f
C3378 XA.XIR[5].XIC[2].icell.SM Vbias 0.00701f
C3379 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00212f
C3380 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.SM 0.00188f
C3381 XA.XIR[10].XIC[11].icell.SM VPWR 0.00158f
C3382 XA.XIR[12].XIC[4].icell.PDM Iout 0.00112f
C3383 XA.XIR[11].XIC[7].icell.PUM VPWR 0.01036f
C3384 XThR.Tn[2] Vbias 3.71826f
C3385 XA.XIR[0].XIC[14].icell.Ien Iout 0.06455f
C3386 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02698f
C3387 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.01406f
C3388 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PUM 0.00209f
C3389 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00529f
C3390 XA.XIR[4].XIC[5].icell.PUM Vbias 0.00347f
C3391 XThR.Tn[2] XA.XIR[3].XIC[1].icell.SM 0.00121f
C3392 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.03982f
C3393 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.01406f
C3394 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.01406f
C3395 XA.XIR[6].XIC[5].icell.SM VPWR 0.00158f
C3396 XA.XIR[10].XIC[8].icell.Ien VPWR 0.19065f
C3397 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Iout 0.00401f
C3398 XA.XIR[15].XIC[9].icell.SM VPWR 0.00158f
C3399 XA.XIR[3].XIC[8].icell.PDM Vbias 0.04058f
C3400 XThR.Tn[2] XA.XIR[2].XIC[5].icell.PDM 0.0033f
C3401 XThR.XTB7.A XThR.Tn[4] 0.02736f
C3402 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PUM 0.00529f
C3403 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04522f
C3404 XA.XIR[10].XIC[5].icell.Ien Iout 0.06483f
C3405 XA.XIR[6].XIC[2].icell.SM Iout 0.00388f
C3406 XA.XIR[5].XIC[8].icell.PUM VPWR 0.01036f
C3407 data[6] data[7] 0.04128f
C3408 XThR.Tn[13] XA.XIR[14].XIC[10].icell.Ien 0.00321f
C3409 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PUM 0.00131f
C3410 XA.XIR[2].XIC[7].icell.SM Vbias 0.00701f
C3411 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00212f
C3412 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C3413 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00529f
C3414 XA.XIR[4].XIC[11].icell.PDM VPWR 0.00863f
C3415 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00212f
C3416 XThR.XTB5.Y a_n997_1803# 0.06458f
C3417 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02698f
C3418 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.03976f
C3419 XA.XIR[12].XIC[11].icell.PDM VPWR 0.00863f
C3420 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00529f
C3421 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00212f
C3422 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.SM 0.00188f
C3423 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.03976f
C3424 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.SM 0.00383f
C3425 XThR.Tn[6] XA.XIR[7].XIC[10].icell.SM 0.00121f
C3426 XA.XIR[3].XIC[11].icell.Ien VPWR 0.19065f
C3427 XA.XIR[4].XIC[8].icell.PDM Iout 0.00112f
C3428 XThC.Tn[5] Iout 0.84073f
C3429 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04522f
C3430 XThC.Tn[8] XThR.Tn[11] 0.28062f
C3431 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12] 0.0033f
C3432 XA.XIR[9].XIC[7].icell.Ien Vbias 0.21238f
C3433 XA.XIR[8].XIC[4].icell.SM VPWR 0.00158f
C3434 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.03424f
C3435 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.SM 0.00188f
C3436 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00212f
C3437 XA.XIR[3].XIC[8].icell.Ien Iout 0.06483f
C3438 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PUM 0.00131f
C3439 VPWR data[0] 0.52929f
C3440 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04522f
C3441 XA.XIR[10].XIC[13].icell.Ien VPWR 0.19065f
C3442 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00529f
C3443 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.SM 0.00383f
C3444 XA.XIR[8].XIC[1].icell.SM Iout 0.00388f
C3445 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[7].icell.Ien 0.00212f
C3446 XA.XIR[14].XIC[0].icell.PDM Iout 0.00112f
C3447 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.SM 0.00188f
C3448 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.SM 0.00188f
C3449 XThR.XTB7.Y a_n997_1803# 0.00571f
C3450 VPWR bias[1] 1.23968f
C3451 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02698f
C3452 XA.XIR[10].XIC[9].icell.Ien Iout 0.06483f
C3453 XA.XIR[15].XIC[11].icell.Ien VPWR 0.32782f
C3454 XA.XIR[13].XIC_15.icell.PDM VPWR 0.06959f
C3455 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.SM 0.00188f
C3456 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.SM 0.00383f
C3457 XA.XIR[2].XIC[12].icell.PUM Vbias 0.00347f
C3458 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C3459 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PUM 0.00529f
C3460 XA.XIR[4].XIC[13].icell.Ien VPWR 0.19065f
C3461 XThC.XTB7.B a_8739_9569# 0.0168f
C3462 XThR.Tn[3] XA.XIR[4].XIC[9].icell.SM 0.00121f
C3463 XA.XIR[9].XIC[8].icell.SM Iout 0.00388f
C3464 XA.XIR[7].XIC[3].icell.SM Vbias 0.00701f
C3465 XThR.Tn[14] XA.XIR[15].XIC[6].icell.Ien 0.00321f
C3466 XA.XIR[14].XIC[10].icell.Ien Vbias 0.21238f
C3467 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.15089f
C3468 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.SM 0.00383f
C3469 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PUM 0.00529f
C3470 XA.XIR[1].XIC[4].icell.SM Vbias 0.00701f
C3471 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04522f
C3472 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00212f
C3473 XA.XIR[15].XIC[2].icell.PUM VPWR 0.01036f
C3474 XA.XIR[3].XIC[11].icell.SM Iout 0.00388f
C3475 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04522f
C3476 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04f
C3477 XA.XIR[12].XIC[2].icell.PDM Vbias 0.04058f
C3478 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02698f
C3479 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.SM 0.00383f
C3480 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.SM 0.00383f
C3481 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02698f
C3482 XThC.XTB3.Y XThC.Tn[7] 0.00819f
C3483 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.15089f
C3484 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04522f
C3485 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02698f
C3486 XThR.XTBN.A a_n997_3755# 0.01939f
C3487 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PUM 0.00529f
C3488 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.SM 0.00383f
C3489 XThC.Tn[8] XThR.Tn[7] 0.28062f
C3490 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00529f
C3491 XA.XIR[0].XIC[7].icell.PDM Vbias 0.04063f
C3492 XA.XIR[2].XIC_15.icell.PDM Iout 0.0013f
C3493 XThR.Tn[13] XA.XIR[14].XIC[1].icell.SM 0.00121f
C3494 XA.XIR[8].XIC[10].icell.SM Vbias 0.00701f
C3495 XA.XIR[7].XIC[9].icell.PUM VPWR 0.01036f
C3496 XThR.Tn[4] XA.XIR[5].XIC[9].icell.SM 0.00121f
C3497 XA.XIR[11].XIC[2].icell.PUM Vbias 0.00347f
C3498 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08017f
C3499 XA.XIR[15].XIC_dummy_right.icell.SM VPWR 0.00123f
C3500 XThC.Tn[13] XThR.Tn[2] 0.28063f
C3501 XThC.Tn[4] XThC.Tn[5] 0.42055f
C3502 XThC.Tn[11] XThR.Tn[12] 0.28062f
C3503 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01897f
C3504 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.01406f
C3505 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04522f
C3506 XThR.Tn[13] XA.XIR[13].XIC[5].icell.PDM 0.0033f
C3507 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.SM 0.00188f
C3508 XA.XIR[1].XIC[10].icell.PUM VPWR 0.01036f
C3509 XThR.Tn[0] XA.XIR[1].XIC[1].icell.SM 0.00121f
C3510 XA.XIR[9].XIC[0].icell.SM VPWR 0.00158f
C3511 XA.XIR[10].XIC[12].icell.PDM Iout 0.00112f
C3512 XA.XIR[13].XIC[1].icell.Ien Iout 0.06483f
C3513 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.SM 0.00383f
C3514 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01776f
C3515 XA.XIR[5].XIC_dummy_left.icell.Ien Vbias 0.00342f
C3516 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.PUM 0.00112f
C3517 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PUM 0.00131f
C3518 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.03976f
C3519 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00212f
C3520 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.SM 0.00188f
C3521 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06536f
C3522 XThR.Tn[0] XA.XIR[0].XIC[4].icell.PDM 0.0033f
C3523 XA.XIR[0].XIC[10].icell.Ien VPWR 0.19003f
C3524 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.15089f
C3525 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.01406f
C3526 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PUM 0.00131f
C3527 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.SM 0.00383f
C3528 XThR.Tn[12] XA.XIR[12].XIC[7].icell.PDM 0.0033f
C3529 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00529f
C3530 XA.XIR[0].XIC[7].icell.Ien Iout 0.06455f
C3531 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C3532 XA.XIR[9].XIC[14].icell.SM Vbias 0.00701f
C3533 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PUM 0.00529f
C3534 XA.XIR[3].XIC_dummy_right.icell.SM VPWR 0.00123f
C3535 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01718f
C3536 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PUM 0.00131f
C3537 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.SM 0.00188f
C3538 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00212f
C3539 XThC.Tn[10] XThR.Tn[10] 0.28062f
C3540 XThR.Tn[9] XA.XIR[10].XIC[3].icell.SM 0.00121f
C3541 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PUM 0.00529f
C3542 XA.XIR[15].XIC[8].icell.PUM Vbias 0.00347f
C3543 XA.XIR[7].XIC[14].icell.PDM VPWR 0.00873f
C3544 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PUM 0.00131f
C3545 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04522f
C3546 XA.XIR[8].XIC[0].icell.Ien Vbias 0.21102f
C3547 XThC.XTB7.B XThC.Tn[11] 0.03903f
C3548 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00212f
C3549 a_n1049_5611# VPWR 0.71844f
C3550 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04522f
C3551 XA.XIR[2].XIC[0].icell.SM Vbias 0.00675f
C3552 XA.XIR[1].XIC_15.icell.PDM VPWR 0.06959f
C3553 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06536f
C3554 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.SM 0.00188f
C3555 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00212f
C3556 XA.XIR[14].XIC[1].icell.SM Vbias 0.00701f
C3557 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.SM 0.00188f
C3558 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10] 0.0033f
C3559 XA.XIR[4].XIC[4].icell.PDM VPWR 0.00863f
C3560 XA.XIR[10].XIC[12].icell.PUM VPWR 0.01036f
C3561 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.SM 0.00383f
C3562 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00529f
C3563 XA.XIR[13].XIC[5].icell.PDM Vbias 0.04058f
C3564 XA.XIR[13].XIC_15.icell.SM Iout 0.0047f
C3565 XThR.Tn[6] XA.XIR[7].XIC[3].icell.SM 0.00121f
C3566 XA.XIR[3].XIC[4].icell.Ien VPWR 0.19065f
C3567 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PUM 0.00529f
C3568 XThR.Tn[12] XA.XIR[12].XIC[11].icell.PDM 0.0033f
C3569 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PUM 0.00529f
C3570 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PDM 0.00594f
C3571 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.SM 0.00188f
C3572 XA.XIR[15].XIC[10].icell.PUM VPWR 0.01036f
C3573 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.01406f
C3574 XA.XIR[12].XIC[6].icell.PDM Vbias 0.04058f
C3575 XA.XIR[3].XIC[1].icell.Ien Iout 0.06483f
C3576 XA.XIR[2].XIC[6].icell.PUM VPWR 0.01036f
C3577 XThC.XTB3.Y a_3773_9615# 0.00124f
C3578 XA.XIR[13].XIC[11].icell.SM VPWR 0.00158f
C3579 XThR.XTBN.A XThR.Tn[11] 0.11968f
C3580 XA.XIR[14].XIC[7].icell.PUM VPWR 0.01036f
C3581 XA.XIR[11].XIC[6].icell.PUM Vbias 0.00347f
C3582 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04522f
C3583 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.03976f
C3584 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.SM 0.00188f
C3585 XThR.XTBN.Y a_n1049_7493# 0.08456f
C3586 a_3773_9615# XThC.Tn[2] 0.01175f
C3587 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00212f
C3588 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.SM 0.00383f
C3589 XThR.Tn[1] XA.XIR[2].XIC[5].icell.Ien 0.00321f
C3590 XA.XIR[13].XIC[8].icell.Ien VPWR 0.19065f
C3591 XThR.XTBN.Y XA.XIR[14].XIC_dummy_left.icell.Iout 0.00119f
C3592 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.SM 0.00188f
C3593 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00212f
C3594 XA.XIR[6].XIC[4].icell.SM Vbias 0.00701f
C3595 XA.XIR[10].XIC[7].icell.Ien Vbias 0.21238f
C3596 XA.XIR[9].XIC[4].icell.SM VPWR 0.00158f
C3597 XA.XIR[13].XIC[5].icell.Ien Iout 0.06483f
C3598 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00529f
C3599 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.15089f
C3600 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PDM 0.00182f
C3601 XA.XIR[9].XIC[1].icell.SM Iout 0.00388f
C3602 XA.XIR[11].XIC[0].icell.PDM VPWR 0.00863f
C3603 XA.XIR[5].XIC[7].icell.PUM Vbias 0.00347f
C3604 XThR.Tn[3] XA.XIR[4].XIC[2].icell.SM 0.00121f
C3605 XThC.Tn[0] VPWR 6.02351f
C3606 XA.XIR[12].XIC[6].icell.Ien Iout 0.06483f
C3607 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04522f
C3608 XThC.XTB1.Y XThC.Tn[7] 0.0045f
C3609 XA.XIR[7].XIC_15.icell.SM Vbias 0.00701f
C3610 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.SM 0.00188f
C3611 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00212f
C3612 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PUM 0.00131f
C3613 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PUM 0.00131f
C3614 XA.XIR[4].XIC[10].icell.PDM Vbias 0.04058f
C3615 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14] 0.0033f
C3616 XThR.XTB6.A data[4] 0.48493f
C3617 XA.XIR[11].XIC[9].icell.PDM Iout 0.00112f
C3618 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00529f
C3619 XA.XIR[6].XIC[10].icell.PUM VPWR 0.01036f
C3620 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.01406f
C3621 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.15089f
C3622 XThC.Tn[8] XThR.Tn[14] 0.28062f
C3623 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PUM 0.00134f
C3624 XA.XIR[3].XIC[10].icell.Ien Vbias 0.21238f
C3625 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PUM 0.00131f
C3626 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04522f
C3627 XThC.XTB7.B data[0] 0.0138f
C3628 XA.XIR[8].XIC[3].icell.SM Vbias 0.00701f
C3629 XA.XIR[7].XIC[2].icell.PUM VPWR 0.01036f
C3630 XA.XIR[5].XIC[13].icell.PDM VPWR 0.00863f
C3631 XThR.Tn[4] XA.XIR[5].XIC[2].icell.SM 0.00121f
C3632 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PUM 0.00487f
C3633 XA.XIR[13].XIC[13].icell.Ien VPWR 0.19065f
C3634 XThR.Tn[8] XA.XIR[8].XIC[7].icell.PDM 0.0033f
C3635 XThC.XTB7.Y a_7875_9569# 0.00476f
C3636 XThR.XTBN.A XThR.Tn[7] 0.01439f
C3637 XA.XIR[1].XIC[3].icell.PUM VPWR 0.01036f
C3638 XA.XIR[5].XIC[10].icell.PDM Iout 0.00112f
C3639 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C3640 XA.XIR[13].XIC[9].icell.Ien Iout 0.06483f
C3641 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C3642 XThR.Tn[7] XA.XIR[8].XIC[6].icell.Ien 0.00321f
C3643 XA.XIR[4].XIC[10].icell.Ien Iout 0.06483f
C3644 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.SM 0.00383f
C3645 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PUM 0.00529f
C3646 XThR.XTB3.Y data[4] 0.03253f
C3647 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PUM 0.00131f
C3648 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.01406f
C3649 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.15089f
C3650 XA.XIR[8].XIC[9].icell.PUM VPWR 0.01036f
C3651 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PUM 0.00529f
C3652 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PUM 0.00209f
C3653 XA.XIR[9].XIC[10].icell.SM Vbias 0.00701f
C3654 XA.XIR[0].XIC[3].icell.Ien VPWR 0.19003f
C3655 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.SM 0.00188f
C3656 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PUM 0.00131f
C3657 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.SM 0.00383f
C3658 XA.XIR[4].XIC[12].icell.Ien Vbias 0.21238f
C3659 a_6243_9615# XThC.Tn[5] 0.00158f
C3660 XA.XIR[12].XIC_15.icell.PDM Vbias 0.04206f
C3661 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.01406f
C3662 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00529f
C3663 XA.XIR[0].XIC[0].icell.Ien Iout 0.06447f
C3664 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.01406f
C3665 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[8].icell.SM 0.00383f
C3666 XA.XIR[10].XIC[0].icell.SM VPWR 0.00158f
C3667 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.01406f
C3668 XA.XIR[6].XIC_15.icell.PDM VPWR 0.06959f
C3669 XThR.Tn[5] XA.XIR[5].XIC[7].icell.PDM 0.0033f
C3670 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.33685f
C3671 XA.XIR[3].XIC[13].icell.SM Vbias 0.00701f
C3672 XA.XIR[10].XIC[14].icell.Ien VPWR 0.1907f
C3673 XA.XIR[15].XIC[1].icell.PUM Vbias 0.00347f
C3674 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02698f
C3675 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.SM 0.00188f
C3676 XA.XIR[10].XIC[10].icell.Ien Iout 0.06483f
C3677 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00529f
C3678 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PUM 0.00529f
C3679 XA.XIR[5].XIC[12].icell.Ien Iout 0.06483f
C3680 XA.XIR[14].XIC[2].icell.PUM Vbias 0.00347f
C3681 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08017f
C3682 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.03976f
C3683 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PUM 0.00487f
C3684 XA.XIR[7].XIC[8].icell.PUM Vbias 0.00347f
C3685 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.SM 0.00188f
C3686 XThC.Tn[6] XThR.Tn[11] 0.28062f
C3687 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00212f
C3688 XA.XIR[4].XIC[13].icell.SM Iout 0.00388f
C3689 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00529f
C3690 XA.XIR[13].XIC[12].icell.PDM Iout 0.00112f
C3691 XA.XIR[1].XIC[9].icell.PUM Vbias 0.00347f
C3692 XA.XIR[8].XIC[14].icell.PDM VPWR 0.00873f
C3693 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.03011f
C3694 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01193f
C3695 XThC.XTB5.Y Vbias 0.0131f
C3696 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.15089f
C3697 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35783f
C3698 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.03976f
C3699 XA.XIR[15].XIC[4].icell.PDM Iout 0.00112f
C3700 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C3701 XA.XIR[0].XIC[9].icell.Ien Vbias 0.21246f
C3702 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PUM 0.00131f
C3703 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PUM 0.00529f
C3704 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.03424f
C3705 XA.XIR[12].XIC_15.icell.PUM Vbias 0.00347f
C3706 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C3707 XThR.Tn[12] XA.XIR[13].XIC[11].icell.SM 0.00121f
C3708 XA.XIR[7].XIC[11].icell.PDM Iout 0.00112f
C3709 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.15089f
C3710 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PUM 0.00131f
C3711 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PUM 0.00504f
C3712 XThC.Tn[10] XThR.Tn[13] 0.28062f
C3713 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PUM 0.00529f
C3714 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.SM 0.00383f
C3715 XThR.Tn[12] XA.XIR[13].XIC[8].icell.Ien 0.00321f
C3716 XA.XIR[1].XIC[12].icell.PDM Iout 0.00112f
C3717 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00529f
C3718 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04522f
C3719 XA.XIR[12].XIC[2].icell.Ien VPWR 0.19065f
C3720 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04522f
C3721 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11595f
C3722 XA.XIR[0].XIC[13].icell.SM VPWR 0.00158f
C3723 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.SM 0.00383f
C3724 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.15089f
C3725 XThC.Tn[12] XThR.Tn[3] 0.28062f
C3726 XA.XIR[5].XIC[0].icell.Ien Vbias 0.21102f
C3727 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.SM 0.00188f
C3728 XA.XIR[1].XIC[14].icell.PDM Vbias 0.04058f
C3729 XA.XIR[0].XIC[10].icell.SM Iout 0.00367f
C3730 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C3731 XA.XIR[11].XIC[5].icell.PDM VPWR 0.00863f
C3732 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.SM 0.00383f
C3733 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01193f
C3734 XThC.XTBN.Y Vbias 0.13985f
C3735 XA.XIR[4].XIC[3].icell.PDM Vbias 0.04058f
C3736 XThC.Tn[2] XThR.Tn[2] 0.28062f
C3737 XThC.Tn[6] XThR.Tn[7] 0.28062f
C3738 XThC.Tn[0] XThR.Tn[12] 0.28064f
C3739 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00212f
C3740 XA.XIR[13].XIC[12].icell.PUM VPWR 0.01036f
C3741 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C3742 XA.XIR[10].XIC[4].icell.SM VPWR 0.00158f
C3743 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.03011f
C3744 XA.XIR[6].XIC[3].icell.PUM VPWR 0.01036f
C3745 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.SM 0.00383f
C3746 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.SM 0.00188f
C3747 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.15119f
C3748 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PUM 0.00131f
C3749 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.01406f
C3750 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Ien 0.00217f
C3751 XA.XIR[3].XIC[3].icell.Ien Vbias 0.21238f
C3752 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PUM 0.00529f
C3753 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.SM 0.00383f
C3754 XA.XIR[10].XIC[1].icell.SM Iout 0.00388f
C3755 XA.XIR[5].XIC[6].icell.PDM VPWR 0.00863f
C3756 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00529f
C3757 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C3758 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00212f
C3759 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.SM 0.00188f
C3760 XA.XIR[8].XIC_15.icell.SM Vbias 0.00701f
C3761 XA.XIR[2].XIC[5].icell.PUM Vbias 0.00347f
C3762 XA.XIR[7].XIC[13].icell.Ien Iout 0.06483f
C3763 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.01406f
C3764 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.01406f
C3765 XA.XIR[14].XIC[6].icell.PUM Vbias 0.00347f
C3766 XThR.Tn[12] XA.XIR[13].XIC[13].icell.Ien 0.00321f
C3767 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.SM 0.00383f
C3768 XA.XIR[5].XIC[3].icell.PDM Iout 0.00112f
C3769 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02698f
C3770 XA.XIR[4].XIC[6].icell.Ien VPWR 0.19065f
C3771 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00529f
C3772 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08027f
C3773 XA.XIR[1].XIC[14].icell.Ien Iout 0.06483f
C3774 XA.XIR[7].XIC_dummy_right.icell.PUM Vbias 0.00248f
C3775 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C3776 XA.XIR[12].XIC[11].icell.SM Vbias 0.00701f
C3777 XA.XIR[13].XIC[7].icell.Ien Vbias 0.21238f
C3778 XA.XIR[4].XIC[3].icell.Ien Iout 0.06483f
C3779 XA.XIR[3].XIC[7].icell.SM VPWR 0.00158f
C3780 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PUM 0.00131f
C3781 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C3782 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.SM 0.00188f
C3783 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00212f
C3784 XThC.Tn[10] Vbias 2.3362f
C3785 XA.XIR[8].XIC[2].icell.PUM VPWR 0.01036f
C3786 XA.XIR[9].XIC[3].icell.SM Vbias 0.00701f
C3787 XA.XIR[0].XIC[14].icell.SM Iout 0.00367f
C3788 XA.XIR[3].XIC[4].icell.SM Iout 0.00388f
C3789 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.03976f
C3790 XA.XIR[12].XIC[8].icell.Ien Vbias 0.21238f
C3791 XThC.XTB7.B XThC.Tn[0] 0.00139f
C3792 XA.XIR[2].XIC[11].icell.PDM VPWR 0.00863f
C3793 XA.XIR[10].XIC[8].icell.SM VPWR 0.00158f
C3794 a_4861_9615# Vbias 0.00521f
C3795 XThR.XTB2.Y a_n1049_5317# 0.00844f
C3796 XA.XIR[2].XIC[8].icell.PDM Iout 0.00112f
C3797 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.SM 0.00383f
C3798 XThC.XTB6.Y XThC.Tn[8] 0.02461f
C3799 XA.XIR[10].XIC[0].icell.PDM Vbias 0.04002f
C3800 XA.XIR[14].XIC[9].icell.PDM Iout 0.00112f
C3801 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.SM 0.00188f
C3802 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PUM 0.00529f
C3803 XThR.Tn[1] XA.XIR[2].XIC[8].icell.SM 0.00121f
C3804 XThC.XTB5.Y XThC.Tn[13] 0.00145f
C3805 XThR.XTB6.Y a_n997_3755# 0.0046f
C3806 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01415f
C3807 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02698f
C3808 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.SM 0.00383f
C3809 XA.XIR[6].XIC[9].icell.PUM Vbias 0.00347f
C3810 XA.XIR[9].XIC[9].icell.PUM VPWR 0.01036f
C3811 XThR.Tn[0] Iout 1.16633f
C3812 XThR.Tn[9] XA.XIR[9].XIC[13].icell.PDM 0.0033f
C3813 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.01406f
C3814 XThR.Tn[5] Vbias 3.71719f
C3815 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04522f
C3816 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04522f
C3817 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.03424f
C3818 XA.XIR[7].XIC[1].icell.PUM Vbias 0.00347f
C3819 XA.XIR[5].XIC[12].icell.PDM Vbias 0.04058f
C3820 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PUM 0.00131f
C3821 XThC.XTB6.A a_7875_9569# 0.00149f
C3822 XThR.Tn[14] XA.XIR[15].XIC[2].icell.SM 0.00121f
C3823 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.SM 0.00383f
C3824 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C3825 XA.XIR[11].XIC[0].icell.PUM VPWR 0.01036f
C3826 XA.XIR[3].XIC[12].icell.PUM VPWR 0.01036f
C3827 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.03976f
C3828 XA.XIR[1].XIC[2].icell.PUM Vbias 0.00347f
C3829 XThC.Tn[0] XA.XIR[10].XIC_dummy_left.icell.Iout 0.00111f
C3830 XThR.Tn[3] XA.XIR[3].XIC[10].icell.PDM 0.0033f
C3831 XA.XIR[12].XIC[13].icell.Ien Vbias 0.21238f
C3832 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00529f
C3833 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00212f
C3834 XA.XIR[2].XIC[13].icell.Ien VPWR 0.19065f
C3835 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02698f
C3836 XA.XIR[0].XIC[2].icell.Ien Vbias 0.21246f
C3837 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.03424f
C3838 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PUM 0.00131f
C3839 XA.XIR[6].XIC[12].icell.PDM Iout 0.00112f
C3840 XA.XIR[7].XIC[7].icell.PDM VPWR 0.00863f
C3841 XA.XIR[8].XIC[8].icell.PUM Vbias 0.00347f
C3842 a_9827_9569# VPWR 0.0017f
C3843 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.15089f
C3844 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PUM 0.00529f
C3845 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PUM 0.00131f
C3846 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.SM 0.00383f
C3847 XA.XIR[13].XIC[0].icell.SM VPWR 0.00158f
C3848 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00212f
C3849 XA.XIR[6].XIC[14].icell.PDM Vbias 0.04058f
C3850 XThC.XTBN.Y XThC.Tn[13] 0.62331f
C3851 XA.XIR[9].XIC[14].icell.PDM VPWR 0.00873f
C3852 XThR.Tn[4] XA.XIR[4].XIC[10].icell.PDM 0.0033f
C3853 XA.XIR[1].XIC[8].icell.PDM VPWR 0.00863f
C3854 XA.XIR[13].XIC[14].icell.Ien VPWR 0.1907f
C3855 XA.XIR[7].XIC[4].icell.PDM Iout 0.00112f
C3856 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9] 0.0033f
C3857 XThR.Tn[7] XA.XIR[8].XIC[9].icell.SM 0.00121f
C3858 XA.XIR[1].XIC[5].icell.PDM Iout 0.00112f
C3859 XThR.Tn[12] VPWR 7.65279f
C3860 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.SM 0.00188f
C3861 XA.XIR[5].XIC[14].icell.Ien Vbias 0.21238f
C3862 XA.XIR[0].XIC[6].icell.SM VPWR 0.00158f
C3863 XA.XIR[13].XIC[10].icell.Ien Iout 0.06483f
C3864 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00529f
C3865 XThC.XTB4.Y XThC.Tn[8] 0.01306f
C3866 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.03976f
C3867 XThR.Tn[2] XA.XIR[3].XIC[13].icell.Ien 0.00321f
C3868 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.15089f
C3869 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.15089f
C3870 XA.XIR[0].XIC[3].icell.SM Iout 0.00367f
C3871 XThC.Tn[6] XThR.Tn[14] 0.28062f
C3872 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00529f
C3873 XA.XIR[8].XIC[11].icell.PDM Iout 0.00112f
C3874 XThC.Tn[4] XThR.Tn[0] 0.28064f
C3875 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.15089f
C3876 XThC.Tn[10] XThR.Tn[6] 0.28062f
C3877 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.03976f
C3878 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.SM 0.00188f
C3879 XThC.Tn[12] XThR.Tn[8] 0.28062f
C3880 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PUM 0.00131f
C3881 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Iout 0.00347f
C3882 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.01406f
C3883 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.SM 0.00188f
C3884 XA.XIR[10].XIC_15.icell.Ien VPWR 0.25675f
C3885 XA.XIR[6].XIC[14].icell.Ien Iout 0.06483f
C3886 XA.XIR[15].XIC[6].icell.PDM Vbias 0.04058f
C3887 XThC.Tn[11] XThC.Tn[12] 0.22638f
C3888 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04522f
C3889 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C3890 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.SM 0.00383f
C3891 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.03424f
C3892 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.03424f
C3893 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.15089f
C3894 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.SM 0.00188f
C3895 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00212f
C3896 XA.XIR[7].XIC[13].icell.PDM Vbias 0.04058f
C3897 XA.XIR[10].XIC[13].icell.PDM VPWR 0.00863f
C3898 XThR.Tn[10] XA.XIR[11].XIC[6].icell.Ien 0.00321f
C3899 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04522f
C3900 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PUM 0.00131f
C3901 XThC.XTB7.B VPWR 1.33463f
C3902 XThR.Tn[5] XThR.Tn[6] 0.08096f
C3903 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.SM 0.00188f
C3904 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.SM 0.00383f
C3905 XThR.XTB3.Y XThR.Tn[8] 0.00178f
C3906 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PUM 0.00131f
C3907 XA.XIR[3].XIC[0].icell.SM VPWR 0.00158f
C3908 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00529f
C3909 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02698f
C3910 bias[1] bias[0] 0.13857f
C3911 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11595f
C3912 XThC.Tn[13] XThR.Tn[5] 0.28063f
C3913 XA.XIR[9].XIC_15.icell.SM Vbias 0.00701f
C3914 XA.XIR[15].XIC[6].icell.Ien Iout 0.06816f
C3915 XA.XIR[8].XIC[13].icell.Ien Iout 0.06483f
C3916 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C3917 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00212f
C3918 XA.XIR[2].XIC[4].icell.PDM VPWR 0.00863f
C3919 XThR.Tn[11] XA.XIR[11].XIC[14].icell.PDM 0.0033f
C3920 XA.XIR[0].XIC[12].icell.SM Vbias 0.00701f
C3921 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.PUM 0.00112f
C3922 XA.XIR[14].XIC[5].icell.PDM VPWR 0.00863f
C3923 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13] 0.0033f
C3924 XA.XIR[6].XIC[1].icell.PDM Iout 0.00112f
C3925 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[1].icell.SM 0.00383f
C3926 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00212f
C3927 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00212f
C3928 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.SM 0.00188f
C3929 XA.XIR[11].XIC[4].icell.PDM Vbias 0.04058f
C3930 XA.XIR[8].XIC_dummy_right.icell.PUM Vbias 0.00248f
C3931 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.03424f
C3932 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.03424f
C3933 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.03976f
C3934 XThR.XTB2.Y a_n1049_6405# 0.00847f
C3935 XThR.Tn[1] XA.XIR[2].XIC[1].icell.SM 0.00121f
C3936 XThR.XTB7.A a_n1049_7493# 0.0127f
C3937 XA.XIR[13].XIC[4].icell.SM VPWR 0.00158f
C3938 XThC.Tn[11] XThR.Tn[1] 0.28063f
C3939 XA.XIR[10].XIC[3].icell.SM Vbias 0.00701f
C3940 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11336f
C3941 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00212f
C3942 XA.XIR[6].XIC[2].icell.PUM Vbias 0.00347f
C3943 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.SM 0.00188f
C3944 XA.XIR[13].XIC[1].icell.SM Iout 0.00388f
C3945 XThR.Tn[9] XA.XIR[9].XIC[6].icell.PDM 0.0033f
C3946 XA.XIR[12].XIC[5].icell.SM VPWR 0.00158f
C3947 XA.XIR[12].XIC[12].icell.PUM Vbias 0.00347f
C3948 XThR.Tn[6] XA.XIR[6].XIC[14].icell.PDM 0.0033f
C3949 XA.XIR[5].XIC[5].icell.PDM Vbias 0.04058f
C3950 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C3951 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02698f
C3952 XA.XIR[12].XIC[2].icell.SM Iout 0.00388f
C3953 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00212f
C3954 XA.XIR[11].XIC[7].icell.Ien VPWR 0.19065f
C3955 XThC.XTB7.Y a_6243_9615# 0.27822f
C3956 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.SM 0.00188f
C3957 a_n997_1803# VPWR 0.01989f
C3958 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.03976f
C3959 XThR.Tn[5] XA.XIR[6].XIC_15.icell.Ien 0.00116f
C3960 XThR.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.0033f
C3961 XA.XIR[4].XIC[5].icell.Ien Vbias 0.21238f
C3962 XA.XIR[11].XIC[4].icell.Ien Iout 0.06483f
C3963 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.01406f
C3964 XA.XIR[6].XIC[8].icell.PDM VPWR 0.00863f
C3965 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00212f
C3966 XA.XIR[3].XIC[6].icell.SM Vbias 0.00701f
C3967 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C3968 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.01406f
C3969 XA.XIR[6].XIC[5].icell.PDM Iout 0.00112f
C3970 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.03424f
C3971 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.SM 0.00383f
C3972 XA.XIR[15].XIC_15.icell.PDM Vbias 0.04206f
C3973 XThR.Tn[4] XA.XIR[5].XIC[0].icell.Ien 0.00321f
C3974 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.SM 0.00188f
C3975 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04522f
C3976 XA.XIR[5].XIC[8].icell.Ien VPWR 0.19065f
C3977 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.SM 0.00188f
C3978 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.15089f
C3979 XThR.XTB7.B data[6] 0.07481f
C3980 XA.XIR[2].XIC[10].icell.PDM Vbias 0.04058f
C3981 XThC.Tn[1] XThR.Tn[3] 0.28062f
C3982 XThR.Tn[0] XA.XIR[1].XIC[13].icell.Ien 0.00321f
C3983 XThC.XTB2.Y XThC.Tn[8] 0.00167f
C3984 XA.XIR[13].XIC[8].icell.SM VPWR 0.00158f
C3985 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00529f
C3986 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.01406f
C3987 XA.XIR[5].XIC[5].icell.Ien Iout 0.06483f
C3988 XThR.Tn[4] XA.XIR[4].XIC[3].icell.PDM 0.0033f
C3989 XA.XIR[4].XIC[9].icell.SM VPWR 0.00158f
C3990 XA.XIR[13].XIC[0].icell.PDM Vbias 0.04002f
C3991 XThR.Tn[12] XA.XIR[13].XIC[0].icell.SM 0.00127f
C3992 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PUM 0.00529f
C3993 XThR.Tn[7] XA.XIR[8].XIC[2].icell.SM 0.00121f
C3994 XThR.Tn[12] XA.XIR[13].XIC[14].icell.Ien 0.00321f
C3995 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.01406f
C3996 XA.XIR[4].XIC[6].icell.SM Iout 0.00388f
C3997 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.03981f
C3998 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04522f
C3999 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11595f
C4000 XThR.XTB7.B a_n997_3755# 0.01174f
C4001 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.SM 0.00383f
C4002 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02698f
C4003 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.03424f
C4004 XA.XIR[9].XIC[8].icell.PUM Vbias 0.00347f
C4005 XA.XIR[8].XIC[7].icell.PDM VPWR 0.00863f
C4006 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00212f
C4007 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.01406f
C4008 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.03976f
C4009 XThR.Tn[8] XA.XIR[9].XIC[9].icell.Ien 0.00321f
C4010 XThC.XTBN.A XThC.Tn[10] 0.12148f
C4011 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02698f
C4012 XA.XIR[8].XIC[4].icell.PDM Iout 0.00112f
C4013 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01734f
C4014 XA.XIR[14].XIC[1].icell.PDM VPWR 0.00863f
C4015 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.15089f
C4016 XA.XIR[2].XIC[10].icell.Ien Iout 0.06483f
C4017 XThC.Tn[0] XA.XIR[13].XIC_dummy_left.icell.Iout 0.00111f
C4018 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.03976f
C4019 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00529f
C4020 XA.XIR[10].XIC[9].icell.SM VPWR 0.00158f
C4021 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04522f
C4022 XA.XIR[5].XIC[11].icell.SM VPWR 0.00158f
C4023 XThC.Tn[10] XThR.Tn[4] 0.28062f
C4024 XA.XIR[2].XIC[12].icell.Ien Vbias 0.21238f
C4025 XA.XIR[15].XIC_15.icell.PUM Vbias 0.00347f
C4026 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00529f
C4027 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.SM 0.00188f
C4028 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.03424f
C4029 XA.XIR[4].XIC[14].icell.PUM VPWR 0.01036f
C4030 XThC.XTB7.B a_9827_9569# 0.00228f
C4031 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.03976f
C4032 XThR.XTB5.A XThR.XTBN.A 0.06303f
C4033 XA.XIR[9].XIC[11].icell.PDM Iout 0.00112f
C4034 XA.XIR[7].XIC[6].icell.PDM Vbias 0.04058f
C4035 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PUM 0.00131f
C4036 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PUM 0.00529f
C4037 a_7651_9569# Vbias 0.00309f
C4038 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C4039 XA.XIR[1].XIC[7].icell.PDM Vbias 0.04058f
C4040 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04522f
C4041 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.01406f
C4042 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00529f
C4043 XA.XIR[15].XIC[2].icell.Ien VPWR 0.32782f
C4044 XThR.Tn[8] XA.XIR[9].XIC[12].icell.SM 0.00121f
C4045 XA.XIR[3].XIC[14].icell.PDM Iout 0.00112f
C4046 XA.XIR[12].XIC[0].icell.SM Vbias 0.00675f
C4047 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.03424f
C4048 XThR.Tn[4] XThR.Tn[5] 0.08835f
C4049 XA.XIR[12].XIC[14].icell.Ien Vbias 0.21238f
C4050 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PUM 0.00487f
C4051 XThC.XTB6.Y XThC.Tn[6] 0.00689f
C4052 XA.XIR[8].XIC[13].icell.PDM Vbias 0.04058f
C4053 XA.XIR[0].XIC[5].icell.SM Vbias 0.00701f
C4054 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06536f
C4055 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.03976f
C4056 XA.XIR[2].XIC[13].icell.SM Iout 0.00388f
C4057 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04522f
C4058 XA.XIR[7].XIC[9].icell.Ien VPWR 0.19065f
C4059 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.03976f
C4060 XA.XIR[3].XIC_15.icell.PUM Vbias 0.00347f
C4061 XA.XIR[1].XIC[0].icell.PDM Iout 0.00112f
C4062 XThR.XTB7.Y a_n1319_5317# 0.01283f
C4063 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.SM 0.00383f
C4064 XA.XIR[14].XIC[2].icell.PDM Iout 0.00112f
C4065 XA.XIR[7].XIC[6].icell.Ien Iout 0.06483f
C4066 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.03976f
C4067 XA.XIR[1].XIC[10].icell.Ien VPWR 0.19065f
C4068 XA.XIR[9].XIC[3].icell.PDM VPWR 0.00863f
C4069 XA.XIR[10].XIC[11].icell.Ien VPWR 0.19065f
C4070 XThC.Tn[8] Iout 0.83888f
C4071 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02698f
C4072 XA.XIR[4].XIC[0].icell.PDM Iout 0.00112f
C4073 XThR.Tn[12] XA.XIR[13].XIC[4].icell.SM 0.00121f
C4074 XA.XIR[13].XIC_15.icell.Ien VPWR 0.25675f
C4075 XA.XIR[1].XIC[7].icell.Ien Iout 0.06483f
C4076 XThR.Tn[3] XA.XIR[4].XIC[14].icell.Ien 0.00321f
C4077 XA.XIR[9].XIC[13].icell.Ien Iout 0.06483f
C4078 XA.XIR[0].XIC[11].icell.PUM VPWR 0.00971f
C4079 XThR.XTB6.Y XThR.Tn[14] 0.00128f
C4080 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04522f
C4081 XThR.Tn[5] XA.XIR[6].XIC[11].icell.Ien 0.00321f
C4082 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02698f
C4083 XThR.XTB7.B XThR.Tn[11] 0.03888f
C4084 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C4085 XA.XIR[13].XIC[13].icell.PDM VPWR 0.00863f
C4086 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.03424f
C4087 XA.XIR[9].XIC_dummy_right.icell.PUM Vbias 0.00248f
C4088 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PUM 0.00529f
C4089 XA.XIR[15].XIC[11].icell.SM Vbias 0.00701f
C4090 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04522f
C4091 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C4092 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.15089f
C4093 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.SM 0.00188f
C4094 XThR.XTBN.A data[5] 0.0148f
C4095 XThR.Tn[11] XA.XIR[12].XIC[7].icell.Ien 0.00321f
C4096 XThR.Tn[12] a_n997_1803# 0.18719f
C4097 XThC.XTBN.Y XThC.Tn[2] 0.64352f
C4098 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.SM 0.00383f
C4099 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.SM 0.00383f
C4100 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00529f
C4101 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00212f
C4102 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.03976f
C4103 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.SM 0.00188f
C4104 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C4105 XA.XIR[7].XIC[12].icell.SM VPWR 0.00158f
C4106 XA.XIR[8].XIC[1].icell.PUM Vbias 0.00347f
C4107 XThR.Tn[4] XA.XIR[5].XIC[14].icell.Ien 0.00321f
C4108 XA.XIR[15].XIC[8].icell.Ien Vbias 0.17911f
C4109 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02698f
C4110 XThR.Tn[11] XA.XIR[11].XIC[10].icell.PDM 0.0033f
C4111 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04522f
C4112 XThR.XTB3.Y a_n1049_5611# 0.009f
C4113 XA.XIR[5].XIC[1].icell.Ien VPWR 0.19065f
C4114 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02698f
C4115 XA.XIR[1].XIC[13].icell.SM VPWR 0.00158f
C4116 XA.XIR[10].XIC_dummy_right.icell.SM VPWR 0.00123f
C4117 XA.XIR[2].XIC[3].icell.PDM Vbias 0.04058f
C4118 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.SM 0.00383f
C4119 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.SM 0.00383f
C4120 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.01406f
C4121 XA.XIR[14].XIC[4].icell.PDM Vbias 0.04058f
C4122 XA.XIR[4].XIC[2].icell.SM VPWR 0.00158f
C4123 XThC.XTB4.Y XThC.Tn[6] 0.00608f
C4124 a_n1049_6699# XThR.Tn[4] 0.00158f
C4125 data[2] data[3] 0.04128f
C4126 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.03976f
C4127 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.01406f
C4128 XThR.Tn[12] XA.XIR[13].XIC[8].icell.SM 0.00121f
C4129 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.SM 0.00188f
C4130 XA.XIR[0].XIC_15.icell.PUM VPWR 0.0169f
C4131 XThC.XTB3.Y XThC.Tn[10] 0.29462f
C4132 XThC.Tn[1] XThR.Tn[8] 0.28062f
C4133 XA.XIR[13].XIC[3].icell.SM Vbias 0.00701f
C4134 XThR.Tn[1] XA.XIR[1].XIC_15.icell.PDM 0.0033f
C4135 XA.XIR[3].XIC[5].icell.PUM VPWR 0.01036f
C4136 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11217f
C4137 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.03976f
C4138 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04522f
C4139 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C4140 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00529f
C4141 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.03424f
C4142 XThR.Tn[8] XA.XIR[9].XIC[2].icell.Ien 0.00321f
C4143 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00529f
C4144 XThC.XTB3.Y a_4861_9615# 0.0093f
C4145 XA.XIR[12].XIC[4].icell.SM Vbias 0.00701f
C4146 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04522f
C4147 XA.XIR[2].XIC[6].icell.Ien VPWR 0.19065f
C4148 XThC.XTB6.A data[1] 0.37233f
C4149 XThR.XTB7.B XThR.Tn[7] 0.07415f
C4150 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00529f
C4151 XA.XIR[14].XIC[7].icell.Ien VPWR 0.19119f
C4152 XA.XIR[15].XIC[13].icell.Ien Vbias 0.17911f
C4153 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.SM 0.00383f
C4154 XA.XIR[11].XIC[6].icell.Ien Vbias 0.21238f
C4155 XA.XIR[2].XIC[3].icell.Ien Iout 0.06483f
C4156 a_n1049_8581# VPWR 0.71705f
C4157 XA.XIR[14].XIC[4].icell.Ien Iout 0.06483f
C4158 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PUM 0.00131f
C4159 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C4160 XA.XIR[10].XIC[8].icell.PUM Vbias 0.00347f
C4161 XA.XIR[6].XIC[7].icell.PDM Vbias 0.04058f
C4162 XA.XIR[9].XIC[7].icell.PDM VPWR 0.00863f
C4163 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04522f
C4164 a_n1049_7493# XThR.Tn[2] 0.26564f
C4165 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.15089f
C4166 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.03976f
C4167 XThC.Tn[2] XThR.Tn[5] 0.28062f
C4168 XThR.XTBN.Y a_n997_3755# 0.229f
C4169 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02698f
C4170 XA.XIR[5].XIC[7].icell.Ien Vbias 0.21238f
C4171 XA.XIR[9].XIC[4].icell.PDM Iout 0.00112f
C4172 XA.XIR[1].XIC[14].icell.SM Iout 0.00388f
C4173 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.01406f
C4174 XA.XIR[0].XIC[0].icell.PUM VPWR 0.00971f
C4175 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00212f
C4176 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.SM 0.00383f
C4177 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10] 0.0033f
C4178 XThR.Tn[2] XA.XIR[3].XIC[6].icell.Ien 0.00321f
C4179 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.15089f
C4180 XA.XIR[4].XIC[8].icell.SM Vbias 0.00701f
C4181 VPWR bias[0] 1.93694f
C4182 XA.XIR[11].XIC[7].icell.SM Iout 0.00388f
C4183 XA.XIR[0].XIC_15.icell.SM Iout 0.00367f
C4184 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PUM 0.00529f
C4185 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04522f
C4186 XA.XIR[6].XIC[10].icell.Ien VPWR 0.19065f
C4187 XA.XIR[12].XIC[8].icell.SM Vbias 0.00701f
C4188 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.38945f
C4189 XThR.XTB5.Y a_n1319_6405# 0.01188f
C4190 XThC.Tn[0] XThR.Tn[1] 0.28072f
C4191 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02698f
C4192 XA.XIR[3].XIC[11].icell.PUM Vbias 0.00347f
C4193 XA.XIR[10].XIC[10].icell.PUM VPWR 0.01036f
C4194 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PDM 0.00182f
C4195 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00529f
C4196 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04522f
C4197 XA.XIR[6].XIC[7].icell.Ien Iout 0.06483f
C4198 XA.XIR[8].XIC[6].icell.PDM Vbias 0.04058f
C4199 XA.XIR[7].XIC[2].icell.Ien VPWR 0.19065f
C4200 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.03976f
C4201 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.01406f
C4202 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.03596f
C4203 XThC.XTB7.Y a_8963_9569# 0.00474f
C4204 XA.XIR[1].XIC[3].icell.Ien VPWR 0.19065f
C4205 XA.XIR[5].XIC[8].icell.SM Iout 0.00388f
C4206 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04522f
C4207 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.15089f
C4208 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C4209 XA.XIR[13].XIC[9].icell.SM VPWR 0.00158f
C4210 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00212f
C4211 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PUM 0.00131f
C4212 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.03424f
C4213 XA.XIR[0].XIC[4].icell.PUM VPWR 0.00976f
C4214 XA.XIR[9].XIC[13].icell.PDM Vbias 0.04058f
C4215 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.03424f
C4216 XA.XIR[8].XIC[9].icell.Ien VPWR 0.19065f
C4217 XThR.Tn[12] XA.XIR[13].XIC_15.icell.Ien 0.00116f
C4218 XA.XIR[11].XIC[2].icell.PDM VPWR 0.00863f
C4219 XThR.Tn[5] XA.XIR[6].XIC[4].icell.Ien 0.00321f
C4220 XA.XIR[4].XIC[13].icell.PUM Vbias 0.00347f
C4221 XA.XIR[11].XIC[12].icell.SM Iout 0.00388f
C4222 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.PDM 0.00589f
C4223 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.01406f
C4224 XA.XIR[8].XIC[6].icell.Ien Iout 0.06483f
C4225 XA.XIR[6].XIC[13].icell.SM VPWR 0.00158f
C4226 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.03981f
C4227 XA.XIR[10].XIC[3].icell.PDM VPWR 0.00863f
C4228 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02698f
C4229 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Ien 0.00234f
C4230 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PUM 0.00529f
C4231 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00212f
C4232 XA.XIR[15].XIC[1].icell.Ien Vbias 0.17911f
C4233 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00212f
C4234 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PUM 0.00209f
C4235 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00212f
C4236 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.SM 0.00188f
C4237 XThR.XTB6.A VPWR 0.68638f
C4238 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.03424f
C4239 XThR.Tn[10] XA.XIR[11].XIC[2].icell.SM 0.00121f
C4240 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.03511f
C4241 XA.XIR[7].XIC[8].icell.Ien Vbias 0.21238f
C4242 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.03011f
C4243 XThC.Tn[12] VPWR 6.9204f
C4244 XThR.XTBN.Y XThR.Tn[11] 0.52265f
C4245 XThR.Tn[6] XA.XIR[6].XIC[7].icell.PDM 0.0033f
C4246 XA.XIR[5].XIC[14].icell.SM Vbias 0.00701f
C4247 XA.XIR[1].XIC[9].icell.Ien Vbias 0.21238f
C4248 XThR.Tn[10] XA.XIR[10].XIC[6].icell.PDM 0.0033f
C4249 XA.XIR[13].XIC[11].icell.Ien VPWR 0.19065f
C4250 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.SM 0.00188f
C4251 XA.XIR[8].XIC[12].icell.SM VPWR 0.00158f
C4252 XA.XIR[9].XIC[2].icell.PDM Vbias 0.04058f
C4253 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C4254 XA.XIR[15].XIC[12].icell.PUM Vbias 0.00347f
C4255 XThC.XTBN.A a_7651_9569# 0.02087f
C4256 XA.XIR[15].XIC[5].icell.SM VPWR 0.00158f
C4257 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04522f
C4258 XThR.Tn[8] XThR.Tn[9] 0.07233f
C4259 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02698f
C4260 XThR.Tn[7] XA.XIR[7].XIC[12].icell.PDM 0.0033f
C4261 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.0275f
C4262 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01834f
C4263 XThC.XTB7.A Vbias 0.0135f
C4264 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PUM 0.00536f
C4265 XA.XIR[15].XIC[2].icell.SM Iout 0.00388f
C4266 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02698f
C4267 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.01406f
C4268 XA.XIR[0].XIC[10].icell.PUM Vbias 0.00347f
C4269 XThR.Tn[13] XA.XIR[14].XIC[6].icell.Ien 0.00321f
C4270 XThC.Tn[11] XThR.Tn[9] 0.28062f
C4271 XA.XIR[12].XIC_15.icell.Ien Vbias 0.21343f
C4272 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PUM 0.00529f
C4273 XThR.XTB3.Y VPWR 1.07975f
C4274 XA.XIR[6].XIC[14].icell.SM Iout 0.00388f
C4275 XA.XIR[7].XIC[9].icell.SM Iout 0.00388f
C4276 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35783f
C4277 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00212f
C4278 XThR.Tn[0] XA.XIR[1].XIC[6].icell.Ien 0.00321f
C4279 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.03545f
C4280 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C4281 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.SM 0.00188f
C4282 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C4283 XA.XIR[12].XIC[13].icell.PDM Vbias 0.04058f
C4284 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Ien 0.00217f
C4285 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.03424f
C4286 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02698f
C4287 XA.XIR[1].XIC[10].icell.SM Iout 0.00388f
C4288 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.SM 0.00383f
C4289 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PUM 0.00529f
C4290 XA.XIR[12].XIC[3].icell.PUM VPWR 0.01036f
C4291 XA.XIR[7].XIC[11].icell.SM Vbias 0.00701f
C4292 XThR.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.0033f
C4293 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.07827f
C4294 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PUM 0.00529f
C4295 XThR.Tn[1] VPWR 6.75088f
C4296 XA.XIR[13].XIC_dummy_right.icell.SM VPWR 0.00123f
C4297 XA.XIR[5].XIC[1].icell.PUM Vbias 0.00347f
C4298 XA.XIR[1].XIC[12].icell.SM Vbias 0.00701f
C4299 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02698f
C4300 XA.XIR[11].XIC[3].icell.SM VPWR 0.00158f
C4301 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.03982f
C4302 XThR.Tn[9] XA.XIR[10].XIC[11].icell.SM 0.00121f
C4303 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.01406f
C4304 XA.XIR[4].XIC[1].icell.SM Vbias 0.00701f
C4305 XThR.XTBN.Y XThR.Tn[7] 0.89982f
C4306 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.15089f
C4307 XA.XIR[10].XIC[7].icell.PDM VPWR 0.00863f
C4308 XA.XIR[6].XIC[3].icell.Ien VPWR 0.19065f
C4309 XThR.Tn[9] XA.XIR[10].XIC[8].icell.Ien 0.00321f
C4310 XA.XIR[3].XIC[4].icell.PUM Vbias 0.00347f
C4311 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02698f
C4312 XThR.XTB4.Y data[6] 0.0086f
C4313 XA.XIR[6].XIC[0].icell.Ien Iout 0.06474f
C4314 XA.XIR[10].XIC[4].icell.PDM Iout 0.00112f
C4315 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.SM 0.00188f
C4316 XA.XIR[5].XIC[4].icell.SM VPWR 0.00158f
C4317 XThC.Tn[6] Iout 0.83989f
C4318 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00212f
C4319 XThC.Tn[9] XThR.Tn[11] 0.28062f
C4320 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PUM 0.00529f
C4321 XA.XIR[2].XIC[5].icell.Ien Vbias 0.21238f
C4322 XA.XIR[5].XIC[1].icell.SM Iout 0.00388f
C4323 XA.XIR[14].XIC[6].icell.Ien Vbias 0.21238f
C4324 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Iout 0.00395f
C4325 XA.XIR[4].XIC[7].icell.PUM VPWR 0.01036f
C4326 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.03976f
C4327 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00529f
C4328 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.01406f
C4329 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04522f
C4330 XA.XIR[13].XIC[8].icell.PUM Vbias 0.00347f
C4331 XThR.XTB4.Y a_n997_3755# 0.00497f
C4332 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00212f
C4333 XThR.Tn[12] XA.XIR[13].XIC[9].icell.SM 0.00121f
C4334 XThR.Tn[6] XA.XIR[7].XIC[8].icell.Ien 0.00321f
C4335 XThR.Tn[10] XA.XIR[10].XIC_15.icell.PDM 0.0033f
C4336 XA.XIR[3].XIC[10].icell.PDM VPWR 0.00863f
C4337 XA.XIR[9].XIC[6].icell.PDM Vbias 0.04058f
C4338 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04522f
C4339 XA.XIR[8].XIC[2].icell.Ien VPWR 0.19065f
C4340 XThR.XTB5.A XThR.XTB6.Y 0.00193f
C4341 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PUM 0.00529f
C4342 XThR.Tn[8] XA.XIR[9].XIC[5].icell.SM 0.00121f
C4343 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01799f
C4344 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04522f
C4345 XA.XIR[2].XIC[9].icell.SM VPWR 0.00158f
C4346 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C4347 XThC.XTBN.Y a_2979_9615# 0.0607f
C4348 XA.XIR[3].XIC[7].icell.PDM Iout 0.00112f
C4349 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PUM 0.00529f
C4350 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02698f
C4351 XA.XIR[10].XIC[11].icell.PDM VPWR 0.00863f
C4352 a_5949_9615# Vbias 0.00582f
C4353 XThR.Tn[9] XA.XIR[10].XIC[13].icell.Ien 0.00321f
C4354 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04522f
C4355 XA.XIR[2].XIC[6].icell.SM Iout 0.00388f
C4356 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00529f
C4357 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.SM 0.00188f
C4358 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00212f
C4359 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.03424f
C4360 XA.XIR[14].XIC[7].icell.SM Iout 0.00388f
C4361 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.15089f
C4362 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.03976f
C4363 XA.XIR[15].XIC[14].icell.Ien Vbias 0.17911f
C4364 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.SM 0.00383f
C4365 XA.XIR[9].XIC[9].icell.Ien VPWR 0.19065f
C4366 XA.XIR[6].XIC[9].icell.Ien Vbias 0.21238f
C4367 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00212f
C4368 XA.XIR[13].XIC[10].icell.PUM VPWR 0.01036f
C4369 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.01406f
C4370 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00529f
C4371 a_9827_9569# XThC.Tn[12] 0.19481f
C4372 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.01406f
C4373 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PUM 0.00529f
C4374 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.SM 0.00383f
C4375 XThC.XTB3.Y a_7651_9569# 0.00604f
C4376 XThR.Tn[3] XA.XIR[4].XIC[7].icell.Ien 0.00321f
C4377 XThC.Tn[0] XThC.Tn[1] 1.15894f
C4378 XA.XIR[5].XIC[10].icell.SM Vbias 0.00701f
C4379 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.03976f
C4380 XA.XIR[9].XIC[6].icell.Ien Iout 0.06483f
C4381 XA.XIR[7].XIC[1].icell.Ien Vbias 0.21238f
C4382 XThC.Tn[9] XThR.Tn[7] 0.28062f
C4383 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PUM 0.00529f
C4384 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02698f
C4385 XThC.XTB5.A Vbias 0.005f
C4386 XThC.Tn[4] XThC.Tn[6] 0.00202f
C4387 XA.XIR[3].XIC[12].icell.Ien VPWR 0.19065f
C4388 XThR.Tn[2] XA.XIR[3].XIC[9].icell.SM 0.00121f
C4389 XThR.Tn[6] XA.XIR[7].XIC[11].icell.SM 0.00121f
C4390 XThC.Tn[14] XThR.Tn[2] 0.28068f
C4391 XA.XIR[1].XIC[2].icell.Ien Vbias 0.21238f
C4392 XThC.Tn[12] XThR.Tn[12] 0.28062f
C4393 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.01406f
C4394 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02698f
C4395 XThR.Tn[12] XA.XIR[13].XIC[11].icell.Ien 0.00321f
C4396 XA.XIR[2].XIC[14].icell.PUM VPWR 0.01036f
C4397 XThR.Tn[7] XA.XIR[7].XIC[5].icell.PDM 0.0033f
C4398 XThR.Tn[2] XA.XIR[2].XIC[13].icell.PDM 0.0033f
C4399 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.SM 0.00188f
C4400 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04522f
C4401 XA.XIR[0].XIC[3].icell.PUM Vbias 0.00347f
C4402 XA.XIR[14].XIC[0].icell.Ien VPWR 0.19119f
C4403 XA.XIR[8].XIC[8].icell.Ien Vbias 0.21238f
C4404 XA.XIR[6].XIC[10].icell.SM Iout 0.00388f
C4405 XA.XIR[12].XIC[9].icell.SM Vbias 0.00701f
C4406 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.SM 0.00188f
C4407 XA.XIR[14].XIC[12].icell.SM Iout 0.00388f
C4408 XA.XIR[7].XIC[5].icell.SM VPWR 0.00158f
C4409 XThR.Tn[4] XA.XIR[5].XIC[7].icell.Ien 0.00321f
C4410 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PUM 0.00529f
C4411 a_10915_9569# VPWR 0.00307f
C4412 XA.XIR[13].XIC[3].icell.PDM VPWR 0.00863f
C4413 XThR.Tn[1] XA.XIR[2].XIC[13].icell.Ien 0.00321f
C4414 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PUM 0.00529f
C4415 XA.XIR[7].XIC[2].icell.SM Iout 0.00388f
C4416 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01674f
C4417 XA.XIR[1].XIC[6].icell.SM VPWR 0.00158f
C4418 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04522f
C4419 XA.XIR[10].XIC[2].icell.PDM Vbias 0.04058f
C4420 XA.XIR[6].XIC[12].icell.SM Vbias 0.00701f
C4421 XA.XIR[9].XIC[12].icell.SM VPWR 0.00158f
C4422 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00529f
C4423 XThR.Tn[8] XThR.Tn[10] 0.00255f
C4424 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02698f
C4425 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.03976f
C4426 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00212f
C4427 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.SM 0.00188f
C4428 XA.XIR[1].XIC[3].icell.SM Iout 0.00388f
C4429 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04522f
C4430 XThC.XTB5.A a_7331_10587# 0.01243f
C4431 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01096f
C4432 XThR.Tn[1] XA.XIR[1].XIC[8].icell.PDM 0.0033f
C4433 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C4434 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04522f
C4435 XThC.Tn[11] XThR.Tn[10] 0.28062f
C4436 XThR.Tn[5] XA.XIR[6].XIC[7].icell.SM 0.00121f
C4437 XThC.XTB7.B XThC.Tn[12] 0.00772f
C4438 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PUM 0.00131f
C4439 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04522f
C4440 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PUM 0.00529f
C4441 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C4442 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.01406f
C4443 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00529f
C4444 XA.XIR[8].XIC[9].icell.SM Iout 0.00388f
C4445 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PUM 0.00529f
C4446 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[11].icell.Ien 0.00212f
C4447 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.SM 0.00188f
C4448 XA.XIR[11].XIC[13].icell.SM Iout 0.00388f
C4449 XThR.Tn[11] XA.XIR[12].XIC[3].icell.SM 0.00121f
C4450 XThR.XTB5.Y XThR.Tn[13] 0.00145f
C4451 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PUM 0.00529f
C4452 XA.XIR[8].XIC[11].icell.SM Vbias 0.00701f
C4453 XA.XIR[15].XIC[4].icell.SM Vbias 0.00701f
C4454 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00212f
C4455 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04522f
C4456 XThR.Tn[8] XA.XIR[8].XIC_15.icell.PDM 0.0033f
C4457 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C4458 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.15089f
C4459 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.SM 0.00383f
C4460 XA.XIR[12].XIC[11].icell.Ien Vbias 0.21238f
C4461 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.PUM 0.00112f
C4462 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.01406f
C4463 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PUM 0.00131f
C4464 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.15089f
C4465 XThR.Tn[7] XA.XIR[8].XIC[14].icell.Ien 0.00321f
C4466 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.15089f
C4467 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.SM 0.00383f
C4468 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35783f
C4469 XThR.Tn[3] XA.XIR[4].XIC[14].icell.SM 0.00121f
C4470 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C4471 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PUM 0.00529f
C4472 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.15089f
C4473 XA.XIR[3].XIC[3].icell.PDM VPWR 0.00863f
C4474 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PUM 0.00131f
C4475 XThR.Tn[14] XA.XIR[14].XIC[10].icell.PDM 0.0033f
C4476 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PUM 0.00131f
C4477 XThR.Tn[6] XA.XIR[7].XIC[1].icell.Ien 0.00321f
C4478 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00529f
C4479 XA.XIR[0].XIC_15.icell.PDM Vbias 0.04213f
C4480 XA.XIR[2].XIC[2].icell.SM VPWR 0.00158f
C4481 XThR.Tn[5] XA.XIR[5].XIC_15.icell.PDM 0.0033f
C4482 XA.XIR[14].XIC[3].icell.SM VPWR 0.00158f
C4483 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C4484 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PUM 0.00529f
C4485 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C4486 XA.XIR[11].XIC[2].icell.SM Vbias 0.00701f
C4487 XThC.XTB7.A XThC.XTBN.A 0.197f
C4488 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04522f
C4489 XThC.Tn[1] VPWR 5.98031f
C4490 XA.XIR[15].XIC[8].icell.SM Vbias 0.00701f
C4491 XThR.XTB7.A data[6] 0.00197f
C4492 XThC.XTB1.Y a_7651_9569# 0.06353f
C4493 XThR.Tn[4] XA.XIR[5].XIC[14].icell.SM 0.00121f
C4494 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.15089f
C4495 XA.XIR[13].XIC[7].icell.PDM VPWR 0.00863f
C4496 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.SM 0.00188f
C4497 XThR.Tn[0] XA.XIR[1].XIC[9].icell.SM 0.00121f
C4498 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04522f
C4499 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.03976f
C4500 XA.XIR[10].XIC[6].icell.PDM Vbias 0.04058f
C4501 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01776f
C4502 XA.XIR[9].XIC[2].icell.Ien VPWR 0.19065f
C4503 XA.XIR[6].XIC[2].icell.Ien Vbias 0.21238f
C4504 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Ien 0.00591f
C4505 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.01406f
C4506 XA.XIR[12].XIC[8].icell.PDM VPWR 0.00863f
C4507 XA.XIR[13].XIC[4].icell.PDM Iout 0.00112f
C4508 XThR.Tn[3] XA.XIR[4].XIC[0].icell.Ien 0.00321f
C4509 XThR.Tn[0] XA.XIR[0].XIC[12].icell.PDM 0.0033f
C4510 XThC.Tn[9] XThR.Tn[14] 0.28062f
C4511 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.15089f
C4512 XA.XIR[5].XIC[3].icell.SM Vbias 0.00701f
C4513 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PUM 0.00131f
C4514 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.01406f
C4515 XA.XIR[11].XIC[8].icell.PUM VPWR 0.01036f
C4516 XThC.Tn[0] XThR.Tn[9] 0.28064f
C4517 XA.XIR[12].XIC[5].icell.PDM Iout 0.00112f
C4518 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04522f
C4519 XThR.Tn[3] Vbias 3.71826f
C4520 XThR.Tn[2] XA.XIR[3].XIC[2].icell.SM 0.00121f
C4521 XA.XIR[4].XIC[6].icell.PUM Vbias 0.00347f
C4522 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PUM 0.00134f
C4523 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00212f
C4524 XA.XIR[6].XIC[6].icell.SM VPWR 0.00158f
C4525 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.SM 0.00188f
C4526 XThR.Tn[2] XA.XIR[2].XIC[6].icell.PDM 0.0033f
C4527 XA.XIR[3].XIC[9].icell.PDM Vbias 0.04058f
C4528 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00212f
C4529 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.SM 0.00188f
C4530 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PUM 0.00131f
C4531 XA.XIR[8].XIC[1].icell.Ien Vbias 0.21238f
C4532 XA.XIR[6].XIC[3].icell.SM Iout 0.00388f
C4533 XA.XIR[10].XIC[6].icell.Ien Iout 0.06483f
C4534 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.SM 0.00383f
C4535 XA.XIR[5].XIC[9].icell.PUM VPWR 0.01036f
C4536 XThR.XTB5.A XThR.XTB7.B 0.30355f
C4537 XA.XIR[2].XIC[8].icell.SM Vbias 0.00701f
C4538 XA.XIR[13].XIC[11].icell.PDM VPWR 0.00863f
C4539 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13] 0.0033f
C4540 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PUM 0.00131f
C4541 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.SM 0.00188f
C4542 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00212f
C4543 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00212f
C4544 XA.XIR[4].XIC[12].icell.PDM VPWR 0.00863f
C4545 a_6243_9615# XThC.Tn[6] 0.26142f
C4546 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.01406f
C4547 XThR.Tn[11] XA.XIR[11].XIC[12].icell.PDM 0.0033f
C4548 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00529f
C4549 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.03976f
C4550 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.03424f
C4551 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.03976f
C4552 XA.XIR[4].XIC[9].icell.PDM Iout 0.00112f
C4553 XA.XIR[1].XIC_15.icell.SM Iout 0.0047f
C4554 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.01406f
C4555 XA.XIR[0].XIC[2].icell.PDM VPWR 0.00806f
C4556 XA.XIR[11].XIC[14].icell.PDM Iout 0.00112f
C4557 XA.XIR[9].XIC[8].icell.Ien Vbias 0.21238f
C4558 XA.XIR[8].XIC[5].icell.SM VPWR 0.00158f
C4559 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PUM 0.00131f
C4560 XThR.Tn[5] XA.XIR[6].XIC[0].icell.SM 0.00121f
C4561 XA.XIR[3].XIC[9].icell.Ien Iout 0.06483f
C4562 a_n1319_5317# VPWR 0.00672f
C4563 XA.XIR[8].XIC[2].icell.SM Iout 0.00388f
C4564 a_n1049_7787# VPWR 0.72179f
C4565 XA.XIR[14].XIC_dummy_left.icell.SM VPWR 0.00269f
C4566 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02698f
C4567 XA.XIR[12].XIC[10].icell.PUM Vbias 0.00347f
C4568 XThR.Tn[9] XA.XIR[10].XIC[0].icell.SM 0.00127f
C4569 XThR.Tn[9] XA.XIR[10].XIC[14].icell.Ien 0.00321f
C4570 XThC.Tn[7] XThR.Tn[11] 0.28062f
C4571 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.SM 0.00383f
C4572 XA.XIR[5].XIC[14].icell.PDM VPWR 0.00873f
C4573 XA.XIR[2].XIC[13].icell.PUM Vbias 0.00347f
C4574 XA.XIR[10].XIC_15.icell.PDM Vbias 0.04206f
C4575 XA.XIR[15].XIC_15.icell.Ien Vbias 0.17893f
C4576 XA.XIR[4].XIC[14].icell.Ien VPWR 0.1907f
C4577 XA.XIR[9].XIC[9].icell.SM Iout 0.00388f
C4578 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.01406f
C4579 XThR.Tn[3] XA.XIR[4].XIC[10].icell.SM 0.00121f
C4580 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00212f
C4581 XA.XIR[7].XIC[4].icell.SM Vbias 0.00701f
C4582 XThR.Tn[14] XA.XIR[15].XIC[7].icell.Ien 0.00321f
C4583 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04522f
C4584 XThR.Tn[0] XA.XIR[0].XIC[1].icell.PDM 0.0033f
C4585 a_8739_9569# Vbias 0.0026f
C4586 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.15089f
C4587 XThR.XTB5.Y XThR.Tn[6] 0.00349f
C4588 XA.XIR[15].XIC[13].icell.PDM Vbias 0.04058f
C4589 XThR.XTB7.B data[5] 0.00593f
C4590 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.SM 0.00383f
C4591 XA.XIR[1].XIC[5].icell.SM Vbias 0.00701f
C4592 XA.XIR[13].XIC[2].icell.PDM Vbias 0.04058f
C4593 XA.XIR[9].XIC[11].icell.SM Vbias 0.00701f
C4594 XA.XIR[15].XIC[3].icell.PUM VPWR 0.01036f
C4595 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02698f
C4596 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00529f
C4597 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00212f
C4598 XThC.XTB5.A XThC.XTBN.A 0.06305f
C4599 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PDM 0.00182f
C4600 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C4601 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02698f
C4602 XA.XIR[3].XIC[12].icell.SM Iout 0.00388f
C4603 XA.XIR[12].XIC[3].icell.PDM Vbias 0.04058f
C4604 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.15089f
C4605 XThC.Tn[11] XThR.Tn[13] 0.28062f
C4606 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PUM 0.00529f
C4607 XA.XIR[0].XIC[8].icell.PDM Vbias 0.04065f
C4608 XThC.XTB7.A XThC.Tn[2] 0.12602f
C4609 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01776f
C4610 XThR.Tn[13] XA.XIR[14].XIC[2].icell.SM 0.00121f
C4611 XThR.Tn[4] XA.XIR[5].XIC[10].icell.SM 0.00121f
C4612 XA.XIR[7].XIC[10].icell.PUM VPWR 0.01036f
C4613 XA.XIR[3].XIC_15.icell.Ien Vbias 0.21343f
C4614 XA.XIR[1].XIC[1].icell.PDM VPWR 0.00863f
C4615 XThC.Tn[13] XThR.Tn[3] 0.28063f
C4616 XThC.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00111f
C4617 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Iout 0.00347f
C4618 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C4619 XA.XIR[14].XIC[13].icell.SM Iout 0.00388f
C4620 XThR.Tn[13] XA.XIR[13].XIC[6].icell.PDM 0.0033f
C4621 XA.XIR[1].XIC[11].icell.PUM VPWR 0.01036f
C4622 XThR.Tn[0] XA.XIR[1].XIC[2].icell.SM 0.00121f
C4623 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C4624 XThR.Tn[9] VPWR 7.62673f
C4625 XThC.Tn[3] XThR.Tn[2] 0.28062f
C4626 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04522f
C4627 XThC.Tn[1] XThR.Tn[12] 0.28062f
C4628 XA.XIR[4].XIC[1].icell.PDM VPWR 0.00863f
C4629 XThC.Tn[7] XThR.Tn[7] 0.28062f
C4630 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.03976f
C4631 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.03976f
C4632 XA.XIR[10].XIC_15.icell.PUM Vbias 0.00347f
C4633 XA.XIR[0].XIC[11].icell.Ien VPWR 0.19108f
C4634 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.SM 0.00188f
C4635 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.01406f
C4636 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.15089f
C4637 XThR.Tn[0] XA.XIR[0].XIC[5].icell.PDM 0.0033f
C4638 XA.XIR[4].XIC_15.icell.Ien Iout 0.06485f
C4639 XA.XIR[5].XIC_15.icell.SM Vbias 0.00701f
C4640 XThR.Tn[12] XA.XIR[12].XIC[8].icell.PDM 0.0033f
C4641 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.01406f
C4642 XA.XIR[0].XIC[8].icell.Ien Iout 0.06455f
C4643 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00529f
C4644 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[12].icell.SM 0.00383f
C4645 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00212f
C4646 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PUM 0.00131f
C4647 XA.XIR[10].XIC[2].icell.Ien VPWR 0.19065f
C4648 XThR.XTB7.A XThR.Tn[7] 0.00182f
C4649 XThR.Tn[9] XA.XIR[10].XIC[4].icell.SM 0.00121f
C4650 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02698f
C4651 XA.XIR[11].XIC[14].icell.SM Iout 0.00388f
C4652 XA.XIR[3].XIC[2].icell.PDM Vbias 0.04058f
C4653 XThR.Tn[8] Vbias 3.71582f
C4654 XA.XIR[7].XIC_15.icell.PDM VPWR 0.06959f
C4655 XA.XIR[12].XIC_dummy_right.icell.Ien Vbias 0.00287f
C4656 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.03976f
C4657 XA.XIR[5].XIC[2].icell.PUM VPWR 0.01036f
C4658 XA.XIR[6].XIC_15.icell.SM Iout 0.0047f
C4659 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08017f
C4660 XThC.Tn[11] Vbias 2.38011f
C4661 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.SM 0.00383f
C4662 XThC.Tn[0] XThR.Tn[10] 0.2806f
C4663 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06536f
C4664 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00213f
C4665 XA.XIR[2].XIC[1].icell.SM Vbias 0.00701f
C4666 XA.XIR[1].XIC[2].icell.PDM Iout 0.00112f
C4667 XA.XIR[4].XIC[5].icell.PDM VPWR 0.00863f
C4668 XThC.XTB7.B XThC.Tn[1] 0.0014f
C4669 XA.XIR[14].XIC[2].icell.SM Vbias 0.00701f
C4670 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.03976f
C4671 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00529f
C4672 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00212f
C4673 XA.XIR[0].XIC_15.icell.Ien VPWR 0.25652f
C4674 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.SM 0.00188f
C4675 XA.XIR[4].XIC[2].icell.PDM Iout 0.00112f
C4676 XA.XIR[13].XIC[6].icell.PDM Vbias 0.04058f
C4677 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.SM 0.00383f
C4678 XA.XIR[3].XIC[5].icell.Ien VPWR 0.19065f
C4679 XThR.Tn[6] XA.XIR[7].XIC[4].icell.SM 0.00121f
C4680 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C4681 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.01406f
C4682 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PUM 0.00529f
C4683 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04522f
C4684 XThR.XTB6.Y a_n1319_5611# 0.01283f
C4685 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04522f
C4686 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.SM 0.00188f
C4687 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00212f
C4688 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PUM 0.00131f
C4689 XA.XIR[12].XIC[7].icell.PDM Vbias 0.04058f
C4690 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C4691 XThC.XTB3.Y a_5949_9615# 0.009f
C4692 XA.XIR[3].XIC[2].icell.Ien Iout 0.06483f
C4693 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.0353f
C4694 XA.XIR[2].XIC[7].icell.PUM VPWR 0.01036f
C4695 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC[14].icell.SM 0.00383f
C4696 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00529f
C4697 XA.XIR[14].XIC[8].icell.PUM VPWR 0.01036f
C4698 XA.XIR[10].XIC[11].icell.SM Vbias 0.00701f
C4699 XThR.XTB5.A XThR.XTBN.Y 0.00282f
C4700 XThR.Tn[9] XA.XIR[10].XIC[8].icell.SM 0.00121f
C4701 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02698f
C4702 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[4].icell.Ien 0.00212f
C4703 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.SM 0.00188f
C4704 XA.XIR[11].XIC[7].icell.PUM Vbias 0.00347f
C4705 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04522f
C4706 a_n1319_6405# VPWR 0.00676f
C4707 XThR.Tn[1] XA.XIR[2].XIC[6].icell.Ien 0.00321f
C4708 XThR.Tn[13] XA.XIR[13].XIC_15.icell.PDM 0.0033f
C4709 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PUM 0.00529f
C4710 XA.XIR[10].XIC[8].icell.Ien Vbias 0.21238f
C4711 XA.XIR[15].XIC[9].icell.SM Vbias 0.00701f
C4712 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.SM 0.00188f
C4713 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.SM 0.00383f
C4714 XA.XIR[9].XIC[5].icell.SM VPWR 0.00158f
C4715 XA.XIR[6].XIC[5].icell.SM Vbias 0.00701f
C4716 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.15089f
C4717 XA.XIR[13].XIC[6].icell.Ien Iout 0.06483f
C4718 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C4719 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C4720 XThR.Tn[3] XA.XIR[4].XIC[3].icell.SM 0.00121f
C4721 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.15089f
C4722 XA.XIR[9].XIC[2].icell.SM Iout 0.00388f
C4723 XThR.Tn[14] XA.XIR[15].XIC[0].icell.Ien 0.00358f
C4724 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Ien 0.00529f
C4725 XA.XIR[5].XIC[8].icell.PUM Vbias 0.00347f
C4726 XA.XIR[11].XIC[12].icell.Ien Iout 0.06483f
C4727 XA.XIR[12].XIC[7].icell.Ien Iout 0.06483f
C4728 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.15089f
C4729 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PUM 0.00131f
C4730 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02698f
C4731 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.15089f
C4732 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01872f
C4733 XA.XIR[4].XIC[11].icell.PDM Vbias 0.04058f
C4734 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.03432f
C4735 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.SM 0.00383f
C4736 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.1192f
C4737 XA.XIR[11].XIC[10].icell.PDM Iout 0.00112f
C4738 XThC.XTBN.Y XThC.Tn[14] 0.50214f
C4739 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.SM 0.00188f
C4740 XA.XIR[12].XIC[11].icell.PDM Vbias 0.04058f
C4741 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C4742 XA.XIR[6].XIC[11].icell.PUM VPWR 0.01036f
C4743 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.SM 0.00383f
C4744 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.15089f
C4745 XA.XIR[14].XIC[14].icell.PDM Iout 0.00112f
C4746 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC[0].icell.Ien 0.00212f
C4747 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.15089f
C4748 XA.XIR[3].XIC[11].icell.Ien Vbias 0.21238f
C4749 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.SM 0.00383f
C4750 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00529f
C4751 XThR.XTB5.Y a_n997_2667# 0.00427f
C4752 XThR.Tn[4] XA.XIR[5].XIC[3].icell.SM 0.00121f
C4753 XA.XIR[8].XIC[4].icell.SM Vbias 0.00701f
C4754 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.SM 0.00383f
C4755 XA.XIR[7].XIC[3].icell.PUM VPWR 0.01036f
C4756 Vbias data[0] 0.0027f
C4757 XThR.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.0033f
C4758 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C4759 XA.XIR[10].XIC[13].icell.Ien Vbias 0.21238f
C4760 XThR.Tn[3] XThR.Tn[4] 0.08415f
C4761 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.01406f
C4762 XThC.XTB7.Y a_10051_9569# 0.013f
C4763 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PUM 0.00529f
C4764 XA.XIR[5].XIC[11].icell.PDM Iout 0.00112f
C4765 XA.XIR[1].XIC[4].icell.PUM VPWR 0.01036f
C4766 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.SM 0.00383f
C4767 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00529f
C4768 XThC.Tn[5] XThR.Tn[0] 0.28068f
C4769 XThR.Tn[9] XA.XIR[9].XIC[14].icell.PDM 0.0033f
C4770 XThC.Tn[7] XThR.Tn[14] 0.28062f
C4771 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02698f
C4772 XThR.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.00321f
C4773 XThC.Tn[11] XThR.Tn[6] 0.28062f
C4774 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.002f
C4775 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.01406f
C4776 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04522f
C4777 XA.XIR[15].XIC[11].icell.Ien Vbias 0.17911f
C4778 XA.XIR[4].XIC[11].icell.Ien Iout 0.06483f
C4779 XThC.Tn[13] XThR.Tn[8] 0.28063f
C4780 bias[1] Vbias 0.04991f
C4781 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PUM 0.00529f
C4782 XA.XIR[13].XIC_15.icell.PDM Vbias 0.04206f
C4783 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00212f
C4784 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.SM 0.00188f
C4785 XThR.XTB7.Y a_n997_2667# 0.00474f
C4786 XA.XIR[0].XIC[4].icell.Ien VPWR 0.19019f
C4787 XA.XIR[8].XIC[10].icell.PUM VPWR 0.01036f
C4788 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.15089f
C4789 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PUM 0.00131f
C4790 XA.XIR[2].XIC[0].icell.PDM VPWR 0.00863f
C4791 XThC.Tn[11] XThC.Tn[13] 0.00226f
C4792 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02698f
C4793 XA.XIR[4].XIC[13].icell.Ien Vbias 0.21238f
C4794 XA.XIR[0].XIC[1].icell.Ien Iout 0.06455f
C4795 XA.XIR[15].XIC[1].icell.PDM Iout 0.00112f
C4796 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02698f
C4797 XThR.Tn[5] XA.XIR[5].XIC[8].icell.PDM 0.0033f
C4798 XThR.Tn[10] VPWR 7.60864f
C4799 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08017f
C4800 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.01406f
C4801 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04522f
C4802 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39096f
C4803 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.01406f
C4804 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.03424f
C4805 XA.XIR[15].XIC[2].icell.PUM Vbias 0.00347f
C4806 a_7331_10587# data[0] 0.00451f
C4807 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PUM 0.00529f
C4808 XThR.Tn[9] XA.XIR[10].XIC_15.icell.Ien 0.00116f
C4809 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.01406f
C4810 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C4811 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.38953f
C4812 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C4813 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.01406f
C4814 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04522f
C4815 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.002f
C4816 XA.XIR[5].XIC[13].icell.Ien Iout 0.06483f
C4817 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.03976f
C4818 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Ien 0.00217f
C4819 XThC.Tn[14] XThR.Tn[5] 0.28068f
C4820 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PUM 0.00529f
C4821 XA.XIR[7].XIC[9].icell.PUM Vbias 0.00347f
C4822 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.03981f
C4823 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02698f
C4824 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.03982f
C4825 XA.XIR[1].XIC[10].icell.PUM Vbias 0.00347f
C4826 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00529f
C4827 XA.XIR[5].XIC_dummy_right.icell.PUM Vbias 0.00248f
C4828 XThR.XTB6.A XThR.Tn[1] 0.00411f
C4829 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01193f
C4830 XA.XIR[9].XIC[0].icell.SM Vbias 0.00675f
C4831 XA.XIR[8].XIC_15.icell.PDM VPWR 0.06959f
C4832 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00212f
C4833 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.15089f
C4834 XThC.XTBN.A a_8739_9569# 0.01719f
C4835 XThC.Tn[12] XThR.Tn[1] 0.28063f
C4836 XA.XIR[13].XIC_15.icell.PUM Vbias 0.00347f
C4837 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.01406f
C4838 XA.XIR[15].XIC[5].icell.PDM Iout 0.00112f
C4839 XA.XIR[0].XIC[10].icell.Ien Vbias 0.21246f
C4840 XA.XIR[6].XIC[0].icell.PUM VPWR 0.01036f
C4841 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.03429f
C4842 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PUM 0.00131f
C4843 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PDM 0.00552f
C4844 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.SM 0.00188f
C4845 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00212f
C4846 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.15089f
C4847 XThR.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.00342f
C4848 XA.XIR[7].XIC[12].icell.PDM Iout 0.00112f
C4849 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C4850 XA.XIR[11].XIC[10].icell.SM Iout 0.00388f
C4851 XA.XIR[13].XIC[2].icell.Ien VPWR 0.19065f
C4852 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00529f
C4853 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PUM 0.00131f
C4854 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.01406f
C4855 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02698f
C4856 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02698f
C4857 XA.XIR[14].XIC[14].icell.SM Iout 0.00388f
C4858 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01785f
C4859 XA.XIR[1].XIC[13].icell.PDM Iout 0.00112f
C4860 XA.XIR[7].XIC[14].icell.PDM Vbias 0.04058f
C4861 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.03424f
C4862 XA.XIR[12].XIC[3].icell.Ien VPWR 0.19065f
C4863 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00529f
C4864 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.15089f
C4865 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.03424f
C4866 XThC.Tn[0] XThR.Tn[13] 0.28069f
C4867 XThR.Tn[7] XA.XIR[8].XIC[14].icell.SM 0.00121f
C4868 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00529f
C4869 XA.XIR[1].XIC_15.icell.PDM Vbias 0.04206f
C4870 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00212f
C4871 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.03424f
C4872 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04522f
C4873 XA.XIR[11].XIC[6].icell.PDM VPWR 0.00863f
C4874 XA.XIR[0].XIC[11].icell.SM Iout 0.00367f
C4875 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00529f
C4876 a_7875_9569# XThC.Tn[9] 0.19329f
C4877 XThC.XTB6.A XThC.Tn[5] 0.00363f
C4878 XThR.Tn[5] XA.XIR[5].XIC[0].icell.PDM 0.00335f
C4879 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00212f
C4880 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.15089f
C4881 XThC.Tn[2] XThR.Tn[3] 0.28062f
C4882 XA.XIR[4].XIC[4].icell.PDM Vbias 0.04058f
C4883 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Iout 0.00347f
C4884 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C4885 XThC.XTB2.Y XThC.Tn[9] 0.292f
C4886 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00529f
C4887 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.01406f
C4888 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00529f
C4889 XA.XIR[10].XIC[5].icell.SM VPWR 0.00158f
C4890 XA.XIR[10].XIC[12].icell.PUM Vbias 0.00347f
C4891 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.01406f
C4892 XA.XIR[6].XIC[4].icell.PUM VPWR 0.01036f
C4893 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.15089f
C4894 XA.XIR[3].XIC[4].icell.Ien Vbias 0.21238f
C4895 XA.XIR[10].XIC[2].icell.SM Iout 0.00388f
C4896 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.03424f
C4897 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C4898 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.15089f
C4899 XA.XIR[5].XIC[7].icell.PDM VPWR 0.00863f
C4900 XA.XIR[15].XIC[10].icell.PUM Vbias 0.00347f
C4901 XA.XIR[2].XIC[6].icell.PUM Vbias 0.00347f
C4902 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PUM 0.00529f
C4903 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.03424f
C4904 XA.XIR[7].XIC[14].icell.Ien Iout 0.06483f
C4905 XA.XIR[13].XIC[11].icell.SM Vbias 0.00701f
C4906 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PUM 0.00134f
C4907 XA.XIR[14].XIC[7].icell.PUM Vbias 0.00347f
C4908 XA.XIR[7].XIC[0].icell.PDM VPWR 0.00863f
C4909 XA.XIR[5].XIC[4].icell.PDM Iout 0.00112f
C4910 XA.XIR[4].XIC[7].icell.Ien VPWR 0.19065f
C4911 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04522f
C4912 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.0171f
C4913 XThC.XTBN.A XThC.Tn[11] 0.12129f
C4914 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.03424f
C4915 XA.XIR[13].XIC[8].icell.Ien Vbias 0.21238f
C4916 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.SM 0.00383f
C4917 XA.XIR[4].XIC[4].icell.Ien Iout 0.06483f
C4918 XA.XIR[3].XIC[8].icell.SM VPWR 0.00158f
C4919 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PUM 0.00131f
C4920 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.01406f
C4921 XA.XIR[9].XIC[4].icell.SM Vbias 0.00701f
C4922 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.SM 0.00383f
C4923 XA.XIR[8].XIC[3].icell.PUM VPWR 0.01036f
C4924 XA.XIR[0].XIC_dummy_right.icell.SM VPWR 0.00123f
C4925 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.SM 0.00383f
C4926 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.03424f
C4927 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C4928 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.03976f
C4929 XA.XIR[3].XIC[5].icell.SM Iout 0.00388f
C4930 XA.XIR[2].XIC[12].icell.PDM VPWR 0.00863f
C4931 XThC.XTBN.Y a_4067_9615# 0.08456f
C4932 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.03424f
C4933 XThC.Tn[11] XThR.Tn[4] 0.28062f
C4934 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.SM 0.00383f
C4935 XA.XIR[11].XIC[0].icell.PDM Vbias 0.04002f
C4936 XA.XIR[14].XIC[12].icell.Ien Iout 0.06483f
C4937 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.03424f
C4938 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00529f
C4939 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.01406f
C4940 XThC.Tn[0] Vbias 1.90273f
C4941 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.03976f
C4942 XThR.Tn[14] XA.XIR[14].XIC[12].icell.PDM 0.0033f
C4943 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[5].icell.SM 0.00383f
C4944 XA.XIR[2].XIC[9].icell.PDM Iout 0.00112f
C4945 XA.XIR[14].XIC[10].icell.PDM Iout 0.00112f
C4946 XThR.Tn[10] XThR.Tn[12] 0.00142f
C4947 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02698f
C4948 XThR.Tn[1] XA.XIR[2].XIC[9].icell.SM 0.00121f
C4949 XThR.Tn[9] XA.XIR[10].XIC[9].icell.SM 0.00121f
C4950 XA.XIR[9].XIC[10].icell.PUM VPWR 0.01036f
C4951 XA.XIR[6].XIC[10].icell.PUM Vbias 0.00347f
C4952 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.03424f
C4953 XA.XIR[12].XIC[0].icell.PDM Iout 0.00112f
C4954 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PUM 0.00131f
C4955 XThC.XTB3.Y a_8739_9569# 0.07285f
C4956 XThR.Tn[14] XA.XIR[15].XIC[3].icell.SM 0.00121f
C4957 XA.XIR[5].XIC[13].icell.PDM Vbias 0.04058f
C4958 XA.XIR[13].XIC[13].icell.Ien Vbias 0.21238f
C4959 XA.XIR[7].XIC[2].icell.PUM Vbias 0.00347f
C4960 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.SM 0.00188f
C4961 XThC.XTB6.Y XThC.Tn[7] 0.01462f
C4962 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00212f
C4963 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.03424f
C4964 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08027f
C4965 XA.XIR[3].XIC[13].icell.PUM VPWR 0.01036f
C4966 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.03976f
C4967 XA.XIR[1].XIC[3].icell.PUM Vbias 0.00347f
C4968 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04f
C4969 XThR.Tn[3] XA.XIR[3].XIC[11].icell.PDM 0.0033f
C4970 XA.XIR[11].XIC_15.icell.PDM VPWR 0.06959f
C4971 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02698f
C4972 a_n1049_5611# XThR.Tn[6] 0.00158f
C4973 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13469f
C4974 XA.XIR[2].XIC[14].icell.Ien VPWR 0.1907f
C4975 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02698f
C4976 XThC.Tn[9] Iout 0.83891f
C4977 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01799f
C4978 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.01406f
C4979 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06536f
C4980 XA.XIR[14].XIC[1].icell.PUM VPWR 0.01036f
C4981 XA.XIR[0].XIC[3].icell.Ien Vbias 0.21246f
C4982 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02698f
C4983 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.01406f
C4984 XA.XIR[8].XIC[9].icell.PUM Vbias 0.00347f
C4985 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PUM 0.00131f
C4986 XA.XIR[6].XIC[13].icell.PDM Iout 0.00112f
C4987 XA.XIR[7].XIC[8].icell.PDM VPWR 0.00863f
C4988 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.03424f
C4989 XThR.Tn[10] XA.XIR[10].XIC[13].icell.PDM 0.0033f
C4990 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.15089f
C4991 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01799f
C4992 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PUM 0.00131f
C4993 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00529f
C4994 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.03424f
C4995 XThR.Tn[13] VPWR 7.6901f
C4996 XThR.Tn[4] XA.XIR[4].XIC[11].icell.PDM 0.0033f
C4997 XA.XIR[1].XIC[9].icell.PDM VPWR 0.00863f
C4998 XA.XIR[7].XIC[5].icell.PDM Iout 0.00112f
C4999 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.SM 0.00383f
C5000 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.PUM 0.00112f
C5001 XA.XIR[9].XIC_15.icell.PDM VPWR 0.06959f
C5002 XA.XIR[10].XIC[0].icell.SM Vbias 0.00675f
C5003 XA.XIR[6].XIC_15.icell.PDM Vbias 0.04206f
C5004 XThC.XTBN.A data[0] 0.02545f
C5005 XA.XIR[10].XIC[14].icell.Ien Vbias 0.21238f
C5006 XThC.XTB6.Y a_5949_10571# 0.01283f
C5007 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9] 0.0033f
C5008 XThR.Tn[9] XA.XIR[10].XIC[11].icell.Ien 0.00321f
C5009 XA.XIR[15].XIC_dummy_right.icell.Ien Vbias 0.00287f
C5010 XThR.Tn[7] XA.XIR[8].XIC[10].icell.SM 0.00121f
C5011 XA.XIR[1].XIC[6].icell.PDM Iout 0.00112f
C5012 XA.XIR[4].XIC[14].icell.SM VPWR 0.00208f
C5013 XThR.Tn[12] XA.XIR[13].XIC[2].icell.Ien 0.00321f
C5014 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.PDM 0.00589f
C5015 XThC.XTBN.Y XThC.Tn[3] 0.62681f
C5016 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02698f
C5017 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.SM 0.00383f
C5018 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C5019 XA.XIR[0].XIC[7].icell.SM VPWR 0.00158f
C5020 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.15119f
C5021 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.03976f
C5022 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02698f
C5023 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.15089f
C5024 XThR.Tn[2] XA.XIR[3].XIC[14].icell.Ien 0.00321f
C5025 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.03424f
C5026 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.15089f
C5027 XA.XIR[0].XIC[4].icell.SM Iout 0.00367f
C5028 XA.XIR[8].XIC[12].icell.PDM Iout 0.00112f
C5029 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.15089f
C5030 XA.XIR[11].XIC[1].icell.Ien Iout 0.06483f
C5031 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.SM 0.00188f
C5032 XA.XIR[2].XIC[1].icell.PDM VPWR 0.00863f
C5033 XThC.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.00111f
C5034 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04522f
C5035 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.03424f
C5036 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01776f
C5037 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.03976f
C5038 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04522f
C5039 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.03424f
C5040 XThC.XTB4.Y XThC.Tn[7] 0.01797f
C5041 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.04037f
C5042 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.SM 0.00383f
C5043 XA.XIR[8].XIC[14].icell.PDM Vbias 0.04058f
C5044 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.01406f
C5045 XA.XIR[3].XIC_dummy_right.icell.Ien Vbias 0.00287f
C5046 XA.XIR[2].XIC_15.icell.Ien Iout 0.06485f
C5047 XA.XIR[15].XIC[7].icell.PDM Vbias 0.04058f
C5048 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02698f
C5049 XA.XIR[1].XIC[0].icell.Ien VPWR 0.19066f
C5050 XThC.Tn[0] XThR.Tn[6] 0.28065f
C5051 XThC.Tn[2] XThR.Tn[8] 0.28062f
C5052 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00529f
C5053 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04522f
C5054 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.15089f
C5055 XThR.Tn[10] XA.XIR[11].XIC[7].icell.Ien 0.00321f
C5056 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02698f
C5057 XThR.XTB2.Y XThR.Tn[2] 0.00271f
C5058 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.SM 0.00383f
C5059 XA.XIR[4].XIC[0].icell.Ien VPWR 0.19066f
C5060 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00212f
C5061 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.SM 0.00188f
C5062 XThR.Tn[7] XA.XIR[8].XIC[0].icell.Ien 0.00321f
C5063 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.03424f
C5064 XA.XIR[14].XIC[10].icell.SM Iout 0.00388f
C5065 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.SM 0.00383f
C5066 VPWR Vbias 0.21627p
C5067 XThR.Tn[5] XA.XIR[6].XIC[12].icell.Ien 0.00321f
C5068 a_4861_9615# XThC.Tn[3] 0.27012f
C5069 XA.XIR[3].XIC[1].icell.SM VPWR 0.00158f
C5070 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PUM 0.00131f
C5071 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.03976f
C5072 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06536f
C5073 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02698f
C5074 XA.XIR[12].XIC[2].icell.Ien Vbias 0.21238f
C5075 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.SM 0.00383f
C5076 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.01406f
C5077 XA.XIR[8].XIC[14].icell.Ien Iout 0.06483f
C5078 XA.XIR[2].XIC[5].icell.PDM VPWR 0.00863f
C5079 XA.XIR[0].XIC[13].icell.SM Vbias 0.00701f
C5080 XA.XIR[15].XIC[7].icell.Ien Iout 0.06816f
C5081 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.03424f
C5082 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02698f
C5083 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.03424f
C5084 XA.XIR[14].XIC[6].icell.PDM VPWR 0.00863f
C5085 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.03424f
C5086 XA.XIR[2].XIC[2].icell.PDM Iout 0.00112f
C5087 XThC.Tn[3] XThR.Tn[5] 0.28062f
C5088 XA.XIR[11].XIC[5].icell.PDM Vbias 0.04058f
C5089 XA.XIR[11].XIC_15.icell.SM Iout 0.0047f
C5090 XThR.XTB5.A XThR.XTB7.A 0.07862f
C5091 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.SM 0.00383f
C5092 XA.XIR[15].XIC[11].icell.PDM Vbias 0.04058f
C5093 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.SM 0.00188f
C5094 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.03976f
C5095 XA.XIR[13].XIC[5].icell.SM VPWR 0.00158f
C5096 XA.XIR[13].XIC[12].icell.PUM Vbias 0.00347f
C5097 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.SM 0.00383f
C5098 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08027f
C5099 XThR.Tn[1] XA.XIR[2].XIC[2].icell.SM 0.00121f
C5100 XA.XIR[10].XIC[4].icell.SM Vbias 0.00701f
C5101 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.SM 0.00383f
C5102 XA.XIR[1].XIC_15.icell.Ien VPWR 0.25675f
C5103 XA.XIR[9].XIC[3].icell.PUM VPWR 0.01036f
C5104 XA.XIR[6].XIC[3].icell.PUM Vbias 0.00347f
C5105 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Iout 0.00347f
C5106 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.01406f
C5107 XThR.Tn[9] XA.XIR[9].XIC[7].icell.PDM 0.0033f
C5108 XA.XIR[11].XIC[11].icell.SM VPWR 0.00158f
C5109 XA.XIR[12].XIC[6].icell.SM VPWR 0.00158f
C5110 XA.XIR[13].XIC[2].icell.SM Iout 0.00388f
C5111 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02698f
C5112 XThC.Tn[1] XThR.Tn[1] 0.28062f
C5113 XThR.Tn[6] XA.XIR[6].XIC_15.icell.PDM 0.0033f
C5114 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00212f
C5115 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PUM 0.00131f
C5116 XA.XIR[5].XIC[6].icell.PDM Vbias 0.04058f
C5117 a_7331_10587# VPWR 0.0063f
C5118 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02698f
C5119 XA.XIR[12].XIC[3].icell.SM Iout 0.00388f
C5120 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04522f
C5121 XA.XIR[11].XIC[8].icell.Ien VPWR 0.19065f
C5122 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35627f
C5123 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.SM 0.00383f
C5124 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.03976f
C5125 XThR.Tn[3] XA.XIR[3].XIC[4].icell.PDM 0.0033f
C5126 XA.XIR[4].XIC[6].icell.Ien Vbias 0.21238f
C5127 XA.XIR[11].XIC[5].icell.Ien Iout 0.06483f
C5128 XA.XIR[6].XIC[9].icell.PDM VPWR 0.00863f
C5129 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00529f
C5130 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.15089f
C5131 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PDM 0.00182f
C5132 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00529f
C5133 XThR.XTB6.A a_n1319_5317# 0.00295f
C5134 XA.XIR[3].XIC[7].icell.SM Vbias 0.00701f
C5135 XThC.XTB3.Y data[0] 0.03253f
C5136 XA.XIR[5].XIC[9].icell.Ien VPWR 0.19065f
C5137 XA.XIR[6].XIC[6].icell.PDM Iout 0.00112f
C5138 XA.XIR[8].XIC[2].icell.PUM Vbias 0.00347f
C5139 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PUM 0.00131f
C5140 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C5141 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.15089f
C5142 XA.XIR[2].XIC[11].icell.PDM Vbias 0.04058f
C5143 XThR.Tn[0] XA.XIR[1].XIC[14].icell.Ien 0.00321f
C5144 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02698f
C5145 XThR.XTB2.Y a_n997_3979# 0.00191f
C5146 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.15089f
C5147 XA.XIR[4].XIC[10].icell.SM VPWR 0.00158f
C5148 XA.XIR[5].XIC[6].icell.Ien Iout 0.06483f
C5149 XThR.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.0033f
C5150 XA.XIR[10].XIC[8].icell.SM Vbias 0.00701f
C5151 XThR.Tn[12] XThR.Tn[13] 0.07749f
C5152 XThR.Tn[7] XA.XIR[8].XIC[3].icell.SM 0.00121f
C5153 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04522f
C5154 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.01406f
C5155 XA.XIR[4].XIC[7].icell.SM Iout 0.00388f
C5156 XThC.Tn[0] XA.XIR[6].XIC_dummy_left.icell.Iout 0.00111f
C5157 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11218f
C5158 XThR.XTB7.A data[5] 0.06538f
C5159 XA.XIR[11].XIC[13].icell.Ien VPWR 0.19065f
C5160 XA.XIR[9].XIC[9].icell.PUM Vbias 0.00347f
C5161 XA.XIR[0].XIC[0].icell.SM VPWR 0.00158f
C5162 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00529f
C5163 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04522f
C5164 XA.XIR[8].XIC[8].icell.PDM VPWR 0.00863f
C5165 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.03976f
C5166 XThR.Tn[8] XA.XIR[9].XIC[10].icell.Ien 0.00321f
C5167 XThR.Tn[6] VPWR 6.65699f
C5168 a_n1049_7787# XThR.XTB3.Y 0.00124f
C5169 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00529f
C5170 XA.XIR[11].XIC[9].icell.Ien Iout 0.06483f
C5171 XA.XIR[8].XIC[5].icell.PDM Iout 0.00112f
C5172 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.15089f
C5173 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00529f
C5174 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00529f
C5175 XA.XIR[14].XIC_15.icell.PDM VPWR 0.06959f
C5176 XA.XIR[2].XIC[11].icell.Ien Iout 0.06483f
C5177 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.15089f
C5178 XA.XIR[3].XIC[12].icell.PUM Vbias 0.00347f
C5179 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.03976f
C5180 XThC.Tn[13] VPWR 6.93877f
C5181 XA.XIR[5].XIC[12].icell.SM VPWR 0.00158f
C5182 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PUM 0.00209f
C5183 XThR.Tn[1] a_n1049_7787# 0.26879f
C5184 XA.XIR[2].XIC[13].icell.Ien Vbias 0.21238f
C5185 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PUM 0.00529f
C5186 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04522f
C5187 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.SM 0.00188f
C5188 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00212f
C5189 XA.XIR[9].XIC[12].icell.PDM Iout 0.00112f
C5190 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.01406f
C5191 XThR.XTB6.A XThR.Tn[9] 0.00838f
C5192 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.04493f
C5193 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.03981f
C5194 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PUM 0.00131f
C5195 XThC.Tn[0] XThR.Tn[4] 0.28067f
C5196 XA.XIR[7].XIC[7].icell.PDM Vbias 0.04058f
C5197 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.SM 0.00383f
C5198 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.01406f
C5199 a_9827_9569# Vbias 0.00395f
C5200 XThC.Tn[12] XThR.Tn[9] 0.28062f
C5201 XA.XIR[13].XIC[0].icell.SM Vbias 0.00675f
C5202 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C5203 XA.XIR[13].XIC[14].icell.Ien Vbias 0.21238f
C5204 XA.XIR[1].XIC[8].icell.PDM Vbias 0.04058f
C5205 XA.XIR[9].XIC[14].icell.PDM Vbias 0.04058f
C5206 XA.XIR[15].XIC[3].icell.Ien VPWR 0.32782f
C5207 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00529f
C5208 XThR.Tn[8] XA.XIR[9].XIC[13].icell.SM 0.00121f
C5209 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.38945f
C5210 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00529f
C5211 XThR.Tn[12] Vbias 3.71742f
C5212 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08017f
C5213 XA.XIR[3].XIC_15.icell.PDM Iout 0.0013f
C5214 XA.XIR[0].XIC[6].icell.SM Vbias 0.00701f
C5215 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04522f
C5216 XA.XIR[15].XIC[0].icell.Ien Iout 0.06808f
C5217 XA.XIR[6].XIC_15.icell.Ien VPWR 0.25675f
C5218 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.03981f
C5219 XA.XIR[7].XIC[10].icell.Ien VPWR 0.19065f
C5220 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00529f
C5221 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.03976f
C5222 XA.XIR[1].XIC_dummy_left.icell.SM VPWR 0.00269f
C5223 XA.XIR[11].XIC[12].icell.PDM Iout 0.00112f
C5224 XA.XIR[14].XIC[1].icell.Ien Iout 0.06483f
C5225 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01776f
C5226 XA.XIR[1].XIC[11].icell.Ien VPWR 0.19065f
C5227 XA.XIR[7].XIC[7].icell.Ien Iout 0.06483f
C5228 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.03976f
C5229 XThR.XTB3.Y XThR.Tn[9] 0.00285f
C5230 XA.XIR[4].XIC_dummy_left.icell.SM VPWR 0.00269f
C5231 XThR.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.0033f
C5232 XA.XIR[1].XIC[8].icell.Ien Iout 0.06483f
C5233 XA.XIR[9].XIC[14].icell.Ien Iout 0.06483f
C5234 XThR.Tn[12] XA.XIR[13].XIC[5].icell.SM 0.00121f
C5235 XA.XIR[10].XIC_15.icell.Ien Vbias 0.21343f
C5236 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00529f
C5237 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PUM 0.00529f
C5238 XA.XIR[0].XIC[12].icell.PUM VPWR 0.00971f
C5239 XThR.Tn[11] XA.XIR[12].XIC[11].icell.SM 0.00121f
C5240 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Ien 0.00217f
C5241 XThR.Tn[13] a_n997_1803# 0.0021f
C5242 XThC.XTB2.Y a_3773_9615# 0.2342f
C5243 XA.XIR[10].XIC[13].icell.PDM Vbias 0.04058f
C5244 XThC.Tn[10] XThR.Tn[11] 0.28062f
C5245 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.01406f
C5246 XThC.XTB1.Y data[0] 0.06453f
C5247 XThC.Tn[7] Iout 0.84146f
C5248 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00529f
C5249 XA.XIR[8].XIC[1].icell.PDM Iout 0.00112f
C5250 XThC.XTB7.B Vbias 0.04962f
C5251 XThR.Tn[11] XA.XIR[12].XIC[8].icell.Ien 0.00321f
C5252 XA.XIR[10].XIC[3].icell.PUM VPWR 0.01036f
C5253 XA.XIR[6].XIC[2].icell.PDM VPWR 0.00863f
C5254 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.SM 0.00188f
C5255 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.03976f
C5256 XA.XIR[3].XIC[0].icell.SM Vbias 0.00675f
C5257 XA.XIR[7].XIC[13].icell.SM VPWR 0.00158f
C5258 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11178f
C5259 XA.XIR[5].XIC[2].icell.Ien VPWR 0.19065f
C5260 XThR.XTB6.A a_n1319_6405# 0.00306f
C5261 XA.XIR[2].XIC[4].icell.PDM Vbias 0.04058f
C5262 XA.XIR[11].XIC[12].icell.PUM VPWR 0.01036f
C5263 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00529f
C5264 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.01406f
C5265 XA.XIR[14].XIC[5].icell.PDM Vbias 0.04058f
C5266 XA.XIR[4].XIC[3].icell.SM VPWR 0.00158f
C5267 XA.XIR[1].XIC[11].icell.SM Iout 0.00388f
C5268 XA.XIR[14].XIC_15.icell.SM Iout 0.0047f
C5269 XA.XIR[13].XIC[4].icell.SM Vbias 0.00701f
C5270 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04522f
C5271 XA.XIR[4].XIC[0].icell.SM Iout 0.00388f
C5272 XA.XIR[3].XIC[6].icell.PUM VPWR 0.01036f
C5273 XA.XIR[14].XIC[11].icell.SM VPWR 0.00158f
C5274 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.03424f
C5275 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.SM 0.00383f
C5276 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.03976f
C5277 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.SM 0.00383f
C5278 XThC.XTBN.A VPWR 0.88811f
C5279 XThR.Tn[8] XA.XIR[9].XIC[3].icell.Ien 0.00321f
C5280 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00529f
C5281 XA.XIR[12].XIC[5].icell.SM Vbias 0.00701f
C5282 XThR.Tn[11] XA.XIR[12].XIC[13].icell.Ien 0.00321f
C5283 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.01406f
C5284 XA.XIR[2].XIC[7].icell.Ien VPWR 0.19065f
C5285 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.03976f
C5286 XA.XIR[14].XIC[8].icell.Ien VPWR 0.19119f
C5287 a_9827_9569# XThC.Tn[13] 0.00173f
C5288 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.03976f
C5289 XA.XIR[11].XIC[7].icell.Ien Vbias 0.21238f
C5290 XA.XIR[2].XIC[4].icell.Ien Iout 0.06483f
C5291 XThC.Tn[0] XThC.Tn[2] 0.1179f
C5292 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04522f
C5293 XThR.Tn[4] VPWR 6.69328f
C5294 XThC.Tn[10] XThR.Tn[7] 0.28062f
C5295 XA.XIR[14].XIC[5].icell.Ien Iout 0.06483f
C5296 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PUM 0.00131f
C5297 XThC.Tn[13] XThR.Tn[12] 0.28063f
C5298 XThC.Tn[5] XThC.Tn[6] 0.31356f
C5299 a_n997_2667# VPWR 0.0165f
C5300 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.03424f
C5301 XA.XIR[6].XIC[8].icell.PDM Vbias 0.04058f
C5302 XA.XIR[9].XIC[8].icell.PDM VPWR 0.00863f
C5303 XA.XIR[7].XIC[14].icell.SM Iout 0.00388f
C5304 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.15089f
C5305 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00529f
C5306 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.03976f
C5307 XA.XIR[9].XIC[5].icell.PDM Iout 0.00112f
C5308 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.03976f
C5309 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00529f
C5310 XA.XIR[1].XIC_dummy_right.icell.SM VPWR 0.00123f
C5311 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PUM 0.00131f
C5312 XA.XIR[5].XIC[8].icell.Ien Vbias 0.21238f
C5313 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04522f
C5314 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PUM 0.00529f
C5315 XA.XIR[13].XIC[8].icell.SM Vbias 0.00701f
C5316 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10] 0.0033f
C5317 XThR.Tn[2] XA.XIR[3].XIC[7].icell.Ien 0.00321f
C5318 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.15089f
C5319 XA.XIR[4].XIC[9].icell.SM Vbias 0.00701f
C5320 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00529f
C5321 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.01406f
C5322 XA.XIR[6].XIC[11].icell.Ien VPWR 0.19065f
C5323 XA.XIR[14].XIC[13].icell.Ien VPWR 0.19119f
C5324 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.002f
C5325 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.01406f
C5326 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04522f
C5327 XA.XIR[7].XIC[3].icell.Ien VPWR 0.19065f
C5328 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.03976f
C5329 XA.XIR[8].XIC[7].icell.PDM Vbias 0.04058f
C5330 XA.XIR[6].XIC[8].icell.Ien Iout 0.06483f
C5331 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00212f
C5332 XThR.Tn[1] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00126f
C5333 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.01406f
C5334 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04522f
C5335 XThC.Tn[12] XThR.Tn[10] 0.28062f
C5336 XA.XIR[14].XIC[9].icell.Ien Iout 0.06483f
C5337 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.SM 0.00188f
C5338 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02698f
C5339 XThC.XTB7.Y XThC.Tn[8] 0.07806f
C5340 XA.XIR[14].XIC[1].icell.PDM Vbias 0.04058f
C5341 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.15089f
C5342 XA.XIR[5].XIC[9].icell.SM Iout 0.00388f
C5343 XThC.XTB7.B XThC.Tn[13] 0.00276f
C5344 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.03011f
C5345 XA.XIR[7].XIC[0].icell.Ien Iout 0.06474f
C5346 XA.XIR[1].XIC[4].icell.Ien VPWR 0.19065f
C5347 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13469f
C5348 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.01406f
C5349 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04522f
C5350 XA.XIR[10].XIC[9].icell.SM Vbias 0.00701f
C5351 XA.XIR[1].XIC[1].icell.Ien Iout 0.06483f
C5352 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PUM 0.00131f
C5353 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C5354 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.03424f
C5355 XA.XIR[5].XIC[11].icell.SM Vbias 0.00701f
C5356 XA.XIR[0].XIC[5].icell.PUM VPWR 0.00971f
C5357 XThR.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.00321f
C5358 XA.XIR[8].XIC[10].icell.Ien VPWR 0.19065f
C5359 XA.XIR[11].XIC[0].icell.SM VPWR 0.00158f
C5360 XThR.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.0033f
C5361 XA.XIR[11].XIC[14].icell.Ien VPWR 0.1907f
C5362 XA.XIR[4].XIC[14].icell.PUM Vbias 0.00347f
C5363 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C5364 XA.XIR[8].XIC[7].icell.Ien Iout 0.06483f
C5365 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PUM 0.00529f
C5366 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02698f
C5367 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04522f
C5368 XA.XIR[2].XIC[14].icell.SM VPWR 0.00208f
C5369 XThR.Tn[2] XA.XIR[2].XIC[14].icell.PDM 0.0033f
C5370 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02698f
C5371 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.03982f
C5372 XA.XIR[11].XIC[10].icell.Ien Iout 0.06483f
C5373 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.SM 0.00188f
C5374 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00212f
C5375 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Iout 0.00347f
C5376 XA.XIR[15].XIC[2].icell.Ien Vbias 0.17911f
C5377 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08017f
C5378 XA.XIR[6].XIC[11].icell.SM Iout 0.00388f
C5379 XThR.Tn[11] XA.XIR[11].XIC[4].icell.PDM 0.0033f
C5380 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.03011f
C5381 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.0171f
C5382 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.03424f
C5383 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.SM 0.00188f
C5384 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.SM 0.00383f
C5385 XThR.Tn[10] XA.XIR[11].XIC[3].icell.SM 0.00121f
C5386 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Iout 0.00347f
C5387 XThC.Tn[6] XA.XIR[0].XIC[7].icell.Ien 0.00194f
C5388 XA.XIR[7].XIC[9].icell.Ien Vbias 0.21238f
C5389 XA.XIR[14].XIC[12].icell.PDM Iout 0.00112f
C5390 XThR.Tn[6] XA.XIR[6].XIC[8].icell.PDM 0.0033f
C5391 XThC.XTB3.Y VPWR 1.07067f
C5392 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PUM 0.00529f
C5393 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PUM 0.00131f
C5394 XA.XIR[4].XIC_15.icell.SM VPWR 0.00276f
C5395 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.01406f
C5396 XThC.XTB1.Y XThC.Tn[0] 0.19116f
C5397 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.SM 0.00383f
C5398 XThR.Tn[10] XA.XIR[10].XIC[7].icell.PDM 0.0033f
C5399 XA.XIR[1].XIC[10].icell.Ien Vbias 0.21238f
C5400 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.01406f
C5401 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.04037f
C5402 XA.XIR[10].XIC[11].icell.Ien Vbias 0.21238f
C5403 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PUM 0.00529f
C5404 XThC.Tn[2] VPWR 6.00305f
C5405 XA.XIR[8].XIC[13].icell.SM VPWR 0.00158f
C5406 XA.XIR[9].XIC[3].icell.PDM Vbias 0.04058f
C5407 XA.XIR[15].XIC[6].icell.SM VPWR 0.00158f
C5408 XThC.XTBN.A a_9827_9569# 0.09118f
C5409 XThC.XTB7.A a_6243_10571# 0.0017f
C5410 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.03424f
C5411 XA.XIR[13].XIC_15.icell.Ien Vbias 0.21343f
C5412 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02698f
C5413 XThR.Tn[2] XA.XIR[3].XIC[14].icell.SM 0.00121f
C5414 XThR.Tn[7] XA.XIR[7].XIC[13].icell.PDM 0.0033f
C5415 XThC.Tn[5] XA.XIR[0].XIC[6].icell.PDM 0.00307f
C5416 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.03982f
C5417 XA.XIR[0].XIC[11].icell.PUM Vbias 0.00347f
C5418 XA.XIR[15].XIC[3].icell.SM Iout 0.00388f
C5419 XA.XIR[2].XIC[0].icell.Ien VPWR 0.19066f
C5420 XThR.Tn[13] XA.XIR[14].XIC[7].icell.Ien 0.00321f
C5421 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.03424f
C5422 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02708f
C5423 XThC.Tn[10] XThR.Tn[14] 0.28062f
C5424 XA.XIR[13].XIC[13].icell.PDM Vbias 0.04058f
C5425 XA.XIR[6].XIC_dummy_right.icell.SM VPWR 0.00123f
C5426 XThC.Tn[8] XThR.Tn[0] 0.28104f
C5427 XA.XIR[7].XIC[10].icell.SM Iout 0.00388f
C5428 XThR.Tn[0] XA.XIR[1].XIC[7].icell.Ien 0.00321f
C5429 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02698f
C5430 XA.XIR[13].XIC[3].icell.PUM VPWR 0.01036f
C5431 XThC.Tn[1] XThR.Tn[9] 0.28062f
C5432 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11595f
C5433 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02698f
C5434 XA.XIR[5].XIC[1].icell.PDM Iout 0.00112f
C5435 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C5436 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.SM 0.00383f
C5437 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C5438 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.15089f
C5439 XA.XIR[12].XIC[4].icell.PUM VPWR 0.01036f
C5440 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C5441 XA.XIR[7].XIC[12].icell.SM Vbias 0.00701f
C5442 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04522f
C5443 XA.XIR[5].XIC[1].icell.Ien Vbias 0.21238f
C5444 XA.XIR[14].XIC[12].icell.PUM VPWR 0.01036f
C5445 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.SM 0.00383f
C5446 XThR.Tn[10] XA.XIR[10].XIC[11].icell.PDM 0.0033f
C5447 XA.XIR[1].XIC[13].icell.SM Vbias 0.00701f
C5448 XThC.XTB5.Y a_5155_9615# 0.24821f
C5449 XA.XIR[11].XIC[4].icell.SM VPWR 0.00158f
C5450 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.01406f
C5451 XThR.Tn[2] XA.XIR[3].XIC[0].icell.Ien 0.00321f
C5452 XA.XIR[4].XIC[2].icell.SM Vbias 0.00701f
C5453 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.01406f
C5454 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Ien 0.00531f
C5455 XThC.XTB7.A a_4067_9615# 0.0127f
C5456 XA.XIR[11].XIC[1].icell.SM Iout 0.00388f
C5457 XA.XIR[10].XIC[8].icell.PDM VPWR 0.00863f
C5458 XA.XIR[8].XIC[14].icell.SM Iout 0.00388f
C5459 XA.XIR[6].XIC[4].icell.Ien VPWR 0.19065f
C5460 XA.XIR[0].XIC_15.icell.PUM Vbias 0.00347f
C5461 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04522f
C5462 XA.XIR[3].XIC[5].icell.PUM Vbias 0.00347f
C5463 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02698f
C5464 XThC.XTBN.A XThC.XTB7.B 0.35142f
C5465 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00529f
C5466 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04522f
C5467 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04522f
C5468 XA.XIR[10].XIC[5].icell.PDM Iout 0.00112f
C5469 XA.XIR[5].XIC[5].icell.SM VPWR 0.00158f
C5470 XA.XIR[6].XIC[1].icell.Ien Iout 0.06483f
C5471 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08027f
C5472 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.SM 0.00383f
C5473 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.SM 0.00188f
C5474 XA.XIR[2].XIC[6].icell.Ien Vbias 0.21238f
C5475 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PUM 0.00529f
C5476 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.03424f
C5477 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.01406f
C5478 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.01406f
C5479 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04522f
C5480 XA.XIR[14].XIC[7].icell.Ien Vbias 0.21238f
C5481 XA.XIR[5].XIC[2].icell.SM Iout 0.00388f
C5482 XA.XIR[4].XIC[8].icell.PUM VPWR 0.01036f
C5483 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.SM 0.00383f
C5484 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35783f
C5485 XThR.Tn[2] Iout 1.16632f
C5486 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01193f
C5487 XThR.Tn[6] XA.XIR[7].XIC[9].icell.Ien 0.00321f
C5488 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.SM 0.00188f
C5489 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00212f
C5490 XA.XIR[3].XIC[11].icell.PDM VPWR 0.00863f
C5491 XA.XIR[9].XIC[7].icell.PDM Vbias 0.04058f
C5492 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02698f
C5493 XA.XIR[8].XIC[3].icell.Ien VPWR 0.19065f
C5494 XA.XIR[11].XIC[8].icell.SM VPWR 0.00158f
C5495 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.01406f
C5496 XThR.Tn[8] XA.XIR[9].XIC[6].icell.SM 0.00121f
C5497 XA.XIR[3].XIC[8].icell.PDM Iout 0.00112f
C5498 XA.XIR[2].XIC[10].icell.SM VPWR 0.00158f
C5499 XThC.XTBN.Y a_5155_9615# 0.07602f
C5500 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.01406f
C5501 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PUM 0.00529f
C5502 XThR.Tn[11] XA.XIR[12].XIC[0].icell.SM 0.00127f
C5503 XA.XIR[0].XIC[0].icell.PUM Vbias 0.00106f
C5504 XThR.Tn[5] XA.XIR[5].XIC[2].icell.PDM 0.0033f
C5505 XThR.Tn[11] XA.XIR[12].XIC[14].icell.Ien 0.00321f
C5506 XA.XIR[2].XIC[7].icell.SM Iout 0.00388f
C5507 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.SM 0.00188f
C5508 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.03976f
C5509 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04522f
C5510 XThC.XTB1.Y VPWR 1.1176f
C5511 Vbias bias[0] 0.1739f
C5512 bias[1] bias[2] 0.03172f
C5513 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.01406f
C5514 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.SM 0.00188f
C5515 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.SM 0.00188f
C5516 XA.XIR[14].XIC_dummy_left.icell.Ien Vbias 0.00342f
C5517 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.SM 0.00188f
C5518 XA.XIR[6].XIC[10].icell.Ien Vbias 0.21238f
C5519 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00212f
C5520 XA.XIR[9].XIC[10].icell.Ien VPWR 0.19065f
C5521 XThR.Tn[0] XA.XIR[1].XIC[14].icell.SM 0.00121f
C5522 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C5523 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Ien 0.00153f
C5524 XA.XIR[12].XIC[1].icell.PDM VPWR 0.00863f
C5525 XA.XIR[10].XIC[10].icell.PUM Vbias 0.00347f
C5526 XThR.Tn[3] XA.XIR[4].XIC[8].icell.Ien 0.00321f
C5527 XA.XIR[9].XIC[7].icell.Ien Iout 0.06483f
C5528 XThC.Tn[12] XThR.Tn[13] 0.28062f
C5529 XThC.Tn[0] XA.XIR[11].XIC_dummy_left.icell.Iout 0.00111f
C5530 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PUM 0.00529f
C5531 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02698f
C5532 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.03976f
C5533 XA.XIR[7].XIC[2].icell.Ien Vbias 0.21238f
C5534 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02698f
C5535 XThC.XTB7.A XThC.Tn[3] 0.03065f
C5536 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.SM 0.00188f
C5537 XThR.XTB2.Y a_n1049_6699# 0.00851f
C5538 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.15089f
C5539 XA.XIR[3].XIC[13].icell.Ien VPWR 0.19065f
C5540 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.01406f
C5541 XThR.Tn[6] XA.XIR[7].XIC[12].icell.SM 0.00121f
C5542 XA.XIR[1].XIC[3].icell.Ien Vbias 0.21238f
C5543 XThC.Tn[14] XThR.Tn[3] 0.28068f
C5544 XThR.Tn[2] XA.XIR[3].XIC[10].icell.SM 0.00121f
C5545 XA.XIR[13].XIC[9].icell.SM Vbias 0.00701f
C5546 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00529f
C5547 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.SM 0.00188f
C5548 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00212f
C5549 XThR.Tn[7] XA.XIR[7].XIC[6].icell.PDM 0.0033f
C5550 a_2979_9615# XThC.Tn[0] 0.28426f
C5551 XThC.Tn[4] XThR.Tn[2] 0.28062f
C5552 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.01406f
C5553 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.PDM 0.00589f
C5554 XThC.Tn[2] XThR.Tn[12] 0.28062f
C5555 XA.XIR[0].XIC[4].icell.PUM Vbias 0.00347f
C5556 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.SM 0.00188f
C5557 XA.XIR[14].XIC[0].icell.SM VPWR 0.00158f
C5558 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00212f
C5559 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8] 0.0033f
C5560 XThR.Tn[4] XA.XIR[5].XIC[8].icell.Ien 0.00321f
C5561 XA.XIR[7].XIC[6].icell.SM VPWR 0.00158f
C5562 XA.XIR[8].XIC[9].icell.Ien Vbias 0.21238f
C5563 XA.XIR[14].XIC[14].icell.Ien VPWR 0.19124f
C5564 XA.XIR[11].XIC[2].icell.PDM Vbias 0.04058f
C5565 XThR.Tn[1] XA.XIR[2].XIC[14].icell.Ien 0.00321f
C5566 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00212f
C5567 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04522f
C5568 XA.XIR[7].XIC[3].icell.SM Iout 0.00388f
C5569 XA.XIR[1].XIC[7].icell.SM VPWR 0.00158f
C5570 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00212f
C5571 XA.XIR[14].XIC[10].icell.Ien Iout 0.06483f
C5572 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06536f
C5573 XA.XIR[9].XIC[13].icell.SM VPWR 0.00158f
C5574 XA.XIR[10].XIC[3].icell.PDM Vbias 0.04058f
C5575 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PUM 0.00529f
C5576 XA.XIR[6].XIC[13].icell.SM Vbias 0.00701f
C5577 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C5578 XA.XIR[1].XIC[4].icell.SM Iout 0.00388f
C5579 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01897f
C5580 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.03981f
C5581 XThR.Tn[3] XA.XIR[4].XIC[11].icell.SM 0.00121f
C5582 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PUM 0.00131f
C5583 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.01406f
C5584 XA.XIR[0].XIC[10].icell.PDM VPWR 0.00806f
C5585 XThR.Tn[1] XA.XIR[1].XIC[9].icell.PDM 0.0033f
C5586 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00529f
C5587 XThR.Tn[5] XA.XIR[6].XIC[8].icell.SM 0.00121f
C5588 XA.XIR[12].XIC[2].icell.PDM Iout 0.00112f
C5589 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C5590 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PUM 0.00529f
C5591 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C5592 XA.XIR[8].XIC[10].icell.SM Iout 0.00388f
C5593 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.PDM 0.00589f
C5594 XA.XIR[2].XIC_dummy_left.icell.SM VPWR 0.00269f
C5595 XThC.Tn[1] XThR.Tn[10] 0.28062f
C5596 XThC.Tn[12] Vbias 2.39712f
C5597 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PUM 0.00209f
C5598 XA.XIR[11].XIC_15.icell.Ien VPWR 0.25675f
C5599 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.SM 0.00383f
C5600 XThR.Tn[11] XA.XIR[12].XIC[4].icell.SM 0.00121f
C5601 XA.XIR[13].XIC[11].icell.Ien Vbias 0.21238f
C5602 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04522f
C5603 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.SM 0.00383f
C5604 XThC.XTB7.B XThC.Tn[2] 0.00273f
C5605 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PUM 0.00529f
C5606 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35783f
C5607 XThR.Tn[9] XA.XIR[10].XIC[2].icell.Ien 0.00321f
C5608 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.03424f
C5609 XA.XIR[15].XIC[5].icell.SM Vbias 0.00701f
C5610 XThR.Tn[4] XA.XIR[5].XIC[11].icell.SM 0.00121f
C5611 XA.XIR[8].XIC[12].icell.SM Vbias 0.00701f
C5612 XThC.XTB7.Y XThC.Tn[6] 0.2144f
C5613 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.15089f
C5614 XA.XIR[11].XIC[13].icell.PDM VPWR 0.00863f
C5615 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.03976f
C5616 XA.XIR[1].XIC[1].icell.PUM VPWR 0.01036f
C5617 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.01406f
C5618 XThC.XTB6.Y XThC.Tn[10] 0.02461f
C5619 XA.XIR[1].XIC[12].icell.PUM VPWR 0.01036f
C5620 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PUM 0.00131f
C5621 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.01406f
C5622 XA.XIR[4].XIC[1].icell.PUM VPWR 0.01036f
C5623 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00529f
C5624 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.15089f
C5625 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04522f
C5626 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.15119f
C5627 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00529f
C5628 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04522f
C5629 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PDM 0.00182f
C5630 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PUM 0.00131f
C5631 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11595f
C5632 XA.XIR[9].XIC[14].icell.SM Iout 0.00388f
C5633 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.SM 0.00188f
C5634 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.01406f
C5635 XA.XIR[10].XIC_dummy_right.icell.Ien Vbias 0.00287f
C5636 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04522f
C5637 XThR.Tn[6] XA.XIR[7].XIC[2].icell.Ien 0.00321f
C5638 XA.XIR[3].XIC[4].icell.PDM VPWR 0.00863f
C5639 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PUM 0.00131f
C5640 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.01406f
C5641 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PUM 0.00202f
C5642 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C5643 XA.XIR[12].XIC[3].icell.PUM Vbias 0.00347f
C5644 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C5645 XA.XIR[2].XIC[3].icell.SM VPWR 0.00158f
C5646 XA.XIR[8].XIC[0].icell.Ien Iout 0.06474f
C5647 XThR.Tn[1] Vbias 3.71829f
C5648 XThR.Tn[11] XA.XIR[12].XIC[8].icell.SM 0.00121f
C5649 XA.XIR[14].XIC[4].icell.SM VPWR 0.00158f
C5650 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04522f
C5651 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PUM 0.00131f
C5652 XA.XIR[2].XIC[0].icell.SM Iout 0.00388f
C5653 XA.XIR[11].XIC[3].icell.SM Vbias 0.00701f
C5654 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.11124f
C5655 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01776f
C5656 XA.XIR[14].XIC[1].icell.SM Iout 0.00388f
C5657 XThR.Tn[0] XA.XIR[1].XIC[10].icell.SM 0.00121f
C5658 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00212f
C5659 XA.XIR[13].XIC[8].icell.PDM VPWR 0.00863f
C5660 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.03976f
C5661 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00529f
C5662 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00529f
C5663 XA.XIR[6].XIC[3].icell.Ien Vbias 0.21238f
C5664 XA.XIR[10].XIC[7].icell.PDM Vbias 0.04058f
C5665 XA.XIR[9].XIC[3].icell.Ien VPWR 0.19065f
C5666 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04522f
C5667 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.SM 0.00188f
C5668 XA.XIR[13].XIC[5].icell.PDM Iout 0.00112f
C5669 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.01406f
C5670 XA.XIR[12].XIC[9].icell.PDM VPWR 0.00863f
C5671 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08064f
C5672 XThR.Tn[0] XA.XIR[0].XIC[13].icell.PDM 0.0033f
C5673 XA.XIR[5].XIC[4].icell.SM Vbias 0.00701f
C5674 XThR.Tn[3] XA.XIR[4].XIC[1].icell.Ien 0.00321f
C5675 a_2979_9615# VPWR 0.70527f
C5676 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.01406f
C5677 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.SM 0.00383f
C5678 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12] 0.0033f
C5679 XA.XIR[12].XIC[6].icell.PDM Iout 0.00112f
C5680 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00529f
C5681 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13469f
C5682 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PUM 0.00487f
C5683 XThR.Tn[2] XA.XIR[3].XIC[3].icell.SM 0.00121f
C5684 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PUM 0.00209f
C5685 XA.XIR[4].XIC[7].icell.PUM Vbias 0.00347f
C5686 XThC.XTB4.Y XThC.Tn[10] 0.01391f
C5687 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.01406f
C5688 XA.XIR[6].XIC[7].icell.SM VPWR 0.00158f
C5689 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04522f
C5690 XThR.Tn[2] XA.XIR[2].XIC[7].icell.PDM 0.0033f
C5691 XA.XIR[3].XIC[10].icell.PDM Vbias 0.04058f
C5692 XThC.Tn[6] XThR.Tn[0] 0.28071f
C5693 XThC.XTB4.Y a_4861_9615# 0.23756f
C5694 XA.XIR[14].XIC[8].icell.SM VPWR 0.00158f
C5695 XThR.Tn[13] XA.XIR[14].XIC[0].icell.Ien 0.00352f
C5696 XA.XIR[10].XIC[7].icell.Ien Iout 0.06483f
C5697 XThC.Tn[12] XThR.Tn[6] 0.28062f
C5698 XA.XIR[6].XIC[4].icell.SM Iout 0.00388f
C5699 XThC.Tn[14] XThR.Tn[8] 0.28068f
C5700 XA.XIR[5].XIC[10].icell.PUM VPWR 0.01036f
C5701 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00529f
C5702 XThR.Tn[4] XA.XIR[5].XIC[1].icell.Ien 0.00321f
C5703 XA.XIR[8].XIC[2].icell.Ien Vbias 0.21238f
C5704 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PUM 0.00529f
C5705 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PUM 0.00529f
C5706 XA.XIR[2].XIC[9].icell.SM Vbias 0.00701f
C5707 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13] 0.0033f
C5708 XThC.XTB5.Y a_7875_9569# 0.00418f
C5709 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00529f
C5710 XThC.Tn[12] XThC.Tn[13] 0.2418f
C5711 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38962f
C5712 XA.XIR[1].XIC[0].icell.SM VPWR 0.00158f
C5713 XA.XIR[4].XIC[13].icell.PDM VPWR 0.00863f
C5714 XA.XIR[10].XIC[11].icell.PDM Vbias 0.04058f
C5715 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.01406f
C5716 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00529f
C5717 XA.XIR[7].XIC_15.icell.SM Iout 0.0047f
C5718 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02698f
C5719 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C5720 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C5721 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Iout 0.00347f
C5722 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.03976f
C5723 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PUM 0.00487f
C5724 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00212f
C5725 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.SM 0.00188f
C5726 XA.XIR[4].XIC[10].icell.PDM Iout 0.00112f
C5727 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.SM 0.00383f
C5728 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00529f
C5729 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04522f
C5730 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.03982f
C5731 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.SM 0.00383f
C5732 XA.XIR[0].XIC[3].icell.PDM VPWR 0.00806f
C5733 XA.XIR[8].XIC[6].icell.SM VPWR 0.00158f
C5734 XA.XIR[9].XIC[9].icell.Ien Vbias 0.21238f
C5735 XA.XIR[13].XIC[10].icell.PUM Vbias 0.00347f
C5736 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00212f
C5737 XA.XIR[15].XIC[0].icell.PUM VPWR 0.01036f
C5738 XThR.Tn[5] XA.XIR[6].XIC[1].icell.SM 0.00121f
C5739 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PUM 0.00131f
C5740 XA.XIR[3].XIC[10].icell.Ien Iout 0.06483f
C5741 XThR.XTB3.Y XThR.Tn[6] 0.00298f
C5742 XThC.Tn[0] XA.XIR[14].XIC_dummy_left.icell.Iout 0.00111f
C5743 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.01406f
C5744 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00529f
C5745 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.04494f
C5746 XA.XIR[11].XIC[9].icell.SM VPWR 0.00158f
C5747 XA.XIR[8].XIC[3].icell.SM Iout 0.00388f
C5748 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.SM 0.00188f
C5749 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[8].icell.Ien 0.00212f
C5750 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.SM 0.00383f
C5751 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.SM 0.00188f
C5752 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PUM 0.00529f
C5753 XA.XIR[6].XIC[12].icell.PUM VPWR 0.01036f
C5754 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C5755 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PUM 0.00487f
C5756 XA.XIR[3].XIC[12].icell.Ien Vbias 0.21238f
C5757 XThR.Tn[9] XThR.Tn[10] 0.0923f
C5758 XThR.Tn[11] XA.XIR[12].XIC_15.icell.Ien 0.00116f
C5759 XA.XIR[5].XIC_15.icell.PDM VPWR 0.06959f
C5760 XThR.Tn[14] XA.XIR[15].XIC[11].icell.SM 0.00121f
C5761 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.SM 0.00188f
C5762 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.SM 0.00383f
C5763 XA.XIR[2].XIC[14].icell.PUM Vbias 0.00347f
C5764 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.03011f
C5765 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.03982f
C5766 XA.XIR[14].XIC[0].icell.Ien Vbias 0.21102f
C5767 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.03981f
C5768 XThC.Tn[13] XThR.Tn[1] 0.28063f
C5769 XA.XIR[7].XIC[5].icell.SM Vbias 0.00701f
C5770 XA.XIR[9].XIC[10].icell.SM Iout 0.00388f
C5771 XThC.XTBN.Y a_7875_9569# 0.229f
C5772 XThR.Tn[14] XA.XIR[15].XIC[8].icell.Ien 0.00321f
C5773 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.15089f
C5774 a_10915_9569# Vbias 0.00836f
C5775 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C5776 XA.XIR[4].XIC[12].icell.Ien Iout 0.06483f
C5777 XA.XIR[12].XIC_15.icell.PDM Iout 0.0013f
C5778 XA.XIR[13].XIC[3].icell.PDM Vbias 0.04058f
C5779 XA.XIR[1].XIC[6].icell.SM Vbias 0.00701f
C5780 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.15089f
C5781 XA.XIR[9].XIC[12].icell.SM Vbias 0.00701f
C5782 XA.XIR[15].XIC[4].icell.PUM VPWR 0.01036f
C5783 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PUM 0.00504f
C5784 XThR.Tn[14] XA.XIR[14].XIC[4].icell.PDM 0.0033f
C5785 XA.XIR[3].XIC[13].icell.SM Iout 0.00388f
C5786 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.002f
C5787 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.01406f
C5788 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.15089f
C5789 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PUM 0.00529f
C5790 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00529f
C5791 XA.XIR[0].XIC[9].icell.PDM Vbias 0.04065f
C5792 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.SM 0.00383f
C5793 XThR.Tn[13] XA.XIR[14].XIC[3].icell.SM 0.00121f
C5794 XA.XIR[2].XIC_15.icell.SM VPWR 0.00276f
C5795 XA.XIR[7].XIC[11].icell.PUM VPWR 0.01036f
C5796 XA.XIR[11].XIC[11].icell.Ien VPWR 0.19065f
C5797 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Ien 0.00217f
C5798 XThC.Tn[1] XThR.Tn[13] 0.28062f
C5799 XA.XIR[14].XIC_15.icell.Ien VPWR 0.25706f
C5800 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04522f
C5801 XThR.Tn[0] XA.XIR[1].XIC[3].icell.SM 0.00121f
C5802 XThR.Tn[13] XA.XIR[13].XIC[7].icell.PDM 0.0033f
C5803 VPWR bias[2] 1.5142f
C5804 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.1239f
C5805 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06536f
C5806 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02491f
C5807 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.01406f
C5808 XThC.Tn[3] XThR.Tn[3] 0.28062f
C5809 XThR.Tn[14] XA.XIR[15].XIC[13].icell.Ien 0.00321f
C5810 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.03976f
C5811 XA.XIR[14].XIC[13].icell.PDM VPWR 0.00863f
C5812 XThC.XTB2.Y XThC.Tn[10] 0.00106f
C5813 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00212f
C5814 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.03011f
C5815 XThR.Tn[0] XA.XIR[0].XIC[6].icell.PDM 0.0033f
C5816 XA.XIR[0].XIC[12].icell.Ien VPWR 0.19251f
C5817 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.SM 0.00188f
C5818 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PUM 0.00529f
C5819 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.15089f
C5820 XThR.Tn[12] XA.XIR[12].XIC[9].icell.PDM 0.0033f
C5821 XThC.XTB2.Y a_4861_9615# 0.00851f
C5822 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C5823 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.01406f
C5824 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01776f
C5825 XA.XIR[0].XIC[9].icell.Ien Iout 0.06455f
C5826 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.01406f
C5827 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02698f
C5828 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.03424f
C5829 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02698f
C5830 XA.XIR[13].XIC_dummy_right.icell.Ien Vbias 0.00287f
C5831 XA.XIR[10].XIC[3].icell.Ien VPWR 0.19065f
C5832 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02698f
C5833 XA.XIR[6].XIC[0].icell.SM VPWR 0.00158f
C5834 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00212f
C5835 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.SM 0.00188f
C5836 XThR.Tn[9] XA.XIR[10].XIC[5].icell.SM 0.00121f
C5837 XThC.XTBN.A XThC.Tn[12] 0.22686f
C5838 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08017f
C5839 XA.XIR[11].XIC_dummy_right.icell.SM VPWR 0.00123f
C5840 XA.XIR[3].XIC[3].icell.PDM Vbias 0.04058f
C5841 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C5842 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00212f
C5843 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.SM 0.00188f
C5844 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.SM 0.00383f
C5845 XA.XIR[5].XIC[3].icell.PUM VPWR 0.01036f
C5846 XThR.Tn[13] XA.XIR[13].XIC[11].icell.PDM 0.0033f
C5847 XA.XIR[2].XIC[2].icell.SM Vbias 0.00701f
C5848 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Iout 0.00347f
C5849 a_n1049_7493# VPWR 0.72111f
C5850 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.SM 0.00188f
C5851 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00212f
C5852 XThC.Tn[12] XThR.Tn[4] 0.28062f
C5853 XA.XIR[5].XIC[0].icell.Ien Iout 0.06474f
C5854 XA.XIR[14].XIC[3].icell.SM Vbias 0.00701f
C5855 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.11124f
C5856 XA.XIR[4].XIC[6].icell.PDM VPWR 0.00863f
C5857 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.01406f
C5858 XA.XIR[1].XIC[14].icell.PDM Iout 0.00112f
C5859 XThC.Tn[1] Vbias 2.36927f
C5860 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00529f
C5861 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01402f
C5862 XA.XIR[13].XIC[7].icell.PDM Vbias 0.04058f
C5863 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.SM 0.00383f
C5864 XA.XIR[4].XIC[3].icell.PDM Iout 0.00112f
C5865 XThR.Tn[6] XA.XIR[7].XIC[5].icell.SM 0.00121f
C5866 XThC.XTBN.Y Iout 0.00178f
C5867 XA.XIR[3].XIC[6].icell.Ien VPWR 0.19065f
C5868 XA.XIR[1].XIC_15.icell.PUM Vbias 0.00347f
C5869 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PUM 0.00529f
C5870 XA.XIR[9].XIC[2].icell.Ien Vbias 0.21238f
C5871 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02698f
C5872 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PUM 0.00131f
C5873 XA.XIR[3].XIC[3].icell.Ien Iout 0.06483f
C5874 XA.XIR[12].XIC[8].icell.PDM Vbias 0.04058f
C5875 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.01406f
C5876 XA.XIR[2].XIC[8].icell.PUM VPWR 0.01036f
C5877 XThC.XTB5.Y XThC.Tn[4] 0.19958f
C5878 XA.XIR[8].XIC_15.icell.SM Iout 0.0047f
C5879 a_10915_9569# XThC.Tn[13] 0.01061f
C5880 XA.XIR[11].XIC[8].icell.PUM Vbias 0.00347f
C5881 XThR.XTB3.Y XThR.Tn[4] 0.00382f
C5882 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00212f
C5883 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.SM 0.00188f
C5884 XThR.Tn[11] XA.XIR[12].XIC[9].icell.SM 0.00121f
C5885 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.SM 0.00383f
C5886 XThC.XTB6.Y a_7651_9569# 0.0046f
C5887 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00212f
C5888 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00212f
C5889 XThR.XTB3.Y a_n997_2667# 0.002f
C5890 XThR.Tn[1] XA.XIR[2].XIC[7].icell.Ien 0.00321f
C5891 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.SM 0.00188f
C5892 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.SM 0.00188f
C5893 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C5894 XA.XIR[6].XIC[6].icell.SM Vbias 0.00701f
C5895 XA.XIR[9].XIC[6].icell.SM VPWR 0.00158f
C5896 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01799f
C5897 XA.XIR[12].XIC[11].icell.SM Iout 0.00388f
C5898 XA.XIR[13].XIC[7].icell.Ien Iout 0.06483f
C5899 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00529f
C5900 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06536f
C5901 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00529f
C5902 XThR.XTB5.Y a_n997_3755# 0.00418f
C5903 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02698f
C5904 XThC.Tn[10] Iout 0.83982f
C5905 XA.XIR[9].XIC[3].icell.SM Iout 0.00388f
C5906 XA.XIR[5].XIC[9].icell.PUM Vbias 0.00347f
C5907 XThR.Tn[3] XA.XIR[4].XIC[4].icell.SM 0.00121f
C5908 XThR.Tn[14] XA.XIR[15].XIC[1].icell.Ien 0.00321f
C5909 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.PDM 0.00588f
C5910 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02698f
C5911 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04522f
C5912 XA.XIR[12].XIC[8].icell.Ien Iout 0.06483f
C5913 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.03424f
C5914 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00212f
C5915 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.SM 0.00383f
C5916 XA.XIR[13].XIC[11].icell.PDM Vbias 0.04058f
C5917 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.SM 0.00188f
C5918 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PUM 0.00131f
C5919 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02698f
C5920 XA.XIR[4].XIC[12].icell.PDM Vbias 0.04058f
C5921 XA.XIR[11].XIC[10].icell.PUM VPWR 0.01036f
C5922 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00529f
C5923 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.01406f
C5924 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11595f
C5925 XA.XIR[10].XIC[0].icell.PDM Iout 0.00112f
C5926 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.15089f
C5927 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.15089f
C5928 XThR.XTB7.Y a_n997_3755# 0.00476f
C5929 XA.XIR[0].XIC[2].icell.PDM Vbias 0.04065f
C5930 XA.XIR[7].XIC[4].icell.PUM VPWR 0.01036f
C5931 XThR.Tn[4] XA.XIR[5].XIC[4].icell.SM 0.00121f
C5932 XThC.XTBN.Y XThC.Tn[4] 0.61061f
C5933 XA.XIR[8].XIC[5].icell.SM Vbias 0.00701f
C5934 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.SM 0.00188f
C5935 XThR.Tn[5] Iout 1.16627f
C5936 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.SM 0.00383f
C5937 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PUM 0.00131f
C5938 XA.XIR[14].XIC[9].icell.SM VPWR 0.00158f
C5939 XThR.Tn[8] XA.XIR[8].XIC[9].icell.PDM 0.0033f
C5940 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02698f
C5941 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.SM 0.00383f
C5942 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.SM 0.00188f
C5943 XA.XIR[5].XIC[12].icell.PDM Iout 0.00112f
C5944 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.PDM 0.00589f
C5945 XA.XIR[1].XIC[5].icell.PUM VPWR 0.01036f
C5946 XThR.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.00321f
C5947 XThR.Tn[9] XA.XIR[9].XIC_15.icell.PDM 0.0033f
C5948 XThR.Tn[7] XA.XIR[8].XIC[8].icell.Ien 0.00321f
C5949 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.SM 0.00383f
C5950 XThR.XTBN.A data[7] 0.07741f
C5951 XA.XIR[12].XIC[0].icell.Ien VPWR 0.19066f
C5952 XA.XIR[8].XIC[0].icell.PDM VPWR 0.00863f
C5953 XA.XIR[12].XIC[13].icell.Ien Iout 0.06483f
C5954 XA.XIR[5].XIC[14].icell.PDM Vbias 0.04058f
C5955 XThC.XTB4.Y a_7651_9569# 0.00497f
C5956 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.01406f
C5957 XA.XIR[0].XIC[5].icell.Ien VPWR 0.19024f
C5958 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.15089f
C5959 XA.XIR[8].XIC[11].icell.PUM VPWR 0.01036f
C5960 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00212f
C5961 XA.XIR[11].XIC[3].icell.PDM VPWR 0.00863f
C5962 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PUM 0.00131f
C5963 XThC.Tn[1] XThR.Tn[6] 0.28062f
C5964 XA.XIR[4].XIC[14].icell.Ien Vbias 0.21238f
C5965 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.03976f
C5966 XThC.Tn[3] XThR.Tn[8] 0.28062f
C5967 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.01406f
C5968 XA.XIR[0].XIC[2].icell.Ien Iout 0.06455f
C5969 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04522f
C5970 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00529f
C5971 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.03424f
C5972 XThR.Tn[5] XA.XIR[5].XIC[9].icell.PDM 0.0033f
C5973 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[9].icell.SM 0.00383f
C5974 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01897f
C5975 XThC.Tn[6] XThC.Tn[8] 0.00105f
C5976 XThR.Tn[14] a_n997_715# 0.1927f
C5977 XA.XIR[6].XIC[14].icell.PDM Iout 0.00112f
C5978 XA.XIR[15].XIC[3].icell.PUM Vbias 0.00347f
C5979 a_4861_9615# XThC.Tn[4] 0.00198f
C5980 XThR.Tn[1] XA.XIR[2].XIC[14].icell.SM 0.00121f
C5981 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.SM 0.00188f
C5982 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02698f
C5983 XA.XIR[5].XIC[14].icell.Ien Iout 0.06483f
C5984 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01776f
C5985 XA.XIR[6].XIC_15.icell.PUM Vbias 0.00347f
C5986 XA.XIR[14].XIC[11].icell.Ien VPWR 0.19119f
C5987 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.03976f
C5988 XA.XIR[7].XIC[10].icell.PUM Vbias 0.00347f
C5989 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C5990 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02698f
C5991 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.03424f
C5992 XA.XIR[1].XIC[1].icell.PDM Vbias 0.04058f
C5993 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00212f
C5994 XThR.Tn[7] XA.XIR[8].XIC[11].icell.SM 0.00121f
C5995 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.01406f
C5996 XThR.Tn[3] XA.XIR[3].XIC[0].icell.PDM 0.00336f
C5997 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00212f
C5998 XThC.Tn[4] XThR.Tn[5] 0.28062f
C5999 XA.XIR[1].XIC[11].icell.PUM Vbias 0.00347f
C6000 XThC.XTB7.A data[2] 0.00198f
C6001 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08017f
C6002 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01193f
C6003 XThR.Tn[9] Vbias 3.71832f
C6004 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.03424f
C6005 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.15089f
C6006 XA.XIR[4].XIC[1].icell.PDM Vbias 0.04058f
C6007 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C6008 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PUM 0.00529f
C6009 XA.XIR[15].XIC[6].icell.PDM Iout 0.00112f
C6010 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.01406f
C6011 XA.XIR[0].XIC[11].icell.Ien Vbias 0.21246f
C6012 XA.XIR[2].XIC[1].icell.PUM VPWR 0.01036f
C6013 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35783f
C6014 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PUM 0.00131f
C6015 XA.XIR[7].XIC[1].icell.PDM VPWR 0.00863f
C6016 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04522f
C6017 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[1].icell.Ien 0.00212f
C6018 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C6019 XThC.Tn[2] XThR.Tn[1] 0.28077f
C6020 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02698f
C6021 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06536f
C6022 XA.XIR[7].XIC[13].icell.PDM Iout 0.00112f
C6023 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PUM 0.00131f
C6024 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13469f
C6025 XThR.Tn[1] XA.XIR[2].XIC[0].icell.Ien 0.00321f
C6026 XA.XIR[13].XIC[3].icell.Ien VPWR 0.19065f
C6027 XA.XIR[10].XIC[2].icell.Ien Vbias 0.21238f
C6028 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02698f
C6029 XA.XIR[14].XIC_dummy_right.icell.SM VPWR 0.00123f
C6030 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.03424f
C6031 XA.XIR[7].XIC_15.icell.PDM Vbias 0.04206f
C6032 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04522f
C6033 XA.XIR[12].XIC[4].icell.Ien VPWR 0.19065f
C6034 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.15089f
C6035 XThR.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.00321f
C6036 XA.XIR[5].XIC[2].icell.PUM Vbias 0.00347f
C6037 XA.XIR[9].XIC_15.icell.SM Iout 0.0047f
C6038 XThC.XTB5.Y a_6243_9615# 0.00907f
C6039 XA.XIR[11].XIC[7].icell.PDM VPWR 0.00863f
C6040 XA.XIR[0].XIC[12].icell.SM Iout 0.00367f
C6041 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PUM 0.00131f
C6042 XA.XIR[4].XIC[5].icell.PDM Vbias 0.04058f
C6043 XThR.XTB5.Y XThR.Tn[7] 0.00912f
C6044 XThC.XTB7.A a_5155_9615# 0.02287f
C6045 XA.XIR[11].XIC[4].icell.PDM Iout 0.00112f
C6046 XA.XIR[10].XIC[6].icell.SM VPWR 0.00158f
C6047 XA.XIR[6].XIC[5].icell.PUM VPWR 0.01036f
C6048 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.SM 0.00383f
C6049 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13469f
C6050 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PUM 0.00529f
C6051 XA.XIR[0].XIC_15.icell.Ien Vbias 0.21351f
C6052 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.15089f
C6053 XA.XIR[3].XIC[5].icell.Ien Vbias 0.21238f
C6054 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PUM 0.00529f
C6055 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PUM 0.00131f
C6056 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Ien 0.00529f
C6057 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02698f
C6058 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.SM 0.00383f
C6059 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.03976f
C6060 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00212f
C6061 XA.XIR[10].XIC[3].icell.SM Iout 0.00388f
C6062 XA.XIR[5].XIC[8].icell.PDM VPWR 0.00863f
C6063 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.03424f
C6064 XA.XIR[2].XIC[7].icell.PUM Vbias 0.00347f
C6065 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.01406f
C6066 XThC.XTB2.Y a_7651_9569# 0.00191f
C6067 XA.XIR[5].XIC[5].icell.PDM Iout 0.00112f
C6068 XA.XIR[14].XIC[8].icell.PUM Vbias 0.00347f
C6069 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.SM 0.00383f
C6070 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PDM 0.00182f
C6071 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C6072 XA.XIR[4].XIC[8].icell.Ien VPWR 0.19065f
C6073 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00529f
C6074 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.01406f
C6075 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.04614f
C6076 XThR.Tn[7] XA.XIR[8].XIC[1].icell.Ien 0.00321f
C6077 XA.XIR[4].XIC[5].icell.Ien Iout 0.06483f
C6078 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04522f
C6079 XA.XIR[3].XIC[9].icell.SM VPWR 0.00158f
C6080 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PUM 0.00131f
C6081 XThC.Tn[14] VPWR 6.92099f
C6082 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00212f
C6083 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.SM 0.00188f
C6084 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.002f
C6085 XA.XIR[11].XIC[11].icell.PDM VPWR 0.00863f
C6086 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.01406f
C6087 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.15089f
C6088 XA.XIR[9].XIC[5].icell.SM Vbias 0.00701f
C6089 XA.XIR[8].XIC[4].icell.PUM VPWR 0.01036f
C6090 XA.XIR[3].XIC[6].icell.SM Iout 0.00388f
C6091 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.03976f
C6092 XThC.XTBN.Y a_6243_9615# 0.07731f
C6093 XThR.XTB2.Y data[4] 0.00267f
C6094 XA.XIR[2].XIC[13].icell.PDM VPWR 0.00863f
C6095 XA.XIR[15].XIC_15.icell.PDM Iout 0.0013f
C6096 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.03424f
C6097 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.03976f
C6098 XA.XIR[2].XIC[10].icell.PDM Iout 0.00112f
C6099 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Ien 0.00212f
C6100 XThC.Tn[1] XThR.Tn[4] 0.28062f
C6101 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.01406f
C6102 XA.XIR[9].XIC[0].icell.PDM VPWR 0.00863f
C6103 XA.XIR[14].XIC[10].icell.PUM VPWR 0.01036f
C6104 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00212f
C6105 XThR.Tn[1] XA.XIR[2].XIC[10].icell.SM 0.00121f
C6106 XThC.Tn[13] XThR.Tn[9] 0.28063f
C6107 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.SM 0.00383f
C6108 XA.XIR[13].XIC[0].icell.PDM Iout 0.00112f
C6109 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.04587f
C6110 XA.XIR[9].XIC[11].icell.PUM VPWR 0.01036f
C6111 XA.XIR[6].XIC[11].icell.PUM Vbias 0.00347f
C6112 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.01406f
C6113 XA.XIR[12].XIC_dummy_left.icell.SM VPWR 0.00269f
C6114 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02698f
C6115 XA.XIR[4].XIC[11].icell.SM VPWR 0.00158f
C6116 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C6117 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04522f
C6118 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08027f
C6119 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.03424f
C6120 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PUM 0.00131f
C6121 XA.XIR[7].XIC[3].icell.PUM Vbias 0.00347f
C6122 XThR.Tn[14] XA.XIR[15].XIC[4].icell.SM 0.00121f
C6123 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PUM 0.00209f
C6124 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PDM 0.00182f
C6125 XThR.Tn[3] XA.XIR[3].XIC[12].icell.PDM 0.0033f
C6126 XA.XIR[3].XIC[14].icell.PUM VPWR 0.01036f
C6127 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.01406f
C6128 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.03981f
C6129 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Ien 0.00217f
C6130 XA.XIR[1].XIC[4].icell.PUM Vbias 0.00347f
C6131 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01193f
C6132 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02698f
C6133 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00212f
C6134 XA.XIR[8].XIC[10].icell.PUM Vbias 0.00347f
C6135 XA.XIR[5].XIC[0].icell.PDM VPWR 0.00863f
C6136 XA.XIR[0].XIC[4].icell.Ien Vbias 0.21244f
C6137 XA.XIR[14].XIC[3].icell.PDM VPWR 0.00863f
C6138 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PUM 0.00131f
C6139 XA.XIR[7].XIC[9].icell.PDM VPWR 0.00863f
C6140 XA.XIR[2].XIC[12].icell.Ien Iout 0.06483f
C6141 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00529f
C6142 XA.XIR[2].XIC[0].icell.PDM Vbias 0.04002f
C6143 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.15089f
C6144 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.01406f
C6145 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00212f
C6146 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.SM 0.00188f
C6147 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02698f
C6148 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00529f
C6149 XA.XIR[7].XIC[6].icell.PDM Iout 0.00112f
C6150 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.15089f
C6151 XA.XIR[1].XIC[10].icell.PDM VPWR 0.00863f
C6152 XThR.Tn[4] XA.XIR[4].XIC[12].icell.PDM 0.0033f
C6153 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08017f
C6154 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.03424f
C6155 XThR.Tn[10] Vbias 3.71587f
C6156 XThC.Tn[11] XThR.Tn[11] 0.28062f
C6157 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.002f
C6158 XA.XIR[1].XIC_dummy_left.icell.Ien Vbias 0.00342f
C6159 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.01406f
C6160 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00529f
C6161 XThR.Tn[12] XA.XIR[13].XIC[3].icell.Ien 0.00321f
C6162 XA.XIR[1].XIC[7].icell.PDM Iout 0.00112f
C6163 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.SM 0.00383f
C6164 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04f
C6165 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00212f
C6166 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PUM 0.00536f
C6167 XA.XIR[0].XIC[8].icell.SM VPWR 0.00158f
C6168 XThR.Tn[14] XA.XIR[15].XIC[8].icell.SM 0.00121f
C6169 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00529f
C6170 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.15089f
C6171 XA.XIR[8].XIC[0].icell.PUM VPWR 0.01036f
C6172 XA.XIR[12].XIC[0].icell.SM Iout 0.00388f
C6173 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.03976f
C6174 XA.XIR[12].XIC[14].icell.Ien Iout 0.06483f
C6175 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.15089f
C6176 XA.XIR[4].XIC_dummy_left.icell.Ien Vbias 0.00342f
C6177 XThC.Tn[0] XA.XIR[7].XIC_dummy_left.icell.Iout 0.00111f
C6178 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.15089f
C6179 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.03424f
C6180 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02698f
C6181 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.03424f
C6182 XA.XIR[0].XIC[5].icell.SM Iout 0.00367f
C6183 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00529f
C6184 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C6185 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.01406f
C6186 XA.XIR[8].XIC[13].icell.PDM Iout 0.00112f
C6187 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.15089f
C6188 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00529f
C6189 XThR.Tn[8] XA.XIR[9].XIC_15.icell.Ien 0.00116f
C6190 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.03976f
C6191 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C6192 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.01406f
C6193 XA.XIR[8].XIC_15.icell.PDM Vbias 0.04206f
C6194 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PUM 0.00131f
C6195 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.01406f
C6196 XA.XIR[15].XIC[8].icell.PDM Vbias 0.04058f
C6197 XThR.Tn[10] XA.XIR[11].XIC[11].icell.SM 0.00121f
C6198 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C6199 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04f
C6200 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C6201 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8] 0.0033f
C6202 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C6203 XA.XIR[1].XIC[12].icell.Ien VPWR 0.19065f
C6204 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35783f
C6205 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.15089f
C6206 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.SM 0.00188f
C6207 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00212f
C6208 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C6209 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.01406f
C6210 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Iout 0.00347f
C6211 XThR.Tn[10] XA.XIR[11].XIC[8].icell.Ien 0.00321f
C6212 a_6243_10571# VPWR 0.00653f
C6213 XA.XIR[4].XIC[1].icell.Ien VPWR 0.19065f
C6214 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04522f
C6215 XThR.Tn[7] XThR.Tn[8] 0.08873f
C6216 XThC.XTB6.Y a_5949_9615# 0.26831f
C6217 XA.XIR[15].XIC[11].icell.SM Iout 0.00388f
C6218 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.SM 0.00383f
C6219 XThC.Tn[1] XThC.Tn[2] 0.72538f
C6220 XA.XIR[13].XIC[2].icell.Ien Vbias 0.21238f
C6221 XThC.Tn[0] XThC.Tn[3] 0.12427f
C6222 XThC.Tn[11] XThR.Tn[7] 0.28062f
C6223 XThR.Tn[5] XA.XIR[6].XIC[13].icell.Ien 0.00321f
C6224 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.03424f
C6225 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C6226 XA.XIR[3].XIC[2].icell.SM VPWR 0.00158f
C6227 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PUM 0.00131f
C6228 XThR.Tn[3] XA.XIR[3].XIC[1].icell.PDM 0.0033f
C6229 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.01406f
C6230 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02698f
C6231 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00212f
C6232 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.SM 0.00383f
C6233 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.03424f
C6234 XThC.Tn[14] XThR.Tn[12] 0.28068f
C6235 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Iout 0.00347f
C6236 XA.XIR[15].XIC[8].icell.Ien Iout 0.06816f
C6237 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00212f
C6238 XA.XIR[12].XIC[3].icell.Ien Vbias 0.21238f
C6239 XA.XIR[2].XIC[6].icell.PDM VPWR 0.00863f
C6240 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00212f
C6241 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.03976f
C6242 XThR.XTBN.A a_n997_2891# 0.01719f
C6243 XA.XIR[14].XIC[7].icell.PDM VPWR 0.00863f
C6244 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.01406f
C6245 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[2].icell.SM 0.00383f
C6246 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00212f
C6247 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.SM 0.00188f
C6248 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01734f
C6249 XA.XIR[11].XIC[6].icell.PDM Vbias 0.04058f
C6250 XA.XIR[2].XIC[3].icell.PDM Iout 0.00112f
C6251 XThC.XTB5.A XThC.XTB6.Y 0.00193f
C6252 XA.XIR[7].XIC_15.icell.Ien VPWR 0.25675f
C6253 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.SM 0.00188f
C6254 XA.XIR[14].XIC[4].icell.PDM Iout 0.00112f
C6255 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.03981f
C6256 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C6257 XA.XIR[13].XIC[6].icell.SM VPWR 0.00158f
C6258 XThR.Tn[1] XA.XIR[2].XIC[3].icell.SM 0.00121f
C6259 XThR.Tn[4] XA.XIR[4].XIC[1].icell.PDM 0.0033f
C6260 XA.XIR[10].XIC[5].icell.SM Vbias 0.00701f
C6261 XA.XIR[6].XIC[4].icell.PUM Vbias 0.00347f
C6262 XA.XIR[9].XIC[4].icell.PUM VPWR 0.01036f
C6263 XThR.Tn[10] XA.XIR[11].XIC[13].icell.Ien 0.00321f
C6264 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.SM 0.00383f
C6265 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06536f
C6266 XA.XIR[13].XIC[3].icell.SM Iout 0.00388f
C6267 XThR.Tn[9] XA.XIR[9].XIC[8].icell.PDM 0.0033f
C6268 XA.XIR[12].XIC[7].icell.SM VPWR 0.00158f
C6269 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PUM 0.00529f
C6270 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PUM 0.00131f
C6271 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PUM 0.00529f
C6272 XA.XIR[5].XIC[7].icell.PDM Vbias 0.04058f
C6273 a_4067_9615# VPWR 0.70649f
C6274 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.SM 0.00188f
C6275 XA.XIR[12].XIC[4].icell.SM Iout 0.00388f
C6276 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00212f
C6277 XThR.Tn[14] XA.XIR[15].XIC_15.icell.Ien 0.00116f
C6278 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.03976f
C6279 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.03534f
C6280 XThR.Tn[3] XA.XIR[3].XIC[5].icell.PDM 0.0033f
C6281 XA.XIR[7].XIC[0].icell.PDM Vbias 0.04002f
C6282 XThC.Tn[13] XThR.Tn[10] 0.28063f
C6283 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.SM 0.00383f
C6284 XA.XIR[4].XIC[7].icell.Ien Vbias 0.21238f
C6285 XA.XIR[15].XIC[13].icell.Ien Iout 0.06816f
C6286 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C6287 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C6288 XA.XIR[11].XIC[6].icell.Ien Iout 0.06483f
C6289 XA.XIR[6].XIC[10].icell.PDM VPWR 0.00863f
C6290 XThC.XTB4.Y a_5949_9615# 0.00465f
C6291 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C6292 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00529f
C6293 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PUM 0.00131f
C6294 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.03981f
C6295 XA.XIR[3].XIC[8].icell.SM Vbias 0.00701f
C6296 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.01406f
C6297 XA.XIR[14].XIC[11].icell.PDM VPWR 0.00863f
C6298 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08027f
C6299 XA.XIR[6].XIC[7].icell.PDM Iout 0.00112f
C6300 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.03424f
C6301 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00212f
C6302 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04522f
C6303 XA.XIR[8].XIC[3].icell.PUM Vbias 0.00347f
C6304 XA.XIR[7].XIC[2].icell.PDM VPWR 0.00863f
C6305 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04522f
C6306 XA.XIR[5].XIC[10].icell.Ien VPWR 0.19065f
C6307 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PUM 0.00131f
C6308 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02752f
C6309 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PUM 0.00529f
C6310 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.15089f
C6311 XA.XIR[2].XIC[12].icell.PDM Vbias 0.04058f
C6312 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.03424f
C6313 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PUM 0.00529f
C6314 XThC.XTB5.Y a_8963_9569# 0.00427f
C6315 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00529f
C6316 XA.XIR[1].XIC[3].icell.PDM VPWR 0.00863f
C6317 XA.XIR[5].XIC[7].icell.Ien Iout 0.06483f
C6318 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.11124f
C6319 XA.XIR[12].XIC[12].icell.SM VPWR 0.00158f
C6320 XThR.Tn[4] XA.XIR[4].XIC[5].icell.PDM 0.0033f
C6321 XThR.Tn[7] XA.XIR[8].XIC[4].icell.SM 0.00121f
C6322 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02698f
C6323 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.SM 0.00188f
C6324 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.0357f
C6325 XA.XIR[4].XIC[8].icell.SM Iout 0.00388f
C6326 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Ien 0.00529f
C6327 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.SM 0.00383f
C6328 XA.XIR[9].XIC[10].icell.PUM Vbias 0.00347f
C6329 XA.XIR[0].XIC[1].icell.SM VPWR 0.00158f
C6330 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C6331 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C6332 XA.XIR[8].XIC[9].icell.PDM VPWR 0.00863f
C6333 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PUM 0.00529f
C6334 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02698f
C6335 XA.XIR[12].XIC[8].icell.SM Iout 0.00388f
C6336 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.03976f
C6337 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.01406f
C6338 XThR.Tn[8] XA.XIR[9].XIC[11].icell.Ien 0.00321f
C6339 XA.XIR[8].XIC[6].icell.PDM Iout 0.00112f
C6340 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.SM 0.00383f
C6341 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.02035f
C6342 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.15089f
C6343 XA.XIR[6].XIC[12].icell.Ien VPWR 0.19065f
C6344 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.03424f
C6345 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.03504f
C6346 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06536f
C6347 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C6348 XA.XIR[3].XIC[13].icell.PUM Vbias 0.00347f
C6349 XA.XIR[11].XIC_15.icell.PDM Vbias 0.04206f
C6350 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04522f
C6351 XThC.XTB1.Y XThC.Tn[1] 0.01447f
C6352 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04522f
C6353 XA.XIR[5].XIC[13].icell.SM VPWR 0.00158f
C6354 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.SM 0.00383f
C6355 XA.XIR[9].XIC[1].icell.PDM VPWR 0.00863f
C6356 XA.XIR[2].XIC[14].icell.Ien Vbias 0.21238f
C6357 XThC.Tn[0] XA.XIR[8].XIC_dummy_left.icell.Iout 0.00111f
C6358 XThC.Tn[3] VPWR 5.96571f
C6359 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00529f
C6360 XThR.XTB6.Y a_n1049_5317# 0.01199f
C6361 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02698f
C6362 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02698f
C6363 XA.XIR[14].XIC[1].icell.PUM Vbias 0.00347f
C6364 XThC.XTBN.Y a_8963_9569# 0.22784f
C6365 XA.XIR[7].XIC[8].icell.PDM Vbias 0.04058f
C6366 XA.XIR[9].XIC[13].icell.PDM Iout 0.00112f
C6367 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.0277f
C6368 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02698f
C6369 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.SM 0.00383f
C6370 XThR.Tn[13] Vbias 3.71832f
C6371 XA.XIR[1].XIC[9].icell.PDM Vbias 0.04058f
C6372 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04522f
C6373 XThR.XTB5.A data[4] 0.14415f
C6374 XA.XIR[9].XIC_15.icell.PDM Vbias 0.04206f
C6375 XThC.Tn[11] XThR.Tn[14] 0.28062f
C6376 XThC.Tn[9] XThR.Tn[0] 0.28107f
C6377 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00529f
C6378 XA.XIR[15].XIC[4].icell.Ien VPWR 0.32782f
C6379 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.03544f
C6380 XThC.Tn[2] XThR.Tn[9] 0.28062f
C6381 XThR.Tn[8] XA.XIR[9].XIC[0].icell.Ien 0.00321f
C6382 XThR.XTB2.Y XThR.Tn[8] 0.00167f
C6383 XA.XIR[4].XIC[14].icell.SM Vbias 0.00701f
C6384 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.SM 0.00188f
C6385 XA.XIR[15].XIC[1].icell.Ien Iout 0.06816f
C6386 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.03981f
C6387 XA.XIR[0].XIC[7].icell.SM Vbias 0.00701f
C6388 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.03976f
C6389 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PUM 0.00529f
C6390 XA.XIR[7].XIC[11].icell.Ien VPWR 0.19065f
C6391 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PUM 0.00131f
C6392 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.01406f
C6393 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.SM 0.00383f
C6394 XA.XIR[5].XIC[0].icell.PUM VPWR 0.01036f
C6395 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.SM 0.00383f
C6396 XA.XIR[7].XIC[8].icell.Ien Iout 0.06483f
C6397 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.02698f
C6398 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.03976f
C6399 XA.XIR[2].XIC[1].icell.PDM Vbias 0.04058f
C6400 XA.XIR[11].XIC_15.icell.PUM Vbias 0.00347f
C6401 XA.XIR[5].XIC[14].icell.SM Iout 0.00388f
C6402 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.03424f
C6403 XThR.Tn[12] XA.XIR[13].XIC[6].icell.SM 0.00121f
C6404 XA.XIR[1].XIC[9].icell.Ien Iout 0.06483f
C6405 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.SM 0.00188f
C6406 XA.XIR[0].XIC[13].icell.PUM VPWR 0.00971f
C6407 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.SM 0.00383f
C6408 XA.XIR[9].XIC[2].icell.PDM Iout 0.00112f
C6409 XA.XIR[1].XIC[0].icell.Ien Vbias 0.21102f
C6410 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01746f
C6411 XThR.Tn[14] XA.XIR[15].XIC[9].icell.SM 0.00121f
C6412 XA.XIR[11].XIC[2].icell.Ien VPWR 0.19065f
C6413 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PUM 0.00529f
C6414 XThC.XTB2.Y a_5949_9615# 0.00844f
C6415 XThC.XTB7.B a_6243_10571# 0.00108f
C6416 XA.XIR[8].XIC_15.icell.Ien VPWR 0.25675f
C6417 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06536f
C6418 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PUM 0.00529f
C6419 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.SM 0.00188f
C6420 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02698f
C6421 XA.XIR[4].XIC[0].icell.Ien Vbias 0.21102f
C6422 XA.XIR[12].XIC_15.icell.Ien Iout 0.06485f
C6423 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04522f
C6424 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PUM 0.00529f
C6425 XThR.Tn[7] XA.XIR[7].XIC[14].icell.PDM 0.0033f
C6426 XA.XIR[10].XIC[4].icell.PUM VPWR 0.01036f
C6427 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11] 0.0033f
C6428 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.SM 0.00188f
C6429 XA.XIR[6].XIC[3].icell.PDM VPWR 0.00863f
C6430 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00529f
C6431 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.03976f
C6432 XThC.Tn[0] XThR.Tn[11] 0.28067f
C6433 data[5] data[4] 0.64735f
C6434 XA.XIR[3].XIC[1].icell.SM Vbias 0.00701f
C6435 XA.XIR[12].XIC[13].icell.PDM Iout 0.00112f
C6436 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PUM 0.00529f
C6437 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01702f
C6438 VPWR data[6] 0.21221f
C6439 XA.XIR[5].XIC[3].icell.Ien VPWR 0.19065f
C6440 XThR.XTB3.Y a_n1049_7493# 0.23056f
C6441 XA.XIR[7].XIC[11].icell.SM Iout 0.00388f
C6442 XA.XIR[2].XIC[5].icell.PDM Vbias 0.04058f
C6443 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PUM 0.00529f
C6444 XThR.XTBN.A a_n997_1579# 0.00199f
C6445 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C6446 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PUM 0.00529f
C6447 XA.XIR[14].XIC[6].icell.PDM Vbias 0.04058f
C6448 XA.XIR[4].XIC[4].icell.SM VPWR 0.00158f
C6449 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PUM 0.00529f
C6450 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.01406f
C6451 XA.XIR[1].XIC[12].icell.SM Iout 0.00388f
C6452 XA.XIR[13].XIC[5].icell.SM Vbias 0.00701f
C6453 XA.XIR[4].XIC[1].icell.SM Iout 0.00388f
C6454 XThR.Tn[1] a_n1049_7493# 0.00444f
C6455 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04522f
C6456 a_n997_3755# VPWR 0.0138f
C6457 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.03976f
C6458 XA.XIR[3].XIC[7].icell.PUM VPWR 0.01036f
C6459 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00529f
C6460 XA.XIR[9].XIC[3].icell.PUM Vbias 0.00347f
C6461 XA.XIR[1].XIC_15.icell.Ien Vbias 0.21343f
C6462 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.03424f
C6463 XThR.Tn[8] XA.XIR[9].XIC[4].icell.Ien 0.00321f
C6464 XA.XIR[11].XIC[11].icell.SM Vbias 0.00701f
C6465 XA.XIR[2].XIC[8].icell.Ien VPWR 0.19065f
C6466 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.01406f
C6467 XA.XIR[12].XIC[6].icell.SM Vbias 0.00701f
C6468 XThR.Tn[14] XA.XIR[15].XIC[11].icell.Ien 0.00321f
C6469 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C6470 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11175f
C6471 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00529f
C6472 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PDM 0.00182f
C6473 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PUM 0.00529f
C6474 XThC.XTB6.A XThC.Tn[9] 0.00838f
C6475 XA.XIR[11].XIC[8].icell.Ien Vbias 0.21238f
C6476 XA.XIR[2].XIC[5].icell.Ien Iout 0.06483f
C6477 XA.XIR[0].XIC_dummy_right.icell.Ien Vbias 0.003f
C6478 XThC.Tn[13] XThR.Tn[13] 0.28063f
C6479 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.0353f
C6480 XThC.XTB6.Y a_8739_9569# 0.00466f
C6481 XThC.XTB7.A XThC.Tn[4] 0.0274f
C6482 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02698f
C6483 XA.XIR[14].XIC[6].icell.Ien Iout 0.06483f
C6484 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PUM 0.00131f
C6485 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04522f
C6486 XA.XIR[7].XIC_dummy_right.icell.SM VPWR 0.00123f
C6487 XA.XIR[12].XIC[13].icell.PUM VPWR 0.01036f
C6488 XA.XIR[9].XIC[9].icell.PDM VPWR 0.00863f
C6489 XA.XIR[6].XIC[9].icell.PDM Vbias 0.04058f
C6490 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04522f
C6491 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.15089f
C6492 XThC.Tn[0] XThR.Tn[7] 0.28063f
C6493 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00212f
C6494 XThR.Tn[10] XA.XIR[11].XIC[0].icell.SM 0.00121f
C6495 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.03976f
C6496 XA.XIR[9].XIC[6].icell.PDM Iout 0.00112f
C6497 XThR.Tn[10] XA.XIR[11].XIC[14].icell.Ien 0.00321f
C6498 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04522f
C6499 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PUM 0.00131f
C6500 XA.XIR[5].XIC[9].icell.Ien Vbias 0.21238f
C6501 XThC.Tn[5] XThR.Tn[2] 0.28062f
C6502 XThR.XTB5.A XThR.XTB7.Y 0.00179f
C6503 XThC.Tn[3] XThR.Tn[12] 0.28062f
C6504 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.SM 0.00383f
C6505 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PUM 0.00529f
C6506 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.15089f
C6507 XThR.Tn[2] XA.XIR[3].XIC[8].icell.Ien 0.00321f
C6508 XA.XIR[4].XIC[10].icell.SM Vbias 0.00701f
C6509 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PUM 0.00529f
C6510 XThR.XTB1.Y a_n997_3979# 0.06353f
C6511 XA.XIR[2].XIC[11].icell.SM VPWR 0.00158f
C6512 XA.XIR[10].XIC[1].icell.PDM VPWR 0.00863f
C6513 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04522f
C6514 XThC.Tn[0] XA.XIR[9].XIC_dummy_left.icell.Iout 0.00111f
C6515 XA.XIR[15].XIC[14].icell.Ien Iout 0.06816f
C6516 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04522f
C6517 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C6518 XA.XIR[11].XIC[13].icell.Ien Vbias 0.21238f
C6519 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.03011f
C6520 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02698f
C6521 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00529f
C6522 XA.XIR[0].XIC[0].icell.SM Vbias 0.00675f
C6523 XA.XIR[6].XIC[9].icell.Ien Iout 0.06483f
C6524 XA.XIR[8].XIC[8].icell.PDM Vbias 0.04058f
C6525 XThC.Tn[2] XA.XIR[0].XIC[4].icell.Ien 0.00185f
C6526 XA.XIR[7].XIC[4].icell.Ien VPWR 0.19065f
C6527 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.03976f
C6528 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PUM 0.00209f
C6529 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38954f
C6530 XThR.Tn[6] Vbias 3.71582f
C6531 a_n1335_4229# data[4] 0.00451f
C6532 XA.XIR[1].XIC[5].icell.Ien VPWR 0.19065f
C6533 XA.XIR[5].XIC[10].icell.SM Iout 0.00388f
C6534 XA.XIR[7].XIC[1].icell.Ien Iout 0.06483f
C6535 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04522f
C6536 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.15089f
C6537 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PUM 0.00529f
C6538 XA.XIR[14].XIC_15.icell.PDM Vbias 0.04206f
C6539 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.SM 0.00383f
C6540 XThC.Tn[13] Vbias 2.35903f
C6541 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04522f
C6542 XThC.Tn[2] XThR.Tn[10] 0.28062f
C6543 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PUM 0.00131f
C6544 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PUM 0.00529f
C6545 XA.XIR[12].XIC[1].icell.PUM VPWR 0.01036f
C6546 XA.XIR[3].XIC[0].icell.PDM VPWR 0.00863f
C6547 XThR.XTB7.B XThR.XTBN.A 0.35142f
C6548 XA.XIR[12].XIC[13].icell.SM VPWR 0.00158f
C6549 XA.XIR[1].XIC[2].icell.Ien Iout 0.06483f
C6550 XThC.XTB7.B XThC.Tn[3] 0.00532f
C6551 XA.XIR[5].XIC[12].icell.SM Vbias 0.00701f
C6552 XThC.XTB4.Y a_8739_9569# 0.00813f
C6553 XA.XIR[0].XIC[6].icell.PUM VPWR 0.00971f
C6554 XA.XIR[8].XIC[11].icell.Ien VPWR 0.19065f
C6555 XThR.Tn[11] VPWR 7.66128f
C6556 XThR.Tn[5] XA.XIR[6].XIC[6].icell.Ien 0.00321f
C6557 XThC.XTB7.Y XThC.Tn[7] 0.0835f
C6558 XThR.Tn[2] XA.XIR[3].XIC[11].icell.SM 0.00121f
C6559 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.SM 0.00383f
C6560 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00529f
C6561 XThR.XTB7.B a_n1049_5317# 0.01743f
C6562 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.SM 0.00188f
C6563 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.01406f
C6564 XThC.XTB6.Y XThC.Tn[11] 0.02513f
C6565 XA.XIR[12].XIC[9].icell.SM Iout 0.00388f
C6566 XA.XIR[8].XIC[8].icell.Ien Iout 0.06483f
C6567 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.PDM 0.00576f
C6568 XThR.Tn[11] XA.XIR[12].XIC[2].icell.Ien 0.00321f
C6569 XThR.Tn[2] XA.XIR[2].XIC_15.icell.PDM 0.0033f
C6570 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00529f
C6571 XA.XIR[6].XIC[12].icell.SM Iout 0.00388f
C6572 XA.XIR[10].XIC[2].icell.PDM Iout 0.00112f
C6573 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PUM 0.00529f
C6574 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00212f
C6575 XA.XIR[15].XIC[3].icell.Ien Vbias 0.17911f
C6576 XThR.Tn[11] XA.XIR[11].XIC[5].icell.PDM 0.0033f
C6577 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.SM 0.00188f
C6578 XA.XIR[2].XIC_dummy_left.icell.Ien Vbias 0.00342f
C6579 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00212f
C6580 XThR.XTB6.Y a_n997_2891# 0.00466f
C6581 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.SM 0.00188f
C6582 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06536f
C6583 XThR.XTB2.Y a_n1049_5611# 0.00844f
C6584 XA.XIR[6].XIC_15.icell.Ien Vbias 0.21343f
C6585 XA.XIR[9].XIC_15.icell.Ien VPWR 0.25675f
C6586 XThR.Tn[10] XA.XIR[11].XIC[4].icell.SM 0.00121f
C6587 XA.XIR[7].XIC[10].icell.Ien Vbias 0.21238f
C6588 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C6589 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.SM 0.00188f
C6590 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04f
C6591 XThR.Tn[6] XA.XIR[6].XIC[9].icell.PDM 0.0033f
C6592 XA.XIR[14].XIC_15.icell.PUM Vbias 0.00347f
C6593 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PUM 0.00131f
C6594 XA.XIR[1].XIC[11].icell.Ien Vbias 0.21238f
C6595 XThR.Tn[10] XA.XIR[10].XIC[8].icell.PDM 0.0033f
C6596 XThR.XTBN.Y XA.XIR[6].XIC_dummy_left.icell.Ien 0.00159f
C6597 XThR.Tn[13] XA.XIR[14].XIC[11].icell.SM 0.00121f
C6598 XA.XIR[15].XIC[7].icell.SM VPWR 0.00158f
C6599 XA.XIR[8].XIC[2].icell.PDM VPWR 0.00863f
C6600 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.03424f
C6601 XA.XIR[8].XIC[11].icell.SM Iout 0.00388f
C6602 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.SM 0.00383f
C6603 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.01406f
C6604 XA.XIR[0].XIC[12].icell.PUM Vbias 0.00347f
C6605 XA.XIR[2].XIC[1].icell.Ien VPWR 0.19065f
C6606 XA.XIR[15].XIC[4].icell.SM Iout 0.00388f
C6607 XThR.Tn[13] XA.XIR[14].XIC[8].icell.Ien 0.00321f
C6608 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00529f
C6609 XA.XIR[14].XIC[2].icell.Ien VPWR 0.19119f
C6610 XA.XIR[12].XIC[11].icell.Ien Iout 0.06483f
C6611 XThR.Tn[7] VPWR 7.05634f
C6612 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.SM 0.00383f
C6613 XThR.Tn[0] XA.XIR[1].XIC[8].icell.Ien 0.00321f
C6614 XA.XIR[13].XIC[4].icell.PUM VPWR 0.01036f
C6615 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00212f
C6616 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PUM 0.00131f
C6617 XA.XIR[10].XIC[3].icell.PUM Vbias 0.00347f
C6618 XThC.XTB4.Y XThC.Tn[11] 0.30582f
C6619 XA.XIR[6].XIC[2].icell.PDM Vbias 0.04058f
C6620 XThC.Tn[0] XThR.Tn[14] 0.28065f
C6621 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C6622 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.15089f
C6623 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00529f
C6624 XA.XIR[7].XIC[13].icell.SM Vbias 0.00701f
C6625 XA.XIR[12].XIC[5].icell.PUM VPWR 0.01036f
C6626 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.03424f
C6627 XThR.Tn[10] XA.XIR[11].XIC[8].icell.SM 0.00121f
C6628 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.SM 0.00383f
C6629 XThC.Tn[7] XThR.Tn[0] 0.28143f
C6630 XA.XIR[5].XIC[2].icell.Ien Vbias 0.21238f
C6631 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.11124f
C6632 XThC.Tn[13] XThR.Tn[6] 0.28063f
C6633 XA.XIR[11].XIC[12].icell.PUM Vbias 0.00347f
C6634 XA.XIR[15].XIC[12].icell.SM VPWR 0.00158f
C6635 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.03424f
C6636 XA.XIR[11].XIC[5].icell.SM VPWR 0.00158f
C6637 XThR.XTB5.A XThR.Tn[8] 0.00204f
C6638 XThC.Tn[8] XThC.Tn[9] 0.05816f
C6639 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00529f
C6640 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.15119f
C6641 XThR.Tn[2] XA.XIR[3].XIC[1].icell.Ien 0.00321f
C6642 XA.XIR[4].XIC[3].icell.SM Vbias 0.00701f
C6643 XThC.XTB7.A a_6243_9615# 0.02018f
C6644 XThC.Tn[12] XThC.Tn[14] 0.03994f
C6645 XA.XIR[11].XIC[2].icell.SM Iout 0.00388f
C6646 XThR.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.00321f
C6647 XA.XIR[8].XIC_dummy_right.icell.SM VPWR 0.00123f
C6648 XA.XIR[10].XIC[9].icell.PDM VPWR 0.00863f
C6649 XA.XIR[6].XIC[5].icell.Ien VPWR 0.19065f
C6650 XA.XIR[15].XIC[8].icell.SM Iout 0.00388f
C6651 XThC.XTB7.A data[1] 0.06544f
C6652 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.03424f
C6653 XA.XIR[3].XIC[6].icell.PUM Vbias 0.00347f
C6654 XA.XIR[14].XIC[11].icell.SM Vbias 0.00701f
C6655 XA.XIR[10].XIC[6].icell.PDM Iout 0.00112f
C6656 XA.XIR[6].XIC[2].icell.Ien Iout 0.06483f
C6657 XA.XIR[5].XIC[6].icell.SM VPWR 0.00158f
C6658 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00212f
C6659 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.SM 0.00188f
C6660 XThC.XTBN.A Vbias 0.01573f
C6661 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35783f
C6662 XA.XIR[12].XIC[14].icell.PDM VPWR 0.00873f
C6663 XA.XIR[2].XIC[7].icell.Ien Vbias 0.21238f
C6664 XThR.Tn[0] XA.XIR[1].XIC[11].icell.SM 0.00121f
C6665 XA.XIR[5].XIC[3].icell.SM Iout 0.00388f
C6666 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.15107f
C6667 XA.XIR[14].XIC[8].icell.Ien Vbias 0.21238f
C6668 XA.XIR[4].XIC[9].icell.PUM VPWR 0.01036f
C6669 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Iout 0.00347f
C6670 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.01406f
C6671 XThR.Tn[3] Iout 1.1663f
C6672 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02698f
C6673 XA.XIR[12].XIC[9].icell.PUM VPWR 0.01036f
C6674 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PUM 0.00131f
C6675 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04522f
C6676 XThR.Tn[4] Vbias 3.71719f
C6677 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13469f
C6678 XA.XIR[3].XIC[12].icell.PDM VPWR 0.00863f
C6679 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.SM 0.00383f
C6680 XThR.Tn[6] XA.XIR[7].XIC[10].icell.Ien 0.00321f
C6681 XA.XIR[9].XIC[8].icell.PDM Vbias 0.04058f
C6682 XA.XIR[8].XIC[4].icell.Ien VPWR 0.19065f
C6683 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04522f
C6684 XThR.Tn[8] XA.XIR[9].XIC[7].icell.SM 0.00121f
C6685 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39047f
C6686 XA.XIR[3].XIC[9].icell.PDM Iout 0.00112f
C6687 XA.XIR[8].XIC[1].icell.Ien Iout 0.06483f
C6688 XThR.Tn[11] XThR.Tn[12] 0.12904f
C6689 XThC.Tn[14] XThR.Tn[1] 0.28068f
C6690 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04522f
C6691 XA.XIR[2].XIC[8].icell.SM Iout 0.00388f
C6692 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.SM 0.00188f
C6693 XThR.XTB7.B a_n1049_6405# 0.00268f
C6694 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00212f
C6695 XA.XIR[13].XIC[1].icell.PDM VPWR 0.00863f
C6696 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.03981f
C6697 XA.XIR[9].XIC[11].icell.Ien VPWR 0.19065f
C6698 XA.XIR[6].XIC[11].icell.Ien Vbias 0.21238f
C6699 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02698f
C6700 XA.XIR[14].XIC[13].icell.Ien Vbias 0.21238f
C6701 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C6702 XA.XIR[4].XIC[14].icell.PDM VPWR 0.00873f
C6703 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02698f
C6704 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08027f
C6705 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.SM 0.00383f
C6706 XA.XIR[9].XIC[8].icell.Ien Iout 0.06483f
C6707 XA.XIR[12].XIC[14].icell.PUM VPWR 0.01036f
C6708 XThR.Tn[3] XA.XIR[4].XIC[9].icell.Ien 0.00321f
C6709 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.03976f
C6710 XA.XIR[7].XIC[3].icell.Ien Vbias 0.21238f
C6711 XThR.Tn[6] XA.XIR[6].XIC[2].icell.PDM 0.0033f
C6712 XA.XIR[3].XIC[14].icell.Ien VPWR 0.1907f
C6713 XThR.XTBN.Y a_n1049_5317# 0.07731f
C6714 XThR.Tn[10] XA.XIR[11].XIC_15.icell.Ien 0.00116f
C6715 XThR.Tn[6] XA.XIR[7].XIC[13].icell.SM 0.00121f
C6716 XA.XIR[1].XIC[4].icell.Ien Vbias 0.21238f
C6717 XThC.Tn[2] XThR.Tn[13] 0.28062f
C6718 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04522f
C6719 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.01406f
C6720 XA.XIR[15].XIC[0].icell.SM VPWR 0.00158f
C6721 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.SM 0.00188f
C6722 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04522f
C6723 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PUM 0.00131f
C6724 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.04433f
C6725 XThR.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.0033f
C6726 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.03981f
C6727 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.SM 0.00188f
C6728 XThR.Tn[14] VPWR 7.88052f
C6729 XA.XIR[0].XIC[5].icell.PUM Vbias 0.00347f
C6730 XThC.Tn[4] XThR.Tn[3] 0.28062f
C6731 XThR.Tn[4] XA.XIR[5].XIC[9].icell.Ien 0.00321f
C6732 XA.XIR[8].XIC[10].icell.Ien Vbias 0.21238f
C6733 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.01406f
C6734 XA.XIR[7].XIC[7].icell.SM VPWR 0.00158f
C6735 XA.XIR[11].XIC[0].icell.SM Vbias 0.00675f
C6736 XA.XIR[11].XIC[14].icell.Ien Vbias 0.21238f
C6737 XA.XIR[15].XIC_15.icell.Ien Iout 0.06819f
C6738 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Iout 0.00347f
C6739 XA.XIR[10].XIC_15.icell.PDM Iout 0.0013f
C6740 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04522f
C6741 XA.XIR[1].XIC[8].icell.SM VPWR 0.00158f
C6742 XA.XIR[7].XIC[4].icell.SM Iout 0.00388f
C6743 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01776f
C6744 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.002f
C6745 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.01406f
C6746 XThR.Tn[0] XA.XIR[1].XIC[1].icell.Ien 0.00321f
C6747 XA.XIR[9].XIC[0].icell.Ien VPWR 0.19066f
C6748 XA.XIR[2].XIC[14].icell.SM Vbias 0.00701f
C6749 XThR.XTB2.Y VPWR 0.98816f
C6750 XA.XIR[15].XIC[13].icell.PDM Iout 0.00112f
C6751 XA.XIR[13].XIC[2].icell.PDM Iout 0.00112f
C6752 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00212f
C6753 XThR.Tn[3] XA.XIR[4].XIC[12].icell.SM 0.00121f
C6754 XA.XIR[1].XIC[5].icell.SM Iout 0.00388f
C6755 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PUM 0.00529f
C6756 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PUM 0.00131f
C6757 XA.XIR[9].XIC[11].icell.SM Iout 0.00388f
C6758 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.03976f
C6759 XThR.XTB6.Y a_n997_1579# 0.07626f
C6760 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.03429f
C6761 XA.XIR[0].XIC[11].icell.PDM VPWR 0.00806f
C6762 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04522f
C6763 XThR.Tn[1] XA.XIR[1].XIC[10].icell.PDM 0.0033f
C6764 XA.XIR[3].XIC[1].icell.PDM VPWR 0.00863f
C6765 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PUM 0.00131f
C6766 XA.XIR[12].XIC[3].icell.PDM Iout 0.00112f
C6767 XThR.Tn[5] XA.XIR[6].XIC[9].icell.SM 0.00121f
C6768 XA.XIR[12].XIC[14].icell.SM VPWR 0.00208f
C6769 XThC.Tn[0] XA.XIR[2].XIC_dummy_left.icell.Iout 0.00111f
C6770 XThC.XTB5.A data[1] 0.11102f
C6771 XThR.XTB7.B a_n997_2891# 0.0168f
C6772 XThC.XTB6.A a_5949_10571# 0.00467f
C6773 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.01406f
C6774 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00529f
C6775 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01763f
C6776 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00529f
C6777 XA.XIR[3].XIC_15.icell.Ien Iout 0.06485f
C6778 XThC.XTB3.Y Vbias 0.01151f
C6779 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[12].icell.Ien 0.00212f
C6780 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.SM 0.00188f
C6781 XA.XIR[4].XIC_15.icell.SM Vbias 0.00701f
C6782 XThR.Tn[11] XA.XIR[12].XIC[5].icell.SM 0.00121f
C6783 XThC.Tn[13] XThR.Tn[4] 0.28063f
C6784 XThR.Tn[9] XA.XIR[10].XIC[3].icell.Ien 0.00321f
C6785 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04522f
C6786 XThR.Tn[4] XA.XIR[5].XIC[12].icell.SM 0.00121f
C6787 XA.XIR[8].XIC[13].icell.SM Vbias 0.00701f
C6788 XA.XIR[15].XIC[6].icell.SM Vbias 0.00701f
C6789 XThC.Tn[2] Vbias 2.4654f
C6790 XA.XIR[7].XIC[12].icell.PUM VPWR 0.01036f
C6791 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.15089f
C6792 XA.XIR[5].XIC[2].icell.PDM VPWR 0.00863f
C6793 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.01406f
C6794 XA.XIR[1].XIC[13].icell.PUM VPWR 0.01036f
C6795 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.01406f
C6796 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PUM 0.00529f
C6797 XA.XIR[2].XIC[0].icell.Ien Vbias 0.21102f
C6798 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.03424f
C6799 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.0353f
C6800 VPWR data[2] 0.21031f
C6801 XA.XIR[4].XIC[2].icell.PUM VPWR 0.01036f
C6802 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04522f
C6803 XThR.Tn[12] XA.XIR[12].XIC[14].icell.PDM 0.0033f
C6804 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.15089f
C6805 XA.XIR[5].XIC_15.icell.SM Iout 0.0047f
C6806 XA.XIR[9].XIC_dummy_right.icell.SM VPWR 0.00123f
C6807 XThC.XTB5.Y XThC.Tn[5] 0.01095f
C6808 a_10915_9569# XThC.Tn[14] 0.20278f
C6809 XA.XIR[15].XIC[13].icell.PUM VPWR 0.01036f
C6810 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.01406f
C6811 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00212f
C6812 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.15089f
C6813 XA.XIR[3].XIC[5].icell.PDM VPWR 0.00863f
C6814 XA.XIR[13].XIC[3].icell.PUM Vbias 0.00347f
C6815 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PUM 0.00131f
C6816 XThR.Tn[6] XA.XIR[7].XIC[3].icell.Ien 0.00321f
C6817 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Iout 0.00347f
C6818 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.03424f
C6819 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35783f
C6820 XA.XIR[12].XIC[4].icell.PUM Vbias 0.00347f
C6821 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PUM 0.00529f
C6822 XThR.Tn[8] Iout 1.16627f
C6823 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00529f
C6824 XA.XIR[2].XIC[4].icell.SM VPWR 0.00158f
C6825 XA.XIR[3].XIC[2].icell.PDM Iout 0.00112f
C6826 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.SM 0.00188f
C6827 XThC.XTB2.Y data[0] 0.00267f
C6828 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.01406f
C6829 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02698f
C6830 XA.XIR[14].XIC[5].icell.SM VPWR 0.00158f
C6831 XA.XIR[14].XIC[12].icell.PUM Vbias 0.00347f
C6832 XA.XIR[11].XIC[4].icell.SM Vbias 0.00701f
C6833 XThC.Tn[11] Iout 0.84418f
C6834 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04522f
C6835 XA.XIR[2].XIC[1].icell.SM Iout 0.00388f
C6836 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.0353f
C6837 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.SM 0.00188f
C6838 XA.XIR[12].XIC[12].icell.Ien VPWR 0.19065f
C6839 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00212f
C6840 XA.XIR[13].XIC[9].icell.PDM VPWR 0.00863f
C6841 XA.XIR[14].XIC[2].icell.SM Iout 0.00388f
C6842 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04522f
C6843 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.03976f
C6844 XA.XIR[10].XIC[8].icell.PDM Vbias 0.04058f
C6845 XA.XIR[6].XIC[4].icell.Ien Vbias 0.21238f
C6846 XA.XIR[9].XIC[4].icell.Ien VPWR 0.19065f
C6847 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.03424f
C6848 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.03976f
C6849 XA.XIR[13].XIC[6].icell.PDM Iout 0.00112f
C6850 XA.XIR[12].XIC[10].icell.PDM VPWR 0.00863f
C6851 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.01406f
C6852 XThR.Tn[3] XA.XIR[4].XIC[2].icell.Ien 0.00321f
C6853 XThR.Tn[0] XA.XIR[0].XIC[14].icell.PDM 0.0033f
C6854 XA.XIR[5].XIC[5].icell.SM Vbias 0.00701f
C6855 XThR.Tn[10] XA.XIR[11].XIC[9].icell.SM 0.00121f
C6856 a_5155_9615# VPWR 0.7051f
C6857 XA.XIR[12].XIC[7].icell.PDM Iout 0.00112f
C6858 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.SM 0.00383f
C6859 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04522f
C6860 XThC.XTBN.Y XThC.Tn[5] 0.60785f
C6861 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C6862 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C6863 XThR.Tn[2] XA.XIR[3].XIC[4].icell.SM 0.00121f
C6864 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01799f
C6865 XA.XIR[4].XIC[8].icell.PUM Vbias 0.00347f
C6866 XA.XIR[1].XIC_dummy_right.icell.Ien Vbias 0.00287f
C6867 XA.XIR[10].XIC[11].icell.SM Iout 0.00388f
C6868 XA.XIR[15].XIC[13].icell.SM VPWR 0.00158f
C6869 XA.XIR[6].XIC[8].icell.SM VPWR 0.00158f
C6870 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00212f
C6871 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.SM 0.00188f
C6872 XThR.XTBN.Y a_n1049_6405# 0.07602f
C6873 XThR.Tn[2] XA.XIR[2].XIC[8].icell.PDM 0.0033f
C6874 XA.XIR[15].XIC[0].icell.PDM Vbias 0.04002f
C6875 XThR.Tn[13] XA.XIR[14].XIC[0].icell.SM 0.00127f
C6876 XA.XIR[3].XIC[11].icell.PDM Vbias 0.04058f
C6877 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02698f
C6878 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.SM 0.00188f
C6879 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00212f
C6880 XA.XIR[10].XIC[8].icell.Ien Iout 0.06483f
C6881 XThR.Tn[13] XA.XIR[14].XIC[14].icell.Ien 0.00321f
C6882 XA.XIR[11].XIC[8].icell.SM Vbias 0.00701f
C6883 XA.XIR[15].XIC[9].icell.SM Iout 0.00388f
C6884 XA.XIR[6].XIC[5].icell.SM Iout 0.00388f
C6885 XA.XIR[8].XIC[3].icell.Ien Vbias 0.21238f
C6886 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39045f
C6887 XThR.Tn[4] XA.XIR[5].XIC[2].icell.Ien 0.00321f
C6888 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PUM 0.00529f
C6889 XA.XIR[5].XIC[11].icell.PUM VPWR 0.01036f
C6890 XA.XIR[7].XIC[0].icell.SM VPWR 0.00158f
C6891 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.SM 0.00383f
C6892 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.03424f
C6893 XA.XIR[2].XIC[10].icell.SM Vbias 0.00701f
C6894 XThR.XTBN.Y XA.XIR[7].XIC_dummy_left.icell.Ien 0.00158f
C6895 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.03424f
C6896 XThR.Tn[0] XThR.Tn[2] 0.00536f
C6897 XThC.XTB5.Y a_10051_9569# 0.00133f
C6898 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.SM 0.00188f
C6899 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00212f
C6900 XThC.Tn[2] XThR.Tn[6] 0.28062f
C6901 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.SM 0.00188f
C6902 XA.XIR[1].XIC[1].icell.SM VPWR 0.00158f
C6903 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00212f
C6904 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00212f
C6905 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.11124f
C6906 XThC.Tn[4] XThR.Tn[8] 0.28062f
C6907 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.01406f
C6908 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00212f
C6909 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04522f
C6910 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C6911 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00529f
C6912 a_9827_9569# XA.XIR[0].XIC[11].icell.PDM 0.00127f
C6913 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.03976f
C6914 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00212f
C6915 XA.XIR[4].XIC[11].icell.PDM Iout 0.00112f
C6916 XThC.Tn[7] XThC.Tn[8] 0.08099f
C6917 XThC.XTB1.Y Vbias 0.0117f
C6918 XA.XIR[9].XIC[10].icell.Ien Vbias 0.21238f
C6919 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.03425f
C6920 XA.XIR[0].XIC[4].icell.PDM VPWR 0.00809f
C6921 XA.XIR[8].XIC[7].icell.SM VPWR 0.00158f
C6922 XA.XIR[12].XIC[11].icell.PDM Iout 0.00112f
C6923 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04522f
C6924 XThR.Tn[1] XA.XIR[1].XIC[3].icell.PDM 0.0033f
C6925 XThR.Tn[5] XA.XIR[6].XIC[2].icell.SM 0.00121f
C6926 XThR.XTB4.Y a_n1049_5317# 0.00463f
C6927 XA.XIR[3].XIC[11].icell.Ien Iout 0.06483f
C6928 XA.XIR[12].XIC[1].icell.PDM Vbias 0.04058f
C6929 a_4861_9615# XThC.Tn[5] 0.00208f
C6930 XThR.Tn[10] XA.XIR[11].XIC[11].icell.Ien 0.00321f
C6931 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00529f
C6932 XA.XIR[8].XIC[4].icell.SM Iout 0.00388f
C6933 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06536f
C6934 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02698f
C6935 XA.XIR[10].XIC[0].icell.Ien VPWR 0.19066f
C6936 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PUM 0.00529f
C6937 XA.XIR[6].XIC[13].icell.PUM VPWR 0.01036f
C6938 XA.XIR[10].XIC[13].icell.Ien Iout 0.06483f
C6939 XA.XIR[3].XIC[13].icell.Ien Vbias 0.21238f
C6940 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02698f
C6941 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.SM 0.00383f
C6942 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08017f
C6943 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.SM 0.00383f
C6944 XThC.XTB6.Y VPWR 1.03149f
C6945 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04522f
C6946 XThC.Tn[5] XThR.Tn[5] 0.28062f
C6947 XA.XIR[9].XIC_dummy_left.icell.SM VPWR 0.00269f
C6948 XA.XIR[15].XIC[11].icell.Ien Iout 0.06816f
C6949 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.SM 0.00383f
C6950 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.SM 0.00383f
C6951 XThC.XTBN.Y a_10051_9569# 0.23006f
C6952 XA.XIR[14].XIC[0].icell.SM Vbias 0.00675f
C6953 XA.XIR[13].XIC_15.icell.PDM Iout 0.0013f
C6954 XA.XIR[14].XIC[14].icell.Ien Vbias 0.21238f
C6955 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.SM 0.00188f
C6956 XA.XIR[7].XIC[6].icell.SM Vbias 0.00701f
C6957 XThR.XTBN.Y a_n997_2891# 0.22804f
C6958 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04522f
C6959 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00212f
C6960 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00529f
C6961 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.39042f
C6962 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.15089f
C6963 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PUM 0.00529f
C6964 XA.XIR[4].XIC[13].icell.Ien Iout 0.06483f
C6965 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.15089f
C6966 XA.XIR[1].XIC[7].icell.SM Vbias 0.00701f
C6967 XThC.Tn[3] XThR.Tn[1] 0.28062f
C6968 XA.XIR[9].XIC[13].icell.SM Vbias 0.00701f
C6969 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00529f
C6970 XA.XIR[15].XIC[5].icell.PUM VPWR 0.01036f
C6971 XA.XIR[8].XIC[12].icell.PUM VPWR 0.01036f
C6972 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.SM 0.00188f
C6973 XThR.Tn[14] XA.XIR[14].XIC[5].icell.PDM 0.0033f
C6974 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.SM 0.00188f
C6975 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PUM 0.00131f
C6976 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.15089f
C6977 XA.XIR[4].XIC_dummy_right.icell.PUM Vbias 0.00248f
C6978 XA.XIR[12].XIC[10].icell.SM VPWR 0.00158f
C6979 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02698f
C6980 XA.XIR[0].XIC[10].icell.PDM Vbias 0.04065f
C6981 XThR.Tn[13] XA.XIR[14].XIC[4].icell.SM 0.00121f
C6982 XThR.XTB7.B a_n997_1579# 0.00209f
C6983 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11595f
C6984 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.03424f
C6985 XThR.Tn[13] XA.XIR[13].XIC[8].icell.PDM 0.0033f
C6986 XThR.Tn[0] XA.XIR[1].XIC[4].icell.SM 0.00121f
C6987 XA.XIR[11].XIC_15.icell.Ien Vbias 0.21343f
C6988 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Iout 0.00347f
C6989 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PUM 0.00529f
C6990 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.15089f
C6991 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35783f
C6992 XA.XIR[6].XIC_dummy_right.icell.Ien Vbias 0.00287f
C6993 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.03976f
C6994 XA.XIR[9].XIC[0].icell.SM Iout 0.00388f
C6995 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01203f
C6996 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02698f
C6997 XThR.Tn[0] XA.XIR[0].XIC[7].icell.PDM 0.0033f
C6998 XA.XIR[0].XIC[13].icell.Ien VPWR 0.19003f
C6999 XA.XIR[1].XIC[1].icell.PUM Vbias 0.00347f
C7000 XA.XIR[11].XIC[13].icell.PDM Vbias 0.04058f
C7001 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00529f
C7002 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02698f
C7003 XThC.XTB7.B data[2] 0.07481f
C7004 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.03424f
C7005 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06536f
C7006 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04522f
C7007 XThC.XTB4.Y VPWR 0.91505f
C7008 XThR.Tn[12] XA.XIR[12].XIC[10].icell.PDM 0.0033f
C7009 XA.XIR[1].XIC[12].icell.PUM Vbias 0.00347f
C7010 XA.XIR[0].XIC[10].icell.Ien Iout 0.06455f
C7011 XA.XIR[11].XIC[3].icell.PUM VPWR 0.01036f
C7012 XThC.XTB2.Y XThC.Tn[0] 0.00125f
C7013 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.03424f
C7014 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.01406f
C7015 XThR.XTB6.A a_n997_3755# 0.00149f
C7016 XA.XIR[15].XIC[9].icell.PUM VPWR 0.01036f
C7017 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00529f
C7018 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PUM 0.00529f
C7019 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.03424f
C7020 XA.XIR[4].XIC[1].icell.PUM Vbias 0.00347f
C7021 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.03424f
C7022 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[13].icell.SM 0.00383f
C7023 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.01406f
C7024 XA.XIR[10].XIC[4].icell.Ien VPWR 0.19065f
C7025 XThR.Tn[9] XA.XIR[10].XIC[6].icell.SM 0.00121f
C7026 XA.XIR[6].XIC[1].icell.SM VPWR 0.00158f
C7027 XThR.Tn[13] XA.XIR[14].XIC[8].icell.SM 0.00121f
C7028 XA.XIR[3].XIC[4].icell.PDM Vbias 0.04058f
C7029 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C7030 XA.XIR[5].XIC[4].icell.PUM VPWR 0.01036f
C7031 XThR.XTB5.A VPWR 0.83112f
C7032 XA.XIR[7].XIC[14].icell.PDM Iout 0.00112f
C7033 XA.XIR[2].XIC[3].icell.SM Vbias 0.00701f
C7034 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.03424f
C7035 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Ien 0.00586f
C7036 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00529f
C7037 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00529f
C7038 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.SM 0.00188f
C7039 XA.XIR[14].XIC[4].icell.SM Vbias 0.00701f
C7040 XA.XIR[4].XIC[7].icell.PDM VPWR 0.00863f
C7041 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.03424f
C7042 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.03424f
C7043 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PUM 0.00131f
C7044 XA.XIR[1].XIC_15.icell.PDM Iout 0.0013f
C7045 XA.XIR[7].XIC_15.icell.PUM Vbias 0.00347f
C7046 XA.XIR[13].XIC[8].icell.PDM Vbias 0.04058f
C7047 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.SM 0.00188f
C7048 XThR.XTB3.Y a_n997_3755# 0.0061f
C7049 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00212f
C7050 XA.XIR[6].XIC[0].icell.PDM VPWR 0.00863f
C7051 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C7052 XA.XIR[3].XIC[7].icell.Ien VPWR 0.19065f
C7053 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.SM 0.00383f
C7054 XA.XIR[4].XIC[4].icell.PDM Iout 0.00112f
C7055 XThC.Tn[2] XThR.Tn[4] 0.28062f
C7056 XThR.Tn[6] XA.XIR[7].XIC[6].icell.SM 0.00121f
C7057 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04522f
C7058 XA.XIR[15].XIC[14].icell.PUM VPWR 0.01036f
C7059 XA.XIR[9].XIC[3].icell.Ien Vbias 0.21238f
C7060 XThC.Tn[14] XThR.Tn[9] 0.28068f
C7061 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.SM 0.00383f
C7062 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14] 0.0033f
C7063 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Iout 0.00347f
C7064 XA.XIR[8].XIC[0].icell.SM VPWR 0.00158f
C7065 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02698f
C7066 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00212f
C7067 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.SM 0.00188f
C7068 XA.XIR[12].XIC[9].icell.PDM Vbias 0.04058f
C7069 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PUM 0.00131f
C7070 XA.XIR[2].XIC[9].icell.PUM VPWR 0.01036f
C7071 XThC.XTB7.B a_5155_9615# 0.00268f
C7072 XA.XIR[3].XIC[4].icell.Ien Iout 0.06483f
C7073 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00529f
C7074 a_2979_9615# Vbias 0.00694f
C7075 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.03424f
C7076 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.SM 0.00188f
C7077 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.03424f
C7078 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01872f
C7079 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[5].icell.Ien 0.00212f
C7080 XThR.XTB4.Y a_n1049_6405# 0.01546f
C7081 XThC.XTB6.Y a_9827_9569# 0.00871f
C7082 XA.XIR[13].XIC[11].icell.SM Iout 0.00388f
C7083 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11] 0.0033f
C7084 XThR.Tn[1] XA.XIR[2].XIC[8].icell.Ien 0.00321f
C7085 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9] 0.0033f
C7086 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.SM 0.00383f
C7087 XA.XIR[6].XIC[7].icell.SM Vbias 0.00701f
C7088 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.SM 0.00383f
C7089 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02698f
C7090 XA.XIR[9].XIC[7].icell.SM VPWR 0.00158f
C7091 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00529f
C7092 XA.XIR[13].XIC[8].icell.Ien Iout 0.06483f
C7093 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.03976f
C7094 XA.XIR[14].XIC[8].icell.SM Vbias 0.00701f
C7095 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02698f
C7096 XThR.XTB7.A XThR.XTBN.A 0.19736f
C7097 XThR.Tn[3] XA.XIR[4].XIC[5].icell.SM 0.00121f
C7098 XA.XIR[9].XIC[4].icell.SM Iout 0.00388f
C7099 a_4067_9615# XThC.Tn[1] 0.00584f
C7100 XThR.Tn[14] XA.XIR[15].XIC[2].icell.Ien 0.00321f
C7101 XA.XIR[5].XIC[10].icell.PUM Vbias 0.00347f
C7102 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02698f
C7103 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04522f
C7104 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.01406f
C7105 VPWR data[5] 0.4402f
C7106 XA.XIR[11].XIC[0].icell.PDM Iout 0.00112f
C7107 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.03424f
C7108 XA.XIR[1].XIC[0].icell.SM Vbias 0.00675f
C7109 XA.XIR[12].XIC_dummy_left.icell.Ien Vbias 0.00342f
C7110 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PUM 0.00131f
C7111 XThR.XTB7.A a_n1049_5317# 0.02018f
C7112 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PUM 0.00529f
C7113 XA.XIR[4].XIC[13].icell.PDM Vbias 0.04058f
C7114 XThC.Tn[0] Iout 0.82722f
C7115 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.03424f
C7116 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.SM 0.00383f
C7117 XA.XIR[2].XIC[14].icell.PDM VPWR 0.00873f
C7118 XA.XIR[10].XIC_dummy_left.icell.SM VPWR 0.00269f
C7119 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.15089f
C7120 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.15089f
C7121 XA.XIR[15].XIC[14].icell.SM VPWR 0.00208f
C7122 XThC.Tn[12] XThR.Tn[11] 0.28062f
C7123 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02698f
C7124 XA.XIR[0].XIC[3].icell.PDM Vbias 0.04065f
C7125 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00529f
C7126 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.SM 0.00383f
C7127 XA.XIR[8].XIC[6].icell.SM Vbias 0.00701f
C7128 XThR.Tn[4] XA.XIR[5].XIC[5].icell.SM 0.00121f
C7129 XA.XIR[7].XIC[5].icell.PUM VPWR 0.01036f
C7130 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02698f
C7131 XThR.Tn[8] XA.XIR[8].XIC[10].icell.PDM 0.0033f
C7132 a_7875_9569# VPWR 0.00643f
C7133 XThR.Tn[13] XA.XIR[14].XIC_15.icell.Ien 0.00116f
C7134 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02698f
C7135 XA.XIR[11].XIC[9].icell.SM Vbias 0.00701f
C7136 XA.XIR[13].XIC[0].icell.Ien VPWR 0.19066f
C7137 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.SM 0.00383f
C7138 XThR.Tn[1] XA.XIR[2].XIC[11].icell.SM 0.00121f
C7139 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.01406f
C7140 XA.XIR[5].XIC[13].icell.PDM Iout 0.00112f
C7141 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.03424f
C7142 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.SM 0.00383f
C7143 XA.XIR[1].XIC[6].icell.PUM VPWR 0.01036f
C7144 XA.XIR[13].XIC[13].icell.Ien Iout 0.06483f
C7145 XA.XIR[6].XIC[12].icell.PUM Vbias 0.00347f
C7146 XA.XIR[9].XIC[12].icell.PUM VPWR 0.01036f
C7147 XThC.XTB2.Y VPWR 0.97669f
C7148 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C7149 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.SM 0.00383f
C7150 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C7151 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.03981f
C7152 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.03424f
C7153 XA.XIR[12].XIC[1].icell.Ien VPWR 0.19065f
C7154 XThR.Tn[7] XA.XIR[8].XIC[9].icell.Ien 0.00321f
C7155 XA.XIR[5].XIC_15.icell.PDM Vbias 0.04206f
C7156 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00212f
C7157 XA.XIR[0].XIC[6].icell.Ien VPWR 0.1901f
C7158 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.SM 0.00188f
C7159 XThR.XTB4.Y a_n997_2891# 0.00813f
C7160 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.15089f
C7161 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PUM 0.00131f
C7162 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11595f
C7163 XA.XIR[3].XIC[14].icell.SM VPWR 0.00208f
C7164 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.SM 0.00383f
C7165 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00212f
C7166 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02698f
C7167 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PUM 0.00209f
C7168 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04f
C7169 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.SM 0.00188f
C7170 XA.XIR[12].XIC[11].icell.PUM VPWR 0.01036f
C7171 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C7172 XA.XIR[0].XIC[3].icell.Ien Iout 0.06455f
C7173 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00212f
C7174 XThR.XTBN.Y a_n997_1579# 0.23006f
C7175 XThR.Tn[5] XA.XIR[5].XIC[10].icell.PDM 0.0033f
C7176 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02698f
C7177 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PUM 0.00131f
C7178 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.01406f
C7179 XThC.XTB3.Y XThC.Tn[2] 0.1864f
C7180 XA.XIR[10].XIC[0].icell.SM Iout 0.00388f
C7181 XA.XIR[6].XIC_15.icell.PDM Iout 0.0013f
C7182 XA.XIR[15].XIC[4].icell.PUM Vbias 0.00347f
C7183 XA.XIR[10].XIC[14].icell.Ien Iout 0.06483f
C7184 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.03424f
C7185 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02698f
C7186 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.15089f
C7187 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.03424f
C7188 XThC.Tn[1] XThC.Tn[3] 0.10977f
C7189 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.01406f
C7190 XThC.Tn[8] XThR.Tn[2] 0.28062f
C7191 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PUM 0.00529f
C7192 data[1] data[0] 0.64735f
C7193 XThC.Tn[12] XThR.Tn[7] 0.28062f
C7194 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04522f
C7195 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.03976f
C7196 XA.XIR[2].XIC_15.icell.SM Vbias 0.00701f
C7197 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.02226f
C7198 XThC.Tn[6] XThC.Tn[7] 0.16385f
C7199 XA.XIR[7].XIC[11].icell.PUM Vbias 0.00347f
C7200 XA.XIR[15].XIC[12].icell.Ien VPWR 0.32782f
C7201 XA.XIR[11].XIC[11].icell.Ien Vbias 0.21238f
C7202 XThR.Tn[7] XA.XIR[8].XIC[12].icell.SM 0.00121f
C7203 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C7204 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00529f
C7205 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02698f
C7206 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04522f
C7207 XA.XIR[14].XIC_15.icell.Ien Vbias 0.21343f
C7208 Vbias bias[2] 0.05684f
C7209 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01193f
C7210 XA.XIR[3].XIC[0].icell.Ien VPWR 0.19066f
C7211 a_n1335_4229# VPWR 0.00633f
C7212 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.15089f
C7213 XA.XIR[12].XIC_15.icell.SM VPWR 0.00276f
C7214 XA.XIR[14].XIC[13].icell.PDM Vbias 0.04058f
C7215 XA.XIR[8].XIC[14].icell.PDM Iout 0.00112f
C7216 XA.XIR[15].XIC[7].icell.PDM Iout 0.00112f
C7217 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C7218 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.15089f
C7219 XA.XIR[0].XIC[12].icell.Ien Vbias 0.21246f
C7220 XA.XIR[2].XIC[2].icell.PUM VPWR 0.01036f
C7221 XThR.XTB3.Y XThR.Tn[7] 0.00819f
C7222 XA.XIR[14].XIC[3].icell.PUM VPWR 0.01036f
C7223 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04522f
C7224 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02698f
C7225 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.SM 0.00188f
C7226 XA.XIR[8].XIC_15.icell.PUM Vbias 0.00347f
C7227 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00212f
C7228 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02698f
C7229 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PUM 0.00131f
C7230 XA.XIR[13].XIC[4].icell.Ien VPWR 0.19065f
C7231 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.SM 0.00383f
C7232 XThR.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.00321f
C7233 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PUM 0.00198f
C7234 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00212f
C7235 XThC.Tn[14] XThR.Tn[10] 0.28068f
C7236 XA.XIR[10].XIC[3].icell.Ien Vbias 0.21238f
C7237 XA.XIR[6].XIC[0].icell.SM Vbias 0.00675f
C7238 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04522f
C7239 XThC.XTB7.Y XThC.Tn[10] 0.07406f
C7240 VPWR Iout 54.3441f
C7241 a_n1049_5611# XA.XIR[5].XIC_dummy_left.icell.Iout 0.001f
C7242 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.03976f
C7243 XA.XIR[12].XIC[5].icell.Ien VPWR 0.19065f
C7244 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08027f
C7245 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.15089f
C7246 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00529f
C7247 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.SM 0.00188f
C7248 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.SM 0.00383f
C7249 XA.XIR[5].XIC[3].icell.PUM Vbias 0.00347f
C7250 XA.XIR[12].XIC[2].icell.Ien Iout 0.06483f
C7251 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04522f
C7252 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01402f
C7253 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C7254 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C7255 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06536f
C7256 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00529f
C7257 XA.XIR[11].XIC[8].icell.PDM VPWR 0.00863f
C7258 XA.XIR[0].XIC[13].icell.SM Iout 0.00367f
C7259 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.SM 0.00188f
C7260 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00212f
C7261 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00212f
C7262 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.SM 0.00188f
C7263 XA.XIR[4].XIC[6].icell.PDM Vbias 0.04058f
C7264 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PUM 0.00131f
C7265 XA.XIR[11].XIC[5].icell.PDM Iout 0.00112f
C7266 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02698f
C7267 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00529f
C7268 XA.XIR[10].XIC[7].icell.SM VPWR 0.00158f
C7269 XA.XIR[6].XIC[6].icell.PUM VPWR 0.01036f
C7270 XA.XIR[15].XIC[11].icell.PDM Iout 0.00112f
C7271 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.01406f
C7272 XA.XIR[3].XIC[6].icell.Ien Vbias 0.21238f
C7273 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C7274 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.15089f
C7275 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04522f
C7276 XA.XIR[10].XIC[4].icell.SM Iout 0.00388f
C7277 XThR.XTB7.A a_n1049_6405# 0.02287f
C7278 XA.XIR[5].XIC[9].icell.PDM VPWR 0.00863f
C7279 XThR.Tn[13] XA.XIR[14].XIC[9].icell.SM 0.00121f
C7280 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04522f
C7281 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04f
C7282 XThR.Tn[8] XA.XIR[8].XIC[3].icell.PDM 0.0033f
C7283 XA.XIR[2].XIC[8].icell.PUM Vbias 0.00347f
C7284 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.SM 0.00383f
C7285 XA.XIR[4].XIC[9].icell.Ien VPWR 0.19065f
C7286 XA.XIR[5].XIC[6].icell.PDM Iout 0.00112f
C7287 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.SM 0.00383f
C7288 XThR.Tn[12] XA.XIR[13].XIC[0].icell.Ien 0.0035f
C7289 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C7290 XA.XIR[12].XIC[9].icell.Ien VPWR 0.19065f
C7291 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.SM 0.00383f
C7292 XThR.Tn[7] XA.XIR[8].XIC[2].icell.Ien 0.00321f
C7293 XA.XIR[3].XIC[10].icell.SM VPWR 0.00158f
C7294 XA.XIR[4].XIC[6].icell.Ien Iout 0.06483f
C7295 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PUM 0.00131f
C7296 XA.XIR[9].XIC[6].icell.SM Vbias 0.00701f
C7297 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.01406f
C7298 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.15089f
C7299 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.SM 0.00383f
C7300 XA.XIR[8].XIC[5].icell.PUM VPWR 0.01036f
C7301 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.03976f
C7302 XA.XIR[3].XIC[7].icell.SM Iout 0.00388f
C7303 XThC.Tn[0] XA.XIR[5].XIC_dummy_left.icell.Iout 0.00111f
C7304 XA.XIR[10].XIC[12].icell.SM VPWR 0.00158f
C7305 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PUM 0.00529f
C7306 XThC.Tn[4] VPWR 5.94691f
C7307 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00529f
C7308 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.01406f
C7309 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04522f
C7310 XThR.Tn[5] XA.XIR[5].XIC[3].icell.PDM 0.0033f
C7311 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[6].icell.SM 0.00383f
C7312 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.01406f
C7313 XA.XIR[2].XIC[11].icell.PDM Iout 0.00112f
C7314 XA.XIR[15].XIC[10].icell.SM VPWR 0.00158f
C7315 XA.XIR[10].XIC[8].icell.SM Iout 0.00388f
C7316 XA.XIR[11].XIC[10].icell.PUM Vbias 0.00347f
C7317 XA.XIR[13].XIC_dummy_left.icell.SM VPWR 0.00269f
C7318 XThC.Tn[10] XThR.Tn[0] 0.28074f
C7319 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11595f
C7320 XThC.Tn[12] XThR.Tn[14] 0.28062f
C7321 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02698f
C7322 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9] 0.0033f
C7323 XThR.Tn[13] XA.XIR[14].XIC[11].icell.Ien 0.00321f
C7324 XA.XIR[4].XIC[12].icell.SM VPWR 0.00158f
C7325 XThC.Tn[3] XThR.Tn[9] 0.28062f
C7326 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PUM 0.00131f
C7327 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00212f
C7328 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C7329 XThC.XTB7.B a_7875_9569# 0.01174f
C7330 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C7331 XA.XIR[7].XIC[4].icell.PUM Vbias 0.00347f
C7332 XThR.Tn[14] XA.XIR[15].XIC[5].icell.SM 0.00121f
C7333 XA.XIR[14].XIC[9].icell.SM Vbias 0.00701f
C7334 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06536f
C7335 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00212f
C7336 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.SM 0.00188f
C7337 XThR.XTB7.A a_n997_2891# 0.00342f
C7338 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C7339 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C7340 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PUM 0.00529f
C7341 XThR.Tn[3] XA.XIR[3].XIC[13].icell.PDM 0.0033f
C7342 a_n1049_7493# XA.XIR[1].XIC_dummy_left.icell.Iout 0.0013f
C7343 XA.XIR[1].XIC[5].icell.PUM Vbias 0.00347f
C7344 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Ien 0.00529f
C7345 XA.XIR[12].XIC[12].icell.PDM VPWR 0.00863f
C7346 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01193f
C7347 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.SM 0.00383f
C7348 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00212f
C7349 XThC.Tn[12] XA.XIR[0].XIC[11].icell.PDM 0.00102f
C7350 XThR.Tn[8] XA.XIR[9].XIC[12].icell.Ien 0.00321f
C7351 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02698f
C7352 a_8963_9569# XThC.Tn[11] 0.19413f
C7353 XA.XIR[12].XIC[0].icell.Ien Vbias 0.21102f
C7354 XA.XIR[8].XIC[0].icell.PDM Vbias 0.04002f
C7355 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.01406f
C7356 XA.XIR[0].XIC[5].icell.Ien Vbias 0.21245f
C7357 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Iout 0.00347f
C7358 XA.XIR[8].XIC[11].icell.PUM Vbias 0.00347f
C7359 XA.XIR[2].XIC[13].icell.Ien Iout 0.06483f
C7360 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PUM 0.00131f
C7361 XA.XIR[7].XIC[10].icell.PDM VPWR 0.00863f
C7362 XA.XIR[11].XIC[3].icell.PDM Vbias 0.04058f
C7363 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PUM 0.00529f
C7364 XA.XIR[5].XIC_15.icell.Ien VPWR 0.25675f
C7365 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00529f
C7366 XThR.Tn[4] XA.XIR[4].XIC[13].icell.PDM 0.0033f
C7367 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PUM 0.00131f
C7368 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C7369 XA.XIR[1].XIC[11].icell.PDM VPWR 0.00863f
C7370 XA.XIR[7].XIC[7].icell.PDM Iout 0.00112f
C7371 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.15089f
C7372 XA.XIR[2].XIC_dummy_right.icell.PUM Vbias 0.00248f
C7373 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PUM 0.00529f
C7374 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00212f
C7375 XA.XIR[9].XIC[1].icell.PUM VPWR 0.01036f
C7376 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PUM 0.00529f
C7377 XA.XIR[13].XIC[0].icell.SM Iout 0.00388f
C7378 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.SM 0.00188f
C7379 XA.XIR[1].XIC[8].icell.PDM Iout 0.00112f
C7380 XA.XIR[13].XIC[14].icell.Ien Iout 0.06483f
C7381 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.03424f
C7382 XThR.Tn[12] XA.XIR[13].XIC[4].icell.Ien 0.00321f
C7383 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PDM 0.00182f
C7384 XA.XIR[9].XIC[14].icell.PDM Iout 0.00112f
C7385 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.SM 0.00383f
C7386 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.15089f
C7387 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PUM 0.00529f
C7388 XA.XIR[0].XIC[9].icell.SM VPWR 0.00158f
C7389 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.SM 0.00188f
C7390 XThR.Tn[12] Iout 1.16627f
C7391 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.03976f
C7392 XThC.Tn[1] XThR.Tn[11] 0.28062f
C7393 XA.XIR[3].XIC_dummy_left.icell.SM VPWR 0.00269f
C7394 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C7395 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01897f
C7396 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.15089f
C7397 XA.XIR[9].XIC_15.icell.PUM Vbias 0.00347f
C7398 XA.XIR[14].XIC[11].icell.Ien Vbias 0.21238f
C7399 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C7400 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Ien 0.00529f
C7401 XA.XIR[0].XIC[6].icell.SM Iout 0.00367f
C7402 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04522f
C7403 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.03976f
C7404 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.SM 0.00383f
C7405 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.01406f
C7406 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04522f
C7407 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PUM 0.00131f
C7408 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.SM 0.00383f
C7409 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PDM 0.00182f
C7410 XA.XIR[7].XIC[12].icell.Ien VPWR 0.19065f
C7411 XA.XIR[15].XIC[9].icell.PDM Vbias 0.04058f
C7412 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.SM 0.00188f
C7413 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.SM 0.00383f
C7414 a_n1319_5611# VPWR 0.00674f
C7415 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.03424f
C7416 XA.XIR[2].XIC[1].icell.PUM Vbias 0.00347f
C7417 XA.XIR[10].XIC_15.icell.Ien Iout 0.06485f
C7418 XA.XIR[1].XIC[13].icell.Ien VPWR 0.19065f
C7419 XA.XIR[11].XIC_dummy_right.icell.Ien Vbias 0.00287f
C7420 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.01406f
C7421 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.03424f
C7422 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.SM 0.00383f
C7423 XA.XIR[4].XIC[2].icell.Ien VPWR 0.19065f
C7424 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00529f
C7425 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11181f
C7426 XA.XIR[7].XIC[1].icell.PDM Vbias 0.04058f
C7427 XThR.XTBN.A a_n997_3979# 0.02087f
C7428 XA.XIR[10].XIC[13].icell.PDM Iout 0.00112f
C7429 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.01406f
C7430 XThC.Tn[14] XThR.Tn[13] 0.28068f
C7431 XA.XIR[13].XIC[3].icell.Ien Vbias 0.21238f
C7432 XThC.XTB7.B Iout 0.01f
C7433 XThR.Tn[5] XA.XIR[6].XIC[14].icell.Ien 0.00321f
C7434 XA.XIR[3].XIC[3].icell.SM VPWR 0.00158f
C7435 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PUM 0.00131f
C7436 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C7437 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00212f
C7438 XThR.Tn[9] a_n997_3755# 0.19352f
C7439 XThC.XTB7.A XThC.Tn[5] 0.02758f
C7440 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.15089f
C7441 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.01406f
C7442 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Ien 0.00529f
C7443 XA.XIR[3].XIC[0].icell.SM Iout 0.00388f
C7444 XA.XIR[12].XIC[4].icell.Ien Vbias 0.21238f
C7445 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00529f
C7446 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.03424f
C7447 XA.XIR[2].XIC[7].icell.PDM VPWR 0.00863f
C7448 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C7449 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.SM 0.00188f
C7450 XA.XIR[14].XIC[8].icell.PDM VPWR 0.00863f
C7451 XThC.Tn[1] XThR.Tn[7] 0.28062f
C7452 XA.XIR[11].XIC[7].icell.PDM Vbias 0.04058f
C7453 XA.XIR[2].XIC[4].icell.PDM Iout 0.00112f
C7454 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PUM 0.00131f
C7455 XThC.Tn[4] XThR.Tn[12] 0.28062f
C7456 XThC.Tn[6] XThR.Tn[2] 0.28062f
C7457 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.SM 0.00383f
C7458 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C7459 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PUM 0.00529f
C7460 XA.XIR[13].XIC[7].icell.SM VPWR 0.00158f
C7461 XA.XIR[14].XIC[5].icell.PDM Iout 0.00112f
C7462 XThR.Tn[1] XA.XIR[2].XIC[4].icell.SM 0.00121f
C7463 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.SM 0.00383f
C7464 XA.XIR[10].XIC[6].icell.SM Vbias 0.00701f
C7465 XA.XIR[9].XIC[5].icell.PUM VPWR 0.01036f
C7466 XA.XIR[6].XIC[5].icell.PUM Vbias 0.00347f
C7467 XA.XIR[13].XIC[4].icell.SM Iout 0.00388f
C7468 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.01406f
C7469 XThR.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.0033f
C7470 XA.XIR[5].XIC[8].icell.PDM Vbias 0.04058f
C7471 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.0353f
C7472 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PUM 0.00131f
C7473 a_6243_9615# VPWR 0.70588f
C7474 XA.XIR[12].XIC[5].icell.SM Iout 0.00388f
C7475 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.03976f
C7476 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04522f
C7477 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.SM 0.00383f
C7478 XThR.Tn[3] XA.XIR[3].XIC[6].icell.PDM 0.0033f
C7479 XA.XIR[4].XIC[8].icell.Ien Vbias 0.21238f
C7480 VPWR data[1] 0.44103f
C7481 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.03976f
C7482 XA.XIR[10].XIC[13].icell.PUM VPWR 0.01036f
C7483 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.15089f
C7484 XA.XIR[11].XIC[7].icell.Ien Iout 0.06483f
C7485 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00529f
C7486 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00529f
C7487 XA.XIR[6].XIC[11].icell.PDM VPWR 0.00863f
C7488 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.01406f
C7489 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.01406f
C7490 XA.XIR[3].XIC[9].icell.SM Vbias 0.00701f
C7491 XThR.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.0033f
C7492 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.03976f
C7493 XThC.Tn[14] Vbias 2.38887f
C7494 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.03976f
C7495 XThC.Tn[3] XThR.Tn[10] 0.28062f
C7496 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PUM 0.00529f
C7497 XA.XIR[15].XIC[11].icell.PUM VPWR 0.01036f
C7498 XA.XIR[11].XIC[11].icell.PDM Vbias 0.04058f
C7499 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.03424f
C7500 XA.XIR[7].XIC[3].icell.PDM VPWR 0.00863f
C7501 XA.XIR[8].XIC[4].icell.PUM Vbias 0.00347f
C7502 XA.XIR[6].XIC[8].icell.PDM Iout 0.00112f
C7503 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PUM 0.00131f
C7504 XA.XIR[5].XIC[11].icell.Ien VPWR 0.19065f
C7505 XA.XIR[13].XIC[12].icell.SM VPWR 0.00158f
C7506 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04522f
C7507 XThC.XTB7.B XThC.Tn[4] 0.00356f
C7508 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.15089f
C7509 XA.XIR[2].XIC[13].icell.PDM Vbias 0.04058f
C7510 XThC.XTB5.Y XThC.Tn[8] 0.01728f
C7511 XThC.XTB7.Y a_7651_9569# 0.00477f
C7512 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01402f
C7513 XA.XIR[5].XIC[8].icell.Ien Iout 0.06483f
C7514 XA.XIR[1].XIC[4].icell.PDM VPWR 0.00863f
C7515 XThR.Tn[4] XA.XIR[4].XIC[6].icell.PDM 0.0033f
C7516 XThR.XTB1.Y data[4] 0.06453f
C7517 XThC.XTB6.Y XThC.Tn[12] 0.02863f
C7518 XA.XIR[13].XIC[8].icell.SM Iout 0.00388f
C7519 XA.XIR[14].XIC[10].icell.PUM Vbias 0.00347f
C7520 XThC.XTB6.A a_5155_10571# 0.00306f
C7521 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PUM 0.00529f
C7522 XThR.Tn[7] XA.XIR[8].XIC[5].icell.SM 0.00121f
C7523 XA.XIR[9].XIC[0].icell.PDM Vbias 0.04002f
C7524 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02698f
C7525 XA.XIR[4].XIC[9].icell.SM Iout 0.00388f
C7526 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00529f
C7527 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.03976f
C7528 XA.XIR[9].XIC[11].icell.PUM Vbias 0.00347f
C7529 XA.XIR[8].XIC[10].icell.PDM VPWR 0.00863f
C7530 XA.XIR[0].XIC[2].icell.SM VPWR 0.00158f
C7531 XA.XIR[12].XIC[10].icell.Ien VPWR 0.19065f
C7532 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01734f
C7533 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.03976f
C7534 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C7535 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.SM 0.00188f
C7536 XA.XIR[4].XIC[11].icell.SM Vbias 0.00701f
C7537 XThR.Tn[9] XThR.Tn[11] 0.00252f
C7538 a_5949_9615# XThC.Tn[5] 0.27124f
C7539 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00529f
C7540 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.SM 0.00188f
C7541 XA.XIR[8].XIC[7].icell.PDM Iout 0.00112f
C7542 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.03424f
C7543 XA.XIR[6].XIC[13].icell.Ien VPWR 0.19065f
C7544 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.15089f
C7545 XA.XIR[10].XIC[1].icell.PUM VPWR 0.01036f
C7546 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PUM 0.00529f
C7547 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00529f
C7548 XA.XIR[15].XIC_15.icell.SM VPWR 0.00276f
C7549 XA.XIR[3].XIC[14].icell.PUM Vbias 0.00347f
C7550 XA.XIR[10].XIC[13].icell.SM VPWR 0.00158f
C7551 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02698f
C7552 XA.XIR[14].XIC[1].icell.PDM Iout 0.00112f
C7553 XA.XIR[15].XIC[2].icell.PDM Vbias 0.04058f
C7554 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00212f
C7555 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.01406f
C7556 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04522f
C7557 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.SM 0.00383f
C7558 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04522f
C7559 XA.XIR[10].XIC[9].icell.SM Iout 0.00388f
C7560 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02698f
C7561 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00212f
C7562 XA.XIR[5].XIC[11].icell.SM Iout 0.00388f
C7563 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.SM 0.00188f
C7564 XA.XIR[14].XIC[3].icell.PDM Vbias 0.04058f
C7565 XA.XIR[5].XIC[0].icell.PDM Vbias 0.04002f
C7566 XThC.XTBN.Y XThC.Tn[8] 0.50311f
C7567 XThR.Tn[10] XA.XIR[11].XIC[2].icell.Ien 0.00321f
C7568 XA.XIR[7].XIC[9].icell.PDM Vbias 0.04058f
C7569 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13469f
C7570 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.01406f
C7571 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.SM 0.00383f
C7572 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.03424f
C7573 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04522f
C7574 XThC.XTB1.Y a_2979_9615# 0.21263f
C7575 XA.XIR[1].XIC[10].icell.PDM Vbias 0.04058f
C7576 XA.XIR[8].XIC[12].icell.Ien VPWR 0.19065f
C7577 XA.XIR[15].XIC[5].icell.Ien VPWR 0.32782f
C7578 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.PUM 0.00137f
C7579 XA.XIR[3].XIC_15.icell.SM VPWR 0.00276f
C7580 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00212f
C7581 XThR.Tn[8] XA.XIR[9].XIC[1].icell.Ien 0.00321f
C7582 XThC.Tn[1] XThR.Tn[14] 0.28062f
C7583 XThC.XTB4.Y XThC.Tn[12] 0.00209f
C7584 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.SM 0.00383f
C7585 XA.XIR[0].XIC[8].icell.SM Vbias 0.00701f
C7586 XA.XIR[15].XIC[2].icell.Ien Iout 0.06816f
C7587 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.03976f
C7588 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04522f
C7589 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04522f
C7590 XThC.Tn[14] XThR.Tn[6] 0.28068f
C7591 XA.XIR[7].XIC[9].icell.Ien Iout 0.06483f
C7592 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.03976f
C7593 XThC.Tn[8] XThC.Tn[10] 0.00465f
C7594 XThR.XTB5.A XThR.XTB6.A 1.80461f
C7595 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.03424f
C7596 XA.XIR[5].XIC_dummy_right.icell.SM VPWR 0.00123f
C7597 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00529f
C7598 XA.XIR[1].XIC[10].icell.Ien Iout 0.06483f
C7599 XThC.Tn[13] XThC.Tn[14] 0.39285f
C7600 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04522f
C7601 XThR.Tn[12] XA.XIR[13].XIC[7].icell.SM 0.00121f
C7602 XA.XIR[12].XIC[1].icell.SM VPWR 0.00158f
C7603 XA.XIR[9].XIC[3].icell.PDM Iout 0.00112f
C7604 XA.XIR[10].XIC[11].icell.Ien Iout 0.06483f
C7605 XA.XIR[0].XIC[14].icell.PUM VPWR 0.00971f
C7606 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02698f
C7607 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00529f
C7608 XA.XIR[13].XIC_15.icell.Ien Iout 0.06485f
C7609 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C7610 XA.XIR[14].XIC_dummy_right.icell.Ien Vbias 0.00287f
C7611 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02698f
C7612 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00212f
C7613 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.04038f
C7614 XA.XIR[1].XIC[12].icell.Ien Vbias 0.21238f
C7615 XA.XIR[11].XIC[3].icell.Ien VPWR 0.19065f
C7616 XA.XIR[15].XIC[9].icell.Ien VPWR 0.32782f
C7617 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.01406f
C7618 XA.XIR[4].XIC[1].icell.Ien Vbias 0.21238f
C7619 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PUM 0.00529f
C7620 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.03424f
C7621 XA.XIR[13].XIC[13].icell.PDM Iout 0.00112f
C7622 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.SM 0.00383f
C7623 XThR.Tn[7] XA.XIR[7].XIC_15.icell.PDM 0.0033f
C7624 XThC.Tn[8] XThR.Tn[5] 0.28062f
C7625 XA.XIR[6].XIC[4].icell.PDM VPWR 0.00863f
C7626 XA.XIR[10].XIC[5].icell.PUM VPWR 0.01036f
C7627 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C7628 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.03976f
C7629 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.03976f
C7630 XA.XIR[3].XIC[2].icell.SM Vbias 0.00701f
C7631 XThR.XTB7.B XThR.XTB7.A 0.35833f
C7632 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.SM 0.00188f
C7633 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C7634 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04522f
C7635 XA.XIR[5].XIC[4].icell.Ien VPWR 0.19065f
C7636 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.SM 0.00383f
C7637 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C7638 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02698f
C7639 XA.XIR[2].XIC[6].icell.PDM Vbias 0.04058f
C7640 XA.XIR[7].XIC[12].icell.SM Iout 0.00388f
C7641 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00529f
C7642 XA.XIR[14].XIC[7].icell.PDM Vbias 0.04058f
C7643 XA.XIR[4].XIC[5].icell.SM VPWR 0.00158f
C7644 XThR.Tn[12] XA.XIR[13].XIC[12].icell.SM 0.00121f
C7645 XA.XIR[5].XIC[1].icell.Ien Iout 0.06483f
C7646 XA.XIR[1].XIC[13].icell.SM Iout 0.00388f
C7647 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.SM 0.00188f
C7648 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PUM 0.00529f
C7649 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.01406f
C7650 XA.XIR[7].XIC_15.icell.Ien Vbias 0.21343f
C7651 XA.XIR[13].XIC[6].icell.SM Vbias 0.00701f
C7652 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10] 0.0033f
C7653 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Ien 0.00217f
C7654 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04522f
C7655 XA.XIR[4].XIC[2].icell.SM Iout 0.00388f
C7656 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.03976f
C7657 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PUM 0.00529f
C7658 XA.XIR[3].XIC[8].icell.PUM VPWR 0.01036f
C7659 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.SM 0.00383f
C7660 XThR.XTB6.A data[5] 0.37233f
C7661 XA.XIR[9].XIC[4].icell.PUM Vbias 0.00347f
C7662 XA.XIR[10].XIC[14].icell.PDM VPWR 0.00873f
C7663 XA.XIR[8].XIC[3].icell.PDM VPWR 0.00863f
C7664 XA.XIR[12].XIC[7].icell.SM Vbias 0.00701f
C7665 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00529f
C7666 XThR.Tn[8] XA.XIR[9].XIC[5].icell.Ien 0.00321f
C7667 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.0353f
C7668 XA.XIR[2].XIC[9].icell.Ien VPWR 0.19065f
C7669 XThC.XTB7.B a_6243_9615# 0.01743f
C7670 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.15089f
C7671 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Ien 0.00714f
C7672 XThR.XTB2.Y a_n1049_7787# 0.2342f
C7673 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01193f
C7674 XThC.XTB7.B data[1] 0.00593f
C7675 a_4067_9615# Vbias 0.00553f
C7676 XA.XIR[10].XIC[9].icell.PUM VPWR 0.01036f
C7677 XA.XIR[2].XIC[6].icell.Ien Iout 0.06483f
C7678 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PUM 0.00529f
C7679 XA.XIR[13].XIC[13].icell.PUM VPWR 0.01036f
C7680 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04522f
C7681 XA.XIR[14].XIC[7].icell.Ien Iout 0.06483f
C7682 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PUM 0.00131f
C7683 XA.XIR[9].XIC[10].icell.PDM VPWR 0.00863f
C7684 XA.XIR[6].XIC[10].icell.PDM Vbias 0.04058f
C7685 XThC.Tn[3] XThR.Tn[13] 0.28062f
C7686 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.15089f
C7687 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00529f
C7688 XThR.Tn[10] XThR.Tn[11] 0.07356f
C7689 XA.XIR[14].XIC[11].icell.PDM Vbias 0.04058f
C7690 XA.XIR[9].XIC[7].icell.PDM Iout 0.00112f
C7691 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.03976f
C7692 XA.XIR[5].XIC[10].icell.Ien Vbias 0.21238f
C7693 XThC.Tn[5] XThR.Tn[3] 0.28062f
C7694 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PUM 0.00131f
C7695 XA.XIR[7].XIC[2].icell.PDM Vbias 0.04058f
C7696 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PUM 0.00529f
C7697 XA.XIR[11].XIC[1].icell.PDM VPWR 0.00863f
C7698 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04522f
C7699 XA.XIR[1].XIC[3].icell.PDM Vbias 0.04058f
C7700 XThR.Tn[2] XA.XIR[3].XIC[9].icell.Ien 0.00321f
C7701 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.15089f
C7702 XA.XIR[12].XIC[12].icell.SM Vbias 0.00701f
C7703 XA.XIR[2].XIC[12].icell.SM VPWR 0.00158f
C7704 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.SM 0.00383f
C7705 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.SM 0.00188f
C7706 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01897f
C7707 XA.XIR[10].XIC[14].icell.PUM VPWR 0.01036f
C7708 XA.XIR[0].XIC[1].icell.SM Vbias 0.00701f
C7709 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00212f
C7710 XA.XIR[6].XIC[10].icell.Ien Iout 0.06483f
C7711 XA.XIR[7].XIC[5].icell.Ien VPWR 0.19065f
C7712 XA.XIR[8].XIC[9].icell.PDM Vbias 0.04058f
C7713 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.03976f
C7714 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04522f
C7715 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.SM 0.00188f
C7716 a_8963_9569# VPWR 0.0033f
C7717 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04f
C7718 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.SM 0.00383f
C7719 XA.XIR[13].XIC[1].icell.PUM VPWR 0.01036f
C7720 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.15089f
C7721 XA.XIR[13].XIC[13].icell.SM VPWR 0.00158f
C7722 XA.XIR[6].XIC[12].icell.Ien Vbias 0.21238f
C7723 XA.XIR[7].XIC[2].icell.Ien Iout 0.06483f
C7724 XA.XIR[1].XIC[6].icell.Ien VPWR 0.19065f
C7725 XA.XIR[9].XIC[12].icell.Ien VPWR 0.19065f
C7726 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.15089f
C7727 XThR.XTB2.Y XThR.Tn[9] 0.292f
C7728 XA.XIR[1].XIC[3].icell.Ien Iout 0.06483f
C7729 XA.XIR[12].XIC[2].icell.PUM VPWR 0.01036f
C7730 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04522f
C7731 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PUM 0.00131f
C7732 XA.XIR[5].XIC[13].icell.SM Vbias 0.00701f
C7733 XThC.Tn[14] XThR.Tn[4] 0.28068f
C7734 XA.XIR[13].XIC[9].icell.SM Iout 0.00388f
C7735 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Iout 0.00347f
C7736 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C7737 XA.XIR[0].XIC[7].icell.PUM VPWR 0.00971f
C7738 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.03011f
C7739 XThR.Tn[5] XA.XIR[6].XIC[7].icell.Ien 0.00321f
C7740 XA.XIR[9].XIC[1].icell.PDM Vbias 0.04058f
C7741 XThC.Tn[3] Vbias 2.38713f
C7742 XThR.Tn[6] XA.XIR[7].XIC_15.icell.Ien 0.00116f
C7743 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01897f
C7744 XThR.XTB6.Y a_n997_3979# 0.0046f
C7745 XThR.Tn[2] XA.XIR[3].XIC[12].icell.SM 0.00121f
C7746 XThR.XTB6.A a_n1335_4229# 0.00304f
C7747 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.01406f
C7748 XA.XIR[8].XIC[9].icell.Ien Iout 0.06483f
C7749 XA.XIR[11].XIC[2].icell.PDM Iout 0.00112f
C7750 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04522f
C7751 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PUM 0.00529f
C7752 XThR.Tn[11] XA.XIR[12].XIC[3].icell.Ien 0.00321f
C7753 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.SM 0.00188f
C7754 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00212f
C7755 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.SM 0.00188f
C7756 XA.XIR[6].XIC[13].icell.SM Iout 0.00388f
C7757 XA.XIR[15].XIC[4].icell.Ien Vbias 0.17911f
C7758 XA.XIR[10].XIC[3].icell.PDM Iout 0.00112f
C7759 XA.XIR[10].XIC[14].icell.SM VPWR 0.00208f
C7760 XThR.Tn[11] XA.XIR[11].XIC[6].icell.PDM 0.0033f
C7761 XThC.XTB5.Y XThC.Tn[6] 0.00352f
C7762 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.SM 0.00188f
C7763 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.03424f
C7764 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00212f
C7765 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04522f
C7766 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35783f
C7767 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.SM 0.00188f
C7768 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.SM 0.00383f
C7769 XThR.Tn[10] XA.XIR[11].XIC[5].icell.SM 0.00121f
C7770 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C7771 XA.XIR[7].XIC[11].icell.Ien Vbias 0.21238f
C7772 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PUM 0.00529f
C7773 XThR.Tn[6] XA.XIR[6].XIC[10].icell.PDM 0.0033f
C7774 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.01406f
C7775 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PDM 0.00182f
C7776 XThR.Tn[5] a_n1049_5317# 0.00158f
C7777 XThR.Tn[10] XA.XIR[10].XIC[9].icell.PDM 0.0033f
C7778 XThC.Tn[12] Iout 0.84582f
C7779 XA.XIR[3].XIC[1].icell.PUM VPWR 0.01036f
C7780 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.03976f
C7781 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00529f
C7782 XA.XIR[13].XIC[11].icell.Ien Iout 0.06483f
C7783 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.002f
C7784 XA.XIR[8].XIC[12].icell.SM Iout 0.00388f
C7785 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.01406f
C7786 XA.XIR[15].XIC[5].icell.SM Iout 0.00388f
C7787 XA.XIR[2].XIC[2].icell.Ien VPWR 0.19065f
C7788 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.03982f
C7789 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01734f
C7790 XA.XIR[0].XIC[13].icell.PUM Vbias 0.00347f
C7791 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.SM 0.00383f
C7792 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00529f
C7793 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C7794 XA.XIR[14].XIC[3].icell.Ien VPWR 0.19119f
C7795 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00529f
C7796 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.SM 0.00383f
C7797 XA.XIR[11].XIC[2].icell.Ien Vbias 0.21238f
C7798 XA.XIR[8].XIC_15.icell.Ien Vbias 0.21343f
C7799 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.03424f
C7800 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00212f
C7801 XThR.Tn[0] XA.XIR[1].XIC[9].icell.Ien 0.00321f
C7802 XA.XIR[13].XIC[5].icell.PUM VPWR 0.01036f
C7803 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PUM 0.00529f
C7804 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PUM 0.00131f
C7805 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PUM 0.00131f
C7806 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PUM 0.00487f
C7807 XThC.XTBN.Y XThC.Tn[6] 0.61358f
C7808 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.SM 0.00383f
C7809 XA.XIR[6].XIC[3].icell.PDM Vbias 0.04058f
C7810 XA.XIR[10].XIC[4].icell.PUM Vbias 0.00347f
C7811 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.15089f
C7812 XA.XIR[12].XIC[6].icell.PUM VPWR 0.01036f
C7813 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.15089f
C7814 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01402f
C7815 XA.XIR[5].XIC[3].icell.Ien Vbias 0.21238f
C7816 XThC.XTB7.Y a_5949_9615# 0.00153f
C7817 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.SM 0.00383f
C7818 XA.XIR[10].XIC[12].icell.Ien VPWR 0.19065f
C7819 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.01406f
C7820 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PUM 0.00529f
C7821 XA.XIR[11].XIC[6].icell.SM VPWR 0.00158f
C7822 XThR.Tn[5] XA.XIR[6].XIC[14].icell.SM 0.00121f
C7823 XThR.Tn[1] Iout 1.16635f
C7824 XThR.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.00321f
C7825 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.15089f
C7826 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PUM 0.00529f
C7827 XA.XIR[4].XIC[4].icell.SM Vbias 0.00701f
C7828 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PUM 0.00202f
C7829 XA.XIR[11].XIC[3].icell.SM Iout 0.00388f
C7830 XThC.Tn[3] XThR.Tn[6] 0.28062f
C7831 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04522f
C7832 XA.XIR[6].XIC[6].icell.Ien VPWR 0.19065f
C7833 XA.XIR[10].XIC[10].icell.PDM VPWR 0.00863f
C7834 XA.XIR[15].XIC[10].icell.Ien VPWR 0.32782f
C7835 XThC.Tn[5] XThR.Tn[8] 0.28062f
C7836 XA.XIR[3].XIC[7].icell.PUM Vbias 0.00347f
C7837 XA.XIR[13].XIC[14].icell.PDM VPWR 0.00873f
C7838 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.SM 0.00383f
C7839 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00529f
C7840 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00529f
C7841 XA.XIR[10].XIC[7].icell.PDM Iout 0.00112f
C7842 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04522f
C7843 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PUM 0.00487f
C7844 XA.XIR[6].XIC[3].icell.Ien Iout 0.06483f
C7845 XThR.Tn[11] XA.XIR[11].XIC_15.icell.PDM 0.0033f
C7846 XA.XIR[5].XIC[7].icell.SM VPWR 0.00158f
C7847 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7] 0.0033f
C7848 a_7651_9569# XThC.Tn[8] 0.1927f
C7849 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.SM 0.00188f
C7850 XA.XIR[2].XIC[8].icell.Ien Vbias 0.21238f
C7851 XThR.Tn[0] XA.XIR[1].XIC[12].icell.SM 0.00121f
C7852 XA.XIR[13].XIC[9].icell.PUM VPWR 0.01036f
C7853 XThC.XTB5.A XThC.XTB7.Y 0.00179f
C7854 XA.XIR[5].XIC[4].icell.SM Iout 0.00388f
C7855 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04522f
C7856 XA.XIR[4].XIC[10].icell.PUM VPWR 0.01036f
C7857 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.01406f
C7858 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.15089f
C7859 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PUM 0.00131f
C7860 XThR.Tn[12] XA.XIR[13].XIC[13].icell.SM 0.00121f
C7861 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PUM 0.00131f
C7862 XThR.Tn[6] XA.XIR[7].XIC[11].icell.Ien 0.00321f
C7863 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38957f
C7864 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00212f
C7865 XA.XIR[3].XIC[13].icell.PDM VPWR 0.00863f
C7866 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.SM 0.00188f
C7867 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.SM 0.00188f
C7868 XA.XIR[12].XIC[13].icell.PUM Vbias 0.00347f
C7869 XA.XIR[9].XIC[9].icell.PDM Vbias 0.04058f
C7870 XThR.Tn[11] XThR.Tn[13] 0.00153f
C7871 XA.XIR[8].XIC[5].icell.Ien VPWR 0.19065f
C7872 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.01406f
C7873 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.SM 0.00383f
C7874 XThR.Tn[5] XA.XIR[6].XIC[0].icell.Ien 0.00321f
C7875 XThC.Tn[6] XThR.Tn[5] 0.28062f
C7876 XA.XIR[3].XIC[10].icell.PDM Iout 0.00112f
C7877 XThR.Tn[8] XA.XIR[9].XIC[8].icell.SM 0.00121f
C7878 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.03011f
C7879 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.01406f
C7880 XA.XIR[8].XIC[2].icell.Ien Iout 0.06483f
C7881 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02698f
C7882 XA.XIR[2].XIC[9].icell.SM Iout 0.00388f
C7883 XThR.XTB2.Y XThR.Tn[10] 0.00106f
C7884 XThR.Tn[9] XA.XIR[10].XIC[0].icell.Ien 0.00352f
C7885 XA.XIR[10].XIC[11].icell.PDM Iout 0.00112f
C7886 XA.XIR[5].XIC[12].icell.PUM VPWR 0.01036f
C7887 XThC.Tn[4] XThR.Tn[1] 0.28063f
C7888 XA.XIR[13].XIC[14].icell.PUM VPWR 0.01036f
C7889 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00212f
C7890 XA.XIR[10].XIC[1].icell.PDM Vbias 0.04058f
C7891 XA.XIR[2].XIC[11].icell.SM Vbias 0.00701f
C7892 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02698f
C7893 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.SM 0.00188f
C7894 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C7895 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PUM 0.00501f
C7896 XA.XIR[4].XIC_15.icell.PDM VPWR 0.06959f
C7897 XThC.XTB7.B a_8963_9569# 0.02071f
C7898 XThR.Tn[3] XA.XIR[4].XIC[10].icell.Ien 0.00321f
C7899 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04522f
C7900 XA.XIR[9].XIC[9].icell.Ien Iout 0.06483f
C7901 XA.XIR[7].XIC[4].icell.Ien Vbias 0.21238f
C7902 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.SM 0.00188f
C7903 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.03976f
C7904 XThR.Tn[6] XA.XIR[6].XIC[3].icell.PDM 0.0033f
C7905 XA.XIR[9].XIC_dummy_left.icell.Ien Vbias 0.00342f
C7906 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.03011f
C7907 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00212f
C7908 XA.XIR[1].XIC[5].icell.Ien Vbias 0.21238f
C7909 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04522f
C7910 XThC.XTB6.A XThC.XTB7.A 0.44014f
C7911 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00529f
C7912 XA.XIR[15].XIC[1].icell.SM VPWR 0.00158f
C7913 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00212f
C7914 XA.XIR[3].XIC[12].icell.Ien Iout 0.06483f
C7915 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PUM 0.00131f
C7916 XA.XIR[12].XIC[1].icell.PUM Vbias 0.00347f
C7917 XThR.Tn[7] XA.XIR[7].XIC[8].icell.PDM 0.0033f
C7918 XA.XIR[3].XIC[0].icell.PDM Vbias 0.04002f
C7919 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00212f
C7920 XA.XIR[12].XIC[13].icell.SM Vbias 0.00701f
C7921 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.01406f
C7922 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00212f
C7923 XA.XIR[0].XIC[6].icell.PUM Vbias 0.00347f
C7924 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.SM 0.00188f
C7925 XThR.Tn[4] XA.XIR[5].XIC[10].icell.Ien 0.00321f
C7926 XA.XIR[7].XIC[8].icell.SM VPWR 0.00158f
C7927 XThR.Tn[13] XA.XIR[14].XIC[2].icell.Ien 0.00321f
C7928 XA.XIR[8].XIC[11].icell.Ien Vbias 0.21238f
C7929 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PUM 0.00529f
C7930 XThR.Tn[11] Vbias 3.71832f
C7931 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.03011f
C7932 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04522f
C7933 XA.XIR[14].XIC[0].icell.Ien Iout 0.06474f
C7934 XThR.XTB7.B a_n997_3979# 0.01152f
C7935 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PUM 0.00529f
C7936 XA.XIR[1].XIC[9].icell.SM VPWR 0.00158f
C7937 XThR.Tn[0] XA.XIR[1].XIC[2].icell.Ien 0.00321f
C7938 XThC.XTB2.Y XThC.Tn[1] 0.17879f
C7939 XA.XIR[7].XIC[5].icell.SM Iout 0.00388f
C7940 XA.XIR[9].XIC[1].icell.Ien VPWR 0.19065f
C7941 XThR.XTB6.A a_n1319_5611# 0.00467f
C7942 XA.XIR[10].XIC[10].icell.SM VPWR 0.00158f
C7943 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.03424f
C7944 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.SM 0.00188f
C7945 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.03424f
C7946 XA.XIR[13].XIC[3].icell.PDM Iout 0.00112f
C7947 XThR.XTBN.Y XA.XIR[8].XIC_dummy_left.icell.Ien 0.00238f
C7948 XA.XIR[13].XIC[14].icell.SM VPWR 0.00208f
C7949 XThC.XTB5.Y data[3] 0.00931f
C7950 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PUM 0.00131f
C7951 XA.XIR[1].XIC[6].icell.SM Iout 0.00388f
C7952 XA.XIR[9].XIC[12].icell.SM Iout 0.00388f
C7953 XThR.Tn[3] XA.XIR[4].XIC[13].icell.SM 0.00121f
C7954 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.03424f
C7955 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02698f
C7956 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04522f
C7957 XThR.Tn[1] XA.XIR[1].XIC[11].icell.PDM 0.0033f
C7958 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01103f
C7959 XThR.Tn[5] XA.XIR[6].XIC[10].icell.SM 0.00121f
C7960 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00212f
C7961 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04522f
C7962 XA.XIR[9].XIC_15.icell.Ien Vbias 0.21343f
C7963 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PUM 0.00529f
C7964 XThR.Tn[11] XA.XIR[12].XIC[6].icell.SM 0.00121f
C7965 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04522f
C7966 XThR.Tn[9] XA.XIR[10].XIC[4].icell.Ien 0.00321f
C7967 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.SM 0.00383f
C7968 XA.XIR[15].XIC[7].icell.SM Vbias 0.00701f
C7969 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C7970 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04522f
C7971 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.03424f
C7972 XA.XIR[8].XIC[2].icell.PDM Vbias 0.04058f
C7973 XThR.Tn[4] XA.XIR[5].XIC[13].icell.SM 0.00121f
C7974 XA.XIR[7].XIC[13].icell.PUM VPWR 0.01036f
C7975 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PUM 0.00529f
C7976 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.SM 0.00383f
C7977 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.15089f
C7978 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04f
C7979 XA.XIR[5].XIC[0].icell.SM VPWR 0.00158f
C7980 XThC.Tn[3] XThR.Tn[4] 0.28062f
C7981 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.01406f
C7982 XA.XIR[1].XIC[14].icell.PUM VPWR 0.01036f
C7983 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PUM 0.00529f
C7984 XA.XIR[2].XIC[1].icell.Ien Vbias 0.21238f
C7985 XA.XIR[14].XIC[2].icell.Ien Vbias 0.21238f
C7986 XThR.Tn[7] Vbias 3.71582f
C7987 XA.XIR[4].XIC[3].icell.PUM VPWR 0.01036f
C7988 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.03424f
C7989 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PUM 0.00131f
C7990 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00529f
C7991 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.01406f
C7992 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00212f
C7993 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04522f
C7994 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00212f
C7995 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.SM 0.00188f
C7996 XA.XIR[13].XIC[4].icell.PUM Vbias 0.00347f
C7997 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.15089f
C7998 XA.XIR[3].XIC[6].icell.PDM VPWR 0.00863f
C7999 XThR.Tn[6] XA.XIR[7].XIC[4].icell.Ien 0.00321f
C8000 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04522f
C8001 XThR.Tn[8] XA.XIR[9].XIC[1].icell.SM 0.00121f
C8002 XA.XIR[12].XIC[5].icell.PUM Vbias 0.00347f
C8003 XThC.XTB3.Y a_4067_9615# 0.23056f
C8004 XA.XIR[3].XIC[3].icell.PDM Iout 0.00112f
C8005 XA.XIR[2].XIC[5].icell.SM VPWR 0.00158f
C8006 XA.XIR[13].XIC[12].icell.Ien VPWR 0.19065f
C8007 XA.XIR[14].XIC[6].icell.SM VPWR 0.00158f
C8008 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04522f
C8009 XA.XIR[15].XIC[12].icell.SM Vbias 0.00701f
C8010 XA.XIR[11].XIC[5].icell.SM Vbias 0.00701f
C8011 XA.XIR[2].XIC[2].icell.SM Iout 0.00388f
C8012 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.15089f
C8013 a_4067_9615# XThC.Tn[2] 0.27699f
C8014 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PUM 0.00131f
C8015 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C8016 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.SM 0.00188f
C8017 XA.XIR[14].XIC[3].icell.SM Iout 0.00388f
C8018 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.03424f
C8019 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13] 0.0033f
C8020 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00212f
C8021 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.03976f
C8022 XA.XIR[13].XIC[10].icell.PDM VPWR 0.00863f
C8023 XA.XIR[9].XIC[5].icell.Ien VPWR 0.19065f
C8024 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00529f
C8025 XA.XIR[10].XIC[9].icell.PDM Vbias 0.04058f
C8026 XA.XIR[6].XIC[5].icell.Ien Vbias 0.21238f
C8027 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04522f
C8028 XThC.Tn[1] Iout 0.84479f
C8029 XA.XIR[13].XIC[7].icell.PDM Iout 0.00112f
C8030 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.01406f
C8031 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PUM 0.00131f
C8032 XThC.XTB5.A XThC.XTB6.A 1.80461f
C8033 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01799f
C8034 XThR.Tn[0] XA.XIR[0].XIC_15.icell.PDM 0.0033f
C8035 XThC.Tn[13] XThR.Tn[11] 0.28063f
C8036 XA.XIR[5].XIC[6].icell.SM Vbias 0.00701f
C8037 XA.XIR[9].XIC[2].icell.Ien Iout 0.06483f
C8038 XThR.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.00321f
C8039 XA.XIR[7].XIC_dummy_right.icell.Ien Vbias 0.00287f
C8040 XA.XIR[0].XIC[1].icell.PDM VPWR 0.00806f
C8041 XA.XIR[12].XIC[14].icell.PDM Vbias 0.04058f
C8042 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02698f
C8043 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.SM 0.00383f
C8044 XA.XIR[12].XIC[8].icell.PDM Iout 0.00112f
C8045 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.SM 0.00188f
C8046 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00529f
C8047 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.15089f
C8048 XThR.Tn[2] XA.XIR[3].XIC[5].icell.SM 0.00121f
C8049 XA.XIR[4].XIC[9].icell.PUM Vbias 0.00347f
C8050 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.01406f
C8051 XA.XIR[12].XIC[9].icell.PUM Vbias 0.00347f
C8052 XA.XIR[6].XIC[9].icell.SM VPWR 0.00158f
C8053 XThR.Tn[2] XA.XIR[2].XIC[9].icell.PDM 0.0033f
C8054 XA.XIR[3].XIC[12].icell.PDM Vbias 0.04058f
C8055 XThR.Tn[13] XThR.Tn[14] 0.16991f
C8056 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.03424f
C8057 XA.XIR[8].XIC[4].icell.Ien Vbias 0.21238f
C8058 XA.XIR[6].XIC[6].icell.SM Iout 0.00388f
C8059 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11595f
C8060 XThR.Tn[4] XA.XIR[5].XIC[3].icell.Ien 0.00321f
C8061 XA.XIR[7].XIC[1].icell.SM VPWR 0.00158f
C8062 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.SM 0.00188f
C8063 XA.XIR[10].XIC_dummy_left.icell.Ien Vbias 0.00342f
C8064 XThC.XTB7.Y a_8739_9569# 0.00474f
C8065 XA.XIR[1].XIC[2].icell.SM VPWR 0.00158f
C8066 XA.XIR[13].XIC[11].icell.PDM Iout 0.00112f
C8067 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.03424f
C8068 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.03976f
C8069 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00212f
C8070 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.SM 0.00188f
C8071 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.SM 0.00383f
C8072 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C8073 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.SM 0.00188f
C8074 XA.XIR[4].XIC[12].icell.PDM Iout 0.00112f
C8075 XThC.XTB3.Y XThC.Tn[3] 0.01287f
C8076 XA.XIR[13].XIC[1].icell.PDM Vbias 0.04058f
C8077 XA.XIR[0].XIC[5].icell.PDM VPWR 0.00929f
C8078 XThR.Tn[6] XThR.Tn[7] 0.08065f
C8079 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04522f
C8080 XA.XIR[8].XIC[8].icell.SM VPWR 0.00158f
C8081 XThR.Tn[1] XA.XIR[1].XIC[4].icell.PDM 0.0033f
C8082 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Ien 0.00529f
C8083 XA.XIR[9].XIC[11].icell.Ien Vbias 0.21238f
C8084 XThR.Tn[12] XA.XIR[13].XIC[14].icell.SM 0.00121f
C8085 XThR.Tn[5] XA.XIR[6].XIC[3].icell.SM 0.00121f
C8086 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00212f
C8087 XA.XIR[11].XIC[0].icell.Ien VPWR 0.19066f
C8088 XThC.Tn[2] XThC.Tn[3] 0.34561f
C8089 XA.XIR[4].XIC[14].icell.PDM Vbias 0.04058f
C8090 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.SM 0.00188f
C8091 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00529f
C8092 XThC.Tn[9] XThR.Tn[2] 0.28062f
C8093 XA.XIR[12].XIC[14].icell.PUM Vbias 0.00347f
C8094 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.01406f
C8095 XThC.Tn[13] XThR.Tn[7] 0.28063f
C8096 XA.XIR[8].XIC[5].icell.SM Iout 0.00388f
C8097 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02698f
C8098 XA.XIR[6].XIC[14].icell.PUM VPWR 0.01036f
C8099 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.SM 0.00188f
C8100 XA.XIR[10].XIC[1].icell.Ien VPWR 0.19065f
C8101 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[9].icell.Ien 0.00212f
C8102 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.03424f
C8103 XThR.XTBN.Y a_n997_3979# 0.23021f
C8104 XA.XIR[3].XIC[14].icell.Ien Vbias 0.21238f
C8105 XA.XIR[15].XIC[0].icell.SM Vbias 0.00675f
C8106 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02698f
C8107 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.SM 0.00383f
C8108 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.SM 0.00383f
C8109 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.SM 0.00188f
C8110 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.SM 0.00383f
C8111 XA.XIR[10].XIC[11].icell.PUM VPWR 0.01036f
C8112 XA.XIR[5].XIC[14].icell.PDM Iout 0.00112f
C8113 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PUM 0.00529f
C8114 XThR.Tn[14] Vbias 3.71851f
C8115 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PUM 0.00131f
C8116 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.01406f
C8117 XA.XIR[7].XIC[7].icell.SM Vbias 0.00701f
C8118 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.15089f
C8119 XA.XIR[4].XIC[14].icell.Ien Iout 0.06483f
C8120 XA.XIR[5].XIC_15.icell.PUM Vbias 0.00347f
C8121 XA.XIR[1].XIC[8].icell.SM Vbias 0.00701f
C8122 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.15089f
C8123 XA.XIR[13].XIC[10].icell.SM VPWR 0.00158f
C8124 XA.XIR[8].XIC[13].icell.PUM VPWR 0.01036f
C8125 XA.XIR[9].XIC[0].icell.Ien Vbias 0.21102f
C8126 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02698f
C8127 XA.XIR[15].XIC[6].icell.PUM VPWR 0.01036f
C8128 XThR.Tn[14] XA.XIR[14].XIC[6].icell.PDM 0.0033f
C8129 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.15089f
C8130 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PUM 0.00131f
C8131 XThR.XTB1.Y VPWR 1.12978f
C8132 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04522f
C8133 XThC.XTB2.Y a_3523_10575# 0.01006f
C8134 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00529f
C8135 XThR.Tn[13] XA.XIR[14].XIC[5].icell.SM 0.00121f
C8136 XA.XIR[0].XIC[11].icell.PDM Vbias 0.04065f
C8137 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13469f
C8138 XA.XIR[3].XIC[1].icell.PDM Vbias 0.04058f
C8139 XThC.XTB7.Y XThC.Tn[11] 0.07471f
C8140 XA.XIR[12].XIC[14].icell.SM Vbias 0.00701f
C8141 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.SM 0.00188f
C8142 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04522f
C8143 XThR.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.00321f
C8144 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PUM 0.00529f
C8145 XThR.Tn[13] XA.XIR[13].XIC[9].icell.PDM 0.0033f
C8146 XA.XIR[10].XIC_15.icell.SM VPWR 0.00276f
C8147 XThR.Tn[0] XA.XIR[1].XIC[5].icell.SM 0.00121f
C8148 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.03424f
C8149 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.SM 0.00383f
C8150 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PUM 0.00529f
C8151 XA.XIR[1].XIC[1].icell.PDM Iout 0.00112f
C8152 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00212f
C8153 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.03976f
C8154 XA.XIR[7].XIC[12].icell.PUM Vbias 0.00347f
C8155 XA.XIR[12].XIC[4].icell.PDM VPWR 0.00863f
C8156 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.SM 0.00383f
C8157 XA.XIR[0].XIC[14].icell.Ien VPWR 0.19008f
C8158 XThR.Tn[9] Iout 1.16627f
C8159 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00212f
C8160 XThR.Tn[0] XA.XIR[0].XIC[8].icell.PDM 0.0033f
C8161 XA.XIR[4].XIC[1].icell.PDM Iout 0.00112f
C8162 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.SM 0.00188f
C8163 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PUM 0.00529f
C8164 XA.XIR[5].XIC[2].icell.PDM Vbias 0.04058f
C8165 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02734f
C8166 XA.XIR[11].XIC[4].icell.PUM VPWR 0.01036f
C8167 XA.XIR[1].XIC[13].icell.PUM Vbias 0.00347f
C8168 XA.XIR[0].XIC[11].icell.Ien Iout 0.06455f
C8169 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00212f
C8170 XThR.Tn[11] a_n997_2667# 0.19413f
C8171 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.03424f
C8172 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.SM 0.00383f
C8173 XA.XIR[4].XIC[2].icell.PUM Vbias 0.00347f
C8174 XA.XIR[10].XIC[5].icell.Ien VPWR 0.19065f
C8175 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00212f
C8176 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.SM 0.00188f
C8177 XA.XIR[15].XIC[13].icell.PUM Vbias 0.00347f
C8178 XA.XIR[6].XIC[2].icell.SM VPWR 0.00158f
C8179 XThR.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.0033f
C8180 XThR.Tn[9] XA.XIR[10].XIC[7].icell.SM 0.00121f
C8181 XA.XIR[3].XIC[5].icell.PDM Vbias 0.04058f
C8182 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01402f
C8183 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.SM 0.00188f
C8184 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00212f
C8185 XA.XIR[10].XIC[2].icell.Ien Iout 0.06483f
C8186 XThC.XTB5.A XThC.Tn[8] 0.00205f
C8187 XA.XIR[5].XIC[5].icell.PUM VPWR 0.01036f
C8188 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.SM 0.00383f
C8189 XA.XIR[8].XIC_dummy_right.icell.Ien Vbias 0.00287f
C8190 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02698f
C8191 XThR.Tn[2] XThR.XTB4.Y 0.0021f
C8192 XA.XIR[2].XIC[4].icell.SM Vbias 0.00701f
C8193 XA.XIR[7].XIC_15.icell.PDM Iout 0.0013f
C8194 XA.XIR[14].XIC[5].icell.SM Vbias 0.00701f
C8195 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00212f
C8196 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.SM 0.00188f
C8197 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.01406f
C8198 XA.XIR[4].XIC[8].icell.PDM VPWR 0.00863f
C8199 XThC.Tn[5] VPWR 5.95818f
C8200 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00529f
C8201 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.03424f
C8202 XA.XIR[12].XIC[12].icell.Ien Vbias 0.21238f
C8203 XA.XIR[13].XIC[9].icell.PDM Vbias 0.04058f
C8204 XA.XIR[4].XIC[5].icell.PDM Iout 0.00112f
C8205 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.SM 0.00383f
C8206 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04522f
C8207 XA.XIR[3].XIC[8].icell.Ien VPWR 0.19065f
C8208 XThR.Tn[6] XA.XIR[7].XIC[7].icell.SM 0.00121f
C8209 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.03424f
C8210 XA.XIR[9].XIC[4].icell.Ien Vbias 0.21238f
C8211 XA.XIR[8].XIC[1].icell.SM VPWR 0.00158f
C8212 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PUM 0.00131f
C8213 XA.XIR[0].XIC_15.icell.Ien Iout 0.06455f
C8214 XThR.Tn[14] XA.XIR[14].XIC_15.icell.PDM 0.0033f
C8215 XA.XIR[3].XIC[5].icell.Ien Iout 0.06483f
C8216 XA.XIR[14].XIC[0].icell.PDM VPWR 0.00863f
C8217 XA.XIR[12].XIC[10].icell.PDM Vbias 0.04058f
C8218 XThC.Tn[13] XThR.Tn[14] 0.28063f
C8219 XThC.Tn[11] XThR.Tn[0] 0.28077f
C8220 XA.XIR[2].XIC[10].icell.PUM VPWR 0.01036f
C8221 data[7] VGND 0.49949f
C8222 data[6] VGND 0.47974f
C8223 data[4] VGND 0.59317f
C8224 data[5] VGND 1.17814f
C8225 Iout VGND 0.31933p
C8226 data[3] VGND 0.49912f
C8227 data[2] VGND 0.48064f
C8228 data[0] VGND 0.59421f
C8229 data[1] VGND 1.17844f
C8230 bias[2] VGND 0.77552f
C8231 bias[0] VGND 1.22004f
C8232 Vbias VGND 0.22928p
C8233 bias[1] VGND 0.62458f
C8234 VPWR VGND 0.33989p
C8235 a_n997_715# VGND 0.5638f
C8236 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.74784f
C8237 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70255f
C8238 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C8239 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64161f
C8240 XA.XIR[15].XIC_15.icell.SM VGND 0.00474f
C8241 XA.XIR[15].XIC_dummy_right.icell.PUM VGND 0.00226f
C8242 XA.XIR[15].XIC_15.icell.Ien VGND 0.43984f
C8243 XA.XIR[15].XIC[14].icell.SM VGND 0.00502f
C8244 XA.XIR[15].XIC_15.icell.PUM VGND 0.00284f
C8245 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.22893f
C8246 XA.XIR[15].XIC[14].icell.Ien VGND 0.44037f
C8247 XA.XIR[15].XIC[13].icell.SM VGND 0.00502f
C8248 XA.XIR[15].XIC[14].icell.PUM VGND 0.00301f
C8249 XA.XIR[15].XIC_15.icell.PDM VGND 0.18566f
C8250 XA.XIR[15].XIC[13].icell.Ien VGND 0.44037f
C8251 XA.XIR[15].XIC[12].icell.SM VGND 0.00502f
C8252 XA.XIR[15].XIC[13].icell.PUM VGND 0.00301f
C8253 XA.XIR[15].XIC[14].icell.PDM VGND 0.18513f
C8254 XA.XIR[15].XIC[12].icell.Ien VGND 0.44037f
C8255 XA.XIR[15].XIC[11].icell.SM VGND 0.00502f
C8256 XA.XIR[15].XIC[12].icell.PUM VGND 0.00301f
C8257 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85333f
C8258 XA.XIR[15].XIC[13].icell.PDM VGND 0.18513f
C8259 XA.XIR[15].XIC[11].icell.Ien VGND 0.44037f
C8260 XA.XIR[15].XIC[10].icell.SM VGND 0.00502f
C8261 XA.XIR[15].XIC[11].icell.PUM VGND 0.00301f
C8262 XA.XIR[15].XIC[12].icell.PDM VGND 0.18513f
C8263 XA.XIR[15].XIC[10].icell.Ien VGND 0.44037f
C8264 XA.XIR[15].XIC[9].icell.SM VGND 0.00502f
C8265 XA.XIR[15].XIC[10].icell.PUM VGND 0.00301f
C8266 XA.XIR[15].XIC[11].icell.PDM VGND 0.18513f
C8267 XA.XIR[15].XIC[9].icell.Ien VGND 0.44037f
C8268 XA.XIR[15].XIC[8].icell.SM VGND 0.00502f
C8269 XA.XIR[15].XIC[9].icell.PUM VGND 0.00301f
C8270 XA.XIR[15].XIC[10].icell.PDM VGND 0.18513f
C8271 XA.XIR[15].XIC[8].icell.Ien VGND 0.44037f
C8272 XA.XIR[15].XIC[7].icell.SM VGND 0.00502f
C8273 XA.XIR[15].XIC[8].icell.PUM VGND 0.00301f
C8274 XA.XIR[15].XIC[9].icell.PDM VGND 0.18513f
C8275 XA.XIR[15].XIC[7].icell.Ien VGND 0.44037f
C8276 XA.XIR[15].XIC[6].icell.SM VGND 0.00502f
C8277 XA.XIR[15].XIC[7].icell.PUM VGND 0.00301f
C8278 XA.XIR[15].XIC[8].icell.PDM VGND 0.18513f
C8279 XA.XIR[15].XIC[6].icell.Ien VGND 0.44037f
C8280 XA.XIR[15].XIC[5].icell.SM VGND 0.00502f
C8281 XA.XIR[15].XIC[6].icell.PUM VGND 0.00301f
C8282 XA.XIR[15].XIC[7].icell.PDM VGND 0.18513f
C8283 XA.XIR[15].XIC[5].icell.Ien VGND 0.44037f
C8284 XA.XIR[15].XIC[4].icell.SM VGND 0.00502f
C8285 XA.XIR[15].XIC[5].icell.PUM VGND 0.00301f
C8286 XA.XIR[15].XIC[6].icell.PDM VGND 0.18513f
C8287 XA.XIR[15].XIC[4].icell.Ien VGND 0.44037f
C8288 XA.XIR[15].XIC[3].icell.SM VGND 0.00502f
C8289 XA.XIR[15].XIC[4].icell.PUM VGND 0.00301f
C8290 XA.XIR[15].XIC[5].icell.PDM VGND 0.18513f
C8291 XA.XIR[15].XIC[3].icell.Ien VGND 0.44037f
C8292 XA.XIR[15].XIC[2].icell.SM VGND 0.00502f
C8293 XA.XIR[15].XIC[3].icell.PUM VGND 0.00301f
C8294 XA.XIR[15].XIC[4].icell.PDM VGND 0.18513f
C8295 XA.XIR[15].XIC[2].icell.Ien VGND 0.44037f
C8296 XA.XIR[15].XIC[1].icell.SM VGND 0.00502f
C8297 XA.XIR[15].XIC[2].icell.PUM VGND 0.00301f
C8298 XA.XIR[15].XIC[3].icell.PDM VGND 0.18513f
C8299 XA.XIR[15].XIC[1].icell.Ien VGND 0.44037f
C8300 XA.XIR[15].XIC[0].icell.SM VGND 0.00502f
C8301 XA.XIR[15].XIC[1].icell.PUM VGND 0.00301f
C8302 XA.XIR[15].XIC[2].icell.PDM VGND 0.18513f
C8303 XA.XIR[15].XIC[0].icell.Ien VGND 0.44058f
C8304 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01043f
C8305 XA.XIR[15].XIC[0].icell.PUM VGND 0.00549f
C8306 XA.XIR[15].XIC[1].icell.PDM VGND 0.18513f
C8307 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.60728f
C8308 XA.XIR[15].XIC_dummy_left.icell.PUM VGND 0.00226f
C8309 XA.XIR[15].XIC[0].icell.PDM VGND 0.18522f
C8310 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22263f
C8311 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80232f
C8312 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C8313 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.6141f
C8314 XA.XIR[14].XIC_15.icell.SM VGND 0.00474f
C8315 XA.XIR[14].XIC_dummy_right.icell.PUM VGND 0.00226f
C8316 XA.XIR[14].XIC_15.icell.Ien VGND 0.37606f
C8317 XA.XIR[14].XIC[14].icell.SM VGND 0.00502f
C8318 XA.XIR[14].XIC_15.icell.PUM VGND 0.00284f
C8319 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23008f
C8320 XA.XIR[14].XIC[14].icell.Ien VGND 0.37698f
C8321 XA.XIR[14].XIC[13].icell.SM VGND 0.00502f
C8322 XA.XIR[14].XIC[14].icell.PUM VGND 0.00301f
C8323 XA.XIR[14].XIC_15.icell.PDM VGND 0.18645f
C8324 XA.XIR[14].XIC[13].icell.Ien VGND 0.37698f
C8325 XA.XIR[14].XIC[12].icell.SM VGND 0.00502f
C8326 XA.XIR[14].XIC[13].icell.PUM VGND 0.00301f
C8327 XA.XIR[14].XIC[14].icell.PDM VGND 0.18592f
C8328 XA.XIR[14].XIC[12].icell.Ien VGND 0.37698f
C8329 XA.XIR[14].XIC[11].icell.SM VGND 0.00502f
C8330 XA.XIR[14].XIC[12].icell.PUM VGND 0.00301f
C8331 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85333f
C8332 XA.XIR[14].XIC[13].icell.PDM VGND 0.18592f
C8333 XA.XIR[14].XIC[11].icell.Ien VGND 0.37698f
C8334 XA.XIR[14].XIC[10].icell.SM VGND 0.00502f
C8335 XA.XIR[14].XIC[11].icell.PUM VGND 0.00301f
C8336 XA.XIR[14].XIC[12].icell.PDM VGND 0.18592f
C8337 XA.XIR[14].XIC[10].icell.Ien VGND 0.37698f
C8338 XA.XIR[14].XIC[9].icell.SM VGND 0.00502f
C8339 XA.XIR[14].XIC[10].icell.PUM VGND 0.00301f
C8340 XA.XIR[14].XIC[11].icell.PDM VGND 0.18592f
C8341 XA.XIR[14].XIC[9].icell.Ien VGND 0.37698f
C8342 XA.XIR[14].XIC[8].icell.SM VGND 0.00502f
C8343 XA.XIR[14].XIC[9].icell.PUM VGND 0.00301f
C8344 XA.XIR[14].XIC[10].icell.PDM VGND 0.18592f
C8345 XA.XIR[14].XIC[8].icell.Ien VGND 0.37698f
C8346 XA.XIR[14].XIC[7].icell.SM VGND 0.00502f
C8347 XA.XIR[14].XIC[8].icell.PUM VGND 0.00301f
C8348 XA.XIR[14].XIC[9].icell.PDM VGND 0.18592f
C8349 XA.XIR[14].XIC[7].icell.Ien VGND 0.37698f
C8350 XA.XIR[14].XIC[6].icell.SM VGND 0.00502f
C8351 XA.XIR[14].XIC[7].icell.PUM VGND 0.00301f
C8352 XA.XIR[14].XIC[8].icell.PDM VGND 0.18592f
C8353 XA.XIR[14].XIC[6].icell.Ien VGND 0.37698f
C8354 XA.XIR[14].XIC[5].icell.SM VGND 0.00502f
C8355 XA.XIR[14].XIC[6].icell.PUM VGND 0.00301f
C8356 XA.XIR[14].XIC[7].icell.PDM VGND 0.18592f
C8357 XA.XIR[14].XIC[5].icell.Ien VGND 0.37698f
C8358 XA.XIR[14].XIC[4].icell.SM VGND 0.00502f
C8359 XA.XIR[14].XIC[5].icell.PUM VGND 0.00301f
C8360 XA.XIR[14].XIC[6].icell.PDM VGND 0.18592f
C8361 XA.XIR[14].XIC[4].icell.Ien VGND 0.37698f
C8362 XA.XIR[14].XIC[3].icell.SM VGND 0.00502f
C8363 XA.XIR[14].XIC[4].icell.PUM VGND 0.00301f
C8364 XA.XIR[14].XIC[5].icell.PDM VGND 0.18592f
C8365 XA.XIR[14].XIC[3].icell.Ien VGND 0.37698f
C8366 XA.XIR[14].XIC[2].icell.SM VGND 0.00502f
C8367 XA.XIR[14].XIC[3].icell.PUM VGND 0.00301f
C8368 XA.XIR[14].XIC[4].icell.PDM VGND 0.18592f
C8369 XA.XIR[14].XIC[2].icell.Ien VGND 0.37698f
C8370 XA.XIR[14].XIC[1].icell.SM VGND 0.00502f
C8371 XThR.Tn[14] VGND 14.00401f
C8372 XA.XIR[14].XIC[2].icell.PUM VGND 0.00301f
C8373 XA.XIR[14].XIC[3].icell.PDM VGND 0.18592f
C8374 XA.XIR[14].XIC[1].icell.Ien VGND 0.37698f
C8375 XA.XIR[14].XIC[0].icell.SM VGND 0.00502f
C8376 a_n997_1579# VGND 0.54776f
C8377 XA.XIR[14].XIC[1].icell.PUM VGND 0.00301f
C8378 XA.XIR[14].XIC[2].icell.PDM VGND 0.18592f
C8379 XA.XIR[14].XIC[0].icell.Ien VGND 0.3772f
C8380 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01043f
C8381 XA.XIR[14].XIC[0].icell.PUM VGND 0.00549f
C8382 XA.XIR[14].XIC[1].icell.PDM VGND 0.18592f
C8383 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.58213f
C8384 XA.XIR[14].XIC_dummy_left.icell.PUM VGND 0.00226f
C8385 XA.XIR[14].XIC[0].icell.PDM VGND 0.18601f
C8386 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22378f
C8387 a_n997_1803# VGND 0.53618f
C8388 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.80236f
C8389 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C8390 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.6141f
C8391 XA.XIR[13].XIC_15.icell.SM VGND 0.00474f
C8392 XA.XIR[13].XIC_dummy_right.icell.PUM VGND 0.00226f
C8393 XA.XIR[13].XIC_15.icell.Ien VGND 0.37606f
C8394 XA.XIR[13].XIC[14].icell.SM VGND 0.00502f
C8395 XA.XIR[13].XIC_15.icell.PUM VGND 0.00284f
C8396 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23008f
C8397 XA.XIR[13].XIC[14].icell.Ien VGND 0.37698f
C8398 XA.XIR[13].XIC[13].icell.SM VGND 0.00502f
C8399 XA.XIR[13].XIC[14].icell.PUM VGND 0.00301f
C8400 XA.XIR[13].XIC_15.icell.PDM VGND 0.18645f
C8401 XA.XIR[13].XIC[13].icell.Ien VGND 0.37698f
C8402 XA.XIR[13].XIC[12].icell.SM VGND 0.00502f
C8403 XA.XIR[13].XIC[13].icell.PUM VGND 0.00301f
C8404 XA.XIR[13].XIC[14].icell.PDM VGND 0.18592f
C8405 XA.XIR[13].XIC[12].icell.Ien VGND 0.37698f
C8406 XA.XIR[13].XIC[11].icell.SM VGND 0.00502f
C8407 XA.XIR[13].XIC[12].icell.PUM VGND 0.00301f
C8408 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85333f
C8409 XA.XIR[13].XIC[13].icell.PDM VGND 0.18592f
C8410 XA.XIR[13].XIC[11].icell.Ien VGND 0.37698f
C8411 XA.XIR[13].XIC[10].icell.SM VGND 0.00502f
C8412 XA.XIR[13].XIC[11].icell.PUM VGND 0.00301f
C8413 XA.XIR[13].XIC[12].icell.PDM VGND 0.18592f
C8414 XA.XIR[13].XIC[10].icell.Ien VGND 0.37698f
C8415 XA.XIR[13].XIC[9].icell.SM VGND 0.00502f
C8416 XA.XIR[13].XIC[10].icell.PUM VGND 0.00301f
C8417 XA.XIR[13].XIC[11].icell.PDM VGND 0.18592f
C8418 XA.XIR[13].XIC[9].icell.Ien VGND 0.37698f
C8419 XA.XIR[13].XIC[8].icell.SM VGND 0.00502f
C8420 XA.XIR[13].XIC[9].icell.PUM VGND 0.00301f
C8421 XA.XIR[13].XIC[10].icell.PDM VGND 0.18592f
C8422 XA.XIR[13].XIC[8].icell.Ien VGND 0.37698f
C8423 XA.XIR[13].XIC[7].icell.SM VGND 0.00502f
C8424 XA.XIR[13].XIC[8].icell.PUM VGND 0.00301f
C8425 XA.XIR[13].XIC[9].icell.PDM VGND 0.18592f
C8426 XA.XIR[13].XIC[7].icell.Ien VGND 0.37698f
C8427 XA.XIR[13].XIC[6].icell.SM VGND 0.00502f
C8428 XA.XIR[13].XIC[7].icell.PUM VGND 0.00301f
C8429 XA.XIR[13].XIC[8].icell.PDM VGND 0.18592f
C8430 XA.XIR[13].XIC[6].icell.Ien VGND 0.37698f
C8431 XA.XIR[13].XIC[5].icell.SM VGND 0.00502f
C8432 XA.XIR[13].XIC[6].icell.PUM VGND 0.00301f
C8433 XA.XIR[13].XIC[7].icell.PDM VGND 0.18592f
C8434 XA.XIR[13].XIC[5].icell.Ien VGND 0.37698f
C8435 XA.XIR[13].XIC[4].icell.SM VGND 0.00502f
C8436 XA.XIR[13].XIC[5].icell.PUM VGND 0.00301f
C8437 XA.XIR[13].XIC[6].icell.PDM VGND 0.18592f
C8438 XA.XIR[13].XIC[4].icell.Ien VGND 0.37698f
C8439 XA.XIR[13].XIC[3].icell.SM VGND 0.00502f
C8440 XA.XIR[13].XIC[4].icell.PUM VGND 0.00301f
C8441 XA.XIR[13].XIC[5].icell.PDM VGND 0.18592f
C8442 XA.XIR[13].XIC[3].icell.Ien VGND 0.37698f
C8443 XA.XIR[13].XIC[2].icell.SM VGND 0.00502f
C8444 XA.XIR[13].XIC[3].icell.PUM VGND 0.00301f
C8445 XA.XIR[13].XIC[4].icell.PDM VGND 0.18592f
C8446 XA.XIR[13].XIC[2].icell.Ien VGND 0.37698f
C8447 XA.XIR[13].XIC[1].icell.SM VGND 0.00502f
C8448 XThR.Tn[13] VGND 13.88476f
C8449 XA.XIR[13].XIC[2].icell.PUM VGND 0.00301f
C8450 XA.XIR[13].XIC[3].icell.PDM VGND 0.18592f
C8451 XA.XIR[13].XIC[1].icell.Ien VGND 0.37698f
C8452 XA.XIR[13].XIC[0].icell.SM VGND 0.00502f
C8453 XA.XIR[13].XIC[1].icell.PUM VGND 0.00301f
C8454 XA.XIR[13].XIC[2].icell.PDM VGND 0.18592f
C8455 XA.XIR[13].XIC[0].icell.Ien VGND 0.3772f
C8456 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01043f
C8457 XA.XIR[13].XIC[0].icell.PUM VGND 0.00549f
C8458 XA.XIR[13].XIC[1].icell.PDM VGND 0.18592f
C8459 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.58069f
C8460 XA.XIR[13].XIC_dummy_left.icell.PUM VGND 0.00226f
C8461 XA.XIR[13].XIC[0].icell.PDM VGND 0.18601f
C8462 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22378f
C8463 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80102f
C8464 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C8465 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.6141f
C8466 XA.XIR[12].XIC_15.icell.SM VGND 0.00474f
C8467 XA.XIR[12].XIC_dummy_right.icell.PUM VGND 0.00226f
C8468 XA.XIR[12].XIC_15.icell.Ien VGND 0.37606f
C8469 XA.XIR[12].XIC[14].icell.SM VGND 0.00502f
C8470 XA.XIR[12].XIC_15.icell.PUM VGND 0.00284f
C8471 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23008f
C8472 XA.XIR[12].XIC[14].icell.Ien VGND 0.37698f
C8473 XA.XIR[12].XIC[13].icell.SM VGND 0.00502f
C8474 XA.XIR[12].XIC[14].icell.PUM VGND 0.00301f
C8475 XA.XIR[12].XIC_15.icell.PDM VGND 0.18645f
C8476 XA.XIR[12].XIC[13].icell.Ien VGND 0.37698f
C8477 XA.XIR[12].XIC[12].icell.SM VGND 0.00502f
C8478 XA.XIR[12].XIC[13].icell.PUM VGND 0.00301f
C8479 XA.XIR[12].XIC[14].icell.PDM VGND 0.18592f
C8480 XA.XIR[12].XIC[12].icell.Ien VGND 0.37698f
C8481 XA.XIR[12].XIC[11].icell.SM VGND 0.00502f
C8482 XA.XIR[12].XIC[12].icell.PUM VGND 0.00301f
C8483 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85333f
C8484 XA.XIR[12].XIC[13].icell.PDM VGND 0.18592f
C8485 XA.XIR[12].XIC[11].icell.Ien VGND 0.37698f
C8486 XA.XIR[12].XIC[10].icell.SM VGND 0.00502f
C8487 XA.XIR[12].XIC[11].icell.PUM VGND 0.00301f
C8488 XA.XIR[12].XIC[12].icell.PDM VGND 0.18592f
C8489 XA.XIR[12].XIC[10].icell.Ien VGND 0.37698f
C8490 XA.XIR[12].XIC[9].icell.SM VGND 0.00502f
C8491 XA.XIR[12].XIC[10].icell.PUM VGND 0.00301f
C8492 XA.XIR[12].XIC[11].icell.PDM VGND 0.18592f
C8493 XA.XIR[12].XIC[9].icell.Ien VGND 0.37698f
C8494 XA.XIR[12].XIC[8].icell.SM VGND 0.00502f
C8495 XA.XIR[12].XIC[9].icell.PUM VGND 0.00301f
C8496 XA.XIR[12].XIC[10].icell.PDM VGND 0.18592f
C8497 XA.XIR[12].XIC[8].icell.Ien VGND 0.37698f
C8498 XA.XIR[12].XIC[7].icell.SM VGND 0.00502f
C8499 XA.XIR[12].XIC[8].icell.PUM VGND 0.00301f
C8500 XA.XIR[12].XIC[9].icell.PDM VGND 0.18592f
C8501 XA.XIR[12].XIC[7].icell.Ien VGND 0.37698f
C8502 XA.XIR[12].XIC[6].icell.SM VGND 0.00502f
C8503 XA.XIR[12].XIC[7].icell.PUM VGND 0.00301f
C8504 XA.XIR[12].XIC[8].icell.PDM VGND 0.18592f
C8505 XA.XIR[12].XIC[6].icell.Ien VGND 0.37698f
C8506 XA.XIR[12].XIC[5].icell.SM VGND 0.00502f
C8507 XA.XIR[12].XIC[6].icell.PUM VGND 0.00301f
C8508 XA.XIR[12].XIC[7].icell.PDM VGND 0.18592f
C8509 XA.XIR[12].XIC[5].icell.Ien VGND 0.37698f
C8510 XA.XIR[12].XIC[4].icell.SM VGND 0.00502f
C8511 XA.XIR[12].XIC[5].icell.PUM VGND 0.00301f
C8512 XA.XIR[12].XIC[6].icell.PDM VGND 0.18592f
C8513 XA.XIR[12].XIC[4].icell.Ien VGND 0.37698f
C8514 XA.XIR[12].XIC[3].icell.SM VGND 0.00502f
C8515 XA.XIR[12].XIC[4].icell.PUM VGND 0.00301f
C8516 XA.XIR[12].XIC[5].icell.PDM VGND 0.18592f
C8517 XA.XIR[12].XIC[3].icell.Ien VGND 0.37698f
C8518 XA.XIR[12].XIC[2].icell.SM VGND 0.00502f
C8519 XA.XIR[12].XIC[3].icell.PUM VGND 0.00301f
C8520 XA.XIR[12].XIC[4].icell.PDM VGND 0.18592f
C8521 XA.XIR[12].XIC[2].icell.Ien VGND 0.37698f
C8522 XA.XIR[12].XIC[1].icell.SM VGND 0.00502f
C8523 XThR.Tn[12] VGND 13.77499f
C8524 XA.XIR[12].XIC[2].icell.PUM VGND 0.00301f
C8525 XA.XIR[12].XIC[3].icell.PDM VGND 0.18592f
C8526 XA.XIR[12].XIC[1].icell.Ien VGND 0.37698f
C8527 XA.XIR[12].XIC[0].icell.SM VGND 0.00502f
C8528 XA.XIR[12].XIC[1].icell.PUM VGND 0.00301f
C8529 XA.XIR[12].XIC[2].icell.PDM VGND 0.18592f
C8530 XA.XIR[12].XIC[0].icell.Ien VGND 0.3772f
C8531 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01043f
C8532 XA.XIR[12].XIC[0].icell.PUM VGND 0.00549f
C8533 XA.XIR[12].XIC[1].icell.PDM VGND 0.18592f
C8534 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.57898f
C8535 XA.XIR[12].XIC_dummy_left.icell.PUM VGND 0.00226f
C8536 XA.XIR[12].XIC[0].icell.PDM VGND 0.18601f
C8537 a_n997_2667# VGND 0.54569f
C8538 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22378f
C8539 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.80337f
C8540 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C8541 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.6141f
C8542 XA.XIR[11].XIC_15.icell.SM VGND 0.00474f
C8543 XA.XIR[11].XIC_dummy_right.icell.PUM VGND 0.00226f
C8544 XA.XIR[11].XIC_15.icell.Ien VGND 0.37606f
C8545 XA.XIR[11].XIC[14].icell.SM VGND 0.00502f
C8546 XA.XIR[11].XIC_15.icell.PUM VGND 0.00284f
C8547 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23008f
C8548 XA.XIR[11].XIC[14].icell.Ien VGND 0.37698f
C8549 XA.XIR[11].XIC[13].icell.SM VGND 0.00502f
C8550 XA.XIR[11].XIC[14].icell.PUM VGND 0.00301f
C8551 XA.XIR[11].XIC_15.icell.PDM VGND 0.18645f
C8552 XA.XIR[11].XIC[13].icell.Ien VGND 0.37698f
C8553 XA.XIR[11].XIC[12].icell.SM VGND 0.00502f
C8554 XA.XIR[11].XIC[13].icell.PUM VGND 0.00301f
C8555 XA.XIR[11].XIC[14].icell.PDM VGND 0.18592f
C8556 XA.XIR[11].XIC[12].icell.Ien VGND 0.37698f
C8557 XA.XIR[11].XIC[11].icell.SM VGND 0.00502f
C8558 XA.XIR[11].XIC[12].icell.PUM VGND 0.00301f
C8559 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85333f
C8560 XA.XIR[11].XIC[13].icell.PDM VGND 0.18592f
C8561 XA.XIR[11].XIC[11].icell.Ien VGND 0.37698f
C8562 XA.XIR[11].XIC[10].icell.SM VGND 0.00502f
C8563 XA.XIR[11].XIC[11].icell.PUM VGND 0.00301f
C8564 XA.XIR[11].XIC[12].icell.PDM VGND 0.18592f
C8565 XA.XIR[11].XIC[10].icell.Ien VGND 0.37698f
C8566 XA.XIR[11].XIC[9].icell.SM VGND 0.00502f
C8567 XA.XIR[11].XIC[10].icell.PUM VGND 0.00301f
C8568 XA.XIR[11].XIC[11].icell.PDM VGND 0.18592f
C8569 XA.XIR[11].XIC[9].icell.Ien VGND 0.37698f
C8570 XA.XIR[11].XIC[8].icell.SM VGND 0.00502f
C8571 XA.XIR[11].XIC[9].icell.PUM VGND 0.00301f
C8572 XA.XIR[11].XIC[10].icell.PDM VGND 0.18592f
C8573 XA.XIR[11].XIC[8].icell.Ien VGND 0.37698f
C8574 XA.XIR[11].XIC[7].icell.SM VGND 0.00502f
C8575 XA.XIR[11].XIC[8].icell.PUM VGND 0.00301f
C8576 XA.XIR[11].XIC[9].icell.PDM VGND 0.18592f
C8577 XA.XIR[11].XIC[7].icell.Ien VGND 0.37698f
C8578 XA.XIR[11].XIC[6].icell.SM VGND 0.00502f
C8579 XA.XIR[11].XIC[7].icell.PUM VGND 0.00301f
C8580 XA.XIR[11].XIC[8].icell.PDM VGND 0.18592f
C8581 XA.XIR[11].XIC[6].icell.Ien VGND 0.37698f
C8582 XA.XIR[11].XIC[5].icell.SM VGND 0.00502f
C8583 XA.XIR[11].XIC[6].icell.PUM VGND 0.00301f
C8584 XA.XIR[11].XIC[7].icell.PDM VGND 0.18592f
C8585 XA.XIR[11].XIC[5].icell.Ien VGND 0.37698f
C8586 XA.XIR[11].XIC[4].icell.SM VGND 0.00502f
C8587 XA.XIR[11].XIC[5].icell.PUM VGND 0.00301f
C8588 XA.XIR[11].XIC[6].icell.PDM VGND 0.18592f
C8589 XA.XIR[11].XIC[4].icell.Ien VGND 0.37698f
C8590 XA.XIR[11].XIC[3].icell.SM VGND 0.00502f
C8591 XA.XIR[11].XIC[4].icell.PUM VGND 0.00301f
C8592 XA.XIR[11].XIC[5].icell.PDM VGND 0.18592f
C8593 XA.XIR[11].XIC[3].icell.Ien VGND 0.37698f
C8594 XA.XIR[11].XIC[2].icell.SM VGND 0.00502f
C8595 XA.XIR[11].XIC[3].icell.PUM VGND 0.00301f
C8596 XA.XIR[11].XIC[4].icell.PDM VGND 0.18592f
C8597 XA.XIR[11].XIC[2].icell.Ien VGND 0.37698f
C8598 XA.XIR[11].XIC[1].icell.SM VGND 0.00502f
C8599 XThR.Tn[11] VGND 13.83609f
C8600 XA.XIR[11].XIC[2].icell.PUM VGND 0.00301f
C8601 XA.XIR[11].XIC[3].icell.PDM VGND 0.18592f
C8602 XA.XIR[11].XIC[1].icell.Ien VGND 0.37698f
C8603 XA.XIR[11].XIC[0].icell.SM VGND 0.00502f
C8604 a_n997_2891# VGND 0.54779f
C8605 a_n1331_2891# VGND 0.00194f
C8606 XA.XIR[11].XIC[1].icell.PUM VGND 0.00301f
C8607 XA.XIR[11].XIC[2].icell.PDM VGND 0.18592f
C8608 XA.XIR[11].XIC[0].icell.Ien VGND 0.3772f
C8609 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01043f
C8610 XA.XIR[11].XIC[0].icell.PUM VGND 0.00549f
C8611 XA.XIR[11].XIC[1].icell.PDM VGND 0.18592f
C8612 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57909f
C8613 XA.XIR[11].XIC_dummy_left.icell.PUM VGND 0.00226f
C8614 XA.XIR[11].XIC[0].icell.PDM VGND 0.18601f
C8615 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22378f
C8616 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80221f
C8617 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C8618 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.6141f
C8619 XA.XIR[10].XIC_15.icell.SM VGND 0.00474f
C8620 XA.XIR[10].XIC_dummy_right.icell.PUM VGND 0.00226f
C8621 XA.XIR[10].XIC_15.icell.Ien VGND 0.37606f
C8622 XA.XIR[10].XIC[14].icell.SM VGND 0.00502f
C8623 XA.XIR[10].XIC_15.icell.PUM VGND 0.00284f
C8624 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23008f
C8625 XA.XIR[10].XIC[14].icell.Ien VGND 0.37698f
C8626 XA.XIR[10].XIC[13].icell.SM VGND 0.00502f
C8627 XA.XIR[10].XIC[14].icell.PUM VGND 0.00301f
C8628 XA.XIR[10].XIC_15.icell.PDM VGND 0.18645f
C8629 XA.XIR[10].XIC[13].icell.Ien VGND 0.37698f
C8630 XA.XIR[10].XIC[12].icell.SM VGND 0.00502f
C8631 XA.XIR[10].XIC[13].icell.PUM VGND 0.00301f
C8632 XA.XIR[10].XIC[14].icell.PDM VGND 0.18592f
C8633 XA.XIR[10].XIC[12].icell.Ien VGND 0.37698f
C8634 XA.XIR[10].XIC[11].icell.SM VGND 0.00502f
C8635 XA.XIR[10].XIC[12].icell.PUM VGND 0.00301f
C8636 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85333f
C8637 XA.XIR[10].XIC[13].icell.PDM VGND 0.18592f
C8638 XA.XIR[10].XIC[11].icell.Ien VGND 0.37698f
C8639 XA.XIR[10].XIC[10].icell.SM VGND 0.00502f
C8640 XA.XIR[10].XIC[11].icell.PUM VGND 0.00301f
C8641 XA.XIR[10].XIC[12].icell.PDM VGND 0.18592f
C8642 XA.XIR[10].XIC[10].icell.Ien VGND 0.37698f
C8643 XA.XIR[10].XIC[9].icell.SM VGND 0.00502f
C8644 XA.XIR[10].XIC[10].icell.PUM VGND 0.00301f
C8645 XA.XIR[10].XIC[11].icell.PDM VGND 0.18592f
C8646 XA.XIR[10].XIC[9].icell.Ien VGND 0.37698f
C8647 XA.XIR[10].XIC[8].icell.SM VGND 0.00502f
C8648 XA.XIR[10].XIC[9].icell.PUM VGND 0.00301f
C8649 XA.XIR[10].XIC[10].icell.PDM VGND 0.18592f
C8650 XA.XIR[10].XIC[8].icell.Ien VGND 0.37698f
C8651 XA.XIR[10].XIC[7].icell.SM VGND 0.00502f
C8652 XA.XIR[10].XIC[8].icell.PUM VGND 0.00301f
C8653 XA.XIR[10].XIC[9].icell.PDM VGND 0.18592f
C8654 XA.XIR[10].XIC[7].icell.Ien VGND 0.37698f
C8655 XA.XIR[10].XIC[6].icell.SM VGND 0.00502f
C8656 XA.XIR[10].XIC[7].icell.PUM VGND 0.00301f
C8657 XA.XIR[10].XIC[8].icell.PDM VGND 0.18592f
C8658 XA.XIR[10].XIC[6].icell.Ien VGND 0.37698f
C8659 XA.XIR[10].XIC[5].icell.SM VGND 0.00502f
C8660 XA.XIR[10].XIC[6].icell.PUM VGND 0.00301f
C8661 XA.XIR[10].XIC[7].icell.PDM VGND 0.18592f
C8662 XA.XIR[10].XIC[5].icell.Ien VGND 0.37698f
C8663 XA.XIR[10].XIC[4].icell.SM VGND 0.00502f
C8664 XA.XIR[10].XIC[5].icell.PUM VGND 0.00301f
C8665 XA.XIR[10].XIC[6].icell.PDM VGND 0.18592f
C8666 XA.XIR[10].XIC[4].icell.Ien VGND 0.37698f
C8667 XA.XIR[10].XIC[3].icell.SM VGND 0.00502f
C8668 XA.XIR[10].XIC[4].icell.PUM VGND 0.00301f
C8669 XA.XIR[10].XIC[5].icell.PDM VGND 0.18592f
C8670 XA.XIR[10].XIC[3].icell.Ien VGND 0.37698f
C8671 XA.XIR[10].XIC[2].icell.SM VGND 0.00502f
C8672 XA.XIR[10].XIC[3].icell.PUM VGND 0.00301f
C8673 XA.XIR[10].XIC[4].icell.PDM VGND 0.18592f
C8674 XA.XIR[10].XIC[2].icell.Ien VGND 0.37698f
C8675 XA.XIR[10].XIC[1].icell.SM VGND 0.00502f
C8676 XThR.Tn[10] VGND 13.77667f
C8677 XA.XIR[10].XIC[2].icell.PUM VGND 0.00301f
C8678 XA.XIR[10].XIC[3].icell.PDM VGND 0.18592f
C8679 XA.XIR[10].XIC[1].icell.Ien VGND 0.37698f
C8680 XA.XIR[10].XIC[0].icell.SM VGND 0.00502f
C8681 XA.XIR[10].XIC[1].icell.PUM VGND 0.00301f
C8682 XA.XIR[10].XIC[2].icell.PDM VGND 0.18592f
C8683 XA.XIR[10].XIC[0].icell.Ien VGND 0.3772f
C8684 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01043f
C8685 XA.XIR[10].XIC[0].icell.PUM VGND 0.00549f
C8686 XA.XIR[10].XIC[1].icell.PDM VGND 0.18592f
C8687 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.58069f
C8688 XA.XIR[10].XIC_dummy_left.icell.PUM VGND 0.00226f
C8689 XA.XIR[10].XIC[0].icell.PDM VGND 0.18601f
C8690 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22378f
C8691 a_n997_3755# VGND 0.54793f
C8692 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.80407f
C8693 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C8694 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.6141f
C8695 XA.XIR[9].XIC_15.icell.SM VGND 0.00474f
C8696 XA.XIR[9].XIC_dummy_right.icell.PUM VGND 0.00226f
C8697 XA.XIR[9].XIC_15.icell.Ien VGND 0.37606f
C8698 XA.XIR[9].XIC[14].icell.SM VGND 0.00502f
C8699 XA.XIR[9].XIC_15.icell.PUM VGND 0.00284f
C8700 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23008f
C8701 XA.XIR[9].XIC[14].icell.Ien VGND 0.37698f
C8702 XA.XIR[9].XIC[13].icell.SM VGND 0.00502f
C8703 XA.XIR[9].XIC[14].icell.PUM VGND 0.00301f
C8704 XA.XIR[9].XIC_15.icell.PDM VGND 0.18645f
C8705 XA.XIR[9].XIC[13].icell.Ien VGND 0.37698f
C8706 XA.XIR[9].XIC[12].icell.SM VGND 0.00502f
C8707 XA.XIR[9].XIC[13].icell.PUM VGND 0.00301f
C8708 XA.XIR[9].XIC[14].icell.PDM VGND 0.18592f
C8709 XA.XIR[9].XIC[12].icell.Ien VGND 0.37698f
C8710 XA.XIR[9].XIC[11].icell.SM VGND 0.00502f
C8711 XA.XIR[9].XIC[12].icell.PUM VGND 0.00301f
C8712 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85333f
C8713 XA.XIR[9].XIC[13].icell.PDM VGND 0.18592f
C8714 XA.XIR[9].XIC[11].icell.Ien VGND 0.37698f
C8715 XA.XIR[9].XIC[10].icell.SM VGND 0.00502f
C8716 XA.XIR[9].XIC[11].icell.PUM VGND 0.00301f
C8717 XA.XIR[9].XIC[12].icell.PDM VGND 0.18592f
C8718 XA.XIR[9].XIC[10].icell.Ien VGND 0.37698f
C8719 XA.XIR[9].XIC[9].icell.SM VGND 0.00502f
C8720 XA.XIR[9].XIC[10].icell.PUM VGND 0.00301f
C8721 XA.XIR[9].XIC[11].icell.PDM VGND 0.18592f
C8722 XA.XIR[9].XIC[9].icell.Ien VGND 0.37698f
C8723 XA.XIR[9].XIC[8].icell.SM VGND 0.00502f
C8724 XA.XIR[9].XIC[9].icell.PUM VGND 0.00301f
C8725 XA.XIR[9].XIC[10].icell.PDM VGND 0.18592f
C8726 XA.XIR[9].XIC[8].icell.Ien VGND 0.37698f
C8727 XA.XIR[9].XIC[7].icell.SM VGND 0.00502f
C8728 XA.XIR[9].XIC[8].icell.PUM VGND 0.00301f
C8729 XA.XIR[9].XIC[9].icell.PDM VGND 0.18592f
C8730 XA.XIR[9].XIC[7].icell.Ien VGND 0.37698f
C8731 XA.XIR[9].XIC[6].icell.SM VGND 0.00502f
C8732 XA.XIR[9].XIC[7].icell.PUM VGND 0.00301f
C8733 XA.XIR[9].XIC[8].icell.PDM VGND 0.18592f
C8734 XA.XIR[9].XIC[6].icell.Ien VGND 0.37698f
C8735 XA.XIR[9].XIC[5].icell.SM VGND 0.00502f
C8736 XA.XIR[9].XIC[6].icell.PUM VGND 0.00301f
C8737 XA.XIR[9].XIC[7].icell.PDM VGND 0.18592f
C8738 XA.XIR[9].XIC[5].icell.Ien VGND 0.37698f
C8739 XA.XIR[9].XIC[4].icell.SM VGND 0.00502f
C8740 XA.XIR[9].XIC[5].icell.PUM VGND 0.00301f
C8741 XA.XIR[9].XIC[6].icell.PDM VGND 0.18592f
C8742 XA.XIR[9].XIC[4].icell.Ien VGND 0.37698f
C8743 XA.XIR[9].XIC[3].icell.SM VGND 0.00502f
C8744 XA.XIR[9].XIC[4].icell.PUM VGND 0.00301f
C8745 XA.XIR[9].XIC[5].icell.PDM VGND 0.18592f
C8746 XA.XIR[9].XIC[3].icell.Ien VGND 0.37698f
C8747 XA.XIR[9].XIC[2].icell.SM VGND 0.00502f
C8748 XA.XIR[9].XIC[3].icell.PUM VGND 0.00301f
C8749 XA.XIR[9].XIC[4].icell.PDM VGND 0.18592f
C8750 XA.XIR[9].XIC[2].icell.Ien VGND 0.37698f
C8751 XA.XIR[9].XIC[1].icell.SM VGND 0.00502f
C8752 XThR.Tn[9] VGND 13.78041f
C8753 XA.XIR[9].XIC[2].icell.PUM VGND 0.00301f
C8754 XA.XIR[9].XIC[3].icell.PDM VGND 0.18592f
C8755 XA.XIR[9].XIC[1].icell.Ien VGND 0.37698f
C8756 XA.XIR[9].XIC[0].icell.SM VGND 0.00502f
C8757 XA.XIR[9].XIC[1].icell.PUM VGND 0.00301f
C8758 XA.XIR[9].XIC[2].icell.PDM VGND 0.18592f
C8759 XA.XIR[9].XIC[0].icell.Ien VGND 0.3772f
C8760 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01043f
C8761 XA.XIR[9].XIC[0].icell.PUM VGND 0.00549f
C8762 XA.XIR[9].XIC[1].icell.PDM VGND 0.18592f
C8763 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.58012f
C8764 a_n997_3979# VGND 0.54721f
C8765 XA.XIR[9].XIC_dummy_left.icell.PUM VGND 0.00226f
C8766 XA.XIR[9].XIC[0].icell.PDM VGND 0.18601f
C8767 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22378f
C8768 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80139f
C8769 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C8770 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.6141f
C8771 XA.XIR[8].XIC_15.icell.SM VGND 0.00474f
C8772 XA.XIR[8].XIC_dummy_right.icell.PUM VGND 0.00226f
C8773 XA.XIR[8].XIC_15.icell.Ien VGND 0.37606f
C8774 XA.XIR[8].XIC[14].icell.SM VGND 0.00502f
C8775 XA.XIR[8].XIC_15.icell.PUM VGND 0.00284f
C8776 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23008f
C8777 XA.XIR[8].XIC[14].icell.Ien VGND 0.37698f
C8778 XA.XIR[8].XIC[13].icell.SM VGND 0.00502f
C8779 XA.XIR[8].XIC[14].icell.PUM VGND 0.00301f
C8780 XA.XIR[8].XIC_15.icell.PDM VGND 0.18645f
C8781 XA.XIR[8].XIC[13].icell.Ien VGND 0.37698f
C8782 XA.XIR[8].XIC[12].icell.SM VGND 0.00502f
C8783 XA.XIR[8].XIC[13].icell.PUM VGND 0.00301f
C8784 XA.XIR[8].XIC[14].icell.PDM VGND 0.18592f
C8785 XA.XIR[8].XIC[12].icell.Ien VGND 0.37698f
C8786 XA.XIR[8].XIC[11].icell.SM VGND 0.00502f
C8787 XA.XIR[8].XIC[12].icell.PUM VGND 0.00301f
C8788 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85333f
C8789 XA.XIR[8].XIC[13].icell.PDM VGND 0.18592f
C8790 XA.XIR[8].XIC[11].icell.Ien VGND 0.37698f
C8791 XA.XIR[8].XIC[10].icell.SM VGND 0.00502f
C8792 XA.XIR[8].XIC[11].icell.PUM VGND 0.00301f
C8793 XA.XIR[8].XIC[12].icell.PDM VGND 0.18592f
C8794 XA.XIR[8].XIC[10].icell.Ien VGND 0.37698f
C8795 XA.XIR[8].XIC[9].icell.SM VGND 0.00502f
C8796 XA.XIR[8].XIC[10].icell.PUM VGND 0.00301f
C8797 XA.XIR[8].XIC[11].icell.PDM VGND 0.18592f
C8798 XA.XIR[8].XIC[9].icell.Ien VGND 0.37698f
C8799 XA.XIR[8].XIC[8].icell.SM VGND 0.00502f
C8800 XA.XIR[8].XIC[9].icell.PUM VGND 0.00301f
C8801 XA.XIR[8].XIC[10].icell.PDM VGND 0.18592f
C8802 XA.XIR[8].XIC[8].icell.Ien VGND 0.37698f
C8803 XA.XIR[8].XIC[7].icell.SM VGND 0.00502f
C8804 XA.XIR[8].XIC[8].icell.PUM VGND 0.00301f
C8805 XA.XIR[8].XIC[9].icell.PDM VGND 0.18592f
C8806 XA.XIR[8].XIC[7].icell.Ien VGND 0.37698f
C8807 XA.XIR[8].XIC[6].icell.SM VGND 0.00502f
C8808 XA.XIR[8].XIC[7].icell.PUM VGND 0.00301f
C8809 XA.XIR[8].XIC[8].icell.PDM VGND 0.18592f
C8810 XA.XIR[8].XIC[6].icell.Ien VGND 0.37698f
C8811 XA.XIR[8].XIC[5].icell.SM VGND 0.00502f
C8812 XA.XIR[8].XIC[6].icell.PUM VGND 0.00301f
C8813 XA.XIR[8].XIC[7].icell.PDM VGND 0.18592f
C8814 XA.XIR[8].XIC[5].icell.Ien VGND 0.37698f
C8815 XA.XIR[8].XIC[4].icell.SM VGND 0.00502f
C8816 XA.XIR[8].XIC[5].icell.PUM VGND 0.00301f
C8817 XA.XIR[8].XIC[6].icell.PDM VGND 0.18592f
C8818 XA.XIR[8].XIC[4].icell.Ien VGND 0.37698f
C8819 XA.XIR[8].XIC[3].icell.SM VGND 0.00502f
C8820 XA.XIR[8].XIC[4].icell.PUM VGND 0.00301f
C8821 XA.XIR[8].XIC[5].icell.PDM VGND 0.18592f
C8822 XA.XIR[8].XIC[3].icell.Ien VGND 0.37698f
C8823 XA.XIR[8].XIC[2].icell.SM VGND 0.00502f
C8824 XA.XIR[8].XIC[3].icell.PUM VGND 0.00301f
C8825 XA.XIR[8].XIC[4].icell.PDM VGND 0.18592f
C8826 XA.XIR[8].XIC[2].icell.Ien VGND 0.37698f
C8827 XA.XIR[8].XIC[1].icell.SM VGND 0.00502f
C8828 XA.XIR[8].XIC[2].icell.PUM VGND 0.00301f
C8829 XA.XIR[8].XIC[3].icell.PDM VGND 0.18592f
C8830 XA.XIR[8].XIC[1].icell.Ien VGND 0.37698f
C8831 XA.XIR[8].XIC[0].icell.SM VGND 0.00502f
C8832 XThR.Tn[8] VGND 13.7628f
C8833 XA.XIR[8].XIC[1].icell.PUM VGND 0.00301f
C8834 XA.XIR[8].XIC[2].icell.PDM VGND 0.18592f
C8835 XA.XIR[8].XIC[0].icell.Ien VGND 0.3772f
C8836 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01043f
C8837 XA.XIR[8].XIC[0].icell.PUM VGND 0.00549f
C8838 XA.XIR[8].XIC[1].icell.PDM VGND 0.18592f
C8839 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57973f
C8840 XA.XIR[8].XIC_dummy_left.icell.PUM VGND 0.00226f
C8841 XA.XIR[8].XIC[0].icell.PDM VGND 0.18601f
C8842 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22378f
C8843 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.8017f
C8844 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C8845 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.6141f
C8846 XA.XIR[7].XIC_15.icell.SM VGND 0.00474f
C8847 XA.XIR[7].XIC_dummy_right.icell.PUM VGND 0.00226f
C8848 XA.XIR[7].XIC_15.icell.Ien VGND 0.37606f
C8849 XA.XIR[7].XIC[14].icell.SM VGND 0.00502f
C8850 XA.XIR[7].XIC_15.icell.PUM VGND 0.00284f
C8851 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23008f
C8852 XA.XIR[7].XIC[14].icell.Ien VGND 0.37698f
C8853 XA.XIR[7].XIC[13].icell.SM VGND 0.00502f
C8854 XA.XIR[7].XIC[14].icell.PUM VGND 0.00301f
C8855 XA.XIR[7].XIC_15.icell.PDM VGND 0.18645f
C8856 XA.XIR[7].XIC[13].icell.Ien VGND 0.37698f
C8857 XA.XIR[7].XIC[12].icell.SM VGND 0.00502f
C8858 XA.XIR[7].XIC[13].icell.PUM VGND 0.00301f
C8859 XA.XIR[7].XIC[14].icell.PDM VGND 0.18592f
C8860 XA.XIR[7].XIC[12].icell.Ien VGND 0.37698f
C8861 XA.XIR[7].XIC[11].icell.SM VGND 0.00502f
C8862 XA.XIR[7].XIC[12].icell.PUM VGND 0.00301f
C8863 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85333f
C8864 XA.XIR[7].XIC[13].icell.PDM VGND 0.18592f
C8865 XA.XIR[7].XIC[11].icell.Ien VGND 0.37698f
C8866 XA.XIR[7].XIC[10].icell.SM VGND 0.00502f
C8867 XA.XIR[7].XIC[11].icell.PUM VGND 0.00301f
C8868 XA.XIR[7].XIC[12].icell.PDM VGND 0.18592f
C8869 XA.XIR[7].XIC[10].icell.Ien VGND 0.37698f
C8870 XA.XIR[7].XIC[9].icell.SM VGND 0.00502f
C8871 XA.XIR[7].XIC[10].icell.PUM VGND 0.00301f
C8872 XA.XIR[7].XIC[11].icell.PDM VGND 0.18592f
C8873 XA.XIR[7].XIC[9].icell.Ien VGND 0.37698f
C8874 XA.XIR[7].XIC[8].icell.SM VGND 0.00502f
C8875 XA.XIR[7].XIC[9].icell.PUM VGND 0.00301f
C8876 XA.XIR[7].XIC[10].icell.PDM VGND 0.18592f
C8877 XA.XIR[7].XIC[8].icell.Ien VGND 0.37698f
C8878 XA.XIR[7].XIC[7].icell.SM VGND 0.00502f
C8879 XA.XIR[7].XIC[8].icell.PUM VGND 0.00301f
C8880 XA.XIR[7].XIC[9].icell.PDM VGND 0.18592f
C8881 XA.XIR[7].XIC[7].icell.Ien VGND 0.37698f
C8882 XA.XIR[7].XIC[6].icell.SM VGND 0.00502f
C8883 XA.XIR[7].XIC[7].icell.PUM VGND 0.00301f
C8884 XA.XIR[7].XIC[8].icell.PDM VGND 0.18592f
C8885 XA.XIR[7].XIC[6].icell.Ien VGND 0.37698f
C8886 XA.XIR[7].XIC[5].icell.SM VGND 0.00502f
C8887 XA.XIR[7].XIC[6].icell.PUM VGND 0.00301f
C8888 XA.XIR[7].XIC[7].icell.PDM VGND 0.18592f
C8889 XA.XIR[7].XIC[5].icell.Ien VGND 0.37698f
C8890 XA.XIR[7].XIC[4].icell.SM VGND 0.00502f
C8891 XA.XIR[7].XIC[5].icell.PUM VGND 0.00301f
C8892 XA.XIR[7].XIC[6].icell.PDM VGND 0.18592f
C8893 XA.XIR[7].XIC[4].icell.Ien VGND 0.37698f
C8894 XA.XIR[7].XIC[3].icell.SM VGND 0.00502f
C8895 XA.XIR[7].XIC[4].icell.PUM VGND 0.00301f
C8896 XA.XIR[7].XIC[5].icell.PDM VGND 0.18592f
C8897 XA.XIR[7].XIC[3].icell.Ien VGND 0.37698f
C8898 XA.XIR[7].XIC[2].icell.SM VGND 0.00502f
C8899 XA.XIR[7].XIC[3].icell.PUM VGND 0.00301f
C8900 XA.XIR[7].XIC[4].icell.PDM VGND 0.18592f
C8901 XA.XIR[7].XIC[2].icell.Ien VGND 0.37698f
C8902 XA.XIR[7].XIC[1].icell.SM VGND 0.00502f
C8903 XA.XIR[7].XIC[2].icell.PUM VGND 0.00301f
C8904 XA.XIR[7].XIC[3].icell.PDM VGND 0.18592f
C8905 XA.XIR[7].XIC[1].icell.Ien VGND 0.37698f
C8906 XA.XIR[7].XIC[0].icell.SM VGND 0.00502f
C8907 XA.XIR[7].XIC[1].icell.PUM VGND 0.00301f
C8908 XA.XIR[7].XIC[2].icell.PDM VGND 0.18592f
C8909 XA.XIR[7].XIC[0].icell.Ien VGND 0.3772f
C8910 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01043f
C8911 XThR.Tn[7] VGND 14.24964f
C8912 XA.XIR[7].XIC[0].icell.PUM VGND 0.00549f
C8913 XA.XIR[7].XIC[1].icell.PDM VGND 0.18592f
C8914 XThR.XTBN.A VGND 1.22815f
C8915 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.58218f
C8916 XA.XIR[7].XIC_dummy_left.icell.PUM VGND 0.00236f
C8917 XA.XIR[7].XIC[0].icell.PDM VGND 0.18601f
C8918 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22378f
C8919 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80266f
C8920 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C8921 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.6141f
C8922 XA.XIR[6].XIC_15.icell.SM VGND 0.00474f
C8923 XA.XIR[6].XIC_dummy_right.icell.PUM VGND 0.00226f
C8924 XA.XIR[6].XIC_15.icell.Ien VGND 0.37606f
C8925 XA.XIR[6].XIC[14].icell.SM VGND 0.00502f
C8926 XA.XIR[6].XIC_15.icell.PUM VGND 0.00284f
C8927 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23008f
C8928 XA.XIR[6].XIC[14].icell.Ien VGND 0.37698f
C8929 XA.XIR[6].XIC[13].icell.SM VGND 0.00502f
C8930 XA.XIR[6].XIC[14].icell.PUM VGND 0.00301f
C8931 XA.XIR[6].XIC_15.icell.PDM VGND 0.18645f
C8932 XA.XIR[6].XIC[13].icell.Ien VGND 0.37698f
C8933 XA.XIR[6].XIC[12].icell.SM VGND 0.00502f
C8934 XA.XIR[6].XIC[13].icell.PUM VGND 0.00301f
C8935 XA.XIR[6].XIC[14].icell.PDM VGND 0.18592f
C8936 XA.XIR[6].XIC[12].icell.Ien VGND 0.37698f
C8937 XA.XIR[6].XIC[11].icell.SM VGND 0.00502f
C8938 XA.XIR[6].XIC[12].icell.PUM VGND 0.00301f
C8939 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85333f
C8940 XA.XIR[6].XIC[13].icell.PDM VGND 0.18592f
C8941 XA.XIR[6].XIC[11].icell.Ien VGND 0.37698f
C8942 XA.XIR[6].XIC[10].icell.SM VGND 0.00502f
C8943 XA.XIR[6].XIC[11].icell.PUM VGND 0.00301f
C8944 XA.XIR[6].XIC[12].icell.PDM VGND 0.18592f
C8945 XA.XIR[6].XIC[10].icell.Ien VGND 0.37698f
C8946 XA.XIR[6].XIC[9].icell.SM VGND 0.00502f
C8947 XA.XIR[6].XIC[10].icell.PUM VGND 0.00301f
C8948 XA.XIR[6].XIC[11].icell.PDM VGND 0.18592f
C8949 XA.XIR[6].XIC[9].icell.Ien VGND 0.37698f
C8950 XA.XIR[6].XIC[8].icell.SM VGND 0.00502f
C8951 XA.XIR[6].XIC[9].icell.PUM VGND 0.00301f
C8952 XA.XIR[6].XIC[10].icell.PDM VGND 0.18592f
C8953 XA.XIR[6].XIC[8].icell.Ien VGND 0.37698f
C8954 XA.XIR[6].XIC[7].icell.SM VGND 0.00502f
C8955 XA.XIR[6].XIC[8].icell.PUM VGND 0.00301f
C8956 XA.XIR[6].XIC[9].icell.PDM VGND 0.18592f
C8957 XA.XIR[6].XIC[7].icell.Ien VGND 0.37698f
C8958 XA.XIR[6].XIC[6].icell.SM VGND 0.00502f
C8959 XA.XIR[6].XIC[7].icell.PUM VGND 0.00301f
C8960 XA.XIR[6].XIC[8].icell.PDM VGND 0.18592f
C8961 XA.XIR[6].XIC[6].icell.Ien VGND 0.37698f
C8962 XA.XIR[6].XIC[5].icell.SM VGND 0.00502f
C8963 XA.XIR[6].XIC[6].icell.PUM VGND 0.00301f
C8964 XA.XIR[6].XIC[7].icell.PDM VGND 0.18592f
C8965 XA.XIR[6].XIC[5].icell.Ien VGND 0.37698f
C8966 XA.XIR[6].XIC[4].icell.SM VGND 0.00502f
C8967 XA.XIR[6].XIC[5].icell.PUM VGND 0.00301f
C8968 XA.XIR[6].XIC[6].icell.PDM VGND 0.18592f
C8969 XA.XIR[6].XIC[4].icell.Ien VGND 0.37698f
C8970 XA.XIR[6].XIC[3].icell.SM VGND 0.00502f
C8971 XA.XIR[6].XIC[4].icell.PUM VGND 0.00301f
C8972 XA.XIR[6].XIC[5].icell.PDM VGND 0.18592f
C8973 XA.XIR[6].XIC[3].icell.Ien VGND 0.37698f
C8974 XA.XIR[6].XIC[2].icell.SM VGND 0.00502f
C8975 XA.XIR[6].XIC[3].icell.PUM VGND 0.00301f
C8976 XA.XIR[6].XIC[4].icell.PDM VGND 0.18592f
C8977 XA.XIR[6].XIC[2].icell.Ien VGND 0.37698f
C8978 XA.XIR[6].XIC[1].icell.SM VGND 0.00502f
C8979 XA.XIR[6].XIC[2].icell.PUM VGND 0.00301f
C8980 XA.XIR[6].XIC[3].icell.PDM VGND 0.18592f
C8981 XA.XIR[6].XIC[1].icell.Ien VGND 0.37698f
C8982 XA.XIR[6].XIC[0].icell.SM VGND 0.00502f
C8983 XA.XIR[6].XIC[1].icell.PUM VGND 0.00301f
C8984 XA.XIR[6].XIC[2].icell.PDM VGND 0.18592f
C8985 XA.XIR[6].XIC[0].icell.Ien VGND 0.3772f
C8986 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01043f
C8987 XA.XIR[6].XIC[0].icell.PUM VGND 0.00549f
C8988 XA.XIR[6].XIC[1].icell.PDM VGND 0.18592f
C8989 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.58069f
C8990 XThR.Tn[6] VGND 13.85326f
C8991 a_n1049_5317# VGND 0.02283f
C8992 XA.XIR[6].XIC_dummy_left.icell.PUM VGND 0.00226f
C8993 XThR.XTB7.Y VGND 1.36132f
C8994 XA.XIR[6].XIC[0].icell.PDM VGND 0.18601f
C8995 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22378f
C8996 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80134f
C8997 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C8998 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.6141f
C8999 XA.XIR[5].XIC_15.icell.SM VGND 0.00474f
C9000 XA.XIR[5].XIC_dummy_right.icell.PUM VGND 0.00226f
C9001 XA.XIR[5].XIC_15.icell.Ien VGND 0.37606f
C9002 XA.XIR[5].XIC[14].icell.SM VGND 0.00502f
C9003 XA.XIR[5].XIC_15.icell.PUM VGND 0.00284f
C9004 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23008f
C9005 XA.XIR[5].XIC[14].icell.Ien VGND 0.37698f
C9006 XA.XIR[5].XIC[13].icell.SM VGND 0.00502f
C9007 XA.XIR[5].XIC[14].icell.PUM VGND 0.00301f
C9008 XA.XIR[5].XIC_15.icell.PDM VGND 0.18645f
C9009 XA.XIR[5].XIC[13].icell.Ien VGND 0.37698f
C9010 XA.XIR[5].XIC[12].icell.SM VGND 0.00502f
C9011 XA.XIR[5].XIC[13].icell.PUM VGND 0.00301f
C9012 XA.XIR[5].XIC[14].icell.PDM VGND 0.18592f
C9013 XA.XIR[5].XIC[12].icell.Ien VGND 0.37698f
C9014 XA.XIR[5].XIC[11].icell.SM VGND 0.00502f
C9015 XA.XIR[5].XIC[12].icell.PUM VGND 0.00301f
C9016 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85333f
C9017 XA.XIR[5].XIC[13].icell.PDM VGND 0.18592f
C9018 XA.XIR[5].XIC[11].icell.Ien VGND 0.37698f
C9019 XA.XIR[5].XIC[10].icell.SM VGND 0.00502f
C9020 XA.XIR[5].XIC[11].icell.PUM VGND 0.00301f
C9021 XA.XIR[5].XIC[12].icell.PDM VGND 0.18592f
C9022 XA.XIR[5].XIC[10].icell.Ien VGND 0.37698f
C9023 XA.XIR[5].XIC[9].icell.SM VGND 0.00502f
C9024 XA.XIR[5].XIC[10].icell.PUM VGND 0.00301f
C9025 XA.XIR[5].XIC[11].icell.PDM VGND 0.18592f
C9026 XA.XIR[5].XIC[9].icell.Ien VGND 0.37698f
C9027 XA.XIR[5].XIC[8].icell.SM VGND 0.00502f
C9028 XA.XIR[5].XIC[9].icell.PUM VGND 0.00301f
C9029 XA.XIR[5].XIC[10].icell.PDM VGND 0.18592f
C9030 XA.XIR[5].XIC[8].icell.Ien VGND 0.37698f
C9031 XA.XIR[5].XIC[7].icell.SM VGND 0.00502f
C9032 XA.XIR[5].XIC[8].icell.PUM VGND 0.00301f
C9033 XA.XIR[5].XIC[9].icell.PDM VGND 0.18592f
C9034 XA.XIR[5].XIC[7].icell.Ien VGND 0.37698f
C9035 XA.XIR[5].XIC[6].icell.SM VGND 0.00502f
C9036 XA.XIR[5].XIC[7].icell.PUM VGND 0.00301f
C9037 XA.XIR[5].XIC[8].icell.PDM VGND 0.18592f
C9038 XA.XIR[5].XIC[6].icell.Ien VGND 0.37698f
C9039 XA.XIR[5].XIC[5].icell.SM VGND 0.00502f
C9040 XA.XIR[5].XIC[6].icell.PUM VGND 0.00301f
C9041 XA.XIR[5].XIC[7].icell.PDM VGND 0.18592f
C9042 XA.XIR[5].XIC[5].icell.Ien VGND 0.37698f
C9043 XA.XIR[5].XIC[4].icell.SM VGND 0.00502f
C9044 XA.XIR[5].XIC[5].icell.PUM VGND 0.00301f
C9045 XA.XIR[5].XIC[6].icell.PDM VGND 0.18592f
C9046 XA.XIR[5].XIC[4].icell.Ien VGND 0.37698f
C9047 XA.XIR[5].XIC[3].icell.SM VGND 0.00502f
C9048 XA.XIR[5].XIC[4].icell.PUM VGND 0.00301f
C9049 XA.XIR[5].XIC[5].icell.PDM VGND 0.18592f
C9050 XA.XIR[5].XIC[3].icell.Ien VGND 0.37698f
C9051 XA.XIR[5].XIC[2].icell.SM VGND 0.00502f
C9052 XA.XIR[5].XIC[3].icell.PUM VGND 0.00301f
C9053 XA.XIR[5].XIC[4].icell.PDM VGND 0.18592f
C9054 XA.XIR[5].XIC[2].icell.Ien VGND 0.37698f
C9055 XA.XIR[5].XIC[1].icell.SM VGND 0.00502f
C9056 XA.XIR[5].XIC[2].icell.PUM VGND 0.00301f
C9057 XA.XIR[5].XIC[3].icell.PDM VGND 0.18592f
C9058 XA.XIR[5].XIC[1].icell.Ien VGND 0.37698f
C9059 XA.XIR[5].XIC[0].icell.SM VGND 0.00502f
C9060 a_n1049_5611# VGND 0.02855f
C9061 XA.XIR[5].XIC[1].icell.PUM VGND 0.00301f
C9062 XA.XIR[5].XIC[2].icell.PDM VGND 0.18592f
C9063 XA.XIR[5].XIC[0].icell.Ien VGND 0.3772f
C9064 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01043f
C9065 XA.XIR[5].XIC[0].icell.PUM VGND 0.00549f
C9066 XA.XIR[5].XIC[1].icell.PDM VGND 0.18592f
C9067 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57955f
C9068 XA.XIR[5].XIC_dummy_left.icell.PUM VGND 0.00226f
C9069 XA.XIR[5].XIC[0].icell.PDM VGND 0.18601f
C9070 XThR.Tn[5] VGND 13.83264f
C9071 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22378f
C9072 XThR.XTB6.Y VGND 1.38212f
C9073 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.80311f
C9074 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C9075 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.6141f
C9076 XA.XIR[4].XIC_15.icell.SM VGND 0.00474f
C9077 XA.XIR[4].XIC_dummy_right.icell.PUM VGND 0.00226f
C9078 XA.XIR[4].XIC_15.icell.Ien VGND 0.37606f
C9079 XA.XIR[4].XIC[14].icell.SM VGND 0.00502f
C9080 XA.XIR[4].XIC_15.icell.PUM VGND 0.00284f
C9081 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23008f
C9082 XA.XIR[4].XIC[14].icell.Ien VGND 0.37698f
C9083 XA.XIR[4].XIC[13].icell.SM VGND 0.00502f
C9084 XA.XIR[4].XIC[14].icell.PUM VGND 0.00301f
C9085 XA.XIR[4].XIC_15.icell.PDM VGND 0.18645f
C9086 XA.XIR[4].XIC[13].icell.Ien VGND 0.37698f
C9087 XA.XIR[4].XIC[12].icell.SM VGND 0.00502f
C9088 XA.XIR[4].XIC[13].icell.PUM VGND 0.00301f
C9089 XA.XIR[4].XIC[14].icell.PDM VGND 0.18592f
C9090 XA.XIR[4].XIC[12].icell.Ien VGND 0.37698f
C9091 XA.XIR[4].XIC[11].icell.SM VGND 0.00502f
C9092 XA.XIR[4].XIC[12].icell.PUM VGND 0.00301f
C9093 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85333f
C9094 XA.XIR[4].XIC[13].icell.PDM VGND 0.18592f
C9095 XA.XIR[4].XIC[11].icell.Ien VGND 0.37698f
C9096 XA.XIR[4].XIC[10].icell.SM VGND 0.00502f
C9097 XA.XIR[4].XIC[11].icell.PUM VGND 0.00301f
C9098 XA.XIR[4].XIC[12].icell.PDM VGND 0.18592f
C9099 XA.XIR[4].XIC[10].icell.Ien VGND 0.37698f
C9100 XA.XIR[4].XIC[9].icell.SM VGND 0.00502f
C9101 XA.XIR[4].XIC[10].icell.PUM VGND 0.00301f
C9102 XA.XIR[4].XIC[11].icell.PDM VGND 0.18592f
C9103 XA.XIR[4].XIC[9].icell.Ien VGND 0.37698f
C9104 XA.XIR[4].XIC[8].icell.SM VGND 0.00502f
C9105 XA.XIR[4].XIC[9].icell.PUM VGND 0.00301f
C9106 XA.XIR[4].XIC[10].icell.PDM VGND 0.18592f
C9107 XA.XIR[4].XIC[8].icell.Ien VGND 0.37698f
C9108 XA.XIR[4].XIC[7].icell.SM VGND 0.00502f
C9109 XA.XIR[4].XIC[8].icell.PUM VGND 0.00301f
C9110 XA.XIR[4].XIC[9].icell.PDM VGND 0.18592f
C9111 XA.XIR[4].XIC[7].icell.Ien VGND 0.37698f
C9112 XA.XIR[4].XIC[6].icell.SM VGND 0.00502f
C9113 XA.XIR[4].XIC[7].icell.PUM VGND 0.00301f
C9114 XA.XIR[4].XIC[8].icell.PDM VGND 0.18592f
C9115 XA.XIR[4].XIC[6].icell.Ien VGND 0.37698f
C9116 XA.XIR[4].XIC[5].icell.SM VGND 0.00502f
C9117 XA.XIR[4].XIC[6].icell.PUM VGND 0.00301f
C9118 XA.XIR[4].XIC[7].icell.PDM VGND 0.18592f
C9119 XA.XIR[4].XIC[5].icell.Ien VGND 0.37698f
C9120 XA.XIR[4].XIC[4].icell.SM VGND 0.00502f
C9121 XA.XIR[4].XIC[5].icell.PUM VGND 0.00301f
C9122 XA.XIR[4].XIC[6].icell.PDM VGND 0.18592f
C9123 XA.XIR[4].XIC[4].icell.Ien VGND 0.37698f
C9124 XA.XIR[4].XIC[3].icell.SM VGND 0.00502f
C9125 XA.XIR[4].XIC[4].icell.PUM VGND 0.00301f
C9126 XA.XIR[4].XIC[5].icell.PDM VGND 0.18592f
C9127 XA.XIR[4].XIC[3].icell.Ien VGND 0.37698f
C9128 XA.XIR[4].XIC[2].icell.SM VGND 0.00502f
C9129 XA.XIR[4].XIC[3].icell.PUM VGND 0.00301f
C9130 XA.XIR[4].XIC[4].icell.PDM VGND 0.18592f
C9131 XA.XIR[4].XIC[2].icell.Ien VGND 0.37698f
C9132 XA.XIR[4].XIC[1].icell.SM VGND 0.00502f
C9133 XA.XIR[4].XIC[2].icell.PUM VGND 0.00301f
C9134 XA.XIR[4].XIC[3].icell.PDM VGND 0.18592f
C9135 XA.XIR[4].XIC[1].icell.Ien VGND 0.37698f
C9136 XA.XIR[4].XIC[0].icell.SM VGND 0.00502f
C9137 XA.XIR[4].XIC[1].icell.PUM VGND 0.00301f
C9138 XA.XIR[4].XIC[2].icell.PDM VGND 0.18592f
C9139 XA.XIR[4].XIC[0].icell.Ien VGND 0.3772f
C9140 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01043f
C9141 XA.XIR[4].XIC[0].icell.PUM VGND 0.00549f
C9142 XA.XIR[4].XIC[1].icell.PDM VGND 0.18592f
C9143 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.58f
C9144 XA.XIR[4].XIC_dummy_left.icell.PUM VGND 0.00226f
C9145 XA.XIR[4].XIC[0].icell.PDM VGND 0.18601f
C9146 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22378f
C9147 XThR.Tn[4] VGND 13.90393f
C9148 a_n1049_6405# VGND 0.02893f
C9149 a_n1319_6405# VGND 0.00166f
C9150 XThR.XTB5.Y VGND 1.32753f
C9151 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80148f
C9152 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C9153 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.6141f
C9154 XA.XIR[3].XIC_15.icell.SM VGND 0.00474f
C9155 XA.XIR[3].XIC_dummy_right.icell.PUM VGND 0.00226f
C9156 XA.XIR[3].XIC_15.icell.Ien VGND 0.37606f
C9157 XA.XIR[3].XIC[14].icell.SM VGND 0.00502f
C9158 XA.XIR[3].XIC_15.icell.PUM VGND 0.00284f
C9159 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23008f
C9160 XA.XIR[3].XIC[14].icell.Ien VGND 0.37698f
C9161 XA.XIR[3].XIC[13].icell.SM VGND 0.00502f
C9162 XA.XIR[3].XIC[14].icell.PUM VGND 0.00301f
C9163 XA.XIR[3].XIC_15.icell.PDM VGND 0.18645f
C9164 XA.XIR[3].XIC[13].icell.Ien VGND 0.37698f
C9165 XA.XIR[3].XIC[12].icell.SM VGND 0.00502f
C9166 XA.XIR[3].XIC[13].icell.PUM VGND 0.00301f
C9167 XA.XIR[3].XIC[14].icell.PDM VGND 0.18592f
C9168 XA.XIR[3].XIC[12].icell.Ien VGND 0.37698f
C9169 XA.XIR[3].XIC[11].icell.SM VGND 0.00502f
C9170 XA.XIR[3].XIC[12].icell.PUM VGND 0.00301f
C9171 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85333f
C9172 XA.XIR[3].XIC[13].icell.PDM VGND 0.18592f
C9173 XA.XIR[3].XIC[11].icell.Ien VGND 0.37698f
C9174 XA.XIR[3].XIC[10].icell.SM VGND 0.00502f
C9175 XA.XIR[3].XIC[11].icell.PUM VGND 0.00301f
C9176 XA.XIR[3].XIC[12].icell.PDM VGND 0.18592f
C9177 XA.XIR[3].XIC[10].icell.Ien VGND 0.37698f
C9178 XA.XIR[3].XIC[9].icell.SM VGND 0.00502f
C9179 XA.XIR[3].XIC[10].icell.PUM VGND 0.00301f
C9180 XA.XIR[3].XIC[11].icell.PDM VGND 0.18592f
C9181 XA.XIR[3].XIC[9].icell.Ien VGND 0.37698f
C9182 XA.XIR[3].XIC[8].icell.SM VGND 0.00502f
C9183 XA.XIR[3].XIC[9].icell.PUM VGND 0.00301f
C9184 XA.XIR[3].XIC[10].icell.PDM VGND 0.18592f
C9185 XA.XIR[3].XIC[8].icell.Ien VGND 0.37698f
C9186 XA.XIR[3].XIC[7].icell.SM VGND 0.00502f
C9187 XA.XIR[3].XIC[8].icell.PUM VGND 0.00301f
C9188 XA.XIR[3].XIC[9].icell.PDM VGND 0.18592f
C9189 XA.XIR[3].XIC[7].icell.Ien VGND 0.37698f
C9190 XA.XIR[3].XIC[6].icell.SM VGND 0.00502f
C9191 XA.XIR[3].XIC[7].icell.PUM VGND 0.00301f
C9192 XA.XIR[3].XIC[8].icell.PDM VGND 0.18592f
C9193 XA.XIR[3].XIC[6].icell.Ien VGND 0.37698f
C9194 XA.XIR[3].XIC[5].icell.SM VGND 0.00502f
C9195 XA.XIR[3].XIC[6].icell.PUM VGND 0.00301f
C9196 XA.XIR[3].XIC[7].icell.PDM VGND 0.18592f
C9197 XA.XIR[3].XIC[5].icell.Ien VGND 0.37698f
C9198 XA.XIR[3].XIC[4].icell.SM VGND 0.00502f
C9199 XA.XIR[3].XIC[5].icell.PUM VGND 0.00301f
C9200 XA.XIR[3].XIC[6].icell.PDM VGND 0.18592f
C9201 XA.XIR[3].XIC[4].icell.Ien VGND 0.37698f
C9202 XA.XIR[3].XIC[3].icell.SM VGND 0.00502f
C9203 XA.XIR[3].XIC[4].icell.PUM VGND 0.00301f
C9204 XA.XIR[3].XIC[5].icell.PDM VGND 0.18592f
C9205 XA.XIR[3].XIC[3].icell.Ien VGND 0.37698f
C9206 XA.XIR[3].XIC[2].icell.SM VGND 0.00502f
C9207 XA.XIR[3].XIC[3].icell.PUM VGND 0.00301f
C9208 XA.XIR[3].XIC[4].icell.PDM VGND 0.18592f
C9209 XA.XIR[3].XIC[2].icell.Ien VGND 0.37698f
C9210 XA.XIR[3].XIC[1].icell.SM VGND 0.00502f
C9211 XA.XIR[3].XIC[2].icell.PUM VGND 0.00301f
C9212 XA.XIR[3].XIC[3].icell.PDM VGND 0.18592f
C9213 XA.XIR[3].XIC[1].icell.Ien VGND 0.37698f
C9214 XA.XIR[3].XIC[0].icell.SM VGND 0.00502f
C9215 XA.XIR[3].XIC[1].icell.PUM VGND 0.00301f
C9216 XA.XIR[3].XIC[2].icell.PDM VGND 0.18592f
C9217 XA.XIR[3].XIC[0].icell.Ien VGND 0.3772f
C9218 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01043f
C9219 XA.XIR[3].XIC[0].icell.PUM VGND 0.00549f
C9220 XA.XIR[3].XIC[1].icell.PDM VGND 0.18592f
C9221 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.58069f
C9222 a_n1049_6699# VGND 0.02979f
C9223 XA.XIR[3].XIC_dummy_left.icell.PUM VGND 0.00226f
C9224 XA.XIR[3].XIC[0].icell.PDM VGND 0.18601f
C9225 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22378f
C9226 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80366f
C9227 XThR.Tn[3] VGND 13.84852f
C9228 XThR.XTB4.Y VGND 1.76953f
C9229 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C9230 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.6141f
C9231 XA.XIR[2].XIC_15.icell.SM VGND 0.00474f
C9232 XA.XIR[2].XIC_dummy_right.icell.PUM VGND 0.00226f
C9233 XA.XIR[2].XIC_15.icell.Ien VGND 0.37606f
C9234 XA.XIR[2].XIC[14].icell.SM VGND 0.00502f
C9235 XA.XIR[2].XIC_15.icell.PUM VGND 0.00284f
C9236 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23008f
C9237 XA.XIR[2].XIC[14].icell.Ien VGND 0.37698f
C9238 XA.XIR[2].XIC[13].icell.SM VGND 0.00502f
C9239 XA.XIR[2].XIC[14].icell.PUM VGND 0.00301f
C9240 XA.XIR[2].XIC_15.icell.PDM VGND 0.18645f
C9241 XA.XIR[2].XIC[13].icell.Ien VGND 0.37698f
C9242 XA.XIR[2].XIC[12].icell.SM VGND 0.00502f
C9243 XA.XIR[2].XIC[13].icell.PUM VGND 0.00301f
C9244 XA.XIR[2].XIC[14].icell.PDM VGND 0.18592f
C9245 XA.XIR[2].XIC[12].icell.Ien VGND 0.37698f
C9246 XA.XIR[2].XIC[11].icell.SM VGND 0.00502f
C9247 XA.XIR[2].XIC[12].icell.PUM VGND 0.00301f
C9248 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85333f
C9249 XA.XIR[2].XIC[13].icell.PDM VGND 0.18592f
C9250 XA.XIR[2].XIC[11].icell.Ien VGND 0.37698f
C9251 XA.XIR[2].XIC[10].icell.SM VGND 0.00502f
C9252 XA.XIR[2].XIC[11].icell.PUM VGND 0.00301f
C9253 XA.XIR[2].XIC[12].icell.PDM VGND 0.18592f
C9254 XA.XIR[2].XIC[10].icell.Ien VGND 0.37698f
C9255 XA.XIR[2].XIC[9].icell.SM VGND 0.00502f
C9256 XA.XIR[2].XIC[10].icell.PUM VGND 0.00301f
C9257 XA.XIR[2].XIC[11].icell.PDM VGND 0.18592f
C9258 XA.XIR[2].XIC[9].icell.Ien VGND 0.37698f
C9259 XA.XIR[2].XIC[8].icell.SM VGND 0.00502f
C9260 XA.XIR[2].XIC[9].icell.PUM VGND 0.00301f
C9261 XA.XIR[2].XIC[10].icell.PDM VGND 0.18592f
C9262 XA.XIR[2].XIC[8].icell.Ien VGND 0.37698f
C9263 XA.XIR[2].XIC[7].icell.SM VGND 0.00502f
C9264 XA.XIR[2].XIC[8].icell.PUM VGND 0.00301f
C9265 XA.XIR[2].XIC[9].icell.PDM VGND 0.18592f
C9266 XA.XIR[2].XIC[7].icell.Ien VGND 0.37698f
C9267 XA.XIR[2].XIC[6].icell.SM VGND 0.00502f
C9268 XA.XIR[2].XIC[7].icell.PUM VGND 0.00301f
C9269 XA.XIR[2].XIC[8].icell.PDM VGND 0.18592f
C9270 XA.XIR[2].XIC[6].icell.Ien VGND 0.37698f
C9271 XA.XIR[2].XIC[5].icell.SM VGND 0.00502f
C9272 XA.XIR[2].XIC[6].icell.PUM VGND 0.00301f
C9273 XA.XIR[2].XIC[7].icell.PDM VGND 0.18592f
C9274 XA.XIR[2].XIC[5].icell.Ien VGND 0.37698f
C9275 XA.XIR[2].XIC[4].icell.SM VGND 0.00502f
C9276 XA.XIR[2].XIC[5].icell.PUM VGND 0.00301f
C9277 XA.XIR[2].XIC[6].icell.PDM VGND 0.18592f
C9278 XA.XIR[2].XIC[4].icell.Ien VGND 0.37698f
C9279 XA.XIR[2].XIC[3].icell.SM VGND 0.00502f
C9280 XA.XIR[2].XIC[4].icell.PUM VGND 0.00301f
C9281 XA.XIR[2].XIC[5].icell.PDM VGND 0.18592f
C9282 XA.XIR[2].XIC[3].icell.Ien VGND 0.37698f
C9283 XA.XIR[2].XIC[2].icell.SM VGND 0.00502f
C9284 XA.XIR[2].XIC[3].icell.PUM VGND 0.00301f
C9285 XA.XIR[2].XIC[4].icell.PDM VGND 0.18592f
C9286 XA.XIR[2].XIC[2].icell.Ien VGND 0.37698f
C9287 XA.XIR[2].XIC[1].icell.SM VGND 0.00502f
C9288 XA.XIR[2].XIC[2].icell.PUM VGND 0.00301f
C9289 XA.XIR[2].XIC[3].icell.PDM VGND 0.18592f
C9290 XA.XIR[2].XIC[1].icell.Ien VGND 0.37698f
C9291 XA.XIR[2].XIC[0].icell.SM VGND 0.00502f
C9292 XA.XIR[2].XIC[1].icell.PUM VGND 0.00301f
C9293 XA.XIR[2].XIC[2].icell.PDM VGND 0.18592f
C9294 XA.XIR[2].XIC[0].icell.Ien VGND 0.3772f
C9295 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01043f
C9296 XA.XIR[2].XIC[0].icell.PUM VGND 0.00549f
C9297 XA.XIR[2].XIC[1].icell.PDM VGND 0.18592f
C9298 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.58205f
C9299 a_n1335_7243# VGND 0.00179f
C9300 XA.XIR[2].XIC_dummy_left.icell.PUM VGND 0.00226f
C9301 XA.XIR[2].XIC[0].icell.PDM VGND 0.18601f
C9302 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22378f
C9303 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80148f
C9304 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C9305 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.6141f
C9306 XA.XIR[1].XIC_15.icell.SM VGND 0.00474f
C9307 XA.XIR[1].XIC_dummy_right.icell.PUM VGND 0.00226f
C9308 XA.XIR[1].XIC_15.icell.Ien VGND 0.37606f
C9309 XA.XIR[1].XIC[14].icell.SM VGND 0.00502f
C9310 XA.XIR[1].XIC_15.icell.PUM VGND 0.00284f
C9311 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23008f
C9312 XA.XIR[1].XIC[14].icell.Ien VGND 0.37698f
C9313 XA.XIR[1].XIC[13].icell.SM VGND 0.00502f
C9314 XA.XIR[1].XIC[14].icell.PUM VGND 0.00301f
C9315 XA.XIR[1].XIC_15.icell.PDM VGND 0.18645f
C9316 XA.XIR[1].XIC[13].icell.Ien VGND 0.37698f
C9317 XA.XIR[1].XIC[12].icell.SM VGND 0.00502f
C9318 XA.XIR[1].XIC[13].icell.PUM VGND 0.00301f
C9319 XA.XIR[1].XIC[14].icell.PDM VGND 0.18592f
C9320 XA.XIR[1].XIC[12].icell.Ien VGND 0.37698f
C9321 XA.XIR[1].XIC[11].icell.SM VGND 0.00502f
C9322 XA.XIR[1].XIC[12].icell.PUM VGND 0.00301f
C9323 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.86947f
C9324 XA.XIR[1].XIC[13].icell.PDM VGND 0.18592f
C9325 XA.XIR[1].XIC[11].icell.Ien VGND 0.37698f
C9326 XA.XIR[1].XIC[10].icell.SM VGND 0.00502f
C9327 XA.XIR[1].XIC[11].icell.PUM VGND 0.00301f
C9328 XA.XIR[1].XIC[12].icell.PDM VGND 0.18592f
C9329 XA.XIR[1].XIC[10].icell.Ien VGND 0.37698f
C9330 XA.XIR[1].XIC[9].icell.SM VGND 0.00502f
C9331 XA.XIR[1].XIC[10].icell.PUM VGND 0.00301f
C9332 XA.XIR[1].XIC[11].icell.PDM VGND 0.18592f
C9333 XA.XIR[1].XIC[9].icell.Ien VGND 0.37698f
C9334 XA.XIR[1].XIC[8].icell.SM VGND 0.00502f
C9335 XA.XIR[1].XIC[9].icell.PUM VGND 0.00301f
C9336 XA.XIR[1].XIC[10].icell.PDM VGND 0.18592f
C9337 XA.XIR[1].XIC[8].icell.Ien VGND 0.37698f
C9338 XA.XIR[1].XIC[7].icell.SM VGND 0.00502f
C9339 XA.XIR[1].XIC[8].icell.PUM VGND 0.00301f
C9340 XA.XIR[1].XIC[9].icell.PDM VGND 0.18592f
C9341 XA.XIR[1].XIC[7].icell.Ien VGND 0.37698f
C9342 XA.XIR[1].XIC[6].icell.SM VGND 0.00502f
C9343 XA.XIR[1].XIC[7].icell.PUM VGND 0.00301f
C9344 XA.XIR[1].XIC[8].icell.PDM VGND 0.18592f
C9345 XA.XIR[1].XIC[6].icell.Ien VGND 0.37698f
C9346 XA.XIR[1].XIC[5].icell.SM VGND 0.00502f
C9347 XA.XIR[1].XIC[6].icell.PUM VGND 0.00301f
C9348 XA.XIR[1].XIC[7].icell.PDM VGND 0.18592f
C9349 XA.XIR[1].XIC[5].icell.Ien VGND 0.37698f
C9350 XA.XIR[1].XIC[4].icell.SM VGND 0.00502f
C9351 XA.XIR[1].XIC[5].icell.PUM VGND 0.00301f
C9352 XA.XIR[1].XIC[6].icell.PDM VGND 0.18592f
C9353 XA.XIR[1].XIC[4].icell.Ien VGND 0.37698f
C9354 XA.XIR[1].XIC[3].icell.SM VGND 0.00502f
C9355 XA.XIR[1].XIC[4].icell.PUM VGND 0.00301f
C9356 XA.XIR[1].XIC[5].icell.PDM VGND 0.18592f
C9357 XA.XIR[1].XIC[3].icell.Ien VGND 0.37698f
C9358 XA.XIR[1].XIC[2].icell.SM VGND 0.00502f
C9359 XA.XIR[1].XIC[3].icell.PUM VGND 0.00301f
C9360 XA.XIR[1].XIC[4].icell.PDM VGND 0.18592f
C9361 XA.XIR[1].XIC[2].icell.Ien VGND 0.37698f
C9362 XA.XIR[1].XIC[1].icell.SM VGND 0.00502f
C9363 XA.XIR[1].XIC[2].icell.PUM VGND 0.00301f
C9364 XA.XIR[1].XIC[3].icell.PDM VGND 0.18592f
C9365 XA.XIR[1].XIC[1].icell.Ien VGND 0.37698f
C9366 XA.XIR[1].XIC[0].icell.SM VGND 0.00502f
C9367 XThR.Tn[2] VGND 13.90118f
C9368 a_n1049_7493# VGND 0.02449f
C9369 XThR.XTB3.Y VGND 2.09162f
C9370 XThR.XTB7.A VGND 1.95536f
C9371 XA.XIR[1].XIC[1].icell.PUM VGND 0.00301f
C9372 XA.XIR[1].XIC[2].icell.PDM VGND 0.18592f
C9373 XA.XIR[1].XIC[0].icell.Ien VGND 0.3772f
C9374 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01043f
C9375 XA.XIR[1].XIC[0].icell.PUM VGND 0.00549f
C9376 XA.XIR[1].XIC[1].icell.PDM VGND 0.18592f
C9377 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.58043f
C9378 XA.XIR[1].XIC_dummy_left.icell.PUM VGND 0.00226f
C9379 XA.XIR[1].XIC[0].icell.PDM VGND 0.18601f
C9380 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22378f
C9381 a_n1049_7787# VGND 0.03396f
C9382 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83642f
C9383 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C9384 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.62341f
C9385 XA.XIR[0].XIC_15.icell.SM VGND 0.00474f
C9386 XA.XIR[0].XIC_dummy_right.icell.PUM VGND 0.00217f
C9387 XA.XIR[0].XIC_15.icell.Ien VGND 0.38171f
C9388 XA.XIR[0].XIC[14].icell.SM VGND 0.00623f
C9389 XA.XIR[0].XIC_15.icell.PUM VGND 0.00493f
C9390 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.2377f
C9391 XA.XIR[0].XIC[14].icell.Ien VGND 0.38923f
C9392 XA.XIR[0].XIC[13].icell.SM VGND 0.00623f
C9393 XA.XIR[0].XIC[14].icell.PUM VGND 0.00432f
C9394 XA.XIR[0].XIC_15.icell.PDM VGND 0.19612f
C9395 XA.XIR[0].XIC[13].icell.Ien VGND 0.38928f
C9396 XA.XIR[0].XIC[12].icell.SM VGND 0.00623f
C9397 XA.XIR[0].XIC[13].icell.PUM VGND 0.00437f
C9398 XA.XIR[0].XIC[14].icell.PDM VGND 0.23377f
C9399 XA.XIR[0].XIC[12].icell.Ien VGND 0.38587f
C9400 XA.XIR[0].XIC[11].icell.SM VGND 0.00623f
C9401 XA.XIR[0].XIC[12].icell.PUM VGND 0.00432f
C9402 XA.XIR[0].XIC[13].icell.PDM VGND 0.23359f
C9403 XA.XIR[0].XIC[11].icell.Ien VGND 0.38655f
C9404 XA.XIR[0].XIC[10].icell.SM VGND 0.00623f
C9405 XA.XIR[0].XIC[11].icell.PUM VGND 0.00432f
C9406 XA.XIR[0].XIC[12].icell.PDM VGND 0.22958f
C9407 XA.XIR[0].XIC[10].icell.Ien VGND 0.38786f
C9408 XA.XIR[0].XIC[9].icell.SM VGND 0.00623f
C9409 XA.XIR[0].XIC[10].icell.PUM VGND 0.00432f
C9410 XA.XIR[0].XIC[11].icell.PDM VGND 0.22995f
C9411 XA.XIR[0].XIC[9].icell.Ien VGND 0.38615f
C9412 XA.XIR[0].XIC[8].icell.SM VGND 0.00623f
C9413 XA.XIR[0].XIC[9].icell.PUM VGND 0.00432f
C9414 XA.XIR[0].XIC[10].icell.PDM VGND 0.22967f
C9415 XA.XIR[0].XIC[8].icell.Ien VGND 0.38663f
C9416 XA.XIR[0].XIC[7].icell.SM VGND 0.00623f
C9417 XA.XIR[0].XIC[8].icell.PUM VGND 0.00432f
C9418 XA.XIR[0].XIC[9].icell.PDM VGND 0.22958f
C9419 XA.XIR[0].XIC[7].icell.Ien VGND 0.38694f
C9420 XA.XIR[0].XIC[6].icell.SM VGND 0.00623f
C9421 XA.XIR[0].XIC[7].icell.PUM VGND 0.00432f
C9422 XA.XIR[0].XIC[8].icell.PDM VGND 0.22958f
C9423 XA.XIR[0].XIC[6].icell.Ien VGND 0.38678f
C9424 XA.XIR[0].XIC[5].icell.SM VGND 0.00623f
C9425 XA.XIR[0].XIC[6].icell.PUM VGND 0.00444f
C9426 XA.XIR[0].XIC[7].icell.PDM VGND 0.2319f
C9427 XA.XIR[0].XIC[5].icell.Ien VGND 0.38578f
C9428 XA.XIR[0].XIC[4].icell.SM VGND 0.00623f
C9429 XA.XIR[0].XIC[5].icell.PUM VGND 0.00432f
C9430 XA.XIR[0].XIC[6].icell.PDM VGND 0.22933f
C9431 XA.XIR[0].XIC[4].icell.Ien VGND 0.38592f
C9432 XA.XIR[0].XIC[3].icell.SM VGND 0.00623f
C9433 XA.XIR[0].XIC[4].icell.PUM VGND 0.00432f
C9434 XA.XIR[0].XIC[5].icell.PDM VGND 0.23123f
C9435 XA.XIR[0].XIC[3].icell.Ien VGND 0.38713f
C9436 XA.XIR[0].XIC[2].icell.SM VGND 0.00623f
C9437 XA.XIR[0].XIC[3].icell.PUM VGND 0.00432f
C9438 XA.XIR[0].XIC[4].icell.PDM VGND 0.22964f
C9439 XA.XIR[0].XIC[2].icell.Ien VGND 0.38923f
C9440 XA.XIR[0].XIC[1].icell.SM VGND 0.00623f
C9441 XA.XIR[0].XIC[2].icell.PUM VGND 0.00432f
C9442 XA.XIR[0].XIC[3].icell.PDM VGND 0.23247f
C9443 XA.XIR[0].XIC[1].icell.Ien VGND 0.38923f
C9444 XA.XIR[0].XIC[0].icell.SM VGND 0.00623f
C9445 XA.XIR[0].XIC[1].icell.PUM VGND 0.00435f
C9446 XA.XIR[0].XIC[2].icell.PDM VGND 0.23353f
C9447 XA.XIR[0].XIC[0].icell.Ien VGND 0.38923f
C9448 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01043f
C9449 XA.XIR[0].XIC[0].icell.PUM VGND 0.00691f
C9450 XA.XIR[0].XIC[1].icell.PDM VGND 0.23353f
C9451 XThR.Tn[1] VGND 13.93526f
C9452 a_n1335_8107# VGND 0.00163f
C9453 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.59317f
C9454 XThR.XTB2.Y VGND 1.47668f
C9455 XThR.XTB6.A VGND 0.95642f
C9456 XA.XIR[0].XIC_dummy_left.icell.PUM VGND 0.00382f
C9457 XA.XIR[0].XIC[0].icell.PDM VGND 0.23275f
C9458 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.23356f
C9459 a_n1335_8331# VGND 0.00203f
C9460 XThR.Tn[0] VGND 14.21229f
C9461 a_n1049_8581# VGND 0.04324f
C9462 XThR.XTBN.Y VGND 7.54169f
C9463 XThR.XTB1.Y VGND 1.81265f
C9464 XThR.XTB7.B VGND 2.61156f
C9465 XThR.XTB5.A VGND 1.76044f
C9466 XThC.Tn[14] VGND 10.05793f
C9467 XThC.Tn[13] VGND 9.88365f
C9468 XThC.Tn[12] VGND 9.70746f
C9469 XThC.Tn[11] VGND 9.53947f
C9470 XThC.Tn[10] VGND 9.38703f
C9471 XThC.Tn[9] VGND 9.36615f
C9472 XThC.Tn[8] VGND 9.3421f
C9473 a_10915_9569# VGND 0.55837f
C9474 a_10051_9569# VGND 0.55761f
C9475 a_9827_9569# VGND 0.54463f
C9476 a_8963_9569# VGND 0.5545f
C9477 a_8739_9569# VGND 0.55288f
C9478 a_7875_9569# VGND 0.55432f
C9479 a_7651_9569# VGND 0.55717f
C9480 XThC.Tn[7] VGND 10.6251f
C9481 XThC.Tn[6] VGND 10.45213f
C9482 XThC.Tn[5] VGND 10.72388f
C9483 XThC.Tn[4] VGND 10.71214f
C9484 XThC.Tn[3] VGND 9.99606f
C9485 XThC.Tn[2] VGND 10.57741f
C9486 XThC.Tn[1] VGND 10.45212f
C9487 XThC.Tn[0] VGND 10.83531f
C9488 a_6243_9615# VGND 0.0299f
C9489 a_5949_9615# VGND 0.03432f
C9490 a_5155_9615# VGND 0.03619f
C9491 a_4861_9615# VGND 0.03649f
C9492 a_4067_9615# VGND 0.03071f
C9493 a_3773_9615# VGND 0.03867f
C9494 a_2979_9615# VGND 0.04107f
C9495 a_8739_10571# VGND 0.00194f
C9496 XThC.XTBN.Y VGND 7.9042f
C9497 XThC.XTB7.Y VGND 1.36247f
C9498 XThC.XTB6.Y VGND 1.3829f
C9499 a_5155_10571# VGND 0.00165f
C9500 XThC.XTB7.B VGND 2.76743f
C9501 XThC.XTB5.Y VGND 1.32591f
C9502 XThC.XTBN.A VGND 1.23171f
C9503 a_4387_10575# VGND 0.00179f
C9504 a_3523_10575# VGND 0.00163f
C9505 a_3299_10575# VGND 0.00202f
C9506 XThC.XTB4.Y VGND 1.69874f
C9507 XThC.XTB3.Y VGND 1.96765f
C9508 XThC.XTB7.A VGND 1.96059f
C9509 XThC.XTB6.A VGND 0.95757f
C9510 XThC.XTB2.Y VGND 1.47588f
C9511 XThC.XTB1.Y VGND 1.77676f
C9512 XThC.XTB5.A VGND 1.75974f
C9513 XThC.Tn[3].t5 VGND 0.01817f
C9514 XThC.Tn[3].t4 VGND 0.01817f
C9515 XThC.Tn[3].n0 VGND 0.03667f
C9516 XThC.Tn[3].t7 VGND 0.01817f
C9517 XThC.Tn[3].t6 VGND 0.01817f
C9518 XThC.Tn[3].n1 VGND 0.0429f
C9519 XThC.Tn[3].n2 VGND 0.12869f
C9520 XThC.Tn[3].t9 VGND 0.01181f
C9521 XThC.Tn[3].t8 VGND 0.01181f
C9522 XThC.Tn[3].n3 VGND 0.02689f
C9523 XThC.Tn[3].t11 VGND 0.01181f
C9524 XThC.Tn[3].t10 VGND 0.01181f
C9525 XThC.Tn[3].n4 VGND 0.02689f
C9526 XThC.Tn[3].t1 VGND 0.01181f
C9527 XThC.Tn[3].t0 VGND 0.01181f
C9528 XThC.Tn[3].n5 VGND 0.02689f
C9529 XThC.Tn[3].t3 VGND 0.01181f
C9530 XThC.Tn[3].t2 VGND 0.01181f
C9531 XThC.Tn[3].n6 VGND 0.0448f
C9532 XThC.Tn[3].n7 VGND 0.12805f
C9533 XThC.Tn[3].n8 VGND 0.07916f
C9534 XThC.Tn[3].n9 VGND 0.08933f
C9535 XThC.Tn[3].t13 VGND 0.01476f
C9536 XThC.Tn[3].t26 VGND 0.01555f
C9537 XThC.Tn[3].n10 VGND 0.03861f
C9538 XThC.Tn[3].n11 VGND 0.02405f
C9539 XThC.Tn[3].n12 VGND 0.07793f
C9540 XThC.Tn[3].t23 VGND 0.01476f
C9541 XThC.Tn[3].t36 VGND 0.01555f
C9542 XThC.Tn[3].n13 VGND 0.03861f
C9543 XThC.Tn[3].n14 VGND 0.02405f
C9544 XThC.Tn[3].n15 VGND 0.07814f
C9545 XThC.Tn[3].n16 VGND 0.13047f
C9546 XThC.Tn[3].t35 VGND 0.01476f
C9547 XThC.Tn[3].t17 VGND 0.01555f
C9548 XThC.Tn[3].n17 VGND 0.03861f
C9549 XThC.Tn[3].n18 VGND 0.02405f
C9550 XThC.Tn[3].n19 VGND 0.07814f
C9551 XThC.Tn[3].n20 VGND 0.13047f
C9552 XThC.Tn[3].t37 VGND 0.01476f
C9553 XThC.Tn[3].t18 VGND 0.01555f
C9554 XThC.Tn[3].n21 VGND 0.03861f
C9555 XThC.Tn[3].n22 VGND 0.02405f
C9556 XThC.Tn[3].n23 VGND 0.07814f
C9557 XThC.Tn[3].n24 VGND 0.13047f
C9558 XThC.Tn[3].t15 VGND 0.01476f
C9559 XThC.Tn[3].t29 VGND 0.01555f
C9560 XThC.Tn[3].n25 VGND 0.03861f
C9561 XThC.Tn[3].n26 VGND 0.02405f
C9562 XThC.Tn[3].n27 VGND 0.07814f
C9563 XThC.Tn[3].n28 VGND 0.13047f
C9564 XThC.Tn[3].t25 VGND 0.01476f
C9565 XThC.Tn[3].t40 VGND 0.01555f
C9566 XThC.Tn[3].n29 VGND 0.03861f
C9567 XThC.Tn[3].n30 VGND 0.02405f
C9568 XThC.Tn[3].n31 VGND 0.07814f
C9569 XThC.Tn[3].n32 VGND 0.13047f
C9570 XThC.Tn[3].t38 VGND 0.01476f
C9571 XThC.Tn[3].t19 VGND 0.01555f
C9572 XThC.Tn[3].n33 VGND 0.03861f
C9573 XThC.Tn[3].n34 VGND 0.02405f
C9574 XThC.Tn[3].n35 VGND 0.07814f
C9575 XThC.Tn[3].n36 VGND 0.13047f
C9576 XThC.Tn[3].t16 VGND 0.01476f
C9577 XThC.Tn[3].t30 VGND 0.01555f
C9578 XThC.Tn[3].n37 VGND 0.03861f
C9579 XThC.Tn[3].n38 VGND 0.02405f
C9580 XThC.Tn[3].n39 VGND 0.07814f
C9581 XThC.Tn[3].n40 VGND 0.13047f
C9582 XThC.Tn[3].t20 VGND 0.01476f
C9583 XThC.Tn[3].t32 VGND 0.01555f
C9584 XThC.Tn[3].n41 VGND 0.03861f
C9585 XThC.Tn[3].n42 VGND 0.02405f
C9586 XThC.Tn[3].n43 VGND 0.07814f
C9587 XThC.Tn[3].n44 VGND 0.13047f
C9588 XThC.Tn[3].t27 VGND 0.01476f
C9589 XThC.Tn[3].t41 VGND 0.01555f
C9590 XThC.Tn[3].n45 VGND 0.03861f
C9591 XThC.Tn[3].n46 VGND 0.02405f
C9592 XThC.Tn[3].n47 VGND 0.07814f
C9593 XThC.Tn[3].n48 VGND 0.13047f
C9594 XThC.Tn[3].t39 VGND 0.01476f
C9595 XThC.Tn[3].t21 VGND 0.01555f
C9596 XThC.Tn[3].n49 VGND 0.03861f
C9597 XThC.Tn[3].n50 VGND 0.02405f
C9598 XThC.Tn[3].n51 VGND 0.07814f
C9599 XThC.Tn[3].n52 VGND 0.13047f
C9600 XThC.Tn[3].t42 VGND 0.01476f
C9601 XThC.Tn[3].t24 VGND 0.01555f
C9602 XThC.Tn[3].n53 VGND 0.03861f
C9603 XThC.Tn[3].n54 VGND 0.02405f
C9604 XThC.Tn[3].n55 VGND 0.07814f
C9605 XThC.Tn[3].n56 VGND 0.13047f
C9606 XThC.Tn[3].t28 VGND 0.01476f
C9607 XThC.Tn[3].t43 VGND 0.01555f
C9608 XThC.Tn[3].n57 VGND 0.03861f
C9609 XThC.Tn[3].n58 VGND 0.02405f
C9610 XThC.Tn[3].n59 VGND 0.07814f
C9611 XThC.Tn[3].n60 VGND 0.13047f
C9612 XThC.Tn[3].t31 VGND 0.01476f
C9613 XThC.Tn[3].t12 VGND 0.01555f
C9614 XThC.Tn[3].n61 VGND 0.03861f
C9615 XThC.Tn[3].n62 VGND 0.02405f
C9616 XThC.Tn[3].n63 VGND 0.07814f
C9617 XThC.Tn[3].n64 VGND 0.13047f
C9618 XThC.Tn[3].t33 VGND 0.01476f
C9619 XThC.Tn[3].t14 VGND 0.01555f
C9620 XThC.Tn[3].n65 VGND 0.03861f
C9621 XThC.Tn[3].n66 VGND 0.02405f
C9622 XThC.Tn[3].n67 VGND 0.07814f
C9623 XThC.Tn[3].n68 VGND 0.13047f
C9624 XThC.Tn[3].t22 VGND 0.01476f
C9625 XThC.Tn[3].t34 VGND 0.01555f
C9626 XThC.Tn[3].n69 VGND 0.03861f
C9627 XThC.Tn[3].n70 VGND 0.02405f
C9628 XThC.Tn[3].n71 VGND 0.07814f
C9629 XThC.Tn[3].n72 VGND 0.13047f
C9630 XThC.Tn[3].n73 VGND 0.76727f
C9631 XThC.Tn[3].n74 VGND 0.11064f
C9632 XThR.XTB3.Y.t1 VGND 0.06176f
C9633 XThR.XTB3.Y.n0 VGND 0.01521f
C9634 XThR.XTB3.Y.t8 VGND 0.04903f
C9635 XThR.XTB3.Y.t15 VGND 0.02889f
C9636 XThR.XTB3.Y.t13 VGND 0.04903f
C9637 XThR.XTB3.Y.t6 VGND 0.02889f
C9638 XThR.XTB3.Y.t9 VGND 0.04903f
C9639 XThR.XTB3.Y.t17 VGND 0.02889f
C9640 XThR.XTB3.Y.n1 VGND 0.08226f
C9641 XThR.XTB3.Y.n2 VGND 0.08688f
C9642 XThR.XTB3.Y.n3 VGND 0.03573f
C9643 XThR.XTB3.Y.n4 VGND 0.0707f
C9644 XThR.XTB3.Y.t12 VGND 0.04903f
C9645 XThR.XTB3.Y.t4 VGND 0.02889f
C9646 XThR.XTB3.Y.n5 VGND 0.06608f
C9647 XThR.XTB3.Y.n6 VGND 0.03236f
C9648 XThR.XTB3.Y.n7 VGND 0.02685f
C9649 XThR.XTB3.Y.t18 VGND 0.04903f
C9650 XThR.XTB3.Y.t5 VGND 0.02889f
C9651 XThR.XTB3.Y.n8 VGND 0.03005f
C9652 XThR.XTB3.Y.t7 VGND 0.04903f
C9653 XThR.XTB3.Y.t10 VGND 0.02889f
C9654 XThR.XTB3.Y.n9 VGND 0.05992f
C9655 XThR.XTB3.Y.t11 VGND 0.04903f
C9656 XThR.XTB3.Y.t16 VGND 0.02889f
C9657 XThR.XTB3.Y.n10 VGND 0.06454f
C9658 XThR.XTB3.Y.n11 VGND 0.03645f
C9659 XThR.XTB3.Y.n12 VGND 0.06034f
C9660 XThR.XTB3.Y.n13 VGND 0.03128f
C9661 XThR.XTB3.Y.n14 VGND 0.02851f
C9662 XThR.XTB3.Y.n15 VGND 0.06454f
C9663 XThR.XTB3.Y.t14 VGND 0.04903f
C9664 XThR.XTB3.Y.t3 VGND 0.02889f
C9665 XThR.XTB3.Y.n16 VGND 0.05838f
C9666 XThR.XTB3.Y.n17 VGND 0.03236f
C9667 XThR.XTB3.Y.n18 VGND 0.04707f
C9668 XThR.XTB3.Y.n19 VGND 1.31347f
C9669 XThR.XTB3.Y.t0 VGND 0.03152f
C9670 XThR.XTB3.Y.t2 VGND 0.03152f
C9671 XThR.XTB3.Y.n20 VGND 0.06766f
C9672 XThR.XTB3.Y.n21 VGND 0.157f
C9673 XThR.XTB3.Y.n22 VGND 0.03296f
C9674 XThR.XTB1.Y.t1 VGND 0.03165f
C9675 XThR.XTB1.Y.n0 VGND 0.0078f
C9676 XThR.XTB1.Y.t8 VGND 0.02512f
C9677 XThR.XTB1.Y.t15 VGND 0.0148f
C9678 XThR.XTB1.Y.t14 VGND 0.02512f
C9679 XThR.XTB1.Y.t7 VGND 0.0148f
C9680 XThR.XTB1.Y.t10 VGND 0.02512f
C9681 XThR.XTB1.Y.t18 VGND 0.0148f
C9682 XThR.XTB1.Y.n1 VGND 0.04215f
C9683 XThR.XTB1.Y.n2 VGND 0.04452f
C9684 XThR.XTB1.Y.n3 VGND 0.01831f
C9685 XThR.XTB1.Y.n4 VGND 0.03623f
C9686 XThR.XTB1.Y.t13 VGND 0.02512f
C9687 XThR.XTB1.Y.t4 VGND 0.0148f
C9688 XThR.XTB1.Y.n5 VGND 0.03386f
C9689 XThR.XTB1.Y.n6 VGND 0.01658f
C9690 XThR.XTB1.Y.n7 VGND 0.01376f
C9691 XThR.XTB1.Y.t6 VGND 0.02512f
C9692 XThR.XTB1.Y.t11 VGND 0.0148f
C9693 XThR.XTB1.Y.n8 VGND 0.0154f
C9694 XThR.XTB1.Y.t12 VGND 0.02512f
C9695 XThR.XTB1.Y.t16 VGND 0.0148f
C9696 XThR.XTB1.Y.n9 VGND 0.0307f
C9697 XThR.XTB1.Y.t17 VGND 0.02512f
C9698 XThR.XTB1.Y.t5 VGND 0.0148f
C9699 XThR.XTB1.Y.n10 VGND 0.03307f
C9700 XThR.XTB1.Y.n11 VGND 0.01868f
C9701 XThR.XTB1.Y.n12 VGND 0.03092f
C9702 XThR.XTB1.Y.n13 VGND 0.01603f
C9703 XThR.XTB1.Y.n14 VGND 0.01461f
C9704 XThR.XTB1.Y.n15 VGND 0.03307f
C9705 XThR.XTB1.Y.t3 VGND 0.02512f
C9706 XThR.XTB1.Y.t9 VGND 0.0148f
C9707 XThR.XTB1.Y.n16 VGND 0.02991f
C9708 XThR.XTB1.Y.n17 VGND 0.01658f
C9709 XThR.XTB1.Y.n18 VGND 0.02412f
C9710 XThR.XTB1.Y.n19 VGND 0.75219f
C9711 XThR.XTB1.Y.t2 VGND 0.01615f
C9712 XThR.XTB1.Y.t0 VGND 0.01615f
C9713 XThR.XTB1.Y.n20 VGND 0.03467f
C9714 XThR.XTB1.Y.n21 VGND 0.08068f
C9715 XThR.XTB1.Y.n22 VGND 0.01689f
C9716 XThR.XTB4.Y.t8 VGND 0.02956f
C9717 XThR.XTB4.Y.t15 VGND 0.05016f
C9718 XThR.XTB4.Y.t16 VGND 0.02956f
C9719 XThR.XTB4.Y.t5 VGND 0.05016f
C9720 XThR.XTB4.Y.t10 VGND 0.02956f
C9721 XThR.XTB4.Y.t17 VGND 0.05016f
C9722 XThR.XTB4.Y.n0 VGND 0.08416f
C9723 XThR.XTB4.Y.n1 VGND 0.08889f
C9724 XThR.XTB4.Y.n2 VGND 0.03656f
C9725 XThR.XTB4.Y.n3 VGND 0.07234f
C9726 XThR.XTB4.Y.t13 VGND 0.02956f
C9727 XThR.XTB4.Y.t4 VGND 0.05016f
C9728 XThR.XTB4.Y.n4 VGND 0.06761f
C9729 XThR.XTB4.Y.n5 VGND 0.0331f
C9730 XThR.XTB4.Y.n6 VGND 0.01685f
C9731 XThR.XTB4.Y.n7 VGND 0.05355f
C9732 XThR.XTB4.Y.n8 VGND 0.64921f
C9733 XThR.XTB4.Y.t14 VGND 0.02956f
C9734 XThR.XTB4.Y.t7 VGND 0.05016f
C9735 XThR.XTB4.Y.n9 VGND 0.03074f
C9736 XThR.XTB4.Y.t3 VGND 0.02956f
C9737 XThR.XTB4.Y.t12 VGND 0.05016f
C9738 XThR.XTB4.Y.n10 VGND 0.0613f
C9739 XThR.XTB4.Y.t9 VGND 0.02956f
C9740 XThR.XTB4.Y.t2 VGND 0.05016f
C9741 XThR.XTB4.Y.n11 VGND 0.06603f
C9742 XThR.XTB4.Y.n12 VGND 0.03729f
C9743 XThR.XTB4.Y.n13 VGND 0.06174f
C9744 XThR.XTB4.Y.n14 VGND 0.03201f
C9745 XThR.XTB4.Y.n15 VGND 0.02916f
C9746 XThR.XTB4.Y.n16 VGND 0.06603f
C9747 XThR.XTB4.Y.t11 VGND 0.02956f
C9748 XThR.XTB4.Y.t6 VGND 0.05016f
C9749 XThR.XTB4.Y.n17 VGND 0.05972f
C9750 XThR.XTB4.Y.n18 VGND 0.0331f
C9751 XThR.XTB4.Y.n19 VGND 0.05647f
C9752 XThR.XTB4.Y.n20 VGND 1.3092f
C9753 XThR.XTB4.Y.t1 VGND 0.06491f
C9754 XThR.XTB4.Y.n21 VGND 0.12281f
C9755 XThR.XTB4.Y.n22 VGND 0.02892f
C9756 XThR.XTB4.Y.t0 VGND 0.11919f
C9757 XThR.Tn[2].t6 VGND 0.02328f
C9758 XThR.Tn[2].t3 VGND 0.02328f
C9759 XThR.Tn[2].n0 VGND 0.04699f
C9760 XThR.Tn[2].t5 VGND 0.02328f
C9761 XThR.Tn[2].t4 VGND 0.02328f
C9762 XThR.Tn[2].n1 VGND 0.05498f
C9763 XThR.Tn[2].n2 VGND 0.16493f
C9764 XThR.Tn[2].t9 VGND 0.01513f
C9765 XThR.Tn[2].t10 VGND 0.01513f
C9766 XThR.Tn[2].n3 VGND 0.03446f
C9767 XThR.Tn[2].t8 VGND 0.01513f
C9768 XThR.Tn[2].t7 VGND 0.01513f
C9769 XThR.Tn[2].n4 VGND 0.03446f
C9770 XThR.Tn[2].t11 VGND 0.01513f
C9771 XThR.Tn[2].t1 VGND 0.01513f
C9772 XThR.Tn[2].n5 VGND 0.03446f
C9773 XThR.Tn[2].t2 VGND 0.01513f
C9774 XThR.Tn[2].t0 VGND 0.01513f
C9775 XThR.Tn[2].n6 VGND 0.05742f
C9776 XThR.Tn[2].n7 VGND 0.16411f
C9777 XThR.Tn[2].n8 VGND 0.10145f
C9778 XThR.Tn[2].n9 VGND 0.11449f
C9779 XThR.Tn[2].t27 VGND 0.01892f
C9780 XThR.Tn[2].t54 VGND 0.01992f
C9781 XThR.Tn[2].n10 VGND 0.04948f
C9782 XThR.Tn[2].n11 VGND 0.09199f
C9783 XThR.Tn[2].t67 VGND 0.01892f
C9784 XThR.Tn[2].t72 VGND 0.01992f
C9785 XThR.Tn[2].n12 VGND 0.04948f
C9786 XThR.Tn[2].t59 VGND 0.01892f
C9787 XThR.Tn[2].t65 VGND 0.01992f
C9788 XThR.Tn[2].n13 VGND 0.04946f
C9789 XThR.Tn[2].n14 VGND 0.03803f
C9790 XThR.Tn[2].n15 VGND 0.00725f
C9791 XThR.Tn[2].n16 VGND 0.11354f
C9792 XThR.Tn[2].t19 VGND 0.01892f
C9793 XThR.Tn[2].t48 VGND 0.01992f
C9794 XThR.Tn[2].n17 VGND 0.04948f
C9795 XThR.Tn[2].t14 VGND 0.01892f
C9796 XThR.Tn[2].t41 VGND 0.01992f
C9797 XThR.Tn[2].n18 VGND 0.04946f
C9798 XThR.Tn[2].n19 VGND 0.03803f
C9799 XThR.Tn[2].n20 VGND 0.00725f
C9800 XThR.Tn[2].n21 VGND 0.11354f
C9801 XThR.Tn[2].t55 VGND 0.01892f
C9802 XThR.Tn[2].t66 VGND 0.01992f
C9803 XThR.Tn[2].n22 VGND 0.04948f
C9804 XThR.Tn[2].t49 VGND 0.01892f
C9805 XThR.Tn[2].t58 VGND 0.01992f
C9806 XThR.Tn[2].n23 VGND 0.04946f
C9807 XThR.Tn[2].n24 VGND 0.03803f
C9808 XThR.Tn[2].n25 VGND 0.00725f
C9809 XThR.Tn[2].n26 VGND 0.11354f
C9810 XThR.Tn[2].t21 VGND 0.01892f
C9811 XThR.Tn[2].t32 VGND 0.01992f
C9812 XThR.Tn[2].n27 VGND 0.04948f
C9813 XThR.Tn[2].t16 VGND 0.01892f
C9814 XThR.Tn[2].t26 VGND 0.01992f
C9815 XThR.Tn[2].n28 VGND 0.04946f
C9816 XThR.Tn[2].n29 VGND 0.03803f
C9817 XThR.Tn[2].n30 VGND 0.00725f
C9818 XThR.Tn[2].n31 VGND 0.11354f
C9819 XThR.Tn[2].t39 VGND 0.01892f
C9820 XThR.Tn[2].t68 VGND 0.01992f
C9821 XThR.Tn[2].n32 VGND 0.04948f
C9822 XThR.Tn[2].t35 VGND 0.01892f
C9823 XThR.Tn[2].t60 VGND 0.01992f
C9824 XThR.Tn[2].n33 VGND 0.04946f
C9825 XThR.Tn[2].n34 VGND 0.03803f
C9826 XThR.Tn[2].n35 VGND 0.00725f
C9827 XThR.Tn[2].n36 VGND 0.11354f
C9828 XThR.Tn[2].t31 VGND 0.01892f
C9829 XThR.Tn[2].t20 VGND 0.01992f
C9830 XThR.Tn[2].n37 VGND 0.04948f
C9831 XThR.Tn[2].t25 VGND 0.01892f
C9832 XThR.Tn[2].t15 VGND 0.01992f
C9833 XThR.Tn[2].n38 VGND 0.04946f
C9834 XThR.Tn[2].n39 VGND 0.03803f
C9835 XThR.Tn[2].n40 VGND 0.00725f
C9836 XThR.Tn[2].n41 VGND 0.11354f
C9837 XThR.Tn[2].t51 VGND 0.01892f
C9838 XThR.Tn[2].t12 VGND 0.01992f
C9839 XThR.Tn[2].n42 VGND 0.04948f
C9840 XThR.Tn[2].t44 VGND 0.01892f
C9841 XThR.Tn[2].t71 VGND 0.01992f
C9842 XThR.Tn[2].n43 VGND 0.04946f
C9843 XThR.Tn[2].n44 VGND 0.03803f
C9844 XThR.Tn[2].n45 VGND 0.00725f
C9845 XThR.Tn[2].n46 VGND 0.11354f
C9846 XThR.Tn[2].t70 VGND 0.01892f
C9847 XThR.Tn[2].t30 VGND 0.01992f
C9848 XThR.Tn[2].n47 VGND 0.04948f
C9849 XThR.Tn[2].t63 VGND 0.01892f
C9850 XThR.Tn[2].t24 VGND 0.01992f
C9851 XThR.Tn[2].n48 VGND 0.04946f
C9852 XThR.Tn[2].n49 VGND 0.03803f
C9853 XThR.Tn[2].n50 VGND 0.00725f
C9854 XThR.Tn[2].n51 VGND 0.11354f
C9855 XThR.Tn[2].t23 VGND 0.01892f
C9856 XThR.Tn[2].t50 VGND 0.01992f
C9857 XThR.Tn[2].n52 VGND 0.04948f
C9858 XThR.Tn[2].t18 VGND 0.01892f
C9859 XThR.Tn[2].t42 VGND 0.01992f
C9860 XThR.Tn[2].n53 VGND 0.04946f
C9861 XThR.Tn[2].n54 VGND 0.03803f
C9862 XThR.Tn[2].n55 VGND 0.00725f
C9863 XThR.Tn[2].n56 VGND 0.11354f
C9864 XThR.Tn[2].t62 VGND 0.01892f
C9865 XThR.Tn[2].t69 VGND 0.01992f
C9866 XThR.Tn[2].n57 VGND 0.04948f
C9867 XThR.Tn[2].t56 VGND 0.01892f
C9868 XThR.Tn[2].t61 VGND 0.01992f
C9869 XThR.Tn[2].n58 VGND 0.04946f
C9870 XThR.Tn[2].n59 VGND 0.03803f
C9871 XThR.Tn[2].n60 VGND 0.00725f
C9872 XThR.Tn[2].n61 VGND 0.11354f
C9873 XThR.Tn[2].t34 VGND 0.01892f
C9874 XThR.Tn[2].t43 VGND 0.01992f
C9875 XThR.Tn[2].n62 VGND 0.04948f
C9876 XThR.Tn[2].t29 VGND 0.01892f
C9877 XThR.Tn[2].t37 VGND 0.01992f
C9878 XThR.Tn[2].n63 VGND 0.04946f
C9879 XThR.Tn[2].n64 VGND 0.03803f
C9880 XThR.Tn[2].n65 VGND 0.00725f
C9881 XThR.Tn[2].n66 VGND 0.11354f
C9882 XThR.Tn[2].t53 VGND 0.01892f
C9883 XThR.Tn[2].t13 VGND 0.01992f
C9884 XThR.Tn[2].n67 VGND 0.04948f
C9885 XThR.Tn[2].t47 VGND 0.01892f
C9886 XThR.Tn[2].t73 VGND 0.01992f
C9887 XThR.Tn[2].n68 VGND 0.04946f
C9888 XThR.Tn[2].n69 VGND 0.03803f
C9889 XThR.Tn[2].n70 VGND 0.00725f
C9890 XThR.Tn[2].n71 VGND 0.11354f
C9891 XThR.Tn[2].t22 VGND 0.01892f
C9892 XThR.Tn[2].t33 VGND 0.01992f
C9893 XThR.Tn[2].n72 VGND 0.04948f
C9894 XThR.Tn[2].t17 VGND 0.01892f
C9895 XThR.Tn[2].t28 VGND 0.01992f
C9896 XThR.Tn[2].n73 VGND 0.04946f
C9897 XThR.Tn[2].n74 VGND 0.03803f
C9898 XThR.Tn[2].n75 VGND 0.00725f
C9899 XThR.Tn[2].n76 VGND 0.11354f
C9900 XThR.Tn[2].t40 VGND 0.01892f
C9901 XThR.Tn[2].t52 VGND 0.01992f
C9902 XThR.Tn[2].n77 VGND 0.04948f
C9903 XThR.Tn[2].t36 VGND 0.01892f
C9904 XThR.Tn[2].t45 VGND 0.01992f
C9905 XThR.Tn[2].n78 VGND 0.04946f
C9906 XThR.Tn[2].n79 VGND 0.03803f
C9907 XThR.Tn[2].n80 VGND 0.00725f
C9908 XThR.Tn[2].n81 VGND 0.11354f
C9909 XThR.Tn[2].t64 VGND 0.01892f
C9910 XThR.Tn[2].t46 VGND 0.01992f
C9911 XThR.Tn[2].n82 VGND 0.04948f
C9912 XThR.Tn[2].t57 VGND 0.01892f
C9913 XThR.Tn[2].t38 VGND 0.01992f
C9914 XThR.Tn[2].n83 VGND 0.04946f
C9915 XThR.Tn[2].n84 VGND 0.03803f
C9916 XThR.Tn[2].n85 VGND 0.00725f
C9917 XThR.Tn[2].n86 VGND 0.11354f
C9918 XThR.Tn[2].n87 VGND 0.10371f
C9919 XThR.Tn[2].n88 VGND 0.22474f
C9920 XThR.Tn[3].t5 VGND 0.0233f
C9921 XThR.Tn[3].t6 VGND 0.0233f
C9922 XThR.Tn[3].n0 VGND 0.04704f
C9923 XThR.Tn[3].t4 VGND 0.0233f
C9924 XThR.Tn[3].t7 VGND 0.0233f
C9925 XThR.Tn[3].n1 VGND 0.05504f
C9926 XThR.Tn[3].n2 VGND 0.15408f
C9927 XThR.Tn[3].t11 VGND 0.01515f
C9928 XThR.Tn[3].t8 VGND 0.01515f
C9929 XThR.Tn[3].n3 VGND 0.03449f
C9930 XThR.Tn[3].t10 VGND 0.01515f
C9931 XThR.Tn[3].t9 VGND 0.01515f
C9932 XThR.Tn[3].n4 VGND 0.03449f
C9933 XThR.Tn[3].t2 VGND 0.01515f
C9934 XThR.Tn[3].t1 VGND 0.01515f
C9935 XThR.Tn[3].n5 VGND 0.05748f
C9936 XThR.Tn[3].t3 VGND 0.01515f
C9937 XThR.Tn[3].t0 VGND 0.01515f
C9938 XThR.Tn[3].n6 VGND 0.03449f
C9939 XThR.Tn[3].n7 VGND 0.16427f
C9940 XThR.Tn[3].n8 VGND 0.10155f
C9941 XThR.Tn[3].n9 VGND 0.11461f
C9942 XThR.Tn[3].t20 VGND 0.01894f
C9943 XThR.Tn[3].t48 VGND 0.01994f
C9944 XThR.Tn[3].n10 VGND 0.04953f
C9945 XThR.Tn[3].n11 VGND 0.09208f
C9946 XThR.Tn[3].t60 VGND 0.01894f
C9947 XThR.Tn[3].t66 VGND 0.01994f
C9948 XThR.Tn[3].n12 VGND 0.04953f
C9949 XThR.Tn[3].t22 VGND 0.01894f
C9950 XThR.Tn[3].t31 VGND 0.01994f
C9951 XThR.Tn[3].n13 VGND 0.04951f
C9952 XThR.Tn[3].n14 VGND 0.03807f
C9953 XThR.Tn[3].n15 VGND 0.00726f
C9954 XThR.Tn[3].n16 VGND 0.11366f
C9955 XThR.Tn[3].t13 VGND 0.01894f
C9956 XThR.Tn[3].t40 VGND 0.01994f
C9957 XThR.Tn[3].n17 VGND 0.04953f
C9958 XThR.Tn[3].t38 VGND 0.01894f
C9959 XThR.Tn[3].t67 VGND 0.01994f
C9960 XThR.Tn[3].n18 VGND 0.04951f
C9961 XThR.Tn[3].n19 VGND 0.03807f
C9962 XThR.Tn[3].n20 VGND 0.00726f
C9963 XThR.Tn[3].n21 VGND 0.11366f
C9964 XThR.Tn[3].t49 VGND 0.01894f
C9965 XThR.Tn[3].t57 VGND 0.01994f
C9966 XThR.Tn[3].n22 VGND 0.04953f
C9967 XThR.Tn[3].t12 VGND 0.01894f
C9968 XThR.Tn[3].t21 VGND 0.01994f
C9969 XThR.Tn[3].n23 VGND 0.04951f
C9970 XThR.Tn[3].n24 VGND 0.03807f
C9971 XThR.Tn[3].n25 VGND 0.00726f
C9972 XThR.Tn[3].n26 VGND 0.11366f
C9973 XThR.Tn[3].t15 VGND 0.01894f
C9974 XThR.Tn[3].t28 VGND 0.01994f
C9975 XThR.Tn[3].n27 VGND 0.04953f
C9976 XThR.Tn[3].t41 VGND 0.01894f
C9977 XThR.Tn[3].t52 VGND 0.01994f
C9978 XThR.Tn[3].n28 VGND 0.04951f
C9979 XThR.Tn[3].n29 VGND 0.03807f
C9980 XThR.Tn[3].n30 VGND 0.00726f
C9981 XThR.Tn[3].n31 VGND 0.11366f
C9982 XThR.Tn[3].t32 VGND 0.01894f
C9983 XThR.Tn[3].t61 VGND 0.01994f
C9984 XThR.Tn[3].n32 VGND 0.04953f
C9985 XThR.Tn[3].t58 VGND 0.01894f
C9986 XThR.Tn[3].t23 VGND 0.01994f
C9987 XThR.Tn[3].n33 VGND 0.04951f
C9988 XThR.Tn[3].n34 VGND 0.03807f
C9989 XThR.Tn[3].n35 VGND 0.00726f
C9990 XThR.Tn[3].n36 VGND 0.11366f
C9991 XThR.Tn[3].t27 VGND 0.01894f
C9992 XThR.Tn[3].t14 VGND 0.01994f
C9993 XThR.Tn[3].n37 VGND 0.04953f
C9994 XThR.Tn[3].t51 VGND 0.01894f
C9995 XThR.Tn[3].t39 VGND 0.01994f
C9996 XThR.Tn[3].n38 VGND 0.04951f
C9997 XThR.Tn[3].n39 VGND 0.03807f
C9998 XThR.Tn[3].n40 VGND 0.00726f
C9999 XThR.Tn[3].n41 VGND 0.11366f
C10000 XThR.Tn[3].t45 VGND 0.01894f
C10001 XThR.Tn[3].t71 VGND 0.01994f
C10002 XThR.Tn[3].n42 VGND 0.04953f
C10003 XThR.Tn[3].t69 VGND 0.01894f
C10004 XThR.Tn[3].t33 VGND 0.01994f
C10005 XThR.Tn[3].n43 VGND 0.04951f
C10006 XThR.Tn[3].n44 VGND 0.03807f
C10007 XThR.Tn[3].n45 VGND 0.00726f
C10008 XThR.Tn[3].n46 VGND 0.11366f
C10009 XThR.Tn[3].t63 VGND 0.01894f
C10010 XThR.Tn[3].t26 VGND 0.01994f
C10011 XThR.Tn[3].n47 VGND 0.04953f
C10012 XThR.Tn[3].t25 VGND 0.01894f
C10013 XThR.Tn[3].t50 VGND 0.01994f
C10014 XThR.Tn[3].n48 VGND 0.04951f
C10015 XThR.Tn[3].n49 VGND 0.03807f
C10016 XThR.Tn[3].n50 VGND 0.00726f
C10017 XThR.Tn[3].n51 VGND 0.11366f
C10018 XThR.Tn[3].t17 VGND 0.01894f
C10019 XThR.Tn[3].t44 VGND 0.01994f
C10020 XThR.Tn[3].n52 VGND 0.04953f
C10021 XThR.Tn[3].t43 VGND 0.01894f
C10022 XThR.Tn[3].t68 VGND 0.01994f
C10023 XThR.Tn[3].n53 VGND 0.04951f
C10024 XThR.Tn[3].n54 VGND 0.03807f
C10025 XThR.Tn[3].n55 VGND 0.00726f
C10026 XThR.Tn[3].n56 VGND 0.11366f
C10027 XThR.Tn[3].t55 VGND 0.01894f
C10028 XThR.Tn[3].t62 VGND 0.01994f
C10029 XThR.Tn[3].n57 VGND 0.04953f
C10030 XThR.Tn[3].t18 VGND 0.01894f
C10031 XThR.Tn[3].t24 VGND 0.01994f
C10032 XThR.Tn[3].n58 VGND 0.04951f
C10033 XThR.Tn[3].n59 VGND 0.03807f
C10034 XThR.Tn[3].n60 VGND 0.00726f
C10035 XThR.Tn[3].n61 VGND 0.11366f
C10036 XThR.Tn[3].t30 VGND 0.01894f
C10037 XThR.Tn[3].t36 VGND 0.01994f
C10038 XThR.Tn[3].n62 VGND 0.04953f
C10039 XThR.Tn[3].t54 VGND 0.01894f
C10040 XThR.Tn[3].t64 VGND 0.01994f
C10041 XThR.Tn[3].n63 VGND 0.04951f
C10042 XThR.Tn[3].n64 VGND 0.03807f
C10043 XThR.Tn[3].n65 VGND 0.00726f
C10044 XThR.Tn[3].n66 VGND 0.11366f
C10045 XThR.Tn[3].t47 VGND 0.01894f
C10046 XThR.Tn[3].t73 VGND 0.01994f
C10047 XThR.Tn[3].n67 VGND 0.04953f
C10048 XThR.Tn[3].t72 VGND 0.01894f
C10049 XThR.Tn[3].t35 VGND 0.01994f
C10050 XThR.Tn[3].n68 VGND 0.04951f
C10051 XThR.Tn[3].n69 VGND 0.03807f
C10052 XThR.Tn[3].n70 VGND 0.00726f
C10053 XThR.Tn[3].n71 VGND 0.11366f
C10054 XThR.Tn[3].t16 VGND 0.01894f
C10055 XThR.Tn[3].t29 VGND 0.01994f
C10056 XThR.Tn[3].n72 VGND 0.04953f
C10057 XThR.Tn[3].t42 VGND 0.01894f
C10058 XThR.Tn[3].t53 VGND 0.01994f
C10059 XThR.Tn[3].n73 VGND 0.04951f
C10060 XThR.Tn[3].n74 VGND 0.03807f
C10061 XThR.Tn[3].n75 VGND 0.00726f
C10062 XThR.Tn[3].n76 VGND 0.11366f
C10063 XThR.Tn[3].t34 VGND 0.01894f
C10064 XThR.Tn[3].t46 VGND 0.01994f
C10065 XThR.Tn[3].n77 VGND 0.04953f
C10066 XThR.Tn[3].t59 VGND 0.01894f
C10067 XThR.Tn[3].t70 VGND 0.01994f
C10068 XThR.Tn[3].n78 VGND 0.04951f
C10069 XThR.Tn[3].n79 VGND 0.03807f
C10070 XThR.Tn[3].n80 VGND 0.00726f
C10071 XThR.Tn[3].n81 VGND 0.11366f
C10072 XThR.Tn[3].t56 VGND 0.01894f
C10073 XThR.Tn[3].t37 VGND 0.01994f
C10074 XThR.Tn[3].n82 VGND 0.04953f
C10075 XThR.Tn[3].t19 VGND 0.01894f
C10076 XThR.Tn[3].t65 VGND 0.01994f
C10077 XThR.Tn[3].n83 VGND 0.04951f
C10078 XThR.Tn[3].n84 VGND 0.03807f
C10079 XThR.Tn[3].n85 VGND 0.00726f
C10080 XThR.Tn[3].n86 VGND 0.11366f
C10081 XThR.Tn[3].n87 VGND 0.10381f
C10082 XThR.Tn[3].n88 VGND 0.22993f
C10083 XThR.Tn[3].n89 VGND 0.04877f
C10084 XThC.Tn[11].t7 VGND 0.01298f
C10085 XThC.Tn[11].t6 VGND 0.01298f
C10086 XThC.Tn[11].n0 VGND 0.03238f
C10087 XThC.Tn[11].t4 VGND 0.01298f
C10088 XThC.Tn[11].t5 VGND 0.01298f
C10089 XThC.Tn[11].n1 VGND 0.02597f
C10090 XThC.Tn[11].n2 VGND 0.05988f
C10091 XThC.Tn[11].t33 VGND 0.01623f
C10092 XThC.Tn[11].t38 VGND 0.01709f
C10093 XThC.Tn[11].n3 VGND 0.04246f
C10094 XThC.Tn[11].n4 VGND 0.02645f
C10095 XThC.Tn[11].n5 VGND 0.08569f
C10096 XThC.Tn[11].t42 VGND 0.01623f
C10097 XThC.Tn[11].t15 VGND 0.01709f
C10098 XThC.Tn[11].n6 VGND 0.04246f
C10099 XThC.Tn[11].n7 VGND 0.02645f
C10100 XThC.Tn[11].n8 VGND 0.08593f
C10101 XThC.Tn[11].n9 VGND 0.14347f
C10102 XThC.Tn[11].t22 VGND 0.01623f
C10103 XThC.Tn[11].t28 VGND 0.01709f
C10104 XThC.Tn[11].n10 VGND 0.04246f
C10105 XThC.Tn[11].n11 VGND 0.02645f
C10106 XThC.Tn[11].n12 VGND 0.08593f
C10107 XThC.Tn[11].n13 VGND 0.14347f
C10108 XThC.Tn[11].t24 VGND 0.01623f
C10109 XThC.Tn[11].t30 VGND 0.01709f
C10110 XThC.Tn[11].n14 VGND 0.04246f
C10111 XThC.Tn[11].n15 VGND 0.02645f
C10112 XThC.Tn[11].n16 VGND 0.08593f
C10113 XThC.Tn[11].n17 VGND 0.14347f
C10114 XThC.Tn[11].t35 VGND 0.01623f
C10115 XThC.Tn[11].t39 VGND 0.01709f
C10116 XThC.Tn[11].n18 VGND 0.04246f
C10117 XThC.Tn[11].n19 VGND 0.02645f
C10118 XThC.Tn[11].n20 VGND 0.08593f
C10119 XThC.Tn[11].n21 VGND 0.14347f
C10120 XThC.Tn[11].t13 VGND 0.01623f
C10121 XThC.Tn[11].t18 VGND 0.01709f
C10122 XThC.Tn[11].n22 VGND 0.04246f
C10123 XThC.Tn[11].n23 VGND 0.02645f
C10124 XThC.Tn[11].n24 VGND 0.08593f
C10125 XThC.Tn[11].n25 VGND 0.14347f
C10126 XThC.Tn[11].t25 VGND 0.01623f
C10127 XThC.Tn[11].t31 VGND 0.01709f
C10128 XThC.Tn[11].n26 VGND 0.04246f
C10129 XThC.Tn[11].n27 VGND 0.02645f
C10130 XThC.Tn[11].n28 VGND 0.08593f
C10131 XThC.Tn[11].n29 VGND 0.14347f
C10132 XThC.Tn[11].t36 VGND 0.01623f
C10133 XThC.Tn[11].t41 VGND 0.01709f
C10134 XThC.Tn[11].n30 VGND 0.04246f
C10135 XThC.Tn[11].n31 VGND 0.02645f
C10136 XThC.Tn[11].n32 VGND 0.08593f
C10137 XThC.Tn[11].n33 VGND 0.14347f
C10138 XThC.Tn[11].t37 VGND 0.01623f
C10139 XThC.Tn[11].t43 VGND 0.01709f
C10140 XThC.Tn[11].n34 VGND 0.04246f
C10141 XThC.Tn[11].n35 VGND 0.02645f
C10142 XThC.Tn[11].n36 VGND 0.08593f
C10143 XThC.Tn[11].n37 VGND 0.14347f
C10144 XThC.Tn[11].t14 VGND 0.01623f
C10145 XThC.Tn[11].t20 VGND 0.01709f
C10146 XThC.Tn[11].n38 VGND 0.04246f
C10147 XThC.Tn[11].n39 VGND 0.02645f
C10148 XThC.Tn[11].n40 VGND 0.08593f
C10149 XThC.Tn[11].n41 VGND 0.14347f
C10150 XThC.Tn[11].t27 VGND 0.01623f
C10151 XThC.Tn[11].t32 VGND 0.01709f
C10152 XThC.Tn[11].n42 VGND 0.04246f
C10153 XThC.Tn[11].n43 VGND 0.02645f
C10154 XThC.Tn[11].n44 VGND 0.08593f
C10155 XThC.Tn[11].n45 VGND 0.14347f
C10156 XThC.Tn[11].t29 VGND 0.01623f
C10157 XThC.Tn[11].t34 VGND 0.01709f
C10158 XThC.Tn[11].n46 VGND 0.04246f
C10159 XThC.Tn[11].n47 VGND 0.02645f
C10160 XThC.Tn[11].n48 VGND 0.08593f
C10161 XThC.Tn[11].n49 VGND 0.14347f
C10162 XThC.Tn[11].t16 VGND 0.01623f
C10163 XThC.Tn[11].t21 VGND 0.01709f
C10164 XThC.Tn[11].n50 VGND 0.04246f
C10165 XThC.Tn[11].n51 VGND 0.02645f
C10166 XThC.Tn[11].n52 VGND 0.08593f
C10167 XThC.Tn[11].n53 VGND 0.14347f
C10168 XThC.Tn[11].t17 VGND 0.01623f
C10169 XThC.Tn[11].t23 VGND 0.01709f
C10170 XThC.Tn[11].n54 VGND 0.04246f
C10171 XThC.Tn[11].n55 VGND 0.02645f
C10172 XThC.Tn[11].n56 VGND 0.08593f
C10173 XThC.Tn[11].n57 VGND 0.14347f
C10174 XThC.Tn[11].t19 VGND 0.01623f
C10175 XThC.Tn[11].t26 VGND 0.01709f
C10176 XThC.Tn[11].n58 VGND 0.04246f
C10177 XThC.Tn[11].n59 VGND 0.02645f
C10178 XThC.Tn[11].n60 VGND 0.08593f
C10179 XThC.Tn[11].n61 VGND 0.14347f
C10180 XThC.Tn[11].t40 VGND 0.01623f
C10181 XThC.Tn[11].t12 VGND 0.01709f
C10182 XThC.Tn[11].n62 VGND 0.04246f
C10183 XThC.Tn[11].n63 VGND 0.02645f
C10184 XThC.Tn[11].n64 VGND 0.08593f
C10185 XThC.Tn[11].n65 VGND 0.14347f
C10186 XThC.Tn[11].n66 VGND 0.66583f
C10187 XThC.Tn[11].n67 VGND 0.26082f
C10188 XThC.Tn[11].t1 VGND 0.01998f
C10189 XThC.Tn[11].t2 VGND 0.01998f
C10190 XThC.Tn[11].n68 VGND 0.04316f
C10191 XThC.Tn[11].t0 VGND 0.01998f
C10192 XThC.Tn[11].t3 VGND 0.01998f
C10193 XThC.Tn[11].n69 VGND 0.06803f
C10194 XThC.Tn[11].n70 VGND 0.18017f
C10195 XThC.Tn[11].n71 VGND 0.01326f
C10196 XThC.Tn[11].t8 VGND 0.01998f
C10197 XThC.Tn[11].t11 VGND 0.01998f
C10198 XThC.Tn[11].n72 VGND 0.06065f
C10199 XThC.Tn[11].t10 VGND 0.01998f
C10200 XThC.Tn[11].t9 VGND 0.01998f
C10201 XThC.Tn[11].n73 VGND 0.0444f
C10202 XThC.Tn[11].n74 VGND 0.19763f
C10203 XThC.XTB3.Y.t1 VGND 0.06296f
C10204 XThC.XTB3.Y.n0 VGND 0.04069f
C10205 XThC.XTB3.Y.n1 VGND 0.05192f
C10206 XThC.XTB3.Y.t2 VGND 0.03159f
C10207 XThC.XTB3.Y.t0 VGND 0.03159f
C10208 XThC.XTB3.Y.n2 VGND 0.06782f
C10209 XThC.XTB3.Y.t10 VGND 0.04914f
C10210 XThC.XTB3.Y.t17 VGND 0.02896f
C10211 XThC.XTB3.Y.n3 VGND 0.05852f
C10212 XThC.XTB3.Y.t14 VGND 0.04914f
C10213 XThC.XTB3.Y.t5 VGND 0.02896f
C10214 XThC.XTB3.Y.n4 VGND 0.03012f
C10215 XThC.XTB3.Y.t15 VGND 0.04914f
C10216 XThC.XTB3.Y.t6 VGND 0.02896f
C10217 XThC.XTB3.Y.n5 VGND 0.06469f
C10218 XThC.XTB3.Y.t3 VGND 0.04914f
C10219 XThC.XTB3.Y.t9 VGND 0.02896f
C10220 XThC.XTB3.Y.n6 VGND 0.06006f
C10221 XThC.XTB3.Y.n7 VGND 0.03654f
C10222 XThC.XTB3.Y.n8 VGND 0.06049f
C10223 XThC.XTB3.Y.n9 VGND 0.0234f
C10224 XThC.XTB3.Y.n10 VGND 0.02857f
C10225 XThC.XTB3.Y.n11 VGND 0.06469f
C10226 XThC.XTB3.Y.n12 VGND 0.03243f
C10227 XThC.XTB3.Y.n13 VGND 0.05514f
C10228 XThC.XTB3.Y.t16 VGND 0.04914f
C10229 XThC.XTB3.Y.t7 VGND 0.02896f
C10230 XThC.XTB3.Y.n14 VGND 0.06624f
C10231 XThC.XTB3.Y.t4 VGND 0.04914f
C10232 XThC.XTB3.Y.t13 VGND 0.02896f
C10233 XThC.XTB3.Y.t12 VGND 0.04914f
C10234 XThC.XTB3.Y.t18 VGND 0.02896f
C10235 XThC.XTB3.Y.t11 VGND 0.04914f
C10236 XThC.XTB3.Y.t8 VGND 0.02896f
C10237 XThC.XTB3.Y.n15 VGND 0.08245f
C10238 XThC.XTB3.Y.n16 VGND 0.08709f
C10239 XThC.XTB3.Y.n17 VGND 0.03356f
C10240 XThC.XTB3.Y.n18 VGND 0.07087f
C10241 XThC.XTB3.Y.n19 VGND 0.03243f
C10242 XThC.XTB3.Y.n20 VGND 0.02691f
C10243 XThC.XTB3.Y.n21 VGND 1.39635f
C10244 XThC.XTB3.Y.n22 VGND 0.14933f
C10245 XThC.Tn[9].t5 VGND 0.01308f
C10246 XThC.Tn[9].t4 VGND 0.01308f
C10247 XThC.Tn[9].n0 VGND 0.03261f
C10248 XThC.Tn[9].t6 VGND 0.01308f
C10249 XThC.Tn[9].t7 VGND 0.01308f
C10250 XThC.Tn[9].n1 VGND 0.02615f
C10251 XThC.Tn[9].n2 VGND 0.0603f
C10252 XThC.Tn[9].t38 VGND 0.01635f
C10253 XThC.Tn[9].t33 VGND 0.01722f
C10254 XThC.Tn[9].n3 VGND 0.04276f
C10255 XThC.Tn[9].n4 VGND 0.02664f
C10256 XThC.Tn[9].n5 VGND 0.08629f
C10257 XThC.Tn[9].t16 VGND 0.01635f
C10258 XThC.Tn[9].t42 VGND 0.01722f
C10259 XThC.Tn[9].n6 VGND 0.04276f
C10260 XThC.Tn[9].n7 VGND 0.02664f
C10261 XThC.Tn[9].n8 VGND 0.08654f
C10262 XThC.Tn[9].n9 VGND 0.14448f
C10263 XThC.Tn[9].t28 VGND 0.01635f
C10264 XThC.Tn[9].t22 VGND 0.01722f
C10265 XThC.Tn[9].n10 VGND 0.04276f
C10266 XThC.Tn[9].n11 VGND 0.02664f
C10267 XThC.Tn[9].n12 VGND 0.08654f
C10268 XThC.Tn[9].n13 VGND 0.14448f
C10269 XThC.Tn[9].t30 VGND 0.01635f
C10270 XThC.Tn[9].t23 VGND 0.01722f
C10271 XThC.Tn[9].n14 VGND 0.04276f
C10272 XThC.Tn[9].n15 VGND 0.02664f
C10273 XThC.Tn[9].n16 VGND 0.08654f
C10274 XThC.Tn[9].n17 VGND 0.14448f
C10275 XThC.Tn[9].t40 VGND 0.01635f
C10276 XThC.Tn[9].t35 VGND 0.01722f
C10277 XThC.Tn[9].n18 VGND 0.04276f
C10278 XThC.Tn[9].n19 VGND 0.02664f
C10279 XThC.Tn[9].n20 VGND 0.08654f
C10280 XThC.Tn[9].n21 VGND 0.14448f
C10281 XThC.Tn[9].t18 VGND 0.01635f
C10282 XThC.Tn[9].t12 VGND 0.01722f
C10283 XThC.Tn[9].n22 VGND 0.04276f
C10284 XThC.Tn[9].n23 VGND 0.02664f
C10285 XThC.Tn[9].n24 VGND 0.08654f
C10286 XThC.Tn[9].n25 VGND 0.14448f
C10287 XThC.Tn[9].t31 VGND 0.01635f
C10288 XThC.Tn[9].t25 VGND 0.01722f
C10289 XThC.Tn[9].n26 VGND 0.04276f
C10290 XThC.Tn[9].n27 VGND 0.02664f
C10291 XThC.Tn[9].n28 VGND 0.08654f
C10292 XThC.Tn[9].n29 VGND 0.14448f
C10293 XThC.Tn[9].t41 VGND 0.01635f
C10294 XThC.Tn[9].t36 VGND 0.01722f
C10295 XThC.Tn[9].n30 VGND 0.04276f
C10296 XThC.Tn[9].n31 VGND 0.02664f
C10297 XThC.Tn[9].n32 VGND 0.08654f
C10298 XThC.Tn[9].n33 VGND 0.14448f
C10299 XThC.Tn[9].t43 VGND 0.01635f
C10300 XThC.Tn[9].t37 VGND 0.01722f
C10301 XThC.Tn[9].n34 VGND 0.04276f
C10302 XThC.Tn[9].n35 VGND 0.02664f
C10303 XThC.Tn[9].n36 VGND 0.08654f
C10304 XThC.Tn[9].n37 VGND 0.14448f
C10305 XThC.Tn[9].t20 VGND 0.01635f
C10306 XThC.Tn[9].t14 VGND 0.01722f
C10307 XThC.Tn[9].n38 VGND 0.04276f
C10308 XThC.Tn[9].n39 VGND 0.02664f
C10309 XThC.Tn[9].n40 VGND 0.08654f
C10310 XThC.Tn[9].n41 VGND 0.14448f
C10311 XThC.Tn[9].t32 VGND 0.01635f
C10312 XThC.Tn[9].t27 VGND 0.01722f
C10313 XThC.Tn[9].n42 VGND 0.04276f
C10314 XThC.Tn[9].n43 VGND 0.02664f
C10315 XThC.Tn[9].n44 VGND 0.08654f
C10316 XThC.Tn[9].n45 VGND 0.14448f
C10317 XThC.Tn[9].t34 VGND 0.01635f
C10318 XThC.Tn[9].t29 VGND 0.01722f
C10319 XThC.Tn[9].n46 VGND 0.04276f
C10320 XThC.Tn[9].n47 VGND 0.02664f
C10321 XThC.Tn[9].n48 VGND 0.08654f
C10322 XThC.Tn[9].n49 VGND 0.14448f
C10323 XThC.Tn[9].t21 VGND 0.01635f
C10324 XThC.Tn[9].t15 VGND 0.01722f
C10325 XThC.Tn[9].n50 VGND 0.04276f
C10326 XThC.Tn[9].n51 VGND 0.02664f
C10327 XThC.Tn[9].n52 VGND 0.08654f
C10328 XThC.Tn[9].n53 VGND 0.14448f
C10329 XThC.Tn[9].t24 VGND 0.01635f
C10330 XThC.Tn[9].t17 VGND 0.01722f
C10331 XThC.Tn[9].n54 VGND 0.04276f
C10332 XThC.Tn[9].n55 VGND 0.02664f
C10333 XThC.Tn[9].n56 VGND 0.08654f
C10334 XThC.Tn[9].n57 VGND 0.14448f
C10335 XThC.Tn[9].t26 VGND 0.01635f
C10336 XThC.Tn[9].t19 VGND 0.01722f
C10337 XThC.Tn[9].n58 VGND 0.04276f
C10338 XThC.Tn[9].n59 VGND 0.02664f
C10339 XThC.Tn[9].n60 VGND 0.08654f
C10340 XThC.Tn[9].n61 VGND 0.14448f
C10341 XThC.Tn[9].t13 VGND 0.01635f
C10342 XThC.Tn[9].t39 VGND 0.01722f
C10343 XThC.Tn[9].n62 VGND 0.04276f
C10344 XThC.Tn[9].n63 VGND 0.02664f
C10345 XThC.Tn[9].n64 VGND 0.08654f
C10346 XThC.Tn[9].n65 VGND 0.14448f
C10347 XThC.Tn[9].n66 VGND 0.62105f
C10348 XThC.Tn[9].n67 VGND 0.26267f
C10349 XThC.Tn[9].t0 VGND 0.02012f
C10350 XThC.Tn[9].t3 VGND 0.02012f
C10351 XThC.Tn[9].n68 VGND 0.04346f
C10352 XThC.Tn[9].t2 VGND 0.02012f
C10353 XThC.Tn[9].t1 VGND 0.02012f
C10354 XThC.Tn[9].n69 VGND 0.06851f
C10355 XThC.Tn[9].n70 VGND 0.18145f
C10356 XThC.Tn[9].n71 VGND 0.01336f
C10357 XThC.Tn[9].t9 VGND 0.02012f
C10358 XThC.Tn[9].t8 VGND 0.02012f
C10359 XThC.Tn[9].n72 VGND 0.06108f
C10360 XThC.Tn[9].t11 VGND 0.02012f
C10361 XThC.Tn[9].t10 VGND 0.02012f
C10362 XThC.Tn[9].n73 VGND 0.04472f
C10363 XThC.Tn[9].n74 VGND 0.19902f
C10364 XThR.Tn[10].t7 VGND 0.02429f
C10365 XThR.Tn[10].t5 VGND 0.02429f
C10366 XThR.Tn[10].n0 VGND 0.07376f
C10367 XThR.Tn[10].t8 VGND 0.02429f
C10368 XThR.Tn[10].t6 VGND 0.02429f
C10369 XThR.Tn[10].n1 VGND 0.054f
C10370 XThR.Tn[10].n2 VGND 0.24556f
C10371 XThR.Tn[10].t9 VGND 0.02429f
C10372 XThR.Tn[10].t11 VGND 0.02429f
C10373 XThR.Tn[10].n3 VGND 0.05249f
C10374 XThR.Tn[10].t1 VGND 0.02429f
C10375 XThR.Tn[10].t10 VGND 0.02429f
C10376 XThR.Tn[10].n4 VGND 0.07989f
C10377 XThR.Tn[10].n5 VGND 0.22183f
C10378 XThR.Tn[10].n6 VGND 0.01093f
C10379 XThR.Tn[10].t20 VGND 0.01974f
C10380 XThR.Tn[10].t48 VGND 0.02079f
C10381 XThR.Tn[10].n7 VGND 0.05163f
C10382 XThR.Tn[10].n8 VGND 0.09599f
C10383 XThR.Tn[10].t60 VGND 0.01974f
C10384 XThR.Tn[10].t64 VGND 0.02079f
C10385 XThR.Tn[10].n9 VGND 0.05163f
C10386 XThR.Tn[10].t37 VGND 0.01974f
C10387 XThR.Tn[10].t44 VGND 0.02079f
C10388 XThR.Tn[10].n10 VGND 0.05161f
C10389 XThR.Tn[10].n11 VGND 0.03969f
C10390 XThR.Tn[10].n12 VGND 0.00757f
C10391 XThR.Tn[10].n13 VGND 0.11849f
C10392 XThR.Tn[10].t12 VGND 0.01974f
C10393 XThR.Tn[10].t42 VGND 0.02079f
C10394 XThR.Tn[10].n14 VGND 0.05163f
C10395 XThR.Tn[10].t53 VGND 0.01974f
C10396 XThR.Tn[10].t19 VGND 0.02079f
C10397 XThR.Tn[10].n15 VGND 0.05161f
C10398 XThR.Tn[10].n16 VGND 0.03969f
C10399 XThR.Tn[10].n17 VGND 0.00757f
C10400 XThR.Tn[10].n18 VGND 0.11849f
C10401 XThR.Tn[10].t50 VGND 0.01974f
C10402 XThR.Tn[10].t59 VGND 0.02079f
C10403 XThR.Tn[10].n19 VGND 0.05163f
C10404 XThR.Tn[10].t30 VGND 0.01974f
C10405 XThR.Tn[10].t36 VGND 0.02079f
C10406 XThR.Tn[10].n20 VGND 0.05161f
C10407 XThR.Tn[10].n21 VGND 0.03969f
C10408 XThR.Tn[10].n22 VGND 0.00757f
C10409 XThR.Tn[10].n23 VGND 0.11849f
C10410 XThR.Tn[10].t14 VGND 0.01974f
C10411 XThR.Tn[10].t27 VGND 0.02079f
C10412 XThR.Tn[10].n24 VGND 0.05163f
C10413 XThR.Tn[10].t55 VGND 0.01974f
C10414 XThR.Tn[10].t67 VGND 0.02079f
C10415 XThR.Tn[10].n25 VGND 0.05161f
C10416 XThR.Tn[10].n26 VGND 0.03969f
C10417 XThR.Tn[10].n27 VGND 0.00757f
C10418 XThR.Tn[10].n28 VGND 0.11849f
C10419 XThR.Tn[10].t31 VGND 0.01974f
C10420 XThR.Tn[10].t61 VGND 0.02079f
C10421 XThR.Tn[10].n29 VGND 0.05163f
C10422 XThR.Tn[10].t72 VGND 0.01974f
C10423 XThR.Tn[10].t39 VGND 0.02079f
C10424 XThR.Tn[10].n30 VGND 0.05161f
C10425 XThR.Tn[10].n31 VGND 0.03969f
C10426 XThR.Tn[10].n32 VGND 0.00757f
C10427 XThR.Tn[10].n33 VGND 0.11849f
C10428 XThR.Tn[10].t26 VGND 0.01974f
C10429 XThR.Tn[10].t13 VGND 0.02079f
C10430 XThR.Tn[10].n34 VGND 0.05163f
C10431 XThR.Tn[10].t66 VGND 0.01974f
C10432 XThR.Tn[10].t54 VGND 0.02079f
C10433 XThR.Tn[10].n35 VGND 0.05161f
C10434 XThR.Tn[10].n36 VGND 0.03969f
C10435 XThR.Tn[10].n37 VGND 0.00757f
C10436 XThR.Tn[10].n38 VGND 0.11849f
C10437 XThR.Tn[10].t45 VGND 0.01974f
C10438 XThR.Tn[10].t70 VGND 0.02079f
C10439 XThR.Tn[10].n39 VGND 0.05163f
C10440 XThR.Tn[10].t22 VGND 0.01974f
C10441 XThR.Tn[10].t49 VGND 0.02079f
C10442 XThR.Tn[10].n40 VGND 0.05161f
C10443 XThR.Tn[10].n41 VGND 0.03969f
C10444 XThR.Tn[10].n42 VGND 0.00757f
C10445 XThR.Tn[10].n43 VGND 0.11849f
C10446 XThR.Tn[10].t63 VGND 0.01974f
C10447 XThR.Tn[10].t25 VGND 0.02079f
C10448 XThR.Tn[10].n44 VGND 0.05163f
C10449 XThR.Tn[10].t41 VGND 0.01974f
C10450 XThR.Tn[10].t65 VGND 0.02079f
C10451 XThR.Tn[10].n45 VGND 0.05161f
C10452 XThR.Tn[10].n46 VGND 0.03969f
C10453 XThR.Tn[10].n47 VGND 0.00757f
C10454 XThR.Tn[10].n48 VGND 0.11849f
C10455 XThR.Tn[10].t18 VGND 0.01974f
C10456 XThR.Tn[10].t43 VGND 0.02079f
C10457 XThR.Tn[10].n49 VGND 0.05163f
C10458 XThR.Tn[10].t58 VGND 0.01974f
C10459 XThR.Tn[10].t21 VGND 0.02079f
C10460 XThR.Tn[10].n50 VGND 0.05161f
C10461 XThR.Tn[10].n51 VGND 0.03969f
C10462 XThR.Tn[10].n52 VGND 0.00757f
C10463 XThR.Tn[10].n53 VGND 0.11849f
C10464 XThR.Tn[10].t52 VGND 0.01974f
C10465 XThR.Tn[10].t62 VGND 0.02079f
C10466 XThR.Tn[10].n54 VGND 0.05163f
C10467 XThR.Tn[10].t33 VGND 0.01974f
C10468 XThR.Tn[10].t40 VGND 0.02079f
C10469 XThR.Tn[10].n55 VGND 0.05161f
C10470 XThR.Tn[10].n56 VGND 0.03969f
C10471 XThR.Tn[10].n57 VGND 0.00757f
C10472 XThR.Tn[10].n58 VGND 0.11849f
C10473 XThR.Tn[10].t29 VGND 0.01974f
C10474 XThR.Tn[10].t35 VGND 0.02079f
C10475 XThR.Tn[10].n59 VGND 0.05163f
C10476 XThR.Tn[10].t69 VGND 0.01974f
C10477 XThR.Tn[10].t15 VGND 0.02079f
C10478 XThR.Tn[10].n60 VGND 0.05161f
C10479 XThR.Tn[10].n61 VGND 0.03969f
C10480 XThR.Tn[10].n62 VGND 0.00757f
C10481 XThR.Tn[10].n63 VGND 0.11849f
C10482 XThR.Tn[10].t47 VGND 0.01974f
C10483 XThR.Tn[10].t71 VGND 0.02079f
C10484 XThR.Tn[10].n64 VGND 0.05163f
C10485 XThR.Tn[10].t24 VGND 0.01974f
C10486 XThR.Tn[10].t51 VGND 0.02079f
C10487 XThR.Tn[10].n65 VGND 0.05161f
C10488 XThR.Tn[10].n66 VGND 0.03969f
C10489 XThR.Tn[10].n67 VGND 0.00757f
C10490 XThR.Tn[10].n68 VGND 0.11849f
C10491 XThR.Tn[10].t16 VGND 0.01974f
C10492 XThR.Tn[10].t28 VGND 0.02079f
C10493 XThR.Tn[10].n69 VGND 0.05163f
C10494 XThR.Tn[10].t57 VGND 0.01974f
C10495 XThR.Tn[10].t68 VGND 0.02079f
C10496 XThR.Tn[10].n70 VGND 0.05161f
C10497 XThR.Tn[10].n71 VGND 0.03969f
C10498 XThR.Tn[10].n72 VGND 0.00757f
C10499 XThR.Tn[10].n73 VGND 0.11849f
C10500 XThR.Tn[10].t32 VGND 0.01974f
C10501 XThR.Tn[10].t46 VGND 0.02079f
C10502 XThR.Tn[10].n74 VGND 0.05163f
C10503 XThR.Tn[10].t73 VGND 0.01974f
C10504 XThR.Tn[10].t23 VGND 0.02079f
C10505 XThR.Tn[10].n75 VGND 0.05161f
C10506 XThR.Tn[10].n76 VGND 0.03969f
C10507 XThR.Tn[10].n77 VGND 0.00757f
C10508 XThR.Tn[10].n78 VGND 0.11849f
C10509 XThR.Tn[10].t56 VGND 0.01974f
C10510 XThR.Tn[10].t38 VGND 0.02079f
C10511 XThR.Tn[10].n79 VGND 0.05163f
C10512 XThR.Tn[10].t34 VGND 0.01974f
C10513 XThR.Tn[10].t17 VGND 0.02079f
C10514 XThR.Tn[10].n80 VGND 0.05161f
C10515 XThR.Tn[10].n81 VGND 0.03969f
C10516 XThR.Tn[10].n82 VGND 0.00757f
C10517 XThR.Tn[10].n83 VGND 0.11849f
C10518 XThR.Tn[10].n84 VGND 0.10822f
C10519 XThR.Tn[10].n85 VGND 0.33317f
C10520 XThR.Tn[10].t2 VGND 0.01579f
C10521 XThR.Tn[10].t4 VGND 0.01579f
C10522 XThR.Tn[10].n86 VGND 0.03938f
C10523 XThR.Tn[10].t3 VGND 0.01579f
C10524 XThR.Tn[10].t0 VGND 0.01579f
C10525 XThR.Tn[10].n87 VGND 0.03158f
C10526 XThR.Tn[10].n88 VGND 0.07282f
C10527 XThR.Tn[1].t4 VGND 0.02319f
C10528 XThR.Tn[1].t5 VGND 0.02319f
C10529 XThR.Tn[1].n0 VGND 0.04681f
C10530 XThR.Tn[1].t7 VGND 0.02319f
C10531 XThR.Tn[1].t6 VGND 0.02319f
C10532 XThR.Tn[1].n1 VGND 0.05477f
C10533 XThR.Tn[1].n2 VGND 0.15332f
C10534 XThR.Tn[1].t11 VGND 0.01507f
C10535 XThR.Tn[1].t8 VGND 0.01507f
C10536 XThR.Tn[1].n3 VGND 0.03432f
C10537 XThR.Tn[1].t10 VGND 0.01507f
C10538 XThR.Tn[1].t9 VGND 0.01507f
C10539 XThR.Tn[1].n4 VGND 0.03432f
C10540 XThR.Tn[1].t2 VGND 0.01507f
C10541 XThR.Tn[1].t1 VGND 0.01507f
C10542 XThR.Tn[1].n5 VGND 0.03432f
C10543 XThR.Tn[1].t3 VGND 0.01507f
C10544 XThR.Tn[1].t0 VGND 0.01507f
C10545 XThR.Tn[1].n6 VGND 0.05719f
C10546 XThR.Tn[1].n7 VGND 0.16346f
C10547 XThR.Tn[1].n8 VGND 0.10105f
C10548 XThR.Tn[1].n9 VGND 0.11404f
C10549 XThR.Tn[1].t27 VGND 0.01884f
C10550 XThR.Tn[1].t57 VGND 0.01984f
C10551 XThR.Tn[1].n10 VGND 0.04928f
C10552 XThR.Tn[1].n11 VGND 0.09162f
C10553 XThR.Tn[1].t69 VGND 0.01884f
C10554 XThR.Tn[1].t12 VGND 0.01984f
C10555 XThR.Tn[1].n12 VGND 0.04928f
C10556 XThR.Tn[1].t64 VGND 0.01884f
C10557 XThR.Tn[1].t73 VGND 0.01984f
C10558 XThR.Tn[1].n13 VGND 0.04927f
C10559 XThR.Tn[1].n14 VGND 0.03788f
C10560 XThR.Tn[1].n15 VGND 0.00722f
C10561 XThR.Tn[1].n16 VGND 0.1131f
C10562 XThR.Tn[1].t22 VGND 0.01884f
C10563 XThR.Tn[1].t50 VGND 0.01984f
C10564 XThR.Tn[1].n17 VGND 0.04928f
C10565 XThR.Tn[1].t17 VGND 0.01884f
C10566 XThR.Tn[1].t46 VGND 0.01984f
C10567 XThR.Tn[1].n18 VGND 0.04927f
C10568 XThR.Tn[1].n19 VGND 0.03788f
C10569 XThR.Tn[1].n20 VGND 0.00722f
C10570 XThR.Tn[1].n21 VGND 0.1131f
C10571 XThR.Tn[1].t58 VGND 0.01884f
C10572 XThR.Tn[1].t68 VGND 0.01984f
C10573 XThR.Tn[1].n22 VGND 0.04928f
C10574 XThR.Tn[1].t56 VGND 0.01884f
C10575 XThR.Tn[1].t62 VGND 0.01984f
C10576 XThR.Tn[1].n23 VGND 0.04927f
C10577 XThR.Tn[1].n24 VGND 0.03788f
C10578 XThR.Tn[1].n25 VGND 0.00722f
C10579 XThR.Tn[1].n26 VGND 0.1131f
C10580 XThR.Tn[1].t24 VGND 0.01884f
C10581 XThR.Tn[1].t35 VGND 0.01984f
C10582 XThR.Tn[1].n27 VGND 0.04928f
C10583 XThR.Tn[1].t19 VGND 0.01884f
C10584 XThR.Tn[1].t30 VGND 0.01984f
C10585 XThR.Tn[1].n28 VGND 0.04927f
C10586 XThR.Tn[1].n29 VGND 0.03788f
C10587 XThR.Tn[1].n30 VGND 0.00722f
C10588 XThR.Tn[1].n31 VGND 0.1131f
C10589 XThR.Tn[1].t40 VGND 0.01884f
C10590 XThR.Tn[1].t70 VGND 0.01984f
C10591 XThR.Tn[1].n32 VGND 0.04928f
C10592 XThR.Tn[1].t38 VGND 0.01884f
C10593 XThR.Tn[1].t65 VGND 0.01984f
C10594 XThR.Tn[1].n33 VGND 0.04927f
C10595 XThR.Tn[1].n34 VGND 0.03788f
C10596 XThR.Tn[1].n35 VGND 0.00722f
C10597 XThR.Tn[1].n36 VGND 0.1131f
C10598 XThR.Tn[1].t34 VGND 0.01884f
C10599 XThR.Tn[1].t23 VGND 0.01984f
C10600 XThR.Tn[1].n37 VGND 0.04928f
C10601 XThR.Tn[1].t29 VGND 0.01884f
C10602 XThR.Tn[1].t18 VGND 0.01984f
C10603 XThR.Tn[1].n38 VGND 0.04927f
C10604 XThR.Tn[1].n39 VGND 0.03788f
C10605 XThR.Tn[1].n40 VGND 0.00722f
C10606 XThR.Tn[1].n41 VGND 0.1131f
C10607 XThR.Tn[1].t53 VGND 0.01884f
C10608 XThR.Tn[1].t15 VGND 0.01984f
C10609 XThR.Tn[1].n42 VGND 0.04928f
C10610 XThR.Tn[1].t48 VGND 0.01884f
C10611 XThR.Tn[1].t13 VGND 0.01984f
C10612 XThR.Tn[1].n43 VGND 0.04927f
C10613 XThR.Tn[1].n44 VGND 0.03788f
C10614 XThR.Tn[1].n45 VGND 0.00722f
C10615 XThR.Tn[1].n46 VGND 0.1131f
C10616 XThR.Tn[1].t72 VGND 0.01884f
C10617 XThR.Tn[1].t33 VGND 0.01984f
C10618 XThR.Tn[1].n47 VGND 0.04928f
C10619 XThR.Tn[1].t67 VGND 0.01884f
C10620 XThR.Tn[1].t28 VGND 0.01984f
C10621 XThR.Tn[1].n48 VGND 0.04927f
C10622 XThR.Tn[1].n49 VGND 0.03788f
C10623 XThR.Tn[1].n50 VGND 0.00722f
C10624 XThR.Tn[1].n51 VGND 0.1131f
C10625 XThR.Tn[1].t26 VGND 0.01884f
C10626 XThR.Tn[1].t52 VGND 0.01984f
C10627 XThR.Tn[1].n52 VGND 0.04928f
C10628 XThR.Tn[1].t21 VGND 0.01884f
C10629 XThR.Tn[1].t47 VGND 0.01984f
C10630 XThR.Tn[1].n53 VGND 0.04927f
C10631 XThR.Tn[1].n54 VGND 0.03788f
C10632 XThR.Tn[1].n55 VGND 0.00722f
C10633 XThR.Tn[1].n56 VGND 0.1131f
C10634 XThR.Tn[1].t61 VGND 0.01884f
C10635 XThR.Tn[1].t71 VGND 0.01984f
C10636 XThR.Tn[1].n57 VGND 0.04928f
C10637 XThR.Tn[1].t59 VGND 0.01884f
C10638 XThR.Tn[1].t66 VGND 0.01984f
C10639 XThR.Tn[1].n58 VGND 0.04927f
C10640 XThR.Tn[1].n59 VGND 0.03788f
C10641 XThR.Tn[1].n60 VGND 0.00722f
C10642 XThR.Tn[1].n61 VGND 0.1131f
C10643 XThR.Tn[1].t37 VGND 0.01884f
C10644 XThR.Tn[1].t44 VGND 0.01984f
C10645 XThR.Tn[1].n62 VGND 0.04928f
C10646 XThR.Tn[1].t32 VGND 0.01884f
C10647 XThR.Tn[1].t42 VGND 0.01984f
C10648 XThR.Tn[1].n63 VGND 0.04927f
C10649 XThR.Tn[1].n64 VGND 0.03788f
C10650 XThR.Tn[1].n65 VGND 0.00722f
C10651 XThR.Tn[1].n66 VGND 0.1131f
C10652 XThR.Tn[1].t55 VGND 0.01884f
C10653 XThR.Tn[1].t16 VGND 0.01984f
C10654 XThR.Tn[1].n67 VGND 0.04928f
C10655 XThR.Tn[1].t51 VGND 0.01884f
C10656 XThR.Tn[1].t14 VGND 0.01984f
C10657 XThR.Tn[1].n68 VGND 0.04927f
C10658 XThR.Tn[1].n69 VGND 0.03788f
C10659 XThR.Tn[1].n70 VGND 0.00722f
C10660 XThR.Tn[1].n71 VGND 0.1131f
C10661 XThR.Tn[1].t25 VGND 0.01884f
C10662 XThR.Tn[1].t36 VGND 0.01984f
C10663 XThR.Tn[1].n72 VGND 0.04928f
C10664 XThR.Tn[1].t20 VGND 0.01884f
C10665 XThR.Tn[1].t31 VGND 0.01984f
C10666 XThR.Tn[1].n73 VGND 0.04927f
C10667 XThR.Tn[1].n74 VGND 0.03788f
C10668 XThR.Tn[1].n75 VGND 0.00722f
C10669 XThR.Tn[1].n76 VGND 0.1131f
C10670 XThR.Tn[1].t41 VGND 0.01884f
C10671 XThR.Tn[1].t54 VGND 0.01984f
C10672 XThR.Tn[1].n77 VGND 0.04928f
C10673 XThR.Tn[1].t39 VGND 0.01884f
C10674 XThR.Tn[1].t49 VGND 0.01984f
C10675 XThR.Tn[1].n78 VGND 0.04927f
C10676 XThR.Tn[1].n79 VGND 0.03788f
C10677 XThR.Tn[1].n80 VGND 0.00722f
C10678 XThR.Tn[1].n81 VGND 0.1131f
C10679 XThR.Tn[1].t63 VGND 0.01884f
C10680 XThR.Tn[1].t45 VGND 0.01984f
C10681 XThR.Tn[1].n82 VGND 0.04928f
C10682 XThR.Tn[1].t60 VGND 0.01884f
C10683 XThR.Tn[1].t43 VGND 0.01984f
C10684 XThR.Tn[1].n83 VGND 0.04927f
C10685 XThR.Tn[1].n84 VGND 0.03788f
C10686 XThR.Tn[1].n85 VGND 0.00722f
C10687 XThR.Tn[1].n86 VGND 0.1131f
C10688 XThR.Tn[1].n87 VGND 0.1033f
C10689 XThR.Tn[1].n88 VGND 0.29735f
C10690 XThR.Tn[1].n89 VGND 0.04852f
C10691 XThC.Tn[14].t4 VGND 0.01243f
C10692 XThC.Tn[14].t6 VGND 0.01243f
C10693 XThC.Tn[14].n0 VGND 0.03099f
C10694 XThC.Tn[14].t5 VGND 0.01243f
C10695 XThC.Tn[14].t7 VGND 0.01243f
C10696 XThC.Tn[14].n1 VGND 0.02485f
C10697 XThC.Tn[14].n2 VGND 0.06252f
C10698 XThC.Tn[14].t23 VGND 0.01553f
C10699 XThC.Tn[14].t26 VGND 0.01636f
C10700 XThC.Tn[14].n3 VGND 0.04063f
C10701 XThC.Tn[14].n4 VGND 0.02531f
C10702 XThC.Tn[14].n5 VGND 0.08201f
C10703 XThC.Tn[14].t32 VGND 0.01553f
C10704 XThC.Tn[14].t34 VGND 0.01636f
C10705 XThC.Tn[14].n6 VGND 0.04063f
C10706 XThC.Tn[14].n7 VGND 0.02531f
C10707 XThC.Tn[14].n8 VGND 0.08223f
C10708 XThC.Tn[14].n9 VGND 0.1373f
C10709 XThC.Tn[14].t13 VGND 0.01553f
C10710 XThC.Tn[14].t16 VGND 0.01636f
C10711 XThC.Tn[14].n10 VGND 0.04063f
C10712 XThC.Tn[14].n11 VGND 0.02531f
C10713 XThC.Tn[14].n12 VGND 0.08223f
C10714 XThC.Tn[14].n13 VGND 0.1373f
C10715 XThC.Tn[14].t14 VGND 0.01553f
C10716 XThC.Tn[14].t18 VGND 0.01636f
C10717 XThC.Tn[14].n14 VGND 0.04063f
C10718 XThC.Tn[14].n15 VGND 0.02531f
C10719 XThC.Tn[14].n16 VGND 0.08223f
C10720 XThC.Tn[14].n17 VGND 0.1373f
C10721 XThC.Tn[14].t24 VGND 0.01553f
C10722 XThC.Tn[14].t27 VGND 0.01636f
C10723 XThC.Tn[14].n18 VGND 0.04063f
C10724 XThC.Tn[14].n19 VGND 0.02531f
C10725 XThC.Tn[14].n20 VGND 0.08223f
C10726 XThC.Tn[14].n21 VGND 0.1373f
C10727 XThC.Tn[14].t35 VGND 0.01553f
C10728 XThC.Tn[14].t38 VGND 0.01636f
C10729 XThC.Tn[14].n22 VGND 0.04063f
C10730 XThC.Tn[14].n23 VGND 0.02531f
C10731 XThC.Tn[14].n24 VGND 0.08223f
C10732 XThC.Tn[14].n25 VGND 0.1373f
C10733 XThC.Tn[14].t15 VGND 0.01553f
C10734 XThC.Tn[14].t19 VGND 0.01636f
C10735 XThC.Tn[14].n26 VGND 0.04063f
C10736 XThC.Tn[14].n27 VGND 0.02531f
C10737 XThC.Tn[14].n28 VGND 0.08223f
C10738 XThC.Tn[14].n29 VGND 0.1373f
C10739 XThC.Tn[14].t25 VGND 0.01553f
C10740 XThC.Tn[14].t28 VGND 0.01636f
C10741 XThC.Tn[14].n30 VGND 0.04063f
C10742 XThC.Tn[14].n31 VGND 0.02531f
C10743 XThC.Tn[14].n32 VGND 0.08223f
C10744 XThC.Tn[14].n33 VGND 0.1373f
C10745 XThC.Tn[14].t29 VGND 0.01553f
C10746 XThC.Tn[14].t31 VGND 0.01636f
C10747 XThC.Tn[14].n34 VGND 0.04063f
C10748 XThC.Tn[14].n35 VGND 0.02531f
C10749 XThC.Tn[14].n36 VGND 0.08223f
C10750 XThC.Tn[14].n37 VGND 0.1373f
C10751 XThC.Tn[14].t36 VGND 0.01553f
C10752 XThC.Tn[14].t39 VGND 0.01636f
C10753 XThC.Tn[14].n38 VGND 0.04063f
C10754 XThC.Tn[14].n39 VGND 0.02531f
C10755 XThC.Tn[14].n40 VGND 0.08223f
C10756 XThC.Tn[14].n41 VGND 0.1373f
C10757 XThC.Tn[14].t17 VGND 0.01553f
C10758 XThC.Tn[14].t20 VGND 0.01636f
C10759 XThC.Tn[14].n42 VGND 0.04063f
C10760 XThC.Tn[14].n43 VGND 0.02531f
C10761 XThC.Tn[14].n44 VGND 0.08223f
C10762 XThC.Tn[14].n45 VGND 0.1373f
C10763 XThC.Tn[14].t21 VGND 0.01553f
C10764 XThC.Tn[14].t22 VGND 0.01636f
C10765 XThC.Tn[14].n46 VGND 0.04063f
C10766 XThC.Tn[14].n47 VGND 0.02531f
C10767 XThC.Tn[14].n48 VGND 0.08223f
C10768 XThC.Tn[14].n49 VGND 0.1373f
C10769 XThC.Tn[14].t37 VGND 0.01553f
C10770 XThC.Tn[14].t40 VGND 0.01636f
C10771 XThC.Tn[14].n50 VGND 0.04063f
C10772 XThC.Tn[14].n51 VGND 0.02531f
C10773 XThC.Tn[14].n52 VGND 0.08223f
C10774 XThC.Tn[14].n53 VGND 0.1373f
C10775 XThC.Tn[14].t41 VGND 0.01553f
C10776 XThC.Tn[14].t43 VGND 0.01636f
C10777 XThC.Tn[14].n54 VGND 0.04063f
C10778 XThC.Tn[14].n55 VGND 0.02531f
C10779 XThC.Tn[14].n56 VGND 0.08223f
C10780 XThC.Tn[14].n57 VGND 0.1373f
C10781 XThC.Tn[14].t42 VGND 0.01553f
C10782 XThC.Tn[14].t12 VGND 0.01636f
C10783 XThC.Tn[14].n58 VGND 0.04063f
C10784 XThC.Tn[14].n59 VGND 0.02531f
C10785 XThC.Tn[14].n60 VGND 0.08223f
C10786 XThC.Tn[14].n61 VGND 0.1373f
C10787 XThC.Tn[14].t30 VGND 0.01553f
C10788 XThC.Tn[14].t33 VGND 0.01636f
C10789 XThC.Tn[14].n62 VGND 0.04063f
C10790 XThC.Tn[14].n63 VGND 0.02531f
C10791 XThC.Tn[14].n64 VGND 0.08223f
C10792 XThC.Tn[14].n65 VGND 0.1373f
C10793 XThC.Tn[14].n66 VGND 0.90052f
C10794 XThC.Tn[14].n67 VGND 0.26491f
C10795 XThC.Tn[14].t0 VGND 0.01912f
C10796 XThC.Tn[14].t1 VGND 0.01912f
C10797 XThC.Tn[14].n68 VGND 0.0413f
C10798 XThC.Tn[14].t3 VGND 0.01912f
C10799 XThC.Tn[14].t2 VGND 0.01912f
C10800 XThC.Tn[14].n69 VGND 0.06286f
C10801 XThC.Tn[14].n70 VGND 0.17467f
C10802 XThC.Tn[14].n71 VGND 0.02746f
C10803 XThC.Tn[14].t11 VGND 0.01912f
C10804 XThC.Tn[14].t10 VGND 0.01912f
C10805 XThC.Tn[14].n72 VGND 0.05804f
C10806 XThC.Tn[14].t9 VGND 0.01912f
C10807 XThC.Tn[14].t8 VGND 0.01912f
C10808 XThC.Tn[14].n73 VGND 0.04249f
C10809 XThC.Tn[14].n74 VGND 0.18913f
C10810 XThR.Tn[13].t2 VGND 0.02411f
C10811 XThR.Tn[13].t0 VGND 0.02411f
C10812 XThR.Tn[13].n0 VGND 0.05359f
C10813 XThR.Tn[13].t1 VGND 0.02411f
C10814 XThR.Tn[13].t3 VGND 0.02411f
C10815 XThR.Tn[13].n1 VGND 0.0732f
C10816 XThR.Tn[13].n2 VGND 0.24367f
C10817 XThR.Tn[13].t11 VGND 0.01567f
C10818 XThR.Tn[13].t9 VGND 0.01567f
C10819 XThR.Tn[13].n3 VGND 0.03908f
C10820 XThR.Tn[13].t10 VGND 0.01567f
C10821 XThR.Tn[13].t8 VGND 0.01567f
C10822 XThR.Tn[13].n4 VGND 0.03134f
C10823 XThR.Tn[13].n5 VGND 0.07884f
C10824 XThR.Tn[13].t39 VGND 0.01959f
C10825 XThR.Tn[13].t65 VGND 0.02063f
C10826 XThR.Tn[13].n6 VGND 0.05124f
C10827 XThR.Tn[13].n7 VGND 0.09525f
C10828 XThR.Tn[13].t13 VGND 0.01959f
C10829 XThR.Tn[13].t21 VGND 0.02063f
C10830 XThR.Tn[13].n8 VGND 0.05124f
C10831 XThR.Tn[13].t51 VGND 0.01959f
C10832 XThR.Tn[13].t57 VGND 0.02063f
C10833 XThR.Tn[13].n9 VGND 0.05122f
C10834 XThR.Tn[13].n10 VGND 0.03939f
C10835 XThR.Tn[13].n11 VGND 0.00751f
C10836 XThR.Tn[13].n12 VGND 0.11758f
C10837 XThR.Tn[13].t29 VGND 0.01959f
C10838 XThR.Tn[13].t58 VGND 0.02063f
C10839 XThR.Tn[13].n13 VGND 0.05124f
C10840 XThR.Tn[13].t67 VGND 0.01959f
C10841 XThR.Tn[13].t33 VGND 0.02063f
C10842 XThR.Tn[13].n14 VGND 0.05122f
C10843 XThR.Tn[13].n15 VGND 0.03939f
C10844 XThR.Tn[13].n16 VGND 0.00751f
C10845 XThR.Tn[13].n17 VGND 0.11758f
C10846 XThR.Tn[13].t66 VGND 0.01959f
C10847 XThR.Tn[13].t12 VGND 0.02063f
C10848 XThR.Tn[13].n18 VGND 0.05124f
C10849 XThR.Tn[13].t40 VGND 0.01959f
C10850 XThR.Tn[13].t50 VGND 0.02063f
C10851 XThR.Tn[13].n19 VGND 0.05122f
C10852 XThR.Tn[13].n20 VGND 0.03939f
C10853 XThR.Tn[13].n21 VGND 0.00751f
C10854 XThR.Tn[13].n22 VGND 0.11758f
C10855 XThR.Tn[13].t31 VGND 0.01959f
C10856 XThR.Tn[13].t43 VGND 0.02063f
C10857 XThR.Tn[13].n23 VGND 0.05124f
C10858 XThR.Tn[13].t69 VGND 0.01959f
C10859 XThR.Tn[13].t19 VGND 0.02063f
C10860 XThR.Tn[13].n24 VGND 0.05122f
C10861 XThR.Tn[13].n25 VGND 0.03939f
C10862 XThR.Tn[13].n26 VGND 0.00751f
C10863 XThR.Tn[13].n27 VGND 0.11758f
C10864 XThR.Tn[13].t48 VGND 0.01959f
C10865 XThR.Tn[13].t14 VGND 0.02063f
C10866 XThR.Tn[13].n28 VGND 0.05124f
C10867 XThR.Tn[13].t24 VGND 0.01959f
C10868 XThR.Tn[13].t52 VGND 0.02063f
C10869 XThR.Tn[13].n29 VGND 0.05122f
C10870 XThR.Tn[13].n30 VGND 0.03939f
C10871 XThR.Tn[13].n31 VGND 0.00751f
C10872 XThR.Tn[13].n32 VGND 0.11758f
C10873 XThR.Tn[13].t42 VGND 0.01959f
C10874 XThR.Tn[13].t30 VGND 0.02063f
C10875 XThR.Tn[13].n33 VGND 0.05124f
C10876 XThR.Tn[13].t18 VGND 0.01959f
C10877 XThR.Tn[13].t68 VGND 0.02063f
C10878 XThR.Tn[13].n34 VGND 0.05122f
C10879 XThR.Tn[13].n35 VGND 0.03939f
C10880 XThR.Tn[13].n36 VGND 0.00751f
C10881 XThR.Tn[13].n37 VGND 0.11758f
C10882 XThR.Tn[13].t60 VGND 0.01959f
C10883 XThR.Tn[13].t23 VGND 0.02063f
C10884 XThR.Tn[13].n38 VGND 0.05124f
C10885 XThR.Tn[13].t36 VGND 0.01959f
C10886 XThR.Tn[13].t63 VGND 0.02063f
C10887 XThR.Tn[13].n39 VGND 0.05122f
C10888 XThR.Tn[13].n40 VGND 0.03939f
C10889 XThR.Tn[13].n41 VGND 0.00751f
C10890 XThR.Tn[13].n42 VGND 0.11758f
C10891 XThR.Tn[13].t16 VGND 0.01959f
C10892 XThR.Tn[13].t41 VGND 0.02063f
C10893 XThR.Tn[13].n43 VGND 0.05124f
C10894 XThR.Tn[13].t54 VGND 0.01959f
C10895 XThR.Tn[13].t17 VGND 0.02063f
C10896 XThR.Tn[13].n44 VGND 0.05122f
C10897 XThR.Tn[13].n45 VGND 0.03939f
C10898 XThR.Tn[13].n46 VGND 0.00751f
C10899 XThR.Tn[13].n47 VGND 0.11758f
C10900 XThR.Tn[13].t34 VGND 0.01959f
C10901 XThR.Tn[13].t59 VGND 0.02063f
C10902 XThR.Tn[13].n48 VGND 0.05124f
C10903 XThR.Tn[13].t71 VGND 0.01959f
C10904 XThR.Tn[13].t35 VGND 0.02063f
C10905 XThR.Tn[13].n49 VGND 0.05122f
C10906 XThR.Tn[13].n50 VGND 0.03939f
C10907 XThR.Tn[13].n51 VGND 0.00751f
C10908 XThR.Tn[13].n52 VGND 0.11758f
C10909 XThR.Tn[13].t72 VGND 0.01959f
C10910 XThR.Tn[13].t15 VGND 0.02063f
C10911 XThR.Tn[13].n53 VGND 0.05124f
C10912 XThR.Tn[13].t46 VGND 0.01959f
C10913 XThR.Tn[13].t53 VGND 0.02063f
C10914 XThR.Tn[13].n54 VGND 0.05122f
C10915 XThR.Tn[13].n55 VGND 0.03939f
C10916 XThR.Tn[13].n56 VGND 0.00751f
C10917 XThR.Tn[13].n57 VGND 0.11758f
C10918 XThR.Tn[13].t45 VGND 0.01959f
C10919 XThR.Tn[13].t55 VGND 0.02063f
C10920 XThR.Tn[13].n58 VGND 0.05124f
C10921 XThR.Tn[13].t22 VGND 0.01959f
C10922 XThR.Tn[13].t27 VGND 0.02063f
C10923 XThR.Tn[13].n59 VGND 0.05122f
C10924 XThR.Tn[13].n60 VGND 0.03939f
C10925 XThR.Tn[13].n61 VGND 0.00751f
C10926 XThR.Tn[13].n62 VGND 0.11758f
C10927 XThR.Tn[13].t62 VGND 0.01959f
C10928 XThR.Tn[13].t25 VGND 0.02063f
C10929 XThR.Tn[13].n63 VGND 0.05124f
C10930 XThR.Tn[13].t38 VGND 0.01959f
C10931 XThR.Tn[13].t64 VGND 0.02063f
C10932 XThR.Tn[13].n64 VGND 0.05122f
C10933 XThR.Tn[13].n65 VGND 0.03939f
C10934 XThR.Tn[13].n66 VGND 0.00751f
C10935 XThR.Tn[13].n67 VGND 0.11758f
C10936 XThR.Tn[13].t32 VGND 0.01959f
C10937 XThR.Tn[13].t44 VGND 0.02063f
C10938 XThR.Tn[13].n68 VGND 0.05124f
C10939 XThR.Tn[13].t70 VGND 0.01959f
C10940 XThR.Tn[13].t20 VGND 0.02063f
C10941 XThR.Tn[13].n69 VGND 0.05122f
C10942 XThR.Tn[13].n70 VGND 0.03939f
C10943 XThR.Tn[13].n71 VGND 0.00751f
C10944 XThR.Tn[13].n72 VGND 0.11758f
C10945 XThR.Tn[13].t49 VGND 0.01959f
C10946 XThR.Tn[13].t61 VGND 0.02063f
C10947 XThR.Tn[13].n73 VGND 0.05124f
C10948 XThR.Tn[13].t26 VGND 0.01959f
C10949 XThR.Tn[13].t37 VGND 0.02063f
C10950 XThR.Tn[13].n74 VGND 0.05122f
C10951 XThR.Tn[13].n75 VGND 0.03939f
C10952 XThR.Tn[13].n76 VGND 0.00751f
C10953 XThR.Tn[13].n77 VGND 0.11758f
C10954 XThR.Tn[13].t73 VGND 0.01959f
C10955 XThR.Tn[13].t56 VGND 0.02063f
C10956 XThR.Tn[13].n78 VGND 0.05124f
C10957 XThR.Tn[13].t47 VGND 0.01959f
C10958 XThR.Tn[13].t28 VGND 0.02063f
C10959 XThR.Tn[13].n79 VGND 0.05122f
C10960 XThR.Tn[13].n80 VGND 0.03939f
C10961 XThR.Tn[13].n81 VGND 0.00751f
C10962 XThR.Tn[13].n82 VGND 0.11758f
C10963 XThR.Tn[13].n83 VGND 0.10739f
C10964 XThR.Tn[13].n84 VGND 0.42105f
C10965 XThR.Tn[13].t6 VGND 0.02411f
C10966 XThR.Tn[13].t4 VGND 0.02411f
C10967 XThR.Tn[13].n85 VGND 0.05209f
C10968 XThR.Tn[13].t7 VGND 0.02411f
C10969 XThR.Tn[13].t5 VGND 0.02411f
C10970 XThR.Tn[13].n86 VGND 0.07928f
C10971 XThR.Tn[13].n87 VGND 0.22013f
C10972 XThR.Tn[13].n88 VGND 0.02947f
C10973 XThR.Tn[11].t7 VGND 0.01576f
C10974 XThR.Tn[11].t1 VGND 0.01576f
C10975 XThR.Tn[11].n0 VGND 0.03931f
C10976 XThR.Tn[11].t0 VGND 0.01576f
C10977 XThR.Tn[11].t3 VGND 0.01576f
C10978 XThR.Tn[11].n1 VGND 0.03152f
C10979 XThR.Tn[11].n2 VGND 0.0793f
C10980 XThR.Tn[11].t8 VGND 0.02425f
C10981 XThR.Tn[11].t10 VGND 0.02425f
C10982 XThR.Tn[11].n3 VGND 0.07362f
C10983 XThR.Tn[11].t9 VGND 0.02425f
C10984 XThR.Tn[11].t11 VGND 0.02425f
C10985 XThR.Tn[11].n4 VGND 0.0539f
C10986 XThR.Tn[11].n5 VGND 0.24509f
C10987 XThR.Tn[11].t4 VGND 0.02425f
C10988 XThR.Tn[11].t6 VGND 0.02425f
C10989 XThR.Tn[11].n6 VGND 0.05239f
C10990 XThR.Tn[11].t2 VGND 0.02425f
C10991 XThR.Tn[11].t5 VGND 0.02425f
C10992 XThR.Tn[11].n7 VGND 0.07974f
C10993 XThR.Tn[11].n8 VGND 0.2214f
C10994 XThR.Tn[11].n9 VGND 0.02964f
C10995 XThR.Tn[11].t60 VGND 0.01971f
C10996 XThR.Tn[11].t25 VGND 0.02075f
C10997 XThR.Tn[11].n10 VGND 0.05153f
C10998 XThR.Tn[11].n11 VGND 0.09581f
C10999 XThR.Tn[11].t38 VGND 0.01971f
C11000 XThR.Tn[11].t43 VGND 0.02075f
C11001 XThR.Tn[11].n12 VGND 0.05153f
C11002 XThR.Tn[11].t30 VGND 0.01971f
C11003 XThR.Tn[11].t36 VGND 0.02075f
C11004 XThR.Tn[11].n13 VGND 0.05152f
C11005 XThR.Tn[11].n14 VGND 0.03961f
C11006 XThR.Tn[11].n15 VGND 0.00755f
C11007 XThR.Tn[11].n16 VGND 0.11826f
C11008 XThR.Tn[11].t52 VGND 0.01971f
C11009 XThR.Tn[11].t19 VGND 0.02075f
C11010 XThR.Tn[11].n17 VGND 0.05153f
C11011 XThR.Tn[11].t47 VGND 0.01971f
C11012 XThR.Tn[11].t12 VGND 0.02075f
C11013 XThR.Tn[11].n18 VGND 0.05152f
C11014 XThR.Tn[11].n19 VGND 0.03961f
C11015 XThR.Tn[11].n20 VGND 0.00755f
C11016 XThR.Tn[11].n21 VGND 0.11826f
C11017 XThR.Tn[11].t26 VGND 0.01971f
C11018 XThR.Tn[11].t37 VGND 0.02075f
C11019 XThR.Tn[11].n22 VGND 0.05153f
C11020 XThR.Tn[11].t20 VGND 0.01971f
C11021 XThR.Tn[11].t29 VGND 0.02075f
C11022 XThR.Tn[11].n23 VGND 0.05152f
C11023 XThR.Tn[11].n24 VGND 0.03961f
C11024 XThR.Tn[11].n25 VGND 0.00755f
C11025 XThR.Tn[11].n26 VGND 0.11826f
C11026 XThR.Tn[11].t54 VGND 0.01971f
C11027 XThR.Tn[11].t65 VGND 0.02075f
C11028 XThR.Tn[11].n27 VGND 0.05153f
C11029 XThR.Tn[11].t49 VGND 0.01971f
C11030 XThR.Tn[11].t59 VGND 0.02075f
C11031 XThR.Tn[11].n28 VGND 0.05152f
C11032 XThR.Tn[11].n29 VGND 0.03961f
C11033 XThR.Tn[11].n30 VGND 0.00755f
C11034 XThR.Tn[11].n31 VGND 0.11826f
C11035 XThR.Tn[11].t72 VGND 0.01971f
C11036 XThR.Tn[11].t39 VGND 0.02075f
C11037 XThR.Tn[11].n32 VGND 0.05153f
C11038 XThR.Tn[11].t68 VGND 0.01971f
C11039 XThR.Tn[11].t31 VGND 0.02075f
C11040 XThR.Tn[11].n33 VGND 0.05152f
C11041 XThR.Tn[11].n34 VGND 0.03961f
C11042 XThR.Tn[11].n35 VGND 0.00755f
C11043 XThR.Tn[11].n36 VGND 0.11826f
C11044 XThR.Tn[11].t64 VGND 0.01971f
C11045 XThR.Tn[11].t53 VGND 0.02075f
C11046 XThR.Tn[11].n37 VGND 0.05153f
C11047 XThR.Tn[11].t58 VGND 0.01971f
C11048 XThR.Tn[11].t48 VGND 0.02075f
C11049 XThR.Tn[11].n38 VGND 0.05152f
C11050 XThR.Tn[11].n39 VGND 0.03961f
C11051 XThR.Tn[11].n40 VGND 0.00755f
C11052 XThR.Tn[11].n41 VGND 0.11826f
C11053 XThR.Tn[11].t22 VGND 0.01971f
C11054 XThR.Tn[11].t45 VGND 0.02075f
C11055 XThR.Tn[11].n42 VGND 0.05153f
C11056 XThR.Tn[11].t15 VGND 0.01971f
C11057 XThR.Tn[11].t42 VGND 0.02075f
C11058 XThR.Tn[11].n43 VGND 0.05152f
C11059 XThR.Tn[11].n44 VGND 0.03961f
C11060 XThR.Tn[11].n45 VGND 0.00755f
C11061 XThR.Tn[11].n46 VGND 0.11826f
C11062 XThR.Tn[11].t41 VGND 0.01971f
C11063 XThR.Tn[11].t63 VGND 0.02075f
C11064 XThR.Tn[11].n47 VGND 0.05153f
C11065 XThR.Tn[11].t33 VGND 0.01971f
C11066 XThR.Tn[11].t57 VGND 0.02075f
C11067 XThR.Tn[11].n48 VGND 0.05152f
C11068 XThR.Tn[11].n49 VGND 0.03961f
C11069 XThR.Tn[11].n50 VGND 0.00755f
C11070 XThR.Tn[11].n51 VGND 0.11826f
C11071 XThR.Tn[11].t56 VGND 0.01971f
C11072 XThR.Tn[11].t21 VGND 0.02075f
C11073 XThR.Tn[11].n52 VGND 0.05153f
C11074 XThR.Tn[11].t51 VGND 0.01971f
C11075 XThR.Tn[11].t13 VGND 0.02075f
C11076 XThR.Tn[11].n53 VGND 0.05152f
C11077 XThR.Tn[11].n54 VGND 0.03961f
C11078 XThR.Tn[11].n55 VGND 0.00755f
C11079 XThR.Tn[11].n56 VGND 0.11826f
C11080 XThR.Tn[11].t34 VGND 0.01971f
C11081 XThR.Tn[11].t40 VGND 0.02075f
C11082 XThR.Tn[11].n57 VGND 0.05153f
C11083 XThR.Tn[11].t27 VGND 0.01971f
C11084 XThR.Tn[11].t32 VGND 0.02075f
C11085 XThR.Tn[11].n58 VGND 0.05152f
C11086 XThR.Tn[11].n59 VGND 0.03961f
C11087 XThR.Tn[11].n60 VGND 0.00755f
C11088 XThR.Tn[11].n61 VGND 0.11826f
C11089 XThR.Tn[11].t67 VGND 0.01971f
C11090 XThR.Tn[11].t14 VGND 0.02075f
C11091 XThR.Tn[11].n62 VGND 0.05153f
C11092 XThR.Tn[11].t62 VGND 0.01971f
C11093 XThR.Tn[11].t70 VGND 0.02075f
C11094 XThR.Tn[11].n63 VGND 0.05152f
C11095 XThR.Tn[11].n64 VGND 0.03961f
C11096 XThR.Tn[11].n65 VGND 0.00755f
C11097 XThR.Tn[11].n66 VGND 0.11826f
C11098 XThR.Tn[11].t24 VGND 0.01971f
C11099 XThR.Tn[11].t46 VGND 0.02075f
C11100 XThR.Tn[11].n67 VGND 0.05153f
C11101 XThR.Tn[11].t18 VGND 0.01971f
C11102 XThR.Tn[11].t44 VGND 0.02075f
C11103 XThR.Tn[11].n68 VGND 0.05152f
C11104 XThR.Tn[11].n69 VGND 0.03961f
C11105 XThR.Tn[11].n70 VGND 0.00755f
C11106 XThR.Tn[11].n71 VGND 0.11826f
C11107 XThR.Tn[11].t55 VGND 0.01971f
C11108 XThR.Tn[11].t66 VGND 0.02075f
C11109 XThR.Tn[11].n72 VGND 0.05153f
C11110 XThR.Tn[11].t50 VGND 0.01971f
C11111 XThR.Tn[11].t61 VGND 0.02075f
C11112 XThR.Tn[11].n73 VGND 0.05152f
C11113 XThR.Tn[11].n74 VGND 0.03961f
C11114 XThR.Tn[11].n75 VGND 0.00755f
C11115 XThR.Tn[11].n76 VGND 0.11826f
C11116 XThR.Tn[11].t73 VGND 0.01971f
C11117 XThR.Tn[11].t23 VGND 0.02075f
C11118 XThR.Tn[11].n77 VGND 0.05153f
C11119 XThR.Tn[11].t69 VGND 0.01971f
C11120 XThR.Tn[11].t16 VGND 0.02075f
C11121 XThR.Tn[11].n78 VGND 0.05152f
C11122 XThR.Tn[11].n79 VGND 0.03961f
C11123 XThR.Tn[11].n80 VGND 0.00755f
C11124 XThR.Tn[11].n81 VGND 0.11826f
C11125 XThR.Tn[11].t35 VGND 0.01971f
C11126 XThR.Tn[11].t17 VGND 0.02075f
C11127 XThR.Tn[11].n82 VGND 0.05153f
C11128 XThR.Tn[11].t28 VGND 0.01971f
C11129 XThR.Tn[11].t71 VGND 0.02075f
C11130 XThR.Tn[11].n83 VGND 0.05152f
C11131 XThR.Tn[11].n84 VGND 0.03961f
C11132 XThR.Tn[11].n85 VGND 0.00755f
C11133 XThR.Tn[11].n86 VGND 0.11826f
C11134 XThR.Tn[11].n87 VGND 0.10802f
C11135 XThR.Tn[11].n88 VGND 0.38713f
C11136 XThR.Tn[6].t7 VGND 0.0235f
C11137 XThR.Tn[6].t4 VGND 0.0235f
C11138 XThR.Tn[6].n0 VGND 0.04743f
C11139 XThR.Tn[6].t6 VGND 0.0235f
C11140 XThR.Tn[6].t5 VGND 0.0235f
C11141 XThR.Tn[6].n1 VGND 0.0555f
C11142 XThR.Tn[6].n2 VGND 0.16647f
C11143 XThR.Tn[6].t8 VGND 0.01527f
C11144 XThR.Tn[6].t9 VGND 0.01527f
C11145 XThR.Tn[6].n3 VGND 0.03478f
C11146 XThR.Tn[6].t11 VGND 0.01527f
C11147 XThR.Tn[6].t10 VGND 0.01527f
C11148 XThR.Tn[6].n4 VGND 0.03478f
C11149 XThR.Tn[6].t0 VGND 0.01527f
C11150 XThR.Tn[6].t1 VGND 0.01527f
C11151 XThR.Tn[6].n5 VGND 0.05796f
C11152 XThR.Tn[6].t3 VGND 0.01527f
C11153 XThR.Tn[6].t2 VGND 0.01527f
C11154 XThR.Tn[6].n6 VGND 0.03478f
C11155 XThR.Tn[6].n7 VGND 0.16564f
C11156 XThR.Tn[6].n8 VGND 0.1024f
C11157 XThR.Tn[6].n9 VGND 0.11556f
C11158 XThR.Tn[6].t20 VGND 0.0191f
C11159 XThR.Tn[6].t50 VGND 0.02011f
C11160 XThR.Tn[6].n10 VGND 0.04994f
C11161 XThR.Tn[6].n11 VGND 0.09285f
C11162 XThR.Tn[6].t59 VGND 0.0191f
C11163 XThR.Tn[6].t66 VGND 0.02011f
C11164 XThR.Tn[6].n12 VGND 0.04994f
C11165 XThR.Tn[6].t41 VGND 0.0191f
C11166 XThR.Tn[6].t49 VGND 0.02011f
C11167 XThR.Tn[6].n13 VGND 0.04993f
C11168 XThR.Tn[6].n14 VGND 0.03839f
C11169 XThR.Tn[6].n15 VGND 0.00732f
C11170 XThR.Tn[6].n16 VGND 0.11461f
C11171 XThR.Tn[6].t12 VGND 0.0191f
C11172 XThR.Tn[6].t40 VGND 0.02011f
C11173 XThR.Tn[6].n17 VGND 0.04994f
C11174 XThR.Tn[6].t57 VGND 0.0191f
C11175 XThR.Tn[6].t22 VGND 0.02011f
C11176 XThR.Tn[6].n18 VGND 0.04993f
C11177 XThR.Tn[6].n19 VGND 0.03839f
C11178 XThR.Tn[6].n20 VGND 0.00732f
C11179 XThR.Tn[6].n21 VGND 0.11461f
C11180 XThR.Tn[6].t51 VGND 0.0191f
C11181 XThR.Tn[6].t56 VGND 0.02011f
C11182 XThR.Tn[6].n22 VGND 0.04994f
C11183 XThR.Tn[6].t32 VGND 0.0191f
C11184 XThR.Tn[6].t39 VGND 0.02011f
C11185 XThR.Tn[6].n23 VGND 0.04993f
C11186 XThR.Tn[6].n24 VGND 0.03839f
C11187 XThR.Tn[6].n25 VGND 0.00732f
C11188 XThR.Tn[6].n26 VGND 0.11461f
C11189 XThR.Tn[6].t15 VGND 0.0191f
C11190 XThR.Tn[6].t27 VGND 0.02011f
C11191 XThR.Tn[6].n27 VGND 0.04994f
C11192 XThR.Tn[6].t61 VGND 0.0191f
C11193 XThR.Tn[6].t70 VGND 0.02011f
C11194 XThR.Tn[6].n28 VGND 0.04993f
C11195 XThR.Tn[6].n29 VGND 0.03839f
C11196 XThR.Tn[6].n30 VGND 0.00732f
C11197 XThR.Tn[6].n31 VGND 0.11461f
C11198 XThR.Tn[6].t33 VGND 0.0191f
C11199 XThR.Tn[6].t60 VGND 0.02011f
C11200 XThR.Tn[6].n32 VGND 0.04994f
C11201 XThR.Tn[6].t14 VGND 0.0191f
C11202 XThR.Tn[6].t42 VGND 0.02011f
C11203 XThR.Tn[6].n33 VGND 0.04993f
C11204 XThR.Tn[6].n34 VGND 0.03839f
C11205 XThR.Tn[6].n35 VGND 0.00732f
C11206 XThR.Tn[6].n36 VGND 0.11461f
C11207 XThR.Tn[6].t26 VGND 0.0191f
C11208 XThR.Tn[6].t13 VGND 0.02011f
C11209 XThR.Tn[6].n37 VGND 0.04994f
C11210 XThR.Tn[6].t69 VGND 0.0191f
C11211 XThR.Tn[6].t58 VGND 0.02011f
C11212 XThR.Tn[6].n38 VGND 0.04993f
C11213 XThR.Tn[6].n39 VGND 0.03839f
C11214 XThR.Tn[6].n40 VGND 0.00732f
C11215 XThR.Tn[6].n41 VGND 0.11461f
C11216 XThR.Tn[6].t45 VGND 0.0191f
C11217 XThR.Tn[6].t68 VGND 0.02011f
C11218 XThR.Tn[6].n42 VGND 0.04994f
C11219 XThR.Tn[6].t25 VGND 0.0191f
C11220 XThR.Tn[6].t52 VGND 0.02011f
C11221 XThR.Tn[6].n43 VGND 0.04993f
C11222 XThR.Tn[6].n44 VGND 0.03839f
C11223 XThR.Tn[6].n45 VGND 0.00732f
C11224 XThR.Tn[6].n46 VGND 0.11461f
C11225 XThR.Tn[6].t65 VGND 0.0191f
C11226 XThR.Tn[6].t24 VGND 0.02011f
C11227 XThR.Tn[6].n47 VGND 0.04994f
C11228 XThR.Tn[6].t46 VGND 0.0191f
C11229 XThR.Tn[6].t67 VGND 0.02011f
C11230 XThR.Tn[6].n48 VGND 0.04993f
C11231 XThR.Tn[6].n49 VGND 0.03839f
C11232 XThR.Tn[6].n50 VGND 0.00732f
C11233 XThR.Tn[6].n51 VGND 0.11461f
C11234 XThR.Tn[6].t18 VGND 0.0191f
C11235 XThR.Tn[6].t43 VGND 0.02011f
C11236 XThR.Tn[6].n52 VGND 0.04994f
C11237 XThR.Tn[6].t64 VGND 0.0191f
C11238 XThR.Tn[6].t23 VGND 0.02011f
C11239 XThR.Tn[6].n53 VGND 0.04993f
C11240 XThR.Tn[6].n54 VGND 0.03839f
C11241 XThR.Tn[6].n55 VGND 0.00732f
C11242 XThR.Tn[6].n56 VGND 0.11461f
C11243 XThR.Tn[6].t54 VGND 0.0191f
C11244 XThR.Tn[6].t63 VGND 0.02011f
C11245 XThR.Tn[6].n57 VGND 0.04994f
C11246 XThR.Tn[6].t36 VGND 0.0191f
C11247 XThR.Tn[6].t44 VGND 0.02011f
C11248 XThR.Tn[6].n58 VGND 0.04993f
C11249 XThR.Tn[6].n59 VGND 0.03839f
C11250 XThR.Tn[6].n60 VGND 0.00732f
C11251 XThR.Tn[6].n61 VGND 0.11461f
C11252 XThR.Tn[6].t31 VGND 0.0191f
C11253 XThR.Tn[6].t35 VGND 0.02011f
C11254 XThR.Tn[6].n62 VGND 0.04994f
C11255 XThR.Tn[6].t73 VGND 0.0191f
C11256 XThR.Tn[6].t19 VGND 0.02011f
C11257 XThR.Tn[6].n63 VGND 0.04993f
C11258 XThR.Tn[6].n64 VGND 0.03839f
C11259 XThR.Tn[6].n65 VGND 0.00732f
C11260 XThR.Tn[6].n66 VGND 0.11461f
C11261 XThR.Tn[6].t48 VGND 0.0191f
C11262 XThR.Tn[6].t72 VGND 0.02011f
C11263 XThR.Tn[6].n67 VGND 0.04994f
C11264 XThR.Tn[6].t30 VGND 0.0191f
C11265 XThR.Tn[6].t53 VGND 0.02011f
C11266 XThR.Tn[6].n68 VGND 0.04993f
C11267 XThR.Tn[6].n69 VGND 0.03839f
C11268 XThR.Tn[6].n70 VGND 0.00732f
C11269 XThR.Tn[6].n71 VGND 0.11461f
C11270 XThR.Tn[6].t17 VGND 0.0191f
C11271 XThR.Tn[6].t29 VGND 0.02011f
C11272 XThR.Tn[6].n72 VGND 0.04994f
C11273 XThR.Tn[6].t62 VGND 0.0191f
C11274 XThR.Tn[6].t71 VGND 0.02011f
C11275 XThR.Tn[6].n73 VGND 0.04993f
C11276 XThR.Tn[6].n74 VGND 0.03839f
C11277 XThR.Tn[6].n75 VGND 0.00732f
C11278 XThR.Tn[6].n76 VGND 0.11461f
C11279 XThR.Tn[6].t34 VGND 0.0191f
C11280 XThR.Tn[6].t47 VGND 0.02011f
C11281 XThR.Tn[6].n77 VGND 0.04994f
C11282 XThR.Tn[6].t16 VGND 0.0191f
C11283 XThR.Tn[6].t28 VGND 0.02011f
C11284 XThR.Tn[6].n78 VGND 0.04993f
C11285 XThR.Tn[6].n79 VGND 0.03839f
C11286 XThR.Tn[6].n80 VGND 0.00732f
C11287 XThR.Tn[6].n81 VGND 0.11461f
C11288 XThR.Tn[6].t55 VGND 0.0191f
C11289 XThR.Tn[6].t37 VGND 0.02011f
C11290 XThR.Tn[6].n82 VGND 0.04994f
C11291 XThR.Tn[6].t38 VGND 0.0191f
C11292 XThR.Tn[6].t21 VGND 0.02011f
C11293 XThR.Tn[6].n83 VGND 0.04993f
C11294 XThR.Tn[6].n84 VGND 0.03839f
C11295 XThR.Tn[6].n85 VGND 0.00732f
C11296 XThR.Tn[6].n86 VGND 0.11461f
C11297 XThR.Tn[6].n87 VGND 0.10468f
C11298 XThR.Tn[6].n88 VGND 0.17425f
C11299 XThC.Tn[7].t6 VGND 0.01222f
C11300 XThC.Tn[7].t5 VGND 0.01222f
C11301 XThC.Tn[7].n0 VGND 0.03772f
C11302 XThC.Tn[7].t4 VGND 0.01222f
C11303 XThC.Tn[7].t7 VGND 0.01222f
C11304 XThC.Tn[7].n1 VGND 0.02699f
C11305 XThC.Tn[7].n2 VGND 0.13349f
C11306 XThC.Tn[7].t0 VGND 0.0188f
C11307 XThC.Tn[7].t3 VGND 0.0188f
C11308 XThC.Tn[7].n3 VGND 0.04049f
C11309 XThC.Tn[7].t2 VGND 0.0188f
C11310 XThC.Tn[7].t1 VGND 0.0188f
C11311 XThC.Tn[7].n4 VGND 0.06147f
C11312 XThC.Tn[7].n5 VGND 0.18074f
C11313 XThC.Tn[7].t19 VGND 0.01528f
C11314 XThC.Tn[7].t32 VGND 0.01609f
C11315 XThC.Tn[7].n6 VGND 0.03996f
C11316 XThC.Tn[7].n7 VGND 0.02489f
C11317 XThC.Tn[7].n8 VGND 0.08065f
C11318 XThC.Tn[7].t29 VGND 0.01528f
C11319 XThC.Tn[7].t10 VGND 0.01609f
C11320 XThC.Tn[7].n9 VGND 0.03996f
C11321 XThC.Tn[7].n10 VGND 0.02489f
C11322 XThC.Tn[7].n11 VGND 0.08087f
C11323 XThC.Tn[7].n12 VGND 0.13503f
C11324 XThC.Tn[7].t9 VGND 0.01528f
C11325 XThC.Tn[7].t23 VGND 0.01609f
C11326 XThC.Tn[7].n13 VGND 0.03996f
C11327 XThC.Tn[7].n14 VGND 0.02489f
C11328 XThC.Tn[7].n15 VGND 0.08087f
C11329 XThC.Tn[7].n16 VGND 0.13503f
C11330 XThC.Tn[7].t11 VGND 0.01528f
C11331 XThC.Tn[7].t24 VGND 0.01609f
C11332 XThC.Tn[7].n17 VGND 0.03996f
C11333 XThC.Tn[7].n18 VGND 0.02489f
C11334 XThC.Tn[7].n19 VGND 0.08087f
C11335 XThC.Tn[7].n20 VGND 0.13503f
C11336 XThC.Tn[7].t21 VGND 0.01528f
C11337 XThC.Tn[7].t35 VGND 0.01609f
C11338 XThC.Tn[7].n21 VGND 0.03996f
C11339 XThC.Tn[7].n22 VGND 0.02489f
C11340 XThC.Tn[7].n23 VGND 0.08087f
C11341 XThC.Tn[7].n24 VGND 0.13503f
C11342 XThC.Tn[7].t31 VGND 0.01528f
C11343 XThC.Tn[7].t14 VGND 0.01609f
C11344 XThC.Tn[7].n25 VGND 0.03996f
C11345 XThC.Tn[7].n26 VGND 0.02489f
C11346 XThC.Tn[7].n27 VGND 0.08087f
C11347 XThC.Tn[7].n28 VGND 0.13503f
C11348 XThC.Tn[7].t12 VGND 0.01528f
C11349 XThC.Tn[7].t25 VGND 0.01609f
C11350 XThC.Tn[7].n29 VGND 0.03996f
C11351 XThC.Tn[7].n30 VGND 0.02489f
C11352 XThC.Tn[7].n31 VGND 0.08087f
C11353 XThC.Tn[7].n32 VGND 0.13503f
C11354 XThC.Tn[7].t22 VGND 0.01528f
C11355 XThC.Tn[7].t36 VGND 0.01609f
C11356 XThC.Tn[7].n33 VGND 0.03996f
C11357 XThC.Tn[7].n34 VGND 0.02489f
C11358 XThC.Tn[7].n35 VGND 0.08087f
C11359 XThC.Tn[7].n36 VGND 0.13503f
C11360 XThC.Tn[7].t26 VGND 0.01528f
C11361 XThC.Tn[7].t38 VGND 0.01609f
C11362 XThC.Tn[7].n37 VGND 0.03996f
C11363 XThC.Tn[7].n38 VGND 0.02489f
C11364 XThC.Tn[7].n39 VGND 0.08087f
C11365 XThC.Tn[7].n40 VGND 0.13503f
C11366 XThC.Tn[7].t33 VGND 0.01528f
C11367 XThC.Tn[7].t15 VGND 0.01609f
C11368 XThC.Tn[7].n41 VGND 0.03996f
C11369 XThC.Tn[7].n42 VGND 0.02489f
C11370 XThC.Tn[7].n43 VGND 0.08087f
C11371 XThC.Tn[7].n44 VGND 0.13503f
C11372 XThC.Tn[7].t13 VGND 0.01528f
C11373 XThC.Tn[7].t27 VGND 0.01609f
C11374 XThC.Tn[7].n45 VGND 0.03996f
C11375 XThC.Tn[7].n46 VGND 0.02489f
C11376 XThC.Tn[7].n47 VGND 0.08087f
C11377 XThC.Tn[7].n48 VGND 0.13503f
C11378 XThC.Tn[7].t17 VGND 0.01528f
C11379 XThC.Tn[7].t30 VGND 0.01609f
C11380 XThC.Tn[7].n49 VGND 0.03996f
C11381 XThC.Tn[7].n50 VGND 0.02489f
C11382 XThC.Tn[7].n51 VGND 0.08087f
C11383 XThC.Tn[7].n52 VGND 0.13503f
C11384 XThC.Tn[7].t34 VGND 0.01528f
C11385 XThC.Tn[7].t16 VGND 0.01609f
C11386 XThC.Tn[7].n53 VGND 0.03996f
C11387 XThC.Tn[7].n54 VGND 0.02489f
C11388 XThC.Tn[7].n55 VGND 0.08087f
C11389 XThC.Tn[7].n56 VGND 0.13503f
C11390 XThC.Tn[7].t37 VGND 0.01528f
C11391 XThC.Tn[7].t18 VGND 0.01609f
C11392 XThC.Tn[7].n57 VGND 0.03996f
C11393 XThC.Tn[7].n58 VGND 0.02489f
C11394 XThC.Tn[7].n59 VGND 0.08087f
C11395 XThC.Tn[7].n60 VGND 0.13503f
C11396 XThC.Tn[7].t39 VGND 0.01528f
C11397 XThC.Tn[7].t20 VGND 0.01609f
C11398 XThC.Tn[7].n61 VGND 0.03996f
C11399 XThC.Tn[7].n62 VGND 0.02489f
C11400 XThC.Tn[7].n63 VGND 0.08087f
C11401 XThC.Tn[7].n64 VGND 0.13503f
C11402 XThC.Tn[7].t28 VGND 0.01528f
C11403 XThC.Tn[7].t8 VGND 0.01609f
C11404 XThC.Tn[7].n65 VGND 0.03996f
C11405 XThC.Tn[7].n66 VGND 0.02489f
C11406 XThC.Tn[7].n67 VGND 0.08087f
C11407 XThC.Tn[7].n68 VGND 0.13503f
C11408 XThC.Tn[7].n69 VGND 0.33911f
C11409 XThC.Tn[7].n70 VGND 0.02249f
C11410 XThC.Tn[13].t6 VGND 0.0194f
C11411 XThC.Tn[13].t5 VGND 0.0194f
C11412 XThC.Tn[13].n0 VGND 0.04192f
C11413 XThC.Tn[13].t4 VGND 0.0194f
C11414 XThC.Tn[13].t7 VGND 0.0194f
C11415 XThC.Tn[13].n1 VGND 0.06609f
C11416 XThC.Tn[13].n2 VGND 0.17502f
C11417 XThC.Tn[13].t9 VGND 0.0194f
C11418 XThC.Tn[13].t8 VGND 0.0194f
C11419 XThC.Tn[13].n3 VGND 0.05892f
C11420 XThC.Tn[13].t11 VGND 0.0194f
C11421 XThC.Tn[13].t10 VGND 0.0194f
C11422 XThC.Tn[13].n4 VGND 0.04313f
C11423 XThC.Tn[13].n5 VGND 0.19198f
C11424 XThC.Tn[13].n6 VGND 0.01289f
C11425 XThC.Tn[13].t32 VGND 0.01577f
C11426 XThC.Tn[13].t13 VGND 0.01661f
C11427 XThC.Tn[13].n7 VGND 0.04124f
C11428 XThC.Tn[13].n8 VGND 0.02569f
C11429 XThC.Tn[13].n9 VGND 0.08324f
C11430 XThC.Tn[13].t42 VGND 0.01577f
C11431 XThC.Tn[13].t23 VGND 0.01661f
C11432 XThC.Tn[13].n10 VGND 0.04124f
C11433 XThC.Tn[13].n11 VGND 0.02569f
C11434 XThC.Tn[13].n12 VGND 0.08347f
C11435 XThC.Tn[13].n13 VGND 0.13936f
C11436 XThC.Tn[13].t22 VGND 0.01577f
C11437 XThC.Tn[13].t36 VGND 0.01661f
C11438 XThC.Tn[13].n14 VGND 0.04124f
C11439 XThC.Tn[13].n15 VGND 0.02569f
C11440 XThC.Tn[13].n16 VGND 0.08347f
C11441 XThC.Tn[13].n17 VGND 0.13936f
C11442 XThC.Tn[13].t24 VGND 0.01577f
C11443 XThC.Tn[13].t37 VGND 0.01661f
C11444 XThC.Tn[13].n18 VGND 0.04124f
C11445 XThC.Tn[13].n19 VGND 0.02569f
C11446 XThC.Tn[13].n20 VGND 0.08347f
C11447 XThC.Tn[13].n21 VGND 0.13936f
C11448 XThC.Tn[13].t34 VGND 0.01577f
C11449 XThC.Tn[13].t16 VGND 0.01661f
C11450 XThC.Tn[13].n22 VGND 0.04124f
C11451 XThC.Tn[13].n23 VGND 0.02569f
C11452 XThC.Tn[13].n24 VGND 0.08347f
C11453 XThC.Tn[13].n25 VGND 0.13936f
C11454 XThC.Tn[13].t12 VGND 0.01577f
C11455 XThC.Tn[13].t27 VGND 0.01661f
C11456 XThC.Tn[13].n26 VGND 0.04124f
C11457 XThC.Tn[13].n27 VGND 0.02569f
C11458 XThC.Tn[13].n28 VGND 0.08347f
C11459 XThC.Tn[13].n29 VGND 0.13936f
C11460 XThC.Tn[13].t25 VGND 0.01577f
C11461 XThC.Tn[13].t38 VGND 0.01661f
C11462 XThC.Tn[13].n30 VGND 0.04124f
C11463 XThC.Tn[13].n31 VGND 0.02569f
C11464 XThC.Tn[13].n32 VGND 0.08347f
C11465 XThC.Tn[13].n33 VGND 0.13936f
C11466 XThC.Tn[13].t35 VGND 0.01577f
C11467 XThC.Tn[13].t17 VGND 0.01661f
C11468 XThC.Tn[13].n34 VGND 0.04124f
C11469 XThC.Tn[13].n35 VGND 0.02569f
C11470 XThC.Tn[13].n36 VGND 0.08347f
C11471 XThC.Tn[13].n37 VGND 0.13936f
C11472 XThC.Tn[13].t39 VGND 0.01577f
C11473 XThC.Tn[13].t19 VGND 0.01661f
C11474 XThC.Tn[13].n38 VGND 0.04124f
C11475 XThC.Tn[13].n39 VGND 0.02569f
C11476 XThC.Tn[13].n40 VGND 0.08347f
C11477 XThC.Tn[13].n41 VGND 0.13936f
C11478 XThC.Tn[13].t14 VGND 0.01577f
C11479 XThC.Tn[13].t28 VGND 0.01661f
C11480 XThC.Tn[13].n42 VGND 0.04124f
C11481 XThC.Tn[13].n43 VGND 0.02569f
C11482 XThC.Tn[13].n44 VGND 0.08347f
C11483 XThC.Tn[13].n45 VGND 0.13936f
C11484 XThC.Tn[13].t26 VGND 0.01577f
C11485 XThC.Tn[13].t40 VGND 0.01661f
C11486 XThC.Tn[13].n46 VGND 0.04124f
C11487 XThC.Tn[13].n47 VGND 0.02569f
C11488 XThC.Tn[13].n48 VGND 0.08347f
C11489 XThC.Tn[13].n49 VGND 0.13936f
C11490 XThC.Tn[13].t29 VGND 0.01577f
C11491 XThC.Tn[13].t43 VGND 0.01661f
C11492 XThC.Tn[13].n50 VGND 0.04124f
C11493 XThC.Tn[13].n51 VGND 0.02569f
C11494 XThC.Tn[13].n52 VGND 0.08347f
C11495 XThC.Tn[13].n53 VGND 0.13936f
C11496 XThC.Tn[13].t15 VGND 0.01577f
C11497 XThC.Tn[13].t30 VGND 0.01661f
C11498 XThC.Tn[13].n54 VGND 0.04124f
C11499 XThC.Tn[13].n55 VGND 0.02569f
C11500 XThC.Tn[13].n56 VGND 0.08347f
C11501 XThC.Tn[13].n57 VGND 0.13936f
C11502 XThC.Tn[13].t18 VGND 0.01577f
C11503 XThC.Tn[13].t31 VGND 0.01661f
C11504 XThC.Tn[13].n58 VGND 0.04124f
C11505 XThC.Tn[13].n59 VGND 0.02569f
C11506 XThC.Tn[13].n60 VGND 0.08347f
C11507 XThC.Tn[13].n61 VGND 0.13936f
C11508 XThC.Tn[13].t20 VGND 0.01577f
C11509 XThC.Tn[13].t33 VGND 0.01661f
C11510 XThC.Tn[13].n62 VGND 0.04124f
C11511 XThC.Tn[13].n63 VGND 0.02569f
C11512 XThC.Tn[13].n64 VGND 0.08347f
C11513 XThC.Tn[13].n65 VGND 0.13936f
C11514 XThC.Tn[13].t41 VGND 0.01577f
C11515 XThC.Tn[13].t21 VGND 0.01661f
C11516 XThC.Tn[13].n66 VGND 0.04124f
C11517 XThC.Tn[13].n67 VGND 0.02569f
C11518 XThC.Tn[13].n68 VGND 0.08347f
C11519 XThC.Tn[13].n69 VGND 0.13936f
C11520 XThC.Tn[13].n70 VGND 0.72276f
C11521 XThC.Tn[13].n71 VGND 0.25416f
C11522 XThC.Tn[13].t0 VGND 0.01261f
C11523 XThC.Tn[13].t2 VGND 0.01261f
C11524 XThC.Tn[13].n72 VGND 0.02523f
C11525 XThC.Tn[13].t3 VGND 0.01261f
C11526 XThC.Tn[13].t1 VGND 0.01261f
C11527 XThC.Tn[13].n73 VGND 0.03146f
C11528 XThC.Tn[13].n74 VGND 0.05816f
C11529 XThC.Tn[8].t9 VGND 0.01312f
C11530 XThC.Tn[8].t8 VGND 0.01312f
C11531 XThC.Tn[8].n0 VGND 0.03271f
C11532 XThC.Tn[8].t11 VGND 0.01312f
C11533 XThC.Tn[8].t10 VGND 0.01312f
C11534 XThC.Tn[8].n1 VGND 0.02623f
C11535 XThC.Tn[8].n2 VGND 0.06599f
C11536 XThC.Tn[8].n3 VGND 0.02467f
C11537 XThC.Tn[8].t13 VGND 0.0164f
C11538 XThC.Tn[8].t26 VGND 0.01727f
C11539 XThC.Tn[8].n4 VGND 0.04289f
C11540 XThC.Tn[8].n5 VGND 0.02672f
C11541 XThC.Tn[8].n6 VGND 0.08657f
C11542 XThC.Tn[8].t23 VGND 0.0164f
C11543 XThC.Tn[8].t36 VGND 0.01727f
C11544 XThC.Tn[8].n7 VGND 0.04289f
C11545 XThC.Tn[8].n8 VGND 0.02672f
C11546 XThC.Tn[8].n9 VGND 0.08681f
C11547 XThC.Tn[8].n10 VGND 0.14494f
C11548 XThC.Tn[8].t35 VGND 0.0164f
C11549 XThC.Tn[8].t17 VGND 0.01727f
C11550 XThC.Tn[8].n11 VGND 0.04289f
C11551 XThC.Tn[8].n12 VGND 0.02672f
C11552 XThC.Tn[8].n13 VGND 0.08681f
C11553 XThC.Tn[8].n14 VGND 0.14494f
C11554 XThC.Tn[8].t37 VGND 0.0164f
C11555 XThC.Tn[8].t18 VGND 0.01727f
C11556 XThC.Tn[8].n15 VGND 0.04289f
C11557 XThC.Tn[8].n16 VGND 0.02672f
C11558 XThC.Tn[8].n17 VGND 0.08681f
C11559 XThC.Tn[8].n18 VGND 0.14494f
C11560 XThC.Tn[8].t15 VGND 0.0164f
C11561 XThC.Tn[8].t29 VGND 0.01727f
C11562 XThC.Tn[8].n19 VGND 0.04289f
C11563 XThC.Tn[8].n20 VGND 0.02672f
C11564 XThC.Tn[8].n21 VGND 0.08681f
C11565 XThC.Tn[8].n22 VGND 0.14494f
C11566 XThC.Tn[8].t25 VGND 0.0164f
C11567 XThC.Tn[8].t40 VGND 0.01727f
C11568 XThC.Tn[8].n23 VGND 0.04289f
C11569 XThC.Tn[8].n24 VGND 0.02672f
C11570 XThC.Tn[8].n25 VGND 0.08681f
C11571 XThC.Tn[8].n26 VGND 0.14494f
C11572 XThC.Tn[8].t38 VGND 0.0164f
C11573 XThC.Tn[8].t19 VGND 0.01727f
C11574 XThC.Tn[8].n27 VGND 0.04289f
C11575 XThC.Tn[8].n28 VGND 0.02672f
C11576 XThC.Tn[8].n29 VGND 0.08681f
C11577 XThC.Tn[8].n30 VGND 0.14494f
C11578 XThC.Tn[8].t16 VGND 0.0164f
C11579 XThC.Tn[8].t30 VGND 0.01727f
C11580 XThC.Tn[8].n31 VGND 0.04289f
C11581 XThC.Tn[8].n32 VGND 0.02672f
C11582 XThC.Tn[8].n33 VGND 0.08681f
C11583 XThC.Tn[8].n34 VGND 0.14494f
C11584 XThC.Tn[8].t20 VGND 0.0164f
C11585 XThC.Tn[8].t32 VGND 0.01727f
C11586 XThC.Tn[8].n35 VGND 0.04289f
C11587 XThC.Tn[8].n36 VGND 0.02672f
C11588 XThC.Tn[8].n37 VGND 0.08681f
C11589 XThC.Tn[8].n38 VGND 0.14494f
C11590 XThC.Tn[8].t27 VGND 0.0164f
C11591 XThC.Tn[8].t41 VGND 0.01727f
C11592 XThC.Tn[8].n39 VGND 0.04289f
C11593 XThC.Tn[8].n40 VGND 0.02672f
C11594 XThC.Tn[8].n41 VGND 0.08681f
C11595 XThC.Tn[8].n42 VGND 0.14494f
C11596 XThC.Tn[8].t39 VGND 0.0164f
C11597 XThC.Tn[8].t21 VGND 0.01727f
C11598 XThC.Tn[8].n43 VGND 0.04289f
C11599 XThC.Tn[8].n44 VGND 0.02672f
C11600 XThC.Tn[8].n45 VGND 0.08681f
C11601 XThC.Tn[8].n46 VGND 0.14494f
C11602 XThC.Tn[8].t42 VGND 0.0164f
C11603 XThC.Tn[8].t24 VGND 0.01727f
C11604 XThC.Tn[8].n47 VGND 0.04289f
C11605 XThC.Tn[8].n48 VGND 0.02672f
C11606 XThC.Tn[8].n49 VGND 0.08681f
C11607 XThC.Tn[8].n50 VGND 0.14494f
C11608 XThC.Tn[8].t28 VGND 0.0164f
C11609 XThC.Tn[8].t43 VGND 0.01727f
C11610 XThC.Tn[8].n51 VGND 0.04289f
C11611 XThC.Tn[8].n52 VGND 0.02672f
C11612 XThC.Tn[8].n53 VGND 0.08681f
C11613 XThC.Tn[8].n54 VGND 0.14494f
C11614 XThC.Tn[8].t31 VGND 0.0164f
C11615 XThC.Tn[8].t12 VGND 0.01727f
C11616 XThC.Tn[8].n55 VGND 0.04289f
C11617 XThC.Tn[8].n56 VGND 0.02672f
C11618 XThC.Tn[8].n57 VGND 0.08681f
C11619 XThC.Tn[8].n58 VGND 0.14494f
C11620 XThC.Tn[8].t33 VGND 0.0164f
C11621 XThC.Tn[8].t14 VGND 0.01727f
C11622 XThC.Tn[8].n59 VGND 0.04289f
C11623 XThC.Tn[8].n60 VGND 0.02672f
C11624 XThC.Tn[8].n61 VGND 0.08681f
C11625 XThC.Tn[8].n62 VGND 0.14494f
C11626 XThC.Tn[8].t22 VGND 0.0164f
C11627 XThC.Tn[8].t34 VGND 0.01727f
C11628 XThC.Tn[8].n63 VGND 0.04289f
C11629 XThC.Tn[8].n64 VGND 0.02672f
C11630 XThC.Tn[8].n65 VGND 0.08681f
C11631 XThC.Tn[8].n66 VGND 0.14494f
C11632 XThC.Tn[8].n67 VGND 0.60695f
C11633 XThC.Tn[8].n68 VGND 0.23755f
C11634 XThC.Tn[8].t5 VGND 0.02018f
C11635 XThC.Tn[8].t6 VGND 0.02018f
C11636 XThC.Tn[8].n69 VGND 0.0436f
C11637 XThC.Tn[8].t4 VGND 0.02018f
C11638 XThC.Tn[8].t7 VGND 0.02018f
C11639 XThC.Tn[8].n70 VGND 0.06636f
C11640 XThC.Tn[8].n71 VGND 0.18439f
C11641 XThC.Tn[8].n72 VGND 0.02899f
C11642 XThC.Tn[8].t2 VGND 0.02018f
C11643 XThC.Tn[8].t1 VGND 0.02018f
C11644 XThC.Tn[8].n73 VGND 0.04486f
C11645 XThC.Tn[8].t0 VGND 0.02018f
C11646 XThC.Tn[8].t3 VGND 0.02018f
C11647 XThC.Tn[8].n74 VGND 0.06127f
C11648 XThC.Tn[8].n75 VGND 0.19965f
C11649 XThC.XTB1.Y.t1 VGND 0.03224f
C11650 XThC.XTB1.Y.n0 VGND 0.02084f
C11651 XThC.XTB1.Y.n1 VGND 0.02659f
C11652 XThC.XTB1.Y.t0 VGND 0.01618f
C11653 XThC.XTB1.Y.t2 VGND 0.01618f
C11654 XThC.XTB1.Y.n2 VGND 0.03473f
C11655 XThC.XTB1.Y.t17 VGND 0.02517f
C11656 XThC.XTB1.Y.t5 VGND 0.01483f
C11657 XThC.XTB1.Y.n3 VGND 0.02997f
C11658 XThC.XTB1.Y.t6 VGND 0.02517f
C11659 XThC.XTB1.Y.t12 VGND 0.01483f
C11660 XThC.XTB1.Y.n4 VGND 0.01542f
C11661 XThC.XTB1.Y.t8 VGND 0.02517f
C11662 XThC.XTB1.Y.t13 VGND 0.01483f
C11663 XThC.XTB1.Y.n5 VGND 0.03313f
C11664 XThC.XTB1.Y.t11 VGND 0.02517f
C11665 XThC.XTB1.Y.t16 VGND 0.01483f
C11666 XThC.XTB1.Y.n6 VGND 0.03076f
C11667 XThC.XTB1.Y.n7 VGND 0.01871f
C11668 XThC.XTB1.Y.n8 VGND 0.03098f
C11669 XThC.XTB1.Y.n9 VGND 0.01198f
C11670 XThC.XTB1.Y.n10 VGND 0.01463f
C11671 XThC.XTB1.Y.n11 VGND 0.03313f
C11672 XThC.XTB1.Y.n12 VGND 0.01661f
C11673 XThC.XTB1.Y.n13 VGND 0.02824f
C11674 XThC.XTB1.Y.t18 VGND 0.02517f
C11675 XThC.XTB1.Y.t9 VGND 0.01483f
C11676 XThC.XTB1.Y.n14 VGND 0.03392f
C11677 XThC.XTB1.Y.t7 VGND 0.02517f
C11678 XThC.XTB1.Y.t15 VGND 0.01483f
C11679 XThC.XTB1.Y.t14 VGND 0.02517f
C11680 XThC.XTB1.Y.t3 VGND 0.01483f
C11681 XThC.XTB1.Y.t10 VGND 0.02517f
C11682 XThC.XTB1.Y.t4 VGND 0.01483f
C11683 XThC.XTB1.Y.n15 VGND 0.04223f
C11684 XThC.XTB1.Y.n16 VGND 0.0446f
C11685 XThC.XTB1.Y.n17 VGND 0.01719f
C11686 XThC.XTB1.Y.n18 VGND 0.0363f
C11687 XThC.XTB1.Y.n19 VGND 0.01661f
C11688 XThC.XTB1.Y.n20 VGND 0.01378f
C11689 XThC.XTB1.Y.n21 VGND 0.77148f
C11690 XThC.XTB1.Y.n22 VGND 0.07634f
C11691 XThR.Tn[12].t11 VGND 0.02439f
C11692 XThR.Tn[12].t9 VGND 0.02439f
C11693 XThR.Tn[12].n0 VGND 0.07405f
C11694 XThR.Tn[12].t8 VGND 0.02439f
C11695 XThR.Tn[12].t10 VGND 0.02439f
C11696 XThR.Tn[12].n1 VGND 0.05422f
C11697 XThR.Tn[12].n2 VGND 0.24652f
C11698 XThR.Tn[12].t7 VGND 0.01585f
C11699 XThR.Tn[12].t5 VGND 0.01585f
C11700 XThR.Tn[12].n3 VGND 0.03954f
C11701 XThR.Tn[12].t6 VGND 0.01585f
C11702 XThR.Tn[12].t4 VGND 0.01585f
C11703 XThR.Tn[12].n4 VGND 0.03171f
C11704 XThR.Tn[12].n5 VGND 0.07311f
C11705 XThR.Tn[12].t40 VGND 0.01982f
C11706 XThR.Tn[12].t70 VGND 0.02087f
C11707 XThR.Tn[12].n6 VGND 0.05184f
C11708 XThR.Tn[12].n7 VGND 0.09637f
C11709 XThR.Tn[12].t20 VGND 0.01982f
C11710 XThR.Tn[12].t25 VGND 0.02087f
C11711 XThR.Tn[12].n8 VGND 0.05184f
C11712 XThR.Tn[12].t14 VGND 0.01982f
C11713 XThR.Tn[12].t24 VGND 0.02087f
C11714 XThR.Tn[12].n9 VGND 0.05182f
C11715 XThR.Tn[12].n10 VGND 0.03985f
C11716 XThR.Tn[12].n11 VGND 0.0076f
C11717 XThR.Tn[12].n12 VGND 0.11895f
C11718 XThR.Tn[12].t35 VGND 0.01982f
C11719 XThR.Tn[12].t63 VGND 0.02087f
C11720 XThR.Tn[12].n13 VGND 0.05184f
C11721 XThR.Tn[12].t30 VGND 0.01982f
C11722 XThR.Tn[12].t59 VGND 0.02087f
C11723 XThR.Tn[12].n14 VGND 0.05182f
C11724 XThR.Tn[12].n15 VGND 0.03985f
C11725 XThR.Tn[12].n16 VGND 0.0076f
C11726 XThR.Tn[12].n17 VGND 0.11895f
C11727 XThR.Tn[12].t71 VGND 0.01982f
C11728 XThR.Tn[12].t19 VGND 0.02087f
C11729 XThR.Tn[12].n18 VGND 0.05184f
C11730 XThR.Tn[12].t69 VGND 0.01982f
C11731 XThR.Tn[12].t13 VGND 0.02087f
C11732 XThR.Tn[12].n19 VGND 0.05182f
C11733 XThR.Tn[12].n20 VGND 0.03985f
C11734 XThR.Tn[12].n21 VGND 0.0076f
C11735 XThR.Tn[12].n22 VGND 0.11895f
C11736 XThR.Tn[12].t37 VGND 0.01982f
C11737 XThR.Tn[12].t48 VGND 0.02087f
C11738 XThR.Tn[12].n23 VGND 0.05184f
C11739 XThR.Tn[12].t32 VGND 0.01982f
C11740 XThR.Tn[12].t43 VGND 0.02087f
C11741 XThR.Tn[12].n24 VGND 0.05182f
C11742 XThR.Tn[12].n25 VGND 0.03985f
C11743 XThR.Tn[12].n26 VGND 0.0076f
C11744 XThR.Tn[12].n27 VGND 0.11895f
C11745 XThR.Tn[12].t53 VGND 0.01982f
C11746 XThR.Tn[12].t21 VGND 0.02087f
C11747 XThR.Tn[12].n28 VGND 0.05184f
C11748 XThR.Tn[12].t51 VGND 0.01982f
C11749 XThR.Tn[12].t16 VGND 0.02087f
C11750 XThR.Tn[12].n29 VGND 0.05182f
C11751 XThR.Tn[12].n30 VGND 0.03985f
C11752 XThR.Tn[12].n31 VGND 0.0076f
C11753 XThR.Tn[12].n32 VGND 0.11895f
C11754 XThR.Tn[12].t47 VGND 0.01982f
C11755 XThR.Tn[12].t36 VGND 0.02087f
C11756 XThR.Tn[12].n33 VGND 0.05184f
C11757 XThR.Tn[12].t42 VGND 0.01982f
C11758 XThR.Tn[12].t31 VGND 0.02087f
C11759 XThR.Tn[12].n34 VGND 0.05182f
C11760 XThR.Tn[12].n35 VGND 0.03985f
C11761 XThR.Tn[12].n36 VGND 0.0076f
C11762 XThR.Tn[12].n37 VGND 0.11895f
C11763 XThR.Tn[12].t66 VGND 0.01982f
C11764 XThR.Tn[12].t28 VGND 0.02087f
C11765 XThR.Tn[12].n38 VGND 0.05184f
C11766 XThR.Tn[12].t61 VGND 0.01982f
C11767 XThR.Tn[12].t26 VGND 0.02087f
C11768 XThR.Tn[12].n39 VGND 0.05182f
C11769 XThR.Tn[12].n40 VGND 0.03985f
C11770 XThR.Tn[12].n41 VGND 0.0076f
C11771 XThR.Tn[12].n42 VGND 0.11895f
C11772 XThR.Tn[12].t23 VGND 0.01982f
C11773 XThR.Tn[12].t46 VGND 0.02087f
C11774 XThR.Tn[12].n43 VGND 0.05184f
C11775 XThR.Tn[12].t18 VGND 0.01982f
C11776 XThR.Tn[12].t41 VGND 0.02087f
C11777 XThR.Tn[12].n44 VGND 0.05182f
C11778 XThR.Tn[12].n45 VGND 0.03985f
C11779 XThR.Tn[12].n46 VGND 0.0076f
C11780 XThR.Tn[12].n47 VGND 0.11895f
C11781 XThR.Tn[12].t39 VGND 0.01982f
C11782 XThR.Tn[12].t65 VGND 0.02087f
C11783 XThR.Tn[12].n48 VGND 0.05184f
C11784 XThR.Tn[12].t34 VGND 0.01982f
C11785 XThR.Tn[12].t60 VGND 0.02087f
C11786 XThR.Tn[12].n49 VGND 0.05182f
C11787 XThR.Tn[12].n50 VGND 0.03985f
C11788 XThR.Tn[12].n51 VGND 0.0076f
C11789 XThR.Tn[12].n52 VGND 0.11895f
C11790 XThR.Tn[12].t12 VGND 0.01982f
C11791 XThR.Tn[12].t22 VGND 0.02087f
C11792 XThR.Tn[12].n53 VGND 0.05184f
C11793 XThR.Tn[12].t72 VGND 0.01982f
C11794 XThR.Tn[12].t17 VGND 0.02087f
C11795 XThR.Tn[12].n54 VGND 0.05182f
C11796 XThR.Tn[12].n55 VGND 0.03985f
C11797 XThR.Tn[12].n56 VGND 0.0076f
C11798 XThR.Tn[12].n57 VGND 0.11895f
C11799 XThR.Tn[12].t50 VGND 0.01982f
C11800 XThR.Tn[12].t57 VGND 0.02087f
C11801 XThR.Tn[12].n58 VGND 0.05184f
C11802 XThR.Tn[12].t45 VGND 0.01982f
C11803 XThR.Tn[12].t55 VGND 0.02087f
C11804 XThR.Tn[12].n59 VGND 0.05182f
C11805 XThR.Tn[12].n60 VGND 0.03985f
C11806 XThR.Tn[12].n61 VGND 0.0076f
C11807 XThR.Tn[12].n62 VGND 0.11895f
C11808 XThR.Tn[12].t68 VGND 0.01982f
C11809 XThR.Tn[12].t29 VGND 0.02087f
C11810 XThR.Tn[12].n63 VGND 0.05184f
C11811 XThR.Tn[12].t64 VGND 0.01982f
C11812 XThR.Tn[12].t27 VGND 0.02087f
C11813 XThR.Tn[12].n64 VGND 0.05182f
C11814 XThR.Tn[12].n65 VGND 0.03985f
C11815 XThR.Tn[12].n66 VGND 0.0076f
C11816 XThR.Tn[12].n67 VGND 0.11895f
C11817 XThR.Tn[12].t38 VGND 0.01982f
C11818 XThR.Tn[12].t49 VGND 0.02087f
C11819 XThR.Tn[12].n68 VGND 0.05184f
C11820 XThR.Tn[12].t33 VGND 0.01982f
C11821 XThR.Tn[12].t44 VGND 0.02087f
C11822 XThR.Tn[12].n69 VGND 0.05182f
C11823 XThR.Tn[12].n70 VGND 0.03985f
C11824 XThR.Tn[12].n71 VGND 0.0076f
C11825 XThR.Tn[12].n72 VGND 0.11895f
C11826 XThR.Tn[12].t54 VGND 0.01982f
C11827 XThR.Tn[12].t67 VGND 0.02087f
C11828 XThR.Tn[12].n73 VGND 0.05184f
C11829 XThR.Tn[12].t52 VGND 0.01982f
C11830 XThR.Tn[12].t62 VGND 0.02087f
C11831 XThR.Tn[12].n74 VGND 0.05182f
C11832 XThR.Tn[12].n75 VGND 0.03985f
C11833 XThR.Tn[12].n76 VGND 0.0076f
C11834 XThR.Tn[12].n77 VGND 0.11895f
C11835 XThR.Tn[12].t15 VGND 0.01982f
C11836 XThR.Tn[12].t58 VGND 0.02087f
C11837 XThR.Tn[12].n78 VGND 0.05184f
C11838 XThR.Tn[12].t73 VGND 0.01982f
C11839 XThR.Tn[12].t56 VGND 0.02087f
C11840 XThR.Tn[12].n79 VGND 0.05182f
C11841 XThR.Tn[12].n80 VGND 0.03985f
C11842 XThR.Tn[12].n81 VGND 0.0076f
C11843 XThR.Tn[12].n82 VGND 0.11895f
C11844 XThR.Tn[12].n83 VGND 0.10865f
C11845 XThR.Tn[12].n84 VGND 0.37056f
C11846 XThR.Tn[12].t2 VGND 0.02439f
C11847 XThR.Tn[12].t0 VGND 0.02439f
C11848 XThR.Tn[12].n85 VGND 0.0527f
C11849 XThR.Tn[12].t3 VGND 0.02439f
C11850 XThR.Tn[12].t1 VGND 0.02439f
C11851 XThR.Tn[12].n86 VGND 0.0802f
C11852 XThR.Tn[12].n87 VGND 0.2227f
C11853 XThR.Tn[12].n88 VGND 0.01098f
C11854 Vbias.t2 VGND 0.31005f
C11855 Vbias.t1 VGND 1.22012f
C11856 Vbias.n0 VGND 2.27946f
C11857 Vbias.t5 VGND 0.06652f
C11858 Vbias.t4 VGND 0.06652f
C11859 Vbias.n1 VGND 0.44817f
C11860 Vbias.t3 VGND 0.06652f
C11861 Vbias.t0 VGND 0.06652f
C11862 Vbias.n2 VGND 0.44817f
C11863 Vbias.n3 VGND 1.34377f
C11864 Vbias.n4 VGND 0.9411f
C11865 Vbias.n5 VGND 0.62914f
C11866 Vbias.t181 VGND 0.32554f
C11867 Vbias.n6 VGND 0.32151f
C11868 Vbias.n7 VGND 0.34218f
C11869 Vbias.t110 VGND 0.32554f
C11870 Vbias.n8 VGND 0.32151f
C11871 Vbias.t210 VGND 0.32554f
C11872 Vbias.n9 VGND 0.32151f
C11873 Vbias.t24 VGND 0.32554f
C11874 Vbias.n10 VGND 0.32151f
C11875 Vbias.n11 VGND 0.04585f
C11876 Vbias.t238 VGND 0.32554f
C11877 Vbias.n12 VGND 0.32151f
C11878 Vbias.n13 VGND 0.09053f
C11879 Vbias.t165 VGND 0.32554f
C11880 Vbias.n14 VGND 0.32151f
C11881 Vbias.n15 VGND 0.09053f
C11882 Vbias.t92 VGND 0.32554f
C11883 Vbias.n16 VGND 0.32151f
C11884 Vbias.n17 VGND 0.09053f
C11885 Vbias.t20 VGND 0.32554f
C11886 Vbias.n18 VGND 0.32151f
C11887 Vbias.n19 VGND 0.09053f
C11888 Vbias.t204 VGND 0.32554f
C11889 Vbias.n20 VGND 0.32151f
C11890 Vbias.n21 VGND 0.09053f
C11891 Vbias.t232 VGND 0.32554f
C11892 Vbias.n22 VGND 0.32151f
C11893 Vbias.n23 VGND 0.09053f
C11894 Vbias.t161 VGND 0.32554f
C11895 Vbias.n24 VGND 0.32151f
C11896 Vbias.n25 VGND 0.09053f
C11897 Vbias.t89 VGND 0.32554f
C11898 Vbias.n26 VGND 0.32151f
C11899 Vbias.n27 VGND 0.09053f
C11900 Vbias.t207 VGND 0.32554f
C11901 Vbias.n28 VGND 0.32151f
C11902 Vbias.n29 VGND 0.09053f
C11903 Vbias.t85 VGND 0.32554f
C11904 Vbias.n30 VGND 0.32151f
C11905 Vbias.n31 VGND 0.09053f
C11906 Vbias.t175 VGND 0.32554f
C11907 Vbias.n32 VGND 0.32151f
C11908 Vbias.n33 VGND 0.09053f
C11909 Vbias.t104 VGND 0.32554f
C11910 Vbias.n34 VGND 0.32151f
C11911 Vbias.n35 VGND 0.09053f
C11912 Vbias.t35 VGND 0.32554f
C11913 Vbias.n36 VGND 0.32151f
C11914 Vbias.n37 VGND 0.09053f
C11915 Vbias.t151 VGND 0.32554f
C11916 Vbias.n38 VGND 0.32151f
C11917 Vbias.t142 VGND 0.32554f
C11918 Vbias.n39 VGND 0.32151f
C11919 Vbias.n40 VGND 0.34218f
C11920 Vbias.t26 VGND 0.32554f
C11921 Vbias.n41 VGND 0.32151f
C11922 Vbias.t259 VGND 0.32554f
C11923 Vbias.n42 VGND 0.32151f
C11924 Vbias.n43 VGND 0.34218f
C11925 Vbias.t114 VGND 0.32554f
C11926 Vbias.n44 VGND 0.32151f
C11927 Vbias.t223 VGND 0.32554f
C11928 Vbias.n45 VGND 0.32151f
C11929 Vbias.n46 VGND 0.34218f
C11930 Vbias.t106 VGND 0.32554f
C11931 Vbias.n47 VGND 0.32151f
C11932 Vbias.t84 VGND 0.32554f
C11933 Vbias.n48 VGND 0.32151f
C11934 Vbias.n49 VGND 0.34218f
C11935 Vbias.t202 VGND 0.32554f
C11936 Vbias.n50 VGND 0.32151f
C11937 Vbias.t111 VGND 0.32554f
C11938 Vbias.n51 VGND 0.32151f
C11939 Vbias.n52 VGND 0.34218f
C11940 Vbias.t254 VGND 0.32554f
C11941 Vbias.n53 VGND 0.32151f
C11942 Vbias.t178 VGND 0.32554f
C11943 Vbias.n54 VGND 0.32151f
C11944 Vbias.n55 VGND 0.34218f
C11945 Vbias.t39 VGND 0.32554f
C11946 Vbias.n56 VGND 0.32151f
C11947 Vbias.t19 VGND 0.32554f
C11948 Vbias.n57 VGND 0.32151f
C11949 Vbias.n58 VGND 0.34218f
C11950 Vbias.t158 VGND 0.32554f
C11951 Vbias.n59 VGND 0.32151f
C11952 Vbias.t72 VGND 0.32554f
C11953 Vbias.n60 VGND 0.32151f
C11954 Vbias.n61 VGND 0.34218f
C11955 Vbias.t184 VGND 0.32554f
C11956 Vbias.n62 VGND 0.32151f
C11957 Vbias.t101 VGND 0.32554f
C11958 Vbias.n63 VGND 0.32151f
C11959 Vbias.n64 VGND 0.34218f
C11960 Vbias.t245 VGND 0.32554f
C11961 Vbias.n65 VGND 0.32151f
C11962 Vbias.t152 VGND 0.32554f
C11963 Vbias.n66 VGND 0.32151f
C11964 Vbias.n67 VGND 0.34218f
C11965 Vbias.t15 VGND 0.32554f
C11966 Vbias.n68 VGND 0.32151f
C11967 Vbias.t182 VGND 0.32554f
C11968 Vbias.n69 VGND 0.32151f
C11969 Vbias.n70 VGND 0.34218f
C11970 Vbias.t67 VGND 0.32554f
C11971 Vbias.n71 VGND 0.32151f
C11972 Vbias.t59 VGND 0.32554f
C11973 Vbias.n72 VGND 0.32151f
C11974 Vbias.n73 VGND 0.34218f
C11975 Vbias.t174 VGND 0.32554f
C11976 Vbias.n74 VGND 0.32151f
C11977 Vbias.t79 VGND 0.32554f
C11978 Vbias.n75 VGND 0.32151f
C11979 Vbias.n76 VGND 0.34218f
C11980 Vbias.t216 VGND 0.32554f
C11981 Vbias.n77 VGND 0.32151f
C11982 Vbias.t140 VGND 0.32554f
C11983 Vbias.n78 VGND 0.32151f
C11984 Vbias.t215 VGND 0.32554f
C11985 Vbias.n79 VGND 0.32151f
C11986 Vbias.n80 VGND 0.08788f
C11987 Vbias.n81 VGND 0.34218f
C11988 Vbias.t30 VGND 0.32554f
C11989 Vbias.n82 VGND 0.32151f
C11990 Vbias.t100 VGND 0.32554f
C11991 Vbias.n83 VGND 0.32151f
C11992 Vbias.n84 VGND 0.34218f
C11993 Vbias.t6 VGND 0.32554f
C11994 Vbias.n85 VGND 0.32151f
C11995 Vbias.t103 VGND 0.32554f
C11996 Vbias.n86 VGND 0.32151f
C11997 Vbias.n87 VGND 0.34218f
C11998 Vbias.t203 VGND 0.32554f
C11999 Vbias.n88 VGND 0.32151f
C12000 Vbias.t214 VGND 0.32554f
C12001 Vbias.n89 VGND 0.32151f
C12002 Vbias.n90 VGND 0.34218f
C12003 Vbias.t115 VGND 0.32554f
C12004 Vbias.n91 VGND 0.32151f
C12005 Vbias.t206 VGND 0.32554f
C12006 Vbias.n92 VGND 0.32151f
C12007 Vbias.n93 VGND 0.34218f
C12008 Vbias.t38 VGND 0.32554f
C12009 Vbias.n94 VGND 0.32151f
C12010 Vbias.t131 VGND 0.32554f
C12011 Vbias.n95 VGND 0.32151f
C12012 Vbias.n96 VGND 0.34218f
C12013 Vbias.t34 VGND 0.32554f
C12014 Vbias.n97 VGND 0.32151f
C12015 Vbias.t116 VGND 0.32554f
C12016 Vbias.n98 VGND 0.32151f
C12017 Vbias.n99 VGND 0.34218f
C12018 Vbias.t218 VGND 0.32554f
C12019 Vbias.n100 VGND 0.32151f
C12020 Vbias.t42 VGND 0.32554f
C12021 Vbias.n101 VGND 0.32151f
C12022 Vbias.n102 VGND 0.34218f
C12023 Vbias.t209 VGND 0.32554f
C12024 Vbias.n103 VGND 0.32151f
C12025 Vbias.t231 VGND 0.32554f
C12026 Vbias.n104 VGND 0.32151f
C12027 Vbias.n105 VGND 0.34218f
C12028 Vbias.t70 VGND 0.32554f
C12029 Vbias.n106 VGND 0.32151f
C12030 Vbias.t143 VGND 0.32554f
C12031 Vbias.n107 VGND 0.32151f
C12032 Vbias.n108 VGND 0.34218f
C12033 Vbias.t43 VGND 0.32554f
C12034 Vbias.n109 VGND 0.32151f
C12035 Vbias.t134 VGND 0.32554f
C12036 Vbias.n110 VGND 0.32151f
C12037 Vbias.n111 VGND 0.34218f
C12038 Vbias.t228 VGND 0.32554f
C12039 Vbias.n112 VGND 0.32151f
C12040 Vbias.t252 VGND 0.32554f
C12041 Vbias.n113 VGND 0.32151f
C12042 Vbias.n114 VGND 0.34218f
C12043 Vbias.t159 VGND 0.32554f
C12044 Vbias.n115 VGND 0.32151f
C12045 Vbias.t47 VGND 0.32554f
C12046 Vbias.n116 VGND 0.32151f
C12047 Vbias.n117 VGND 0.34218f
C12048 Vbias.t148 VGND 0.32554f
C12049 Vbias.n118 VGND 0.32151f
C12050 Vbias.t170 VGND 0.32554f
C12051 Vbias.n119 VGND 0.32151f
C12052 Vbias.n120 VGND 0.34218f
C12053 Vbias.t78 VGND 0.32554f
C12054 Vbias.n121 VGND 0.32151f
C12055 Vbias.t249 VGND 0.32554f
C12056 Vbias.n122 VGND 0.32151f
C12057 Vbias.n123 VGND 0.34218f
C12058 Vbias.n124 VGND 0.34218f
C12059 Vbias.t86 VGND 0.32554f
C12060 Vbias.n125 VGND 0.32151f
C12061 Vbias.n126 VGND 0.61282f
C12062 Vbias.n127 VGND 0.19121f
C12063 Vbias.t194 VGND 0.32554f
C12064 Vbias.n128 VGND 0.32151f
C12065 Vbias.t61 VGND 0.32554f
C12066 Vbias.n129 VGND 0.32151f
C12067 Vbias.n130 VGND 0.19121f
C12068 Vbias.n131 VGND 0.26094f
C12069 Vbias.n132 VGND 0.35295f
C12070 Vbias.n133 VGND 0.09053f
C12071 Vbias.n134 VGND 0.19121f
C12072 Vbias.n135 VGND 0.62914f
C12073 Vbias.t31 VGND 0.32554f
C12074 Vbias.n136 VGND 0.32151f
C12075 Vbias.n137 VGND 0.09053f
C12076 Vbias.n138 VGND 0.19121f
C12077 Vbias.t132 VGND 0.32554f
C12078 Vbias.n139 VGND 0.32151f
C12079 Vbias.n140 VGND 0.09053f
C12080 Vbias.n141 VGND 0.19121f
C12081 Vbias.t139 VGND 0.32554f
C12082 Vbias.n142 VGND 0.32151f
C12083 Vbias.n143 VGND 0.09053f
C12084 Vbias.n144 VGND 0.19121f
C12085 Vbias.t224 VGND 0.32554f
C12086 Vbias.n145 VGND 0.32151f
C12087 Vbias.n146 VGND 0.09053f
C12088 Vbias.n147 VGND 0.19121f
C12089 Vbias.t58 VGND 0.32554f
C12090 Vbias.n148 VGND 0.32151f
C12091 Vbias.n149 VGND 0.09053f
C12092 Vbias.n150 VGND 0.19121f
C12093 Vbias.t145 VGND 0.32554f
C12094 Vbias.n151 VGND 0.32151f
C12095 Vbias.n152 VGND 0.09053f
C12096 Vbias.n153 VGND 0.19121f
C12097 Vbias.t230 VGND 0.32554f
C12098 Vbias.n154 VGND 0.32151f
C12099 Vbias.n155 VGND 0.09053f
C12100 Vbias.n156 VGND 0.19121f
C12101 Vbias.t253 VGND 0.32554f
C12102 Vbias.n157 VGND 0.32151f
C12103 Vbias.n158 VGND 0.09053f
C12104 Vbias.n159 VGND 0.19121f
C12105 Vbias.t71 VGND 0.32554f
C12106 Vbias.n160 VGND 0.32151f
C12107 Vbias.n161 VGND 0.09053f
C12108 Vbias.n162 VGND 0.19121f
C12109 Vbias.t157 VGND 0.32554f
C12110 Vbias.n163 VGND 0.32151f
C12111 Vbias.n164 VGND 0.09053f
C12112 Vbias.n165 VGND 0.19121f
C12113 Vbias.t177 VGND 0.32554f
C12114 Vbias.n166 VGND 0.32151f
C12115 Vbias.n167 VGND 0.09053f
C12116 Vbias.n168 VGND 0.19121f
C12117 Vbias.t77 VGND 0.32554f
C12118 Vbias.n169 VGND 0.32151f
C12119 Vbias.n170 VGND 0.09053f
C12120 Vbias.n171 VGND 0.19121f
C12121 Vbias.t97 VGND 0.32554f
C12122 Vbias.n172 VGND 0.32151f
C12123 Vbias.n173 VGND 0.09053f
C12124 Vbias.n174 VGND 0.19121f
C12125 Vbias.n175 VGND 0.19121f
C12126 Vbias.t13 VGND 0.32554f
C12127 Vbias.n176 VGND 0.32151f
C12128 Vbias.n177 VGND 0.09053f
C12129 Vbias.n178 VGND 0.19121f
C12130 Vbias.n179 VGND 0.62914f
C12131 Vbias.n180 VGND 0.62914f
C12132 Vbias.t55 VGND 0.32554f
C12133 Vbias.n181 VGND 0.32151f
C12134 Vbias.t189 VGND 0.32554f
C12135 Vbias.n182 VGND 0.32151f
C12136 Vbias.n183 VGND 0.08788f
C12137 Vbias.n184 VGND 0.34218f
C12138 Vbias.t9 VGND 0.32554f
C12139 Vbias.n185 VGND 0.32151f
C12140 Vbias.t83 VGND 0.32554f
C12141 Vbias.n186 VGND 0.32151f
C12142 Vbias.n187 VGND 0.34218f
C12143 Vbias.t10 VGND 0.32554f
C12144 Vbias.n188 VGND 0.32151f
C12145 Vbias.t108 VGND 0.32554f
C12146 Vbias.n189 VGND 0.32151f
C12147 Vbias.n190 VGND 0.34218f
C12148 Vbias.t180 VGND 0.32554f
C12149 Vbias.n191 VGND 0.32151f
C12150 Vbias.t188 VGND 0.32554f
C12151 Vbias.n192 VGND 0.32151f
C12152 Vbias.n193 VGND 0.34218f
C12153 Vbias.t117 VGND 0.32554f
C12154 Vbias.n194 VGND 0.32151f
C12155 Vbias.t208 VGND 0.32554f
C12156 Vbias.n195 VGND 0.32151f
C12157 Vbias.n196 VGND 0.34218f
C12158 Vbias.t23 VGND 0.32554f
C12159 Vbias.n197 VGND 0.32151f
C12160 Vbias.t107 VGND 0.32554f
C12161 Vbias.n198 VGND 0.32151f
C12162 Vbias.n199 VGND 0.34218f
C12163 Vbias.t36 VGND 0.32554f
C12164 Vbias.n200 VGND 0.32151f
C12165 Vbias.t120 VGND 0.32554f
C12166 Vbias.n201 VGND 0.32151f
C12167 Vbias.n202 VGND 0.34218f
C12168 Vbias.t192 VGND 0.32554f
C12169 Vbias.n203 VGND 0.32151f
C12170 Vbias.t28 VGND 0.32554f
C12171 Vbias.n204 VGND 0.32151f
C12172 Vbias.n205 VGND 0.34218f
C12173 Vbias.t212 VGND 0.32554f
C12174 Vbias.n206 VGND 0.32151f
C12175 Vbias.t234 VGND 0.32554f
C12176 Vbias.n207 VGND 0.32151f
C12177 Vbias.n208 VGND 0.34218f
C12178 Vbias.t45 VGND 0.32554f
C12179 Vbias.n209 VGND 0.32151f
C12180 Vbias.t119 VGND 0.32554f
C12181 Vbias.n210 VGND 0.32151f
C12182 Vbias.n211 VGND 0.34218f
C12183 Vbias.t46 VGND 0.32554f
C12184 Vbias.n212 VGND 0.32151f
C12185 Vbias.t136 VGND 0.32554f
C12186 Vbias.n213 VGND 0.32151f
C12187 Vbias.n214 VGND 0.34218f
C12188 Vbias.t211 VGND 0.32554f
C12189 Vbias.n215 VGND 0.32151f
C12190 Vbias.t233 VGND 0.32554f
C12191 Vbias.n216 VGND 0.32151f
C12192 Vbias.n217 VGND 0.34218f
C12193 Vbias.t162 VGND 0.32554f
C12194 Vbias.n218 VGND 0.32151f
C12195 Vbias.t51 VGND 0.32554f
C12196 Vbias.n219 VGND 0.32151f
C12197 Vbias.n220 VGND 0.34218f
C12198 Vbias.t123 VGND 0.32554f
C12199 Vbias.n221 VGND 0.32151f
C12200 Vbias.t149 VGND 0.32554f
C12201 Vbias.n222 VGND 0.32151f
C12202 Vbias.n223 VGND 0.34218f
C12203 Vbias.t80 VGND 0.32554f
C12204 Vbias.n224 VGND 0.32151f
C12205 Vbias.t250 VGND 0.32554f
C12206 Vbias.n225 VGND 0.32151f
C12207 Vbias.t64 VGND 0.32554f
C12208 Vbias.n226 VGND 0.32151f
C12209 Vbias.n227 VGND 0.09053f
C12210 Vbias.n228 VGND 0.34218f
C12211 Vbias.t137 VGND 0.32554f
C12212 Vbias.n229 VGND 0.32151f
C12213 Vbias.n230 VGND 0.19121f
C12214 Vbias.n231 VGND 0.19121f
C12215 Vbias.n232 VGND 0.62914f
C12216 Vbias.n233 VGND 0.62914f
C12217 Vbias.t187 VGND 0.32554f
C12218 Vbias.n234 VGND 0.32151f
C12219 Vbias.n235 VGND 0.34218f
C12220 Vbias.t7 VGND 0.32554f
C12221 Vbias.n236 VGND 0.32151f
C12222 Vbias.t243 VGND 0.32554f
C12223 Vbias.n237 VGND 0.32151f
C12224 Vbias.n238 VGND 0.34218f
C12225 Vbias.t168 VGND 0.32554f
C12226 Vbias.n239 VGND 0.32151f
C12227 Vbias.t21 VGND 0.32554f
C12228 Vbias.n240 VGND 0.32151f
C12229 Vbias.n241 VGND 0.34218f
C12230 Vbias.t90 VGND 0.32554f
C12231 Vbias.n242 VGND 0.32151f
C12232 Vbias.t65 VGND 0.32554f
C12233 Vbias.n243 VGND 0.32151f
C12234 Vbias.n244 VGND 0.34218f
C12235 Vbias.t251 VGND 0.32554f
C12236 Vbias.n245 VGND 0.32151f
C12237 Vbias.t164 VGND 0.32554f
C12238 Vbias.n246 VGND 0.32151f
C12239 Vbias.n247 VGND 0.34218f
C12240 Vbias.t236 VGND 0.32554f
C12241 Vbias.n248 VGND 0.32151f
C12242 Vbias.t163 VGND 0.32554f
C12243 Vbias.n249 VGND 0.32151f
C12244 Vbias.n250 VGND 0.34218f
C12245 Vbias.t91 VGND 0.32554f
C12246 Vbias.n251 VGND 0.32151f
C12247 Vbias.t68 VGND 0.32554f
C12248 Vbias.n252 VGND 0.32151f
C12249 Vbias.n253 VGND 0.34218f
C12250 Vbias.t138 VGND 0.32554f
C12251 Vbias.n254 VGND 0.32151f
C12252 Vbias.t50 VGND 0.32554f
C12253 Vbias.n255 VGND 0.32151f
C12254 Vbias.n256 VGND 0.34218f
C12255 Vbias.t237 VGND 0.32554f
C12256 Vbias.n257 VGND 0.32151f
C12257 Vbias.t150 VGND 0.32554f
C12258 Vbias.n258 VGND 0.32151f
C12259 Vbias.n259 VGND 0.34218f
C12260 Vbias.t221 VGND 0.32554f
C12261 Vbias.n260 VGND 0.32151f
C12262 Vbias.t135 VGND 0.32554f
C12263 Vbias.n261 VGND 0.32151f
C12264 Vbias.n262 VGND 0.34218f
C12265 Vbias.t63 VGND 0.32554f
C12266 Vbias.n263 VGND 0.32151f
C12267 Vbias.t235 VGND 0.32554f
C12268 Vbias.n264 VGND 0.32151f
C12269 Vbias.n265 VGND 0.34218f
C12270 Vbias.t48 VGND 0.32554f
C12271 Vbias.n266 VGND 0.32151f
C12272 Vbias.t37 VGND 0.32554f
C12273 Vbias.n267 VGND 0.32151f
C12274 Vbias.n268 VGND 0.34218f
C12275 Vbias.t222 VGND 0.32554f
C12276 Vbias.n269 VGND 0.32151f
C12277 Vbias.t122 VGND 0.32554f
C12278 Vbias.n270 VGND 0.32151f
C12279 Vbias.n271 VGND 0.34218f
C12280 Vbias.t195 VGND 0.32554f
C12281 Vbias.n272 VGND 0.32151f
C12282 Vbias.t121 VGND 0.32554f
C12283 Vbias.n273 VGND 0.32151f
C12284 Vbias.t49 VGND 0.32554f
C12285 Vbias.n274 VGND 0.32151f
C12286 Vbias.n275 VGND 0.08788f
C12287 Vbias.n276 VGND 0.34218f
C12288 Vbias.n277 VGND 0.34218f
C12289 Vbias.t198 VGND 0.32554f
C12290 Vbias.n278 VGND 0.32151f
C12291 Vbias.t255 VGND 0.32554f
C12292 Vbias.n279 VGND 0.32151f
C12293 Vbias.t176 VGND 0.32554f
C12294 Vbias.n280 VGND 0.32151f
C12295 Vbias.n281 VGND 0.19121f
C12296 Vbias.n282 VGND 0.19121f
C12297 Vbias.n283 VGND 0.09053f
C12298 Vbias.n284 VGND 0.34218f
C12299 Vbias.t73 VGND 0.32554f
C12300 Vbias.n285 VGND 0.32151f
C12301 Vbias.t153 VGND 0.32554f
C12302 Vbias.n286 VGND 0.32151f
C12303 Vbias.n287 VGND 0.33936f
C12304 Vbias.t225 VGND 0.32554f
C12305 Vbias.n288 VGND 0.32151f
C12306 Vbias.n289 VGND 0.62914f
C12307 Vbias.n290 VGND 0.62914f
C12308 Vbias.n291 VGND 0.62914f
C12309 Vbias.t146 VGND 0.32554f
C12310 Vbias.n292 VGND 0.32151f
C12311 Vbias.n293 VGND 0.09053f
C12312 Vbias.n294 VGND 0.19121f
C12313 Vbias.n295 VGND 0.19121f
C12314 Vbias.t205 VGND 0.32554f
C12315 Vbias.n296 VGND 0.32151f
C12316 Vbias.n297 VGND 0.33936f
C12317 Vbias.t133 VGND 0.32554f
C12318 Vbias.n298 VGND 0.32151f
C12319 Vbias.t239 VGND 0.32554f
C12320 Vbias.n299 VGND 0.32151f
C12321 Vbias.n300 VGND 0.33936f
C12322 Vbias.t52 VGND 0.32554f
C12323 Vbias.n301 VGND 0.32151f
C12324 Vbias.t32 VGND 0.32554f
C12325 Vbias.n302 VGND 0.32151f
C12326 Vbias.n303 VGND 0.33936f
C12327 Vbias.t217 VGND 0.32554f
C12328 Vbias.n304 VGND 0.32151f
C12329 Vbias.t126 VGND 0.32554f
C12330 Vbias.n305 VGND 0.32151f
C12331 Vbias.n306 VGND 0.33936f
C12332 Vbias.t199 VGND 0.32554f
C12333 Vbias.n307 VGND 0.32151f
C12334 Vbias.t125 VGND 0.32554f
C12335 Vbias.n308 VGND 0.32151f
C12336 Vbias.n309 VGND 0.33936f
C12337 Vbias.t53 VGND 0.32554f
C12338 Vbias.n310 VGND 0.32151f
C12339 Vbias.t33 VGND 0.32554f
C12340 Vbias.n311 VGND 0.32151f
C12341 Vbias.n312 VGND 0.33936f
C12342 Vbias.t102 VGND 0.32554f
C12343 Vbias.n313 VGND 0.32151f
C12344 Vbias.t18 VGND 0.32554f
C12345 Vbias.n314 VGND 0.32151f
C12346 Vbias.n315 VGND 0.33936f
C12347 Vbias.t200 VGND 0.32554f
C12348 Vbias.n316 VGND 0.32151f
C12349 Vbias.t112 VGND 0.32554f
C12350 Vbias.n317 VGND 0.32151f
C12351 Vbias.n318 VGND 0.33936f
C12352 Vbias.t183 VGND 0.32554f
C12353 Vbias.n319 VGND 0.32151f
C12354 Vbias.t99 VGND 0.32554f
C12355 Vbias.n320 VGND 0.32151f
C12356 Vbias.n321 VGND 0.33936f
C12357 Vbias.t29 VGND 0.32554f
C12358 Vbias.n322 VGND 0.32151f
C12359 Vbias.t196 VGND 0.32554f
C12360 Vbias.n323 VGND 0.32151f
C12361 Vbias.n324 VGND 0.33936f
C12362 Vbias.t14 VGND 0.32554f
C12363 Vbias.n325 VGND 0.32151f
C12364 Vbias.t261 VGND 0.32554f
C12365 Vbias.n326 VGND 0.32151f
C12366 Vbias.n327 VGND 0.33936f
C12367 Vbias.t185 VGND 0.32554f
C12368 Vbias.n328 VGND 0.32151f
C12369 Vbias.t16 VGND 0.32554f
C12370 Vbias.n329 VGND 0.32151f
C12371 Vbias.n330 VGND 0.08788f
C12372 Vbias.t88 VGND 0.32554f
C12373 Vbias.n331 VGND 0.32151f
C12374 Vbias.n332 VGND 0.33936f
C12375 Vbias.t160 VGND 0.32554f
C12376 Vbias.n333 VGND 0.32151f
C12377 Vbias.t87 VGND 0.32554f
C12378 Vbias.n334 VGND 0.32151f
C12379 Vbias.t57 VGND 0.32554f
C12380 Vbias.n335 VGND 0.32151f
C12381 Vbias.t193 VGND 0.32554f
C12382 Vbias.n336 VGND 0.32151f
C12383 Vbias.n337 VGND 0.09053f
C12384 Vbias.n338 VGND 0.19121f
C12385 Vbias.t173 VGND 0.32554f
C12386 Vbias.n339 VGND 0.32151f
C12387 Vbias.n340 VGND 0.09053f
C12388 Vbias.n341 VGND 0.19121f
C12389 Vbias.t25 VGND 0.32554f
C12390 Vbias.n342 VGND 0.32151f
C12391 Vbias.n343 VGND 0.09053f
C12392 Vbias.n344 VGND 0.19121f
C12393 Vbias.t258 VGND 0.32554f
C12394 Vbias.n345 VGND 0.32151f
C12395 Vbias.n346 VGND 0.09053f
C12396 Vbias.n347 VGND 0.19121f
C12397 Vbias.t171 VGND 0.32554f
C12398 Vbias.n348 VGND 0.32151f
C12399 Vbias.n349 VGND 0.09053f
C12400 Vbias.n350 VGND 0.19121f
C12401 Vbias.t96 VGND 0.32554f
C12402 Vbias.n351 VGND 0.32151f
C12403 Vbias.n352 VGND 0.09053f
C12404 Vbias.n353 VGND 0.19121f
C12405 Vbias.t76 VGND 0.32554f
C12406 Vbias.n354 VGND 0.32151f
C12407 Vbias.n355 VGND 0.09053f
C12408 Vbias.n356 VGND 0.19121f
C12409 Vbias.t247 VGND 0.32554f
C12410 Vbias.n357 VGND 0.32151f
C12411 Vbias.n358 VGND 0.09053f
C12412 Vbias.n359 VGND 0.19121f
C12413 Vbias.t156 VGND 0.32554f
C12414 Vbias.n360 VGND 0.32151f
C12415 Vbias.n361 VGND 0.09053f
C12416 Vbias.n362 VGND 0.19121f
C12417 Vbias.t69 VGND 0.32554f
C12418 Vbias.n363 VGND 0.32151f
C12419 Vbias.n364 VGND 0.09053f
C12420 Vbias.n365 VGND 0.19121f
C12421 Vbias.t242 VGND 0.32554f
C12422 Vbias.n366 VGND 0.32151f
C12423 Vbias.n367 VGND 0.09053f
C12424 Vbias.n368 VGND 0.19121f
C12425 Vbias.t229 VGND 0.32554f
C12426 Vbias.n369 VGND 0.32151f
C12427 Vbias.n370 VGND 0.09053f
C12428 Vbias.n371 VGND 0.19121f
C12429 Vbias.t130 VGND 0.32554f
C12430 Vbias.n372 VGND 0.32151f
C12431 Vbias.n373 VGND 0.09053f
C12432 Vbias.n374 VGND 0.19121f
C12433 Vbias.n375 VGND 0.08788f
C12434 Vbias.t129 VGND 0.32554f
C12435 Vbias.n376 VGND 0.32151f
C12436 Vbias.n377 VGND 0.19121f
C12437 Vbias.t12 VGND 0.32554f
C12438 Vbias.n378 VGND 0.32151f
C12439 Vbias.n379 VGND 0.04585f
C12440 Vbias.n380 VGND 0.19121f
C12441 Vbias.t248 VGND 0.32554f
C12442 Vbias.n381 VGND 0.32151f
C12443 Vbias.n382 VGND 0.04585f
C12444 Vbias.n383 VGND 0.19121f
C12445 Vbias.t95 VGND 0.32554f
C12446 Vbias.n384 VGND 0.32151f
C12447 Vbias.n385 VGND 0.04585f
C12448 Vbias.n386 VGND 0.19121f
C12449 Vbias.t75 VGND 0.32554f
C12450 Vbias.n387 VGND 0.32151f
C12451 Vbias.n388 VGND 0.04585f
C12452 Vbias.n389 VGND 0.19121f
C12453 Vbias.t246 VGND 0.32554f
C12454 Vbias.n390 VGND 0.32151f
C12455 Vbias.n391 VGND 0.04585f
C12456 Vbias.n392 VGND 0.19121f
C12457 Vbias.t169 VGND 0.32554f
C12458 Vbias.n393 VGND 0.32151f
C12459 Vbias.n394 VGND 0.04585f
C12460 Vbias.n395 VGND 0.19121f
C12461 Vbias.t147 VGND 0.32554f
C12462 Vbias.n396 VGND 0.32151f
C12463 Vbias.n397 VGND 0.04585f
C12464 Vbias.n398 VGND 0.19121f
C12465 Vbias.t60 VGND 0.32554f
C12466 Vbias.n399 VGND 0.32151f
C12467 Vbias.n400 VGND 0.04585f
C12468 Vbias.n401 VGND 0.19121f
C12469 Vbias.t227 VGND 0.32554f
C12470 Vbias.n402 VGND 0.32151f
C12471 Vbias.n403 VGND 0.04585f
C12472 Vbias.n404 VGND 0.19121f
C12473 Vbias.t141 VGND 0.32554f
C12474 Vbias.n405 VGND 0.32151f
C12475 Vbias.n406 VGND 0.04585f
C12476 Vbias.n407 VGND 0.19121f
C12477 Vbias.t56 VGND 0.32554f
C12478 Vbias.n408 VGND 0.32151f
C12479 Vbias.n409 VGND 0.04585f
C12480 Vbias.n410 VGND 0.19121f
C12481 Vbias.t41 VGND 0.32554f
C12482 Vbias.n411 VGND 0.32151f
C12483 Vbias.n412 VGND 0.04585f
C12484 Vbias.n413 VGND 0.19121f
C12485 Vbias.t201 VGND 0.32554f
C12486 Vbias.n414 VGND 0.32151f
C12487 Vbias.n415 VGND 0.04585f
C12488 Vbias.n416 VGND 0.19121f
C12489 Vbias.n417 VGND 0.04319f
C12490 Vbias.n418 VGND 0.33936f
C12491 Vbias.n419 VGND 0.34218f
C12492 Vbias.n420 VGND 0.08788f
C12493 Vbias.n421 VGND 0.19121f
C12494 Vbias.n422 VGND 0.09053f
C12495 Vbias.n423 VGND 0.34218f
C12496 Vbias.n424 VGND 0.34218f
C12497 Vbias.n425 VGND 0.09053f
C12498 Vbias.n426 VGND 0.19121f
C12499 Vbias.n427 VGND 0.19121f
C12500 Vbias.n428 VGND 0.09053f
C12501 Vbias.n429 VGND 0.34218f
C12502 Vbias.n430 VGND 0.34218f
C12503 Vbias.n431 VGND 0.09053f
C12504 Vbias.n432 VGND 0.19121f
C12505 Vbias.n433 VGND 0.19121f
C12506 Vbias.n434 VGND 0.09053f
C12507 Vbias.n435 VGND 0.34218f
C12508 Vbias.n436 VGND 0.34218f
C12509 Vbias.n437 VGND 0.09053f
C12510 Vbias.n438 VGND 0.19121f
C12511 Vbias.n439 VGND 0.19121f
C12512 Vbias.n440 VGND 0.09053f
C12513 Vbias.n441 VGND 0.34218f
C12514 Vbias.n442 VGND 0.34218f
C12515 Vbias.n443 VGND 0.09053f
C12516 Vbias.n444 VGND 0.19121f
C12517 Vbias.n445 VGND 0.19121f
C12518 Vbias.n446 VGND 0.09053f
C12519 Vbias.n447 VGND 0.34218f
C12520 Vbias.n448 VGND 0.34218f
C12521 Vbias.n449 VGND 0.09053f
C12522 Vbias.n450 VGND 0.19121f
C12523 Vbias.n451 VGND 0.19121f
C12524 Vbias.n452 VGND 0.09053f
C12525 Vbias.n453 VGND 0.34218f
C12526 Vbias.n454 VGND 0.34218f
C12527 Vbias.n455 VGND 0.09053f
C12528 Vbias.n456 VGND 0.19121f
C12529 Vbias.n457 VGND 0.19121f
C12530 Vbias.n458 VGND 0.09053f
C12531 Vbias.n459 VGND 0.34218f
C12532 Vbias.n460 VGND 0.34218f
C12533 Vbias.n461 VGND 0.09053f
C12534 Vbias.n462 VGND 0.19121f
C12535 Vbias.n463 VGND 0.19121f
C12536 Vbias.n464 VGND 0.09053f
C12537 Vbias.n465 VGND 0.34218f
C12538 Vbias.n466 VGND 0.34218f
C12539 Vbias.n467 VGND 0.09053f
C12540 Vbias.n468 VGND 0.19121f
C12541 Vbias.n469 VGND 0.19121f
C12542 Vbias.n470 VGND 0.09053f
C12543 Vbias.n471 VGND 0.34218f
C12544 Vbias.n472 VGND 0.34218f
C12545 Vbias.n473 VGND 0.09053f
C12546 Vbias.n474 VGND 0.19121f
C12547 Vbias.n475 VGND 0.19121f
C12548 Vbias.n476 VGND 0.09053f
C12549 Vbias.n477 VGND 0.34218f
C12550 Vbias.n478 VGND 0.34218f
C12551 Vbias.n479 VGND 0.09053f
C12552 Vbias.n480 VGND 0.19121f
C12553 Vbias.n481 VGND 0.19121f
C12554 Vbias.n482 VGND 0.09053f
C12555 Vbias.n483 VGND 0.34218f
C12556 Vbias.n484 VGND 0.34218f
C12557 Vbias.n485 VGND 0.09053f
C12558 Vbias.n486 VGND 0.19121f
C12559 Vbias.n487 VGND 0.19121f
C12560 Vbias.n488 VGND 0.09053f
C12561 Vbias.n489 VGND 0.34218f
C12562 Vbias.n490 VGND 0.34218f
C12563 Vbias.n491 VGND 0.09053f
C12564 Vbias.n492 VGND 0.19121f
C12565 Vbias.n493 VGND 0.19121f
C12566 Vbias.n494 VGND 0.09053f
C12567 Vbias.n495 VGND 0.34218f
C12568 Vbias.n496 VGND 0.34218f
C12569 Vbias.n497 VGND 0.09053f
C12570 Vbias.n498 VGND 0.19121f
C12571 Vbias.n499 VGND 0.19121f
C12572 Vbias.n500 VGND 0.19121f
C12573 Vbias.n501 VGND 0.09053f
C12574 Vbias.n502 VGND 0.34218f
C12575 Vbias.n503 VGND 0.34218f
C12576 Vbias.n504 VGND 0.09053f
C12577 Vbias.n505 VGND 0.19121f
C12578 Vbias.n506 VGND 0.19121f
C12579 Vbias.t81 VGND 0.32554f
C12580 Vbias.n507 VGND 0.32151f
C12581 Vbias.n508 VGND 0.09053f
C12582 Vbias.n509 VGND 0.19121f
C12583 Vbias.t62 VGND 0.32554f
C12584 Vbias.n510 VGND 0.32151f
C12585 Vbias.n511 VGND 0.09053f
C12586 Vbias.n512 VGND 0.19121f
C12587 Vbias.t166 VGND 0.32554f
C12588 Vbias.n513 VGND 0.32151f
C12589 Vbias.n514 VGND 0.09053f
C12590 Vbias.n515 VGND 0.19121f
C12591 Vbias.t144 VGND 0.32554f
C12592 Vbias.n516 VGND 0.32151f
C12593 Vbias.n517 VGND 0.09053f
C12594 Vbias.n518 VGND 0.19121f
C12595 Vbias.t54 VGND 0.32554f
C12596 Vbias.n519 VGND 0.32151f
C12597 Vbias.n520 VGND 0.09053f
C12598 Vbias.n521 VGND 0.19121f
C12599 Vbias.t240 VGND 0.32554f
C12600 Vbias.n522 VGND 0.32151f
C12601 Vbias.n523 VGND 0.09053f
C12602 Vbias.n524 VGND 0.19121f
C12603 Vbias.t219 VGND 0.32554f
C12604 Vbias.n525 VGND 0.32151f
C12605 Vbias.n526 VGND 0.09053f
C12606 Vbias.n527 VGND 0.19121f
C12607 Vbias.t127 VGND 0.32554f
C12608 Vbias.n528 VGND 0.32151f
C12609 Vbias.n529 VGND 0.09053f
C12610 Vbias.n530 VGND 0.19121f
C12611 Vbias.t40 VGND 0.32554f
C12612 Vbias.n531 VGND 0.32151f
C12613 Vbias.n532 VGND 0.09053f
C12614 Vbias.n533 VGND 0.19121f
C12615 Vbias.t213 VGND 0.32554f
C12616 Vbias.n534 VGND 0.32151f
C12617 Vbias.n535 VGND 0.09053f
C12618 Vbias.n536 VGND 0.19121f
C12619 Vbias.t124 VGND 0.32554f
C12620 Vbias.n537 VGND 0.32151f
C12621 Vbias.n538 VGND 0.09053f
C12622 Vbias.n539 VGND 0.19121f
C12623 Vbias.t113 VGND 0.32554f
C12624 Vbias.n540 VGND 0.32151f
C12625 Vbias.n541 VGND 0.09053f
C12626 Vbias.n542 VGND 0.19121f
C12627 Vbias.t17 VGND 0.32554f
C12628 Vbias.n543 VGND 0.32151f
C12629 Vbias.n544 VGND 0.09053f
C12630 Vbias.n545 VGND 0.19121f
C12631 Vbias.n546 VGND 0.08788f
C12632 Vbias.n547 VGND 0.34218f
C12633 Vbias.n548 VGND 0.34218f
C12634 Vbias.n549 VGND 0.08788f
C12635 Vbias.n550 VGND 0.19121f
C12636 Vbias.n551 VGND 0.09053f
C12637 Vbias.n552 VGND 0.34218f
C12638 Vbias.n553 VGND 0.34218f
C12639 Vbias.n554 VGND 0.09053f
C12640 Vbias.n555 VGND 0.19121f
C12641 Vbias.n556 VGND 0.19121f
C12642 Vbias.n557 VGND 0.09053f
C12643 Vbias.n558 VGND 0.34218f
C12644 Vbias.n559 VGND 0.34218f
C12645 Vbias.n560 VGND 0.09053f
C12646 Vbias.n561 VGND 0.19121f
C12647 Vbias.n562 VGND 0.19121f
C12648 Vbias.n563 VGND 0.09053f
C12649 Vbias.n564 VGND 0.34218f
C12650 Vbias.n565 VGND 0.34218f
C12651 Vbias.n566 VGND 0.09053f
C12652 Vbias.n567 VGND 0.19121f
C12653 Vbias.n568 VGND 0.19121f
C12654 Vbias.n569 VGND 0.09053f
C12655 Vbias.n570 VGND 0.34218f
C12656 Vbias.n571 VGND 0.34218f
C12657 Vbias.n572 VGND 0.09053f
C12658 Vbias.n573 VGND 0.19121f
C12659 Vbias.n574 VGND 0.19121f
C12660 Vbias.n575 VGND 0.09053f
C12661 Vbias.n576 VGND 0.34218f
C12662 Vbias.n577 VGND 0.34218f
C12663 Vbias.n578 VGND 0.09053f
C12664 Vbias.n579 VGND 0.19121f
C12665 Vbias.n580 VGND 0.19121f
C12666 Vbias.n581 VGND 0.09053f
C12667 Vbias.n582 VGND 0.34218f
C12668 Vbias.n583 VGND 0.34218f
C12669 Vbias.n584 VGND 0.09053f
C12670 Vbias.n585 VGND 0.19121f
C12671 Vbias.n586 VGND 0.19121f
C12672 Vbias.n587 VGND 0.09053f
C12673 Vbias.n588 VGND 0.34218f
C12674 Vbias.n589 VGND 0.34218f
C12675 Vbias.n590 VGND 0.09053f
C12676 Vbias.n591 VGND 0.19121f
C12677 Vbias.n592 VGND 0.19121f
C12678 Vbias.n593 VGND 0.09053f
C12679 Vbias.n594 VGND 0.34218f
C12680 Vbias.n595 VGND 0.34218f
C12681 Vbias.n596 VGND 0.09053f
C12682 Vbias.n597 VGND 0.19121f
C12683 Vbias.n598 VGND 0.19121f
C12684 Vbias.n599 VGND 0.09053f
C12685 Vbias.n600 VGND 0.34218f
C12686 Vbias.n601 VGND 0.34218f
C12687 Vbias.n602 VGND 0.09053f
C12688 Vbias.n603 VGND 0.19121f
C12689 Vbias.n604 VGND 0.19121f
C12690 Vbias.n605 VGND 0.09053f
C12691 Vbias.n606 VGND 0.34218f
C12692 Vbias.n607 VGND 0.34218f
C12693 Vbias.n608 VGND 0.09053f
C12694 Vbias.n609 VGND 0.19121f
C12695 Vbias.n610 VGND 0.19121f
C12696 Vbias.n611 VGND 0.09053f
C12697 Vbias.n612 VGND 0.34218f
C12698 Vbias.n613 VGND 0.34218f
C12699 Vbias.n614 VGND 0.09053f
C12700 Vbias.n615 VGND 0.19121f
C12701 Vbias.n616 VGND 0.19121f
C12702 Vbias.n617 VGND 0.09053f
C12703 Vbias.n618 VGND 0.34218f
C12704 Vbias.n619 VGND 0.34218f
C12705 Vbias.n620 VGND 0.09053f
C12706 Vbias.n621 VGND 0.19121f
C12707 Vbias.n622 VGND 0.19121f
C12708 Vbias.n623 VGND 0.09053f
C12709 Vbias.n624 VGND 0.34218f
C12710 Vbias.n625 VGND 0.34218f
C12711 Vbias.n626 VGND 0.09053f
C12712 Vbias.n627 VGND 0.19121f
C12713 Vbias.n628 VGND 0.19121f
C12714 Vbias.t105 VGND 0.32554f
C12715 Vbias.n629 VGND 0.32151f
C12716 Vbias.n630 VGND 0.09053f
C12717 Vbias.n631 VGND 0.19121f
C12718 Vbias.n632 VGND 0.62914f
C12719 Vbias.n633 VGND 0.62914f
C12720 Vbias.t82 VGND 0.32554f
C12721 Vbias.n634 VGND 0.32151f
C12722 Vbias.n635 VGND 0.08788f
C12723 Vbias.t154 VGND 0.32554f
C12724 Vbias.n636 VGND 0.32151f
C12725 Vbias.n637 VGND 0.09053f
C12726 Vbias.n638 VGND 0.19121f
C12727 Vbias.t257 VGND 0.32554f
C12728 Vbias.n639 VGND 0.32151f
C12729 Vbias.n640 VGND 0.09053f
C12730 Vbias.n641 VGND 0.19121f
C12731 Vbias.t8 VGND 0.32554f
C12732 Vbias.n642 VGND 0.32151f
C12733 Vbias.n643 VGND 0.09053f
C12734 Vbias.n644 VGND 0.19121f
C12735 Vbias.t93 VGND 0.32554f
C12736 Vbias.n645 VGND 0.32151f
C12737 Vbias.n646 VGND 0.09053f
C12738 Vbias.n647 VGND 0.19121f
C12739 Vbias.t179 VGND 0.32554f
C12740 Vbias.n648 VGND 0.32151f
C12741 Vbias.n649 VGND 0.09053f
C12742 Vbias.n650 VGND 0.19121f
C12743 Vbias.t11 VGND 0.32554f
C12744 Vbias.n651 VGND 0.32151f
C12745 Vbias.n652 VGND 0.09053f
C12746 Vbias.n653 VGND 0.19121f
C12747 Vbias.t98 VGND 0.32554f
C12748 Vbias.n654 VGND 0.32151f
C12749 Vbias.n655 VGND 0.09053f
C12750 Vbias.n656 VGND 0.19121f
C12751 Vbias.t118 VGND 0.32554f
C12752 Vbias.n657 VGND 0.32151f
C12753 Vbias.n658 VGND 0.09053f
C12754 Vbias.n659 VGND 0.19121f
C12755 Vbias.t190 VGND 0.32554f
C12756 Vbias.n660 VGND 0.32151f
C12757 Vbias.n661 VGND 0.09053f
C12758 Vbias.n662 VGND 0.19121f
C12759 Vbias.t27 VGND 0.32554f
C12760 Vbias.n663 VGND 0.32151f
C12761 Vbias.n664 VGND 0.09053f
C12762 Vbias.n665 VGND 0.19121f
C12763 Vbias.t44 VGND 0.32554f
C12764 Vbias.n666 VGND 0.32151f
C12765 Vbias.n667 VGND 0.09053f
C12766 Vbias.n668 VGND 0.19121f
C12767 Vbias.t197 VGND 0.32554f
C12768 Vbias.n669 VGND 0.32151f
C12769 Vbias.n670 VGND 0.09053f
C12770 Vbias.n671 VGND 0.19121f
C12771 Vbias.t220 VGND 0.32554f
C12772 Vbias.n672 VGND 0.32151f
C12773 Vbias.n673 VGND 0.09053f
C12774 Vbias.n674 VGND 0.19121f
C12775 Vbias.n675 VGND 0.19121f
C12776 Vbias.n676 VGND 0.19121f
C12777 Vbias.n677 VGND 0.09053f
C12778 Vbias.n678 VGND 0.34218f
C12779 Vbias.n679 VGND 0.34218f
C12780 Vbias.n680 VGND 0.34218f
C12781 Vbias.n681 VGND 0.09053f
C12782 Vbias.n682 VGND 0.19121f
C12783 Vbias.n683 VGND 0.19121f
C12784 Vbias.n684 VGND 0.19121f
C12785 Vbias.n685 VGND 0.09053f
C12786 Vbias.n686 VGND 0.34218f
C12787 Vbias.n687 VGND 0.34218f
C12788 Vbias.n688 VGND 0.09053f
C12789 Vbias.n689 VGND 0.19121f
C12790 Vbias.n690 VGND 0.19121f
C12791 Vbias.n691 VGND 0.09053f
C12792 Vbias.n692 VGND 0.34218f
C12793 Vbias.n693 VGND 0.34218f
C12794 Vbias.n694 VGND 0.09053f
C12795 Vbias.n695 VGND 0.19121f
C12796 Vbias.n696 VGND 0.19121f
C12797 Vbias.n697 VGND 0.09053f
C12798 Vbias.n698 VGND 0.34218f
C12799 Vbias.n699 VGND 0.34218f
C12800 Vbias.n700 VGND 0.09053f
C12801 Vbias.n701 VGND 0.19121f
C12802 Vbias.n702 VGND 0.19121f
C12803 Vbias.n703 VGND 0.09053f
C12804 Vbias.n704 VGND 0.34218f
C12805 Vbias.n705 VGND 0.34218f
C12806 Vbias.n706 VGND 0.09053f
C12807 Vbias.n707 VGND 0.19121f
C12808 Vbias.n708 VGND 0.19121f
C12809 Vbias.n709 VGND 0.09053f
C12810 Vbias.n710 VGND 0.34218f
C12811 Vbias.n711 VGND 0.34218f
C12812 Vbias.n712 VGND 0.09053f
C12813 Vbias.n713 VGND 0.19121f
C12814 Vbias.n714 VGND 0.19121f
C12815 Vbias.n715 VGND 0.09053f
C12816 Vbias.n716 VGND 0.34218f
C12817 Vbias.n717 VGND 0.34218f
C12818 Vbias.n718 VGND 0.09053f
C12819 Vbias.n719 VGND 0.19121f
C12820 Vbias.n720 VGND 0.19121f
C12821 Vbias.n721 VGND 0.09053f
C12822 Vbias.n722 VGND 0.34218f
C12823 Vbias.n723 VGND 0.34218f
C12824 Vbias.n724 VGND 0.09053f
C12825 Vbias.n725 VGND 0.19121f
C12826 Vbias.n726 VGND 0.19121f
C12827 Vbias.n727 VGND 0.09053f
C12828 Vbias.n728 VGND 0.34218f
C12829 Vbias.n729 VGND 0.34218f
C12830 Vbias.n730 VGND 0.09053f
C12831 Vbias.n731 VGND 0.19121f
C12832 Vbias.n732 VGND 0.19121f
C12833 Vbias.n733 VGND 0.09053f
C12834 Vbias.n734 VGND 0.34218f
C12835 Vbias.n735 VGND 0.34218f
C12836 Vbias.n736 VGND 0.09053f
C12837 Vbias.n737 VGND 0.19121f
C12838 Vbias.n738 VGND 0.19121f
C12839 Vbias.n739 VGND 0.09053f
C12840 Vbias.n740 VGND 0.34218f
C12841 Vbias.n741 VGND 0.34218f
C12842 Vbias.n742 VGND 0.09053f
C12843 Vbias.n743 VGND 0.19121f
C12844 Vbias.n744 VGND 0.19121f
C12845 Vbias.n745 VGND 0.09053f
C12846 Vbias.n746 VGND 0.34218f
C12847 Vbias.n747 VGND 0.34218f
C12848 Vbias.n748 VGND 0.09053f
C12849 Vbias.n749 VGND 0.19121f
C12850 Vbias.n750 VGND 0.19121f
C12851 Vbias.n751 VGND 0.09053f
C12852 Vbias.n752 VGND 0.34218f
C12853 Vbias.n753 VGND 0.34218f
C12854 Vbias.n754 VGND 0.09053f
C12855 Vbias.n755 VGND 0.19121f
C12856 Vbias.n756 VGND 0.19121f
C12857 Vbias.n757 VGND 0.09053f
C12858 Vbias.n758 VGND 0.34218f
C12859 Vbias.n759 VGND 0.34218f
C12860 Vbias.n760 VGND 0.09053f
C12861 Vbias.n761 VGND 0.19121f
C12862 Vbias.n762 VGND 0.08788f
C12863 Vbias.n763 VGND 0.34218f
C12864 Vbias.n764 VGND 0.34218f
C12865 Vbias.n765 VGND 0.34218f
C12866 Vbias.n766 VGND 0.08788f
C12867 Vbias.t128 VGND 0.32554f
C12868 Vbias.n767 VGND 0.32151f
C12869 Vbias.n768 VGND 0.09053f
C12870 Vbias.n769 VGND 0.19121f
C12871 Vbias.t226 VGND 0.32554f
C12872 Vbias.n770 VGND 0.32151f
C12873 Vbias.n771 VGND 0.09053f
C12874 Vbias.n772 VGND 0.19121f
C12875 Vbias.t241 VGND 0.32554f
C12876 Vbias.n773 VGND 0.32151f
C12877 Vbias.n774 VGND 0.09053f
C12878 Vbias.n775 VGND 0.19121f
C12879 Vbias.t66 VGND 0.32554f
C12880 Vbias.n776 VGND 0.32151f
C12881 Vbias.n777 VGND 0.09053f
C12882 Vbias.n778 VGND 0.19121f
C12883 Vbias.t155 VGND 0.32554f
C12884 Vbias.n779 VGND 0.32151f
C12885 Vbias.n780 VGND 0.09053f
C12886 Vbias.n781 VGND 0.19121f
C12887 Vbias.t244 VGND 0.32554f
C12888 Vbias.n782 VGND 0.32151f
C12889 Vbias.n783 VGND 0.09053f
C12890 Vbias.n784 VGND 0.19121f
C12891 Vbias.t74 VGND 0.32554f
C12892 Vbias.n785 VGND 0.32151f
C12893 Vbias.n786 VGND 0.09053f
C12894 Vbias.n787 VGND 0.19121f
C12895 Vbias.t94 VGND 0.32554f
C12896 Vbias.n788 VGND 0.32151f
C12897 Vbias.n789 VGND 0.09053f
C12898 Vbias.n790 VGND 0.19121f
C12899 Vbias.t167 VGND 0.32554f
C12900 Vbias.n791 VGND 0.32151f
C12901 Vbias.n792 VGND 0.09053f
C12902 Vbias.n793 VGND 0.19121f
C12903 Vbias.t256 VGND 0.32554f
C12904 Vbias.n794 VGND 0.32151f
C12905 Vbias.n795 VGND 0.09053f
C12906 Vbias.n796 VGND 0.19121f
C12907 Vbias.t22 VGND 0.32554f
C12908 Vbias.n797 VGND 0.32151f
C12909 Vbias.n798 VGND 0.09053f
C12910 Vbias.n799 VGND 0.19121f
C12911 Vbias.t172 VGND 0.32554f
C12912 Vbias.n800 VGND 0.32151f
C12913 Vbias.n801 VGND 0.09053f
C12914 Vbias.n802 VGND 0.19121f
C12915 Vbias.t191 VGND 0.32554f
C12916 Vbias.n803 VGND 0.32151f
C12917 Vbias.n804 VGND 0.09053f
C12918 Vbias.n805 VGND 0.19121f
C12919 Vbias.n806 VGND 0.19121f
C12920 Vbias.t109 VGND 0.32554f
C12921 Vbias.n807 VGND 0.32151f
C12922 Vbias.n808 VGND 0.09053f
C12923 Vbias.n809 VGND 0.19121f
C12924 Vbias.n810 VGND 0.62914f
C12925 Vbias.n811 VGND 0.62914f
C12926 Vbias.n812 VGND 0.62914f
C12927 Vbias.n813 VGND 0.19121f
C12928 Vbias.n814 VGND 0.19121f
C12929 Vbias.n815 VGND 0.09053f
C12930 Vbias.n816 VGND 0.34218f
C12931 Vbias.n817 VGND 0.34218f
C12932 Vbias.n818 VGND 0.09053f
C12933 Vbias.n819 VGND 0.19121f
C12934 Vbias.n820 VGND 0.19121f
C12935 Vbias.n821 VGND 0.19121f
C12936 Vbias.n822 VGND 0.09053f
C12937 Vbias.n823 VGND 0.34218f
C12938 Vbias.n824 VGND 0.34218f
C12939 Vbias.n825 VGND 0.09053f
C12940 Vbias.n826 VGND 0.19121f
C12941 Vbias.n827 VGND 0.19121f
C12942 Vbias.n828 VGND 0.09053f
C12943 Vbias.n829 VGND 0.34218f
C12944 Vbias.n830 VGND 0.34218f
C12945 Vbias.n831 VGND 0.09053f
C12946 Vbias.n832 VGND 0.19121f
C12947 Vbias.n833 VGND 0.19121f
C12948 Vbias.n834 VGND 0.09053f
C12949 Vbias.n835 VGND 0.34218f
C12950 Vbias.n836 VGND 0.34218f
C12951 Vbias.n837 VGND 0.09053f
C12952 Vbias.n838 VGND 0.19121f
C12953 Vbias.n839 VGND 0.19121f
C12954 Vbias.n840 VGND 0.09053f
C12955 Vbias.n841 VGND 0.34218f
C12956 Vbias.n842 VGND 0.34218f
C12957 Vbias.n843 VGND 0.09053f
C12958 Vbias.n844 VGND 0.19121f
C12959 Vbias.n845 VGND 0.19121f
C12960 Vbias.n846 VGND 0.09053f
C12961 Vbias.n847 VGND 0.34218f
C12962 Vbias.n848 VGND 0.34218f
C12963 Vbias.n849 VGND 0.09053f
C12964 Vbias.n850 VGND 0.19121f
C12965 Vbias.n851 VGND 0.19121f
C12966 Vbias.n852 VGND 0.09053f
C12967 Vbias.n853 VGND 0.34218f
C12968 Vbias.n854 VGND 0.34218f
C12969 Vbias.n855 VGND 0.09053f
C12970 Vbias.n856 VGND 0.19121f
C12971 Vbias.n857 VGND 0.19121f
C12972 Vbias.n858 VGND 0.09053f
C12973 Vbias.n859 VGND 0.34218f
C12974 Vbias.n860 VGND 0.34218f
C12975 Vbias.n861 VGND 0.09053f
C12976 Vbias.n862 VGND 0.19121f
C12977 Vbias.n863 VGND 0.19121f
C12978 Vbias.n864 VGND 0.09053f
C12979 Vbias.n865 VGND 0.34218f
C12980 Vbias.n866 VGND 0.34218f
C12981 Vbias.n867 VGND 0.09053f
C12982 Vbias.n868 VGND 0.19121f
C12983 Vbias.n869 VGND 0.19121f
C12984 Vbias.n870 VGND 0.09053f
C12985 Vbias.n871 VGND 0.34218f
C12986 Vbias.n872 VGND 0.34218f
C12987 Vbias.n873 VGND 0.09053f
C12988 Vbias.n874 VGND 0.19121f
C12989 Vbias.n875 VGND 0.19121f
C12990 Vbias.n876 VGND 0.09053f
C12991 Vbias.n877 VGND 0.34218f
C12992 Vbias.n878 VGND 0.34218f
C12993 Vbias.n879 VGND 0.09053f
C12994 Vbias.n880 VGND 0.19121f
C12995 Vbias.n881 VGND 0.19121f
C12996 Vbias.n882 VGND 0.09053f
C12997 Vbias.n883 VGND 0.34218f
C12998 Vbias.n884 VGND 0.34218f
C12999 Vbias.n885 VGND 0.09053f
C13000 Vbias.n886 VGND 0.19121f
C13001 Vbias.n887 VGND 0.19121f
C13002 Vbias.n888 VGND 0.09053f
C13003 Vbias.n889 VGND 0.34218f
C13004 Vbias.n890 VGND 0.34218f
C13005 Vbias.n891 VGND 0.09053f
C13006 Vbias.n892 VGND 0.19121f
C13007 Vbias.t186 VGND 0.32554f
C13008 Vbias.n893 VGND 0.32151f
C13009 Vbias.n894 VGND 0.08788f
C13010 Vbias.n895 VGND 0.19121f
C13011 Vbias.n896 VGND 0.09053f
C13012 Vbias.n897 VGND 0.34218f
C13013 Vbias.n898 VGND 0.34218f
C13014 Vbias.n899 VGND 0.09053f
C13015 Vbias.n900 VGND 0.19121f
C13016 Vbias.n901 VGND 0.08788f
C13017 Vbias.n902 VGND 0.34218f
C13018 Vbias.n903 VGND 0.34218f
C13019 Vbias.t260 VGND 0.32554f
C13020 Vbias.n904 VGND 0.32151f
C13021 Vbias.n905 VGND 0.25829f
C13022 Vbias.n906 VGND 0.35295f
C13023 Vbias.n907 VGND 0.08788f
C13024 Vbias.n908 VGND 0.19121f
C13025 Vbias.n909 VGND 0.09053f
C13026 Vbias.n910 VGND 0.35295f
C13027 Vbias.n911 VGND 0.26094f
C13028 Vbias.n912 VGND 0.19121f
C13029 Vbias.n913 VGND 0.19121f
C13030 Vbias.n914 VGND 0.26094f
C13031 Vbias.n915 VGND 0.35295f
C13032 Vbias.n916 VGND 0.09053f
C13033 Vbias.n917 VGND 0.19121f
C13034 Vbias.n918 VGND 0.19121f
C13035 Vbias.n919 VGND 0.09053f
C13036 Vbias.n920 VGND 0.35295f
C13037 Vbias.n921 VGND 0.26094f
C13038 Vbias.n922 VGND 0.19121f
C13039 Vbias.n923 VGND 0.19121f
C13040 Vbias.n924 VGND 0.26094f
C13041 Vbias.n925 VGND 0.35295f
C13042 Vbias.n926 VGND 0.09053f
C13043 Vbias.n927 VGND 0.19121f
C13044 Vbias.n928 VGND 0.19121f
C13045 Vbias.n929 VGND 0.09053f
C13046 Vbias.n930 VGND 0.35295f
C13047 Vbias.n931 VGND 0.26094f
C13048 Vbias.n932 VGND 0.19121f
C13049 Vbias.n933 VGND 0.19121f
C13050 Vbias.n934 VGND 0.26094f
C13051 Vbias.n935 VGND 0.35295f
C13052 Vbias.n936 VGND 0.09053f
C13053 Vbias.n937 VGND 0.19121f
C13054 Vbias.n938 VGND 0.19121f
C13055 Vbias.n939 VGND 0.09053f
C13056 Vbias.n940 VGND 0.35295f
C13057 Vbias.n941 VGND 0.26094f
C13058 Vbias.n942 VGND 0.19121f
C13059 Vbias.n943 VGND 0.19121f
C13060 Vbias.n944 VGND 0.26094f
C13061 Vbias.n945 VGND 0.35295f
C13062 Vbias.n946 VGND 0.09053f
C13063 Vbias.n947 VGND 0.19121f
C13064 Vbias.n948 VGND 0.19121f
C13065 Vbias.n949 VGND 0.09053f
C13066 Vbias.n950 VGND 0.35295f
C13067 Vbias.n951 VGND 0.26094f
C13068 Vbias.n952 VGND 0.19121f
C13069 Vbias.n953 VGND 0.19121f
C13070 Vbias.n954 VGND 0.26094f
C13071 Vbias.n955 VGND 0.35295f
C13072 Vbias.n956 VGND 0.09053f
C13073 Vbias.n957 VGND 0.19121f
C13074 Vbias.n958 VGND 0.19121f
C13075 Vbias.n959 VGND 0.09053f
C13076 Vbias.n960 VGND 0.35295f
C13077 Vbias.n961 VGND 0.26094f
C13078 Vbias.n962 VGND 0.19121f
C13079 Vbias.n963 VGND 0.19121f
C13080 Vbias.n964 VGND 0.26094f
C13081 Vbias.n965 VGND 0.35295f
C13082 Vbias.n966 VGND 0.09053f
C13083 Vbias.n967 VGND 0.19121f
C13084 Vbias.n968 VGND 0.19121f
C13085 Vbias.n969 VGND 0.09053f
C13086 Vbias.n970 VGND 0.35295f
C13087 Vbias.n971 VGND 0.26094f
C13088 Vbias.n972 VGND 0.19121f
C13089 Vbias.n973 VGND 0.19121f
C13090 Vbias.n974 VGND 0.26094f
C13091 Vbias.n975 VGND 0.35295f
C13092 Vbias.n976 VGND 0.34218f
C13093 Vbias.n977 VGND 0.34218f
C13094 Vbias.n978 VGND 0.34218f
C13095 Vbias.n979 VGND 0.34218f
C13096 Vbias.n980 VGND 0.34218f
C13097 Vbias.n981 VGND 0.34218f
C13098 Vbias.n982 VGND 0.34218f
C13099 Vbias.n983 VGND 0.34218f
C13100 Vbias.n984 VGND 0.34218f
C13101 Vbias.n985 VGND 0.34218f
C13102 Vbias.n986 VGND 0.34218f
C13103 Vbias.n987 VGND 0.34218f
C13104 Vbias.n988 VGND 0.33936f
C13105 Vbias.n989 VGND 0.09053f
C13106 Vbias.n990 VGND 0.19121f
C13107 Vbias.n991 VGND 0.19121f
C13108 Vbias.n992 VGND 0.09053f
C13109 Vbias.n993 VGND 0.33936f
C13110 Vbias.n994 VGND 0.04585f
C13111 Vbias.n995 VGND 0.19121f
C13112 Vbias.n996 VGND 0.57705f
C13113 Vbias.n997 VGND 1.84902f
C13114 XThR.Tn[4].t9 VGND 0.0234f
C13115 XThR.Tn[4].t10 VGND 0.0234f
C13116 XThR.Tn[4].n0 VGND 0.04724f
C13117 XThR.Tn[4].t8 VGND 0.0234f
C13118 XThR.Tn[4].t11 VGND 0.0234f
C13119 XThR.Tn[4].n1 VGND 0.05528f
C13120 XThR.Tn[4].n2 VGND 0.1658f
C13121 XThR.Tn[4].t7 VGND 0.01521f
C13122 XThR.Tn[4].t4 VGND 0.01521f
C13123 XThR.Tn[4].n3 VGND 0.03464f
C13124 XThR.Tn[4].t6 VGND 0.01521f
C13125 XThR.Tn[4].t5 VGND 0.01521f
C13126 XThR.Tn[4].n4 VGND 0.03464f
C13127 XThR.Tn[4].t0 VGND 0.01521f
C13128 XThR.Tn[4].t1 VGND 0.01521f
C13129 XThR.Tn[4].n5 VGND 0.05772f
C13130 XThR.Tn[4].t3 VGND 0.01521f
C13131 XThR.Tn[4].t2 VGND 0.01521f
C13132 XThR.Tn[4].n6 VGND 0.03464f
C13133 XThR.Tn[4].n7 VGND 0.16498f
C13134 XThR.Tn[4].n8 VGND 0.10199f
C13135 XThR.Tn[4].n9 VGND 0.1151f
C13136 XThR.Tn[4].t45 VGND 0.01902f
C13137 XThR.Tn[4].t13 VGND 0.02003f
C13138 XThR.Tn[4].n10 VGND 0.04974f
C13139 XThR.Tn[4].n11 VGND 0.09248f
C13140 XThR.Tn[4].t25 VGND 0.01902f
C13141 XThR.Tn[4].t30 VGND 0.02003f
C13142 XThR.Tn[4].n12 VGND 0.04974f
C13143 XThR.Tn[4].t20 VGND 0.01902f
C13144 XThR.Tn[4].t29 VGND 0.02003f
C13145 XThR.Tn[4].n13 VGND 0.04973f
C13146 XThR.Tn[4].n14 VGND 0.03824f
C13147 XThR.Tn[4].n15 VGND 0.00729f
C13148 XThR.Tn[4].n16 VGND 0.11415f
C13149 XThR.Tn[4].t40 VGND 0.01902f
C13150 XThR.Tn[4].t68 VGND 0.02003f
C13151 XThR.Tn[4].n17 VGND 0.04974f
C13152 XThR.Tn[4].t35 VGND 0.01902f
C13153 XThR.Tn[4].t64 VGND 0.02003f
C13154 XThR.Tn[4].n18 VGND 0.04973f
C13155 XThR.Tn[4].n19 VGND 0.03824f
C13156 XThR.Tn[4].n20 VGND 0.00729f
C13157 XThR.Tn[4].n21 VGND 0.11415f
C13158 XThR.Tn[4].t14 VGND 0.01902f
C13159 XThR.Tn[4].t24 VGND 0.02003f
C13160 XThR.Tn[4].n22 VGND 0.04974f
C13161 XThR.Tn[4].t12 VGND 0.01902f
C13162 XThR.Tn[4].t18 VGND 0.02003f
C13163 XThR.Tn[4].n23 VGND 0.04973f
C13164 XThR.Tn[4].n24 VGND 0.03824f
C13165 XThR.Tn[4].n25 VGND 0.00729f
C13166 XThR.Tn[4].n26 VGND 0.11415f
C13167 XThR.Tn[4].t42 VGND 0.01902f
C13168 XThR.Tn[4].t53 VGND 0.02003f
C13169 XThR.Tn[4].n27 VGND 0.04974f
C13170 XThR.Tn[4].t37 VGND 0.01902f
C13171 XThR.Tn[4].t48 VGND 0.02003f
C13172 XThR.Tn[4].n28 VGND 0.04973f
C13173 XThR.Tn[4].n29 VGND 0.03824f
C13174 XThR.Tn[4].n30 VGND 0.00729f
C13175 XThR.Tn[4].n31 VGND 0.11415f
C13176 XThR.Tn[4].t58 VGND 0.01902f
C13177 XThR.Tn[4].t26 VGND 0.02003f
C13178 XThR.Tn[4].n32 VGND 0.04974f
C13179 XThR.Tn[4].t56 VGND 0.01902f
C13180 XThR.Tn[4].t21 VGND 0.02003f
C13181 XThR.Tn[4].n33 VGND 0.04973f
C13182 XThR.Tn[4].n34 VGND 0.03824f
C13183 XThR.Tn[4].n35 VGND 0.00729f
C13184 XThR.Tn[4].n36 VGND 0.11415f
C13185 XThR.Tn[4].t52 VGND 0.01902f
C13186 XThR.Tn[4].t41 VGND 0.02003f
C13187 XThR.Tn[4].n37 VGND 0.04974f
C13188 XThR.Tn[4].t47 VGND 0.01902f
C13189 XThR.Tn[4].t36 VGND 0.02003f
C13190 XThR.Tn[4].n38 VGND 0.04973f
C13191 XThR.Tn[4].n39 VGND 0.03824f
C13192 XThR.Tn[4].n40 VGND 0.00729f
C13193 XThR.Tn[4].n41 VGND 0.11415f
C13194 XThR.Tn[4].t71 VGND 0.01902f
C13195 XThR.Tn[4].t33 VGND 0.02003f
C13196 XThR.Tn[4].n42 VGND 0.04974f
C13197 XThR.Tn[4].t66 VGND 0.01902f
C13198 XThR.Tn[4].t31 VGND 0.02003f
C13199 XThR.Tn[4].n43 VGND 0.04973f
C13200 XThR.Tn[4].n44 VGND 0.03824f
C13201 XThR.Tn[4].n45 VGND 0.00729f
C13202 XThR.Tn[4].n46 VGND 0.11415f
C13203 XThR.Tn[4].t28 VGND 0.01902f
C13204 XThR.Tn[4].t51 VGND 0.02003f
C13205 XThR.Tn[4].n47 VGND 0.04974f
C13206 XThR.Tn[4].t23 VGND 0.01902f
C13207 XThR.Tn[4].t46 VGND 0.02003f
C13208 XThR.Tn[4].n48 VGND 0.04973f
C13209 XThR.Tn[4].n49 VGND 0.03824f
C13210 XThR.Tn[4].n50 VGND 0.00729f
C13211 XThR.Tn[4].n51 VGND 0.11415f
C13212 XThR.Tn[4].t44 VGND 0.01902f
C13213 XThR.Tn[4].t70 VGND 0.02003f
C13214 XThR.Tn[4].n52 VGND 0.04974f
C13215 XThR.Tn[4].t39 VGND 0.01902f
C13216 XThR.Tn[4].t65 VGND 0.02003f
C13217 XThR.Tn[4].n53 VGND 0.04973f
C13218 XThR.Tn[4].n54 VGND 0.03824f
C13219 XThR.Tn[4].n55 VGND 0.00729f
C13220 XThR.Tn[4].n56 VGND 0.11415f
C13221 XThR.Tn[4].t17 VGND 0.01902f
C13222 XThR.Tn[4].t27 VGND 0.02003f
C13223 XThR.Tn[4].n57 VGND 0.04974f
C13224 XThR.Tn[4].t15 VGND 0.01902f
C13225 XThR.Tn[4].t22 VGND 0.02003f
C13226 XThR.Tn[4].n58 VGND 0.04973f
C13227 XThR.Tn[4].n59 VGND 0.03824f
C13228 XThR.Tn[4].n60 VGND 0.00729f
C13229 XThR.Tn[4].n61 VGND 0.11415f
C13230 XThR.Tn[4].t55 VGND 0.01902f
C13231 XThR.Tn[4].t62 VGND 0.02003f
C13232 XThR.Tn[4].n62 VGND 0.04974f
C13233 XThR.Tn[4].t50 VGND 0.01902f
C13234 XThR.Tn[4].t60 VGND 0.02003f
C13235 XThR.Tn[4].n63 VGND 0.04973f
C13236 XThR.Tn[4].n64 VGND 0.03824f
C13237 XThR.Tn[4].n65 VGND 0.00729f
C13238 XThR.Tn[4].n66 VGND 0.11415f
C13239 XThR.Tn[4].t73 VGND 0.01902f
C13240 XThR.Tn[4].t34 VGND 0.02003f
C13241 XThR.Tn[4].n67 VGND 0.04974f
C13242 XThR.Tn[4].t69 VGND 0.01902f
C13243 XThR.Tn[4].t32 VGND 0.02003f
C13244 XThR.Tn[4].n68 VGND 0.04973f
C13245 XThR.Tn[4].n69 VGND 0.03824f
C13246 XThR.Tn[4].n70 VGND 0.00729f
C13247 XThR.Tn[4].n71 VGND 0.11415f
C13248 XThR.Tn[4].t43 VGND 0.01902f
C13249 XThR.Tn[4].t54 VGND 0.02003f
C13250 XThR.Tn[4].n72 VGND 0.04974f
C13251 XThR.Tn[4].t38 VGND 0.01902f
C13252 XThR.Tn[4].t49 VGND 0.02003f
C13253 XThR.Tn[4].n73 VGND 0.04973f
C13254 XThR.Tn[4].n74 VGND 0.03824f
C13255 XThR.Tn[4].n75 VGND 0.00729f
C13256 XThR.Tn[4].n76 VGND 0.11415f
C13257 XThR.Tn[4].t59 VGND 0.01902f
C13258 XThR.Tn[4].t72 VGND 0.02003f
C13259 XThR.Tn[4].n77 VGND 0.04974f
C13260 XThR.Tn[4].t57 VGND 0.01902f
C13261 XThR.Tn[4].t67 VGND 0.02003f
C13262 XThR.Tn[4].n78 VGND 0.04973f
C13263 XThR.Tn[4].n79 VGND 0.03824f
C13264 XThR.Tn[4].n80 VGND 0.00729f
C13265 XThR.Tn[4].n81 VGND 0.11415f
C13266 XThR.Tn[4].t19 VGND 0.01902f
C13267 XThR.Tn[4].t63 VGND 0.02003f
C13268 XThR.Tn[4].n82 VGND 0.04974f
C13269 XThR.Tn[4].t16 VGND 0.01902f
C13270 XThR.Tn[4].t61 VGND 0.02003f
C13271 XThR.Tn[4].n83 VGND 0.04973f
C13272 XThR.Tn[4].n84 VGND 0.03824f
C13273 XThR.Tn[4].n85 VGND 0.00729f
C13274 XThR.Tn[4].n86 VGND 0.11415f
C13275 XThR.Tn[4].n87 VGND 0.10426f
C13276 XThR.Tn[4].n88 VGND 0.19698f
C13277 XThR.Tn[9].t10 VGND 0.02417f
C13278 XThR.Tn[9].t8 VGND 0.02417f
C13279 XThR.Tn[9].n0 VGND 0.0734f
C13280 XThR.Tn[9].t11 VGND 0.02417f
C13281 XThR.Tn[9].t9 VGND 0.02417f
C13282 XThR.Tn[9].n1 VGND 0.05374f
C13283 XThR.Tn[9].n2 VGND 0.24436f
C13284 XThR.Tn[9].t5 VGND 0.01571f
C13285 XThR.Tn[9].t7 VGND 0.01571f
C13286 XThR.Tn[9].n3 VGND 0.03919f
C13287 XThR.Tn[9].t4 VGND 0.01571f
C13288 XThR.Tn[9].t6 VGND 0.01571f
C13289 XThR.Tn[9].n4 VGND 0.03143f
C13290 XThR.Tn[9].n5 VGND 0.07906f
C13291 XThR.Tn[9].t27 VGND 0.01965f
C13292 XThR.Tn[9].t54 VGND 0.02069f
C13293 XThR.Tn[9].n6 VGND 0.05138f
C13294 XThR.Tn[9].n7 VGND 0.09552f
C13295 XThR.Tn[9].t67 VGND 0.01965f
C13296 XThR.Tn[9].t72 VGND 0.02069f
C13297 XThR.Tn[9].n8 VGND 0.05138f
C13298 XThR.Tn[9].t59 VGND 0.01965f
C13299 XThR.Tn[9].t65 VGND 0.02069f
C13300 XThR.Tn[9].n9 VGND 0.05136f
C13301 XThR.Tn[9].n10 VGND 0.0395f
C13302 XThR.Tn[9].n11 VGND 0.00753f
C13303 XThR.Tn[9].n12 VGND 0.1179f
C13304 XThR.Tn[9].t19 VGND 0.01965f
C13305 XThR.Tn[9].t48 VGND 0.02069f
C13306 XThR.Tn[9].n13 VGND 0.05138f
C13307 XThR.Tn[9].t14 VGND 0.01965f
C13308 XThR.Tn[9].t41 VGND 0.02069f
C13309 XThR.Tn[9].n14 VGND 0.05136f
C13310 XThR.Tn[9].n15 VGND 0.0395f
C13311 XThR.Tn[9].n16 VGND 0.00753f
C13312 XThR.Tn[9].n17 VGND 0.1179f
C13313 XThR.Tn[9].t55 VGND 0.01965f
C13314 XThR.Tn[9].t66 VGND 0.02069f
C13315 XThR.Tn[9].n18 VGND 0.05138f
C13316 XThR.Tn[9].t49 VGND 0.01965f
C13317 XThR.Tn[9].t58 VGND 0.02069f
C13318 XThR.Tn[9].n19 VGND 0.05136f
C13319 XThR.Tn[9].n20 VGND 0.0395f
C13320 XThR.Tn[9].n21 VGND 0.00753f
C13321 XThR.Tn[9].n22 VGND 0.1179f
C13322 XThR.Tn[9].t21 VGND 0.01965f
C13323 XThR.Tn[9].t32 VGND 0.02069f
C13324 XThR.Tn[9].n23 VGND 0.05138f
C13325 XThR.Tn[9].t16 VGND 0.01965f
C13326 XThR.Tn[9].t26 VGND 0.02069f
C13327 XThR.Tn[9].n24 VGND 0.05136f
C13328 XThR.Tn[9].n25 VGND 0.0395f
C13329 XThR.Tn[9].n26 VGND 0.00753f
C13330 XThR.Tn[9].n27 VGND 0.1179f
C13331 XThR.Tn[9].t39 VGND 0.01965f
C13332 XThR.Tn[9].t68 VGND 0.02069f
C13333 XThR.Tn[9].n28 VGND 0.05138f
C13334 XThR.Tn[9].t35 VGND 0.01965f
C13335 XThR.Tn[9].t60 VGND 0.02069f
C13336 XThR.Tn[9].n29 VGND 0.05136f
C13337 XThR.Tn[9].n30 VGND 0.0395f
C13338 XThR.Tn[9].n31 VGND 0.00753f
C13339 XThR.Tn[9].n32 VGND 0.1179f
C13340 XThR.Tn[9].t31 VGND 0.01965f
C13341 XThR.Tn[9].t20 VGND 0.02069f
C13342 XThR.Tn[9].n33 VGND 0.05138f
C13343 XThR.Tn[9].t25 VGND 0.01965f
C13344 XThR.Tn[9].t15 VGND 0.02069f
C13345 XThR.Tn[9].n34 VGND 0.05136f
C13346 XThR.Tn[9].n35 VGND 0.0395f
C13347 XThR.Tn[9].n36 VGND 0.00753f
C13348 XThR.Tn[9].n37 VGND 0.1179f
C13349 XThR.Tn[9].t51 VGND 0.01965f
C13350 XThR.Tn[9].t12 VGND 0.02069f
C13351 XThR.Tn[9].n38 VGND 0.05138f
C13352 XThR.Tn[9].t44 VGND 0.01965f
C13353 XThR.Tn[9].t71 VGND 0.02069f
C13354 XThR.Tn[9].n39 VGND 0.05136f
C13355 XThR.Tn[9].n40 VGND 0.0395f
C13356 XThR.Tn[9].n41 VGND 0.00753f
C13357 XThR.Tn[9].n42 VGND 0.1179f
C13358 XThR.Tn[9].t70 VGND 0.01965f
C13359 XThR.Tn[9].t30 VGND 0.02069f
C13360 XThR.Tn[9].n43 VGND 0.05138f
C13361 XThR.Tn[9].t62 VGND 0.01965f
C13362 XThR.Tn[9].t24 VGND 0.02069f
C13363 XThR.Tn[9].n44 VGND 0.05136f
C13364 XThR.Tn[9].n45 VGND 0.0395f
C13365 XThR.Tn[9].n46 VGND 0.00753f
C13366 XThR.Tn[9].n47 VGND 0.1179f
C13367 XThR.Tn[9].t23 VGND 0.01965f
C13368 XThR.Tn[9].t50 VGND 0.02069f
C13369 XThR.Tn[9].n48 VGND 0.05138f
C13370 XThR.Tn[9].t18 VGND 0.01965f
C13371 XThR.Tn[9].t42 VGND 0.02069f
C13372 XThR.Tn[9].n49 VGND 0.05136f
C13373 XThR.Tn[9].n50 VGND 0.0395f
C13374 XThR.Tn[9].n51 VGND 0.00753f
C13375 XThR.Tn[9].n52 VGND 0.1179f
C13376 XThR.Tn[9].t63 VGND 0.01965f
C13377 XThR.Tn[9].t69 VGND 0.02069f
C13378 XThR.Tn[9].n53 VGND 0.05138f
C13379 XThR.Tn[9].t56 VGND 0.01965f
C13380 XThR.Tn[9].t61 VGND 0.02069f
C13381 XThR.Tn[9].n54 VGND 0.05136f
C13382 XThR.Tn[9].n55 VGND 0.0395f
C13383 XThR.Tn[9].n56 VGND 0.00753f
C13384 XThR.Tn[9].n57 VGND 0.1179f
C13385 XThR.Tn[9].t34 VGND 0.01965f
C13386 XThR.Tn[9].t43 VGND 0.02069f
C13387 XThR.Tn[9].n58 VGND 0.05138f
C13388 XThR.Tn[9].t29 VGND 0.01965f
C13389 XThR.Tn[9].t37 VGND 0.02069f
C13390 XThR.Tn[9].n59 VGND 0.05136f
C13391 XThR.Tn[9].n60 VGND 0.0395f
C13392 XThR.Tn[9].n61 VGND 0.00753f
C13393 XThR.Tn[9].n62 VGND 0.1179f
C13394 XThR.Tn[9].t53 VGND 0.01965f
C13395 XThR.Tn[9].t13 VGND 0.02069f
C13396 XThR.Tn[9].n63 VGND 0.05138f
C13397 XThR.Tn[9].t47 VGND 0.01965f
C13398 XThR.Tn[9].t73 VGND 0.02069f
C13399 XThR.Tn[9].n64 VGND 0.05136f
C13400 XThR.Tn[9].n65 VGND 0.0395f
C13401 XThR.Tn[9].n66 VGND 0.00753f
C13402 XThR.Tn[9].n67 VGND 0.1179f
C13403 XThR.Tn[9].t22 VGND 0.01965f
C13404 XThR.Tn[9].t33 VGND 0.02069f
C13405 XThR.Tn[9].n68 VGND 0.05138f
C13406 XThR.Tn[9].t17 VGND 0.01965f
C13407 XThR.Tn[9].t28 VGND 0.02069f
C13408 XThR.Tn[9].n69 VGND 0.05136f
C13409 XThR.Tn[9].n70 VGND 0.0395f
C13410 XThR.Tn[9].n71 VGND 0.00753f
C13411 XThR.Tn[9].n72 VGND 0.1179f
C13412 XThR.Tn[9].t40 VGND 0.01965f
C13413 XThR.Tn[9].t52 VGND 0.02069f
C13414 XThR.Tn[9].n73 VGND 0.05138f
C13415 XThR.Tn[9].t36 VGND 0.01965f
C13416 XThR.Tn[9].t45 VGND 0.02069f
C13417 XThR.Tn[9].n74 VGND 0.05136f
C13418 XThR.Tn[9].n75 VGND 0.0395f
C13419 XThR.Tn[9].n76 VGND 0.00753f
C13420 XThR.Tn[9].n77 VGND 0.1179f
C13421 XThR.Tn[9].t64 VGND 0.01965f
C13422 XThR.Tn[9].t46 VGND 0.02069f
C13423 XThR.Tn[9].n78 VGND 0.05138f
C13424 XThR.Tn[9].t57 VGND 0.01965f
C13425 XThR.Tn[9].t38 VGND 0.02069f
C13426 XThR.Tn[9].n79 VGND 0.05136f
C13427 XThR.Tn[9].n80 VGND 0.0395f
C13428 XThR.Tn[9].n81 VGND 0.00753f
C13429 XThR.Tn[9].n82 VGND 0.1179f
C13430 XThR.Tn[9].n83 VGND 0.10769f
C13431 XThR.Tn[9].n84 VGND 0.34936f
C13432 XThR.Tn[9].t2 VGND 0.02417f
C13433 XThR.Tn[9].t0 VGND 0.02417f
C13434 XThR.Tn[9].n85 VGND 0.05223f
C13435 XThR.Tn[9].t3 VGND 0.02417f
C13436 XThR.Tn[9].t1 VGND 0.02417f
C13437 XThR.Tn[9].n86 VGND 0.0795f
C13438 XThR.Tn[9].n87 VGND 0.22074f
C13439 XThR.Tn[9].n88 VGND 0.02956f
C13440 XThR.Tn[0].t6 VGND 0.02264f
C13441 XThR.Tn[0].t7 VGND 0.02264f
C13442 XThR.Tn[0].n0 VGND 0.04571f
C13443 XThR.Tn[0].t5 VGND 0.02264f
C13444 XThR.Tn[0].t4 VGND 0.02264f
C13445 XThR.Tn[0].n1 VGND 0.05348f
C13446 XThR.Tn[0].n2 VGND 0.16042f
C13447 XThR.Tn[0].t9 VGND 0.01472f
C13448 XThR.Tn[0].t10 VGND 0.01472f
C13449 XThR.Tn[0].n3 VGND 0.03352f
C13450 XThR.Tn[0].t8 VGND 0.01472f
C13451 XThR.Tn[0].t11 VGND 0.01472f
C13452 XThR.Tn[0].n4 VGND 0.03352f
C13453 XThR.Tn[0].t2 VGND 0.01472f
C13454 XThR.Tn[0].t3 VGND 0.01472f
C13455 XThR.Tn[0].n5 VGND 0.03352f
C13456 XThR.Tn[0].t1 VGND 0.01472f
C13457 XThR.Tn[0].t0 VGND 0.01472f
C13458 XThR.Tn[0].n6 VGND 0.05585f
C13459 XThR.Tn[0].n7 VGND 0.15962f
C13460 XThR.Tn[0].n8 VGND 0.09867f
C13461 XThR.Tn[0].n9 VGND 0.11136f
C13462 XThR.Tn[0].t73 VGND 0.0184f
C13463 XThR.Tn[0].t37 VGND 0.01938f
C13464 XThR.Tn[0].n10 VGND 0.04813f
C13465 XThR.Tn[0].n11 VGND 0.08947f
C13466 XThR.Tn[0].t47 VGND 0.0184f
C13467 XThR.Tn[0].t55 VGND 0.01938f
C13468 XThR.Tn[0].n12 VGND 0.04813f
C13469 XThR.Tn[0].t23 VGND 0.0184f
C13470 XThR.Tn[0].t29 VGND 0.01938f
C13471 XThR.Tn[0].n13 VGND 0.04811f
C13472 XThR.Tn[0].n14 VGND 0.037f
C13473 XThR.Tn[0].n15 VGND 0.00705f
C13474 XThR.Tn[0].n16 VGND 0.11044f
C13475 XThR.Tn[0].t63 VGND 0.0184f
C13476 XThR.Tn[0].t30 VGND 0.01938f
C13477 XThR.Tn[0].n17 VGND 0.04813f
C13478 XThR.Tn[0].t39 VGND 0.0184f
C13479 XThR.Tn[0].t68 VGND 0.01938f
C13480 XThR.Tn[0].n18 VGND 0.04811f
C13481 XThR.Tn[0].n19 VGND 0.037f
C13482 XThR.Tn[0].n20 VGND 0.00705f
C13483 XThR.Tn[0].n21 VGND 0.11044f
C13484 XThR.Tn[0].t38 VGND 0.0184f
C13485 XThR.Tn[0].t46 VGND 0.01938f
C13486 XThR.Tn[0].n22 VGND 0.04813f
C13487 XThR.Tn[0].t12 VGND 0.0184f
C13488 XThR.Tn[0].t22 VGND 0.01938f
C13489 XThR.Tn[0].n23 VGND 0.04811f
C13490 XThR.Tn[0].n24 VGND 0.037f
C13491 XThR.Tn[0].n25 VGND 0.00705f
C13492 XThR.Tn[0].n26 VGND 0.11044f
C13493 XThR.Tn[0].t65 VGND 0.0184f
C13494 XThR.Tn[0].t15 VGND 0.01938f
C13495 XThR.Tn[0].n27 VGND 0.04813f
C13496 XThR.Tn[0].t41 VGND 0.0184f
C13497 XThR.Tn[0].t53 VGND 0.01938f
C13498 XThR.Tn[0].n28 VGND 0.04811f
C13499 XThR.Tn[0].n29 VGND 0.037f
C13500 XThR.Tn[0].n30 VGND 0.00705f
C13501 XThR.Tn[0].n31 VGND 0.11044f
C13502 XThR.Tn[0].t20 VGND 0.0184f
C13503 XThR.Tn[0].t48 VGND 0.01938f
C13504 XThR.Tn[0].n32 VGND 0.04813f
C13505 XThR.Tn[0].t58 VGND 0.0184f
C13506 XThR.Tn[0].t24 VGND 0.01938f
C13507 XThR.Tn[0].n33 VGND 0.04811f
C13508 XThR.Tn[0].n34 VGND 0.037f
C13509 XThR.Tn[0].n35 VGND 0.00705f
C13510 XThR.Tn[0].n36 VGND 0.11044f
C13511 XThR.Tn[0].t14 VGND 0.0184f
C13512 XThR.Tn[0].t64 VGND 0.01938f
C13513 XThR.Tn[0].n37 VGND 0.04813f
C13514 XThR.Tn[0].t52 VGND 0.0184f
C13515 XThR.Tn[0].t40 VGND 0.01938f
C13516 XThR.Tn[0].n38 VGND 0.04811f
C13517 XThR.Tn[0].n39 VGND 0.037f
C13518 XThR.Tn[0].n40 VGND 0.00705f
C13519 XThR.Tn[0].n41 VGND 0.11044f
C13520 XThR.Tn[0].t32 VGND 0.0184f
C13521 XThR.Tn[0].t57 VGND 0.01938f
C13522 XThR.Tn[0].n42 VGND 0.04813f
C13523 XThR.Tn[0].t70 VGND 0.0184f
C13524 XThR.Tn[0].t35 VGND 0.01938f
C13525 XThR.Tn[0].n43 VGND 0.04811f
C13526 XThR.Tn[0].n44 VGND 0.037f
C13527 XThR.Tn[0].n45 VGND 0.00705f
C13528 XThR.Tn[0].n46 VGND 0.11044f
C13529 XThR.Tn[0].t50 VGND 0.0184f
C13530 XThR.Tn[0].t13 VGND 0.01938f
C13531 XThR.Tn[0].n47 VGND 0.04813f
C13532 XThR.Tn[0].t26 VGND 0.0184f
C13533 XThR.Tn[0].t51 VGND 0.01938f
C13534 XThR.Tn[0].n48 VGND 0.04811f
C13535 XThR.Tn[0].n49 VGND 0.037f
C13536 XThR.Tn[0].n50 VGND 0.00705f
C13537 XThR.Tn[0].n51 VGND 0.11044f
C13538 XThR.Tn[0].t67 VGND 0.0184f
C13539 XThR.Tn[0].t31 VGND 0.01938f
C13540 XThR.Tn[0].n52 VGND 0.04813f
C13541 XThR.Tn[0].t43 VGND 0.0184f
C13542 XThR.Tn[0].t69 VGND 0.01938f
C13543 XThR.Tn[0].n53 VGND 0.04811f
C13544 XThR.Tn[0].n54 VGND 0.037f
C13545 XThR.Tn[0].n55 VGND 0.00705f
C13546 XThR.Tn[0].n56 VGND 0.11044f
C13547 XThR.Tn[0].t44 VGND 0.0184f
C13548 XThR.Tn[0].t49 VGND 0.01938f
C13549 XThR.Tn[0].n57 VGND 0.04813f
C13550 XThR.Tn[0].t18 VGND 0.0184f
C13551 XThR.Tn[0].t25 VGND 0.01938f
C13552 XThR.Tn[0].n58 VGND 0.04811f
C13553 XThR.Tn[0].n59 VGND 0.037f
C13554 XThR.Tn[0].n60 VGND 0.00705f
C13555 XThR.Tn[0].n61 VGND 0.11044f
C13556 XThR.Tn[0].t17 VGND 0.0184f
C13557 XThR.Tn[0].t27 VGND 0.01938f
C13558 XThR.Tn[0].n62 VGND 0.04813f
C13559 XThR.Tn[0].t56 VGND 0.0184f
C13560 XThR.Tn[0].t61 VGND 0.01938f
C13561 XThR.Tn[0].n63 VGND 0.04811f
C13562 XThR.Tn[0].n64 VGND 0.037f
C13563 XThR.Tn[0].n65 VGND 0.00705f
C13564 XThR.Tn[0].n66 VGND 0.11044f
C13565 XThR.Tn[0].t34 VGND 0.0184f
C13566 XThR.Tn[0].t59 VGND 0.01938f
C13567 XThR.Tn[0].n67 VGND 0.04813f
C13568 XThR.Tn[0].t72 VGND 0.0184f
C13569 XThR.Tn[0].t36 VGND 0.01938f
C13570 XThR.Tn[0].n68 VGND 0.04811f
C13571 XThR.Tn[0].n69 VGND 0.037f
C13572 XThR.Tn[0].n70 VGND 0.00705f
C13573 XThR.Tn[0].n71 VGND 0.11044f
C13574 XThR.Tn[0].t66 VGND 0.0184f
C13575 XThR.Tn[0].t16 VGND 0.01938f
C13576 XThR.Tn[0].n72 VGND 0.04813f
C13577 XThR.Tn[0].t42 VGND 0.0184f
C13578 XThR.Tn[0].t54 VGND 0.01938f
C13579 XThR.Tn[0].n73 VGND 0.04811f
C13580 XThR.Tn[0].n74 VGND 0.037f
C13581 XThR.Tn[0].n75 VGND 0.00705f
C13582 XThR.Tn[0].n76 VGND 0.11044f
C13583 XThR.Tn[0].t21 VGND 0.0184f
C13584 XThR.Tn[0].t33 VGND 0.01938f
C13585 XThR.Tn[0].n77 VGND 0.04813f
C13586 XThR.Tn[0].t60 VGND 0.0184f
C13587 XThR.Tn[0].t71 VGND 0.01938f
C13588 XThR.Tn[0].n78 VGND 0.04811f
C13589 XThR.Tn[0].n79 VGND 0.037f
C13590 XThR.Tn[0].n80 VGND 0.00705f
C13591 XThR.Tn[0].n81 VGND 0.11044f
C13592 XThR.Tn[0].t45 VGND 0.0184f
C13593 XThR.Tn[0].t28 VGND 0.01938f
C13594 XThR.Tn[0].n82 VGND 0.04813f
C13595 XThR.Tn[0].t19 VGND 0.0184f
C13596 XThR.Tn[0].t62 VGND 0.01938f
C13597 XThR.Tn[0].n83 VGND 0.04811f
C13598 XThR.Tn[0].n84 VGND 0.037f
C13599 XThR.Tn[0].n85 VGND 0.00705f
C13600 XThR.Tn[0].n86 VGND 0.11044f
C13601 XThR.Tn[0].n87 VGND 0.10088f
C13602 XThR.Tn[0].n88 VGND 0.28884f
C13603 XThC.Tn[2].t7 VGND 0.01791f
C13604 XThC.Tn[2].t6 VGND 0.01791f
C13605 XThC.Tn[2].n0 VGND 0.03615f
C13606 XThC.Tn[2].t5 VGND 0.01791f
C13607 XThC.Tn[2].t4 VGND 0.01791f
C13608 XThC.Tn[2].n1 VGND 0.0423f
C13609 XThC.Tn[2].n2 VGND 0.11841f
C13610 XThC.Tn[2].t11 VGND 0.01164f
C13611 XThC.Tn[2].t10 VGND 0.01164f
C13612 XThC.Tn[2].n3 VGND 0.02651f
C13613 XThC.Tn[2].t9 VGND 0.01164f
C13614 XThC.Tn[2].t8 VGND 0.01164f
C13615 XThC.Tn[2].n4 VGND 0.02651f
C13616 XThC.Tn[2].t1 VGND 0.01164f
C13617 XThC.Tn[2].t2 VGND 0.01164f
C13618 XThC.Tn[2].n5 VGND 0.02651f
C13619 XThC.Tn[2].t3 VGND 0.01164f
C13620 XThC.Tn[2].t0 VGND 0.01164f
C13621 XThC.Tn[2].n6 VGND 0.04417f
C13622 XThC.Tn[2].n7 VGND 0.12625f
C13623 XThC.Tn[2].n8 VGND 0.07804f
C13624 XThC.Tn[2].n9 VGND 0.08808f
C13625 XThC.Tn[2].t33 VGND 0.01455f
C13626 XThC.Tn[2].t38 VGND 0.01533f
C13627 XThC.Tn[2].n10 VGND 0.03807f
C13628 XThC.Tn[2].n11 VGND 0.02371f
C13629 XThC.Tn[2].n12 VGND 0.07683f
C13630 XThC.Tn[2].t42 VGND 0.01455f
C13631 XThC.Tn[2].t15 VGND 0.01533f
C13632 XThC.Tn[2].n13 VGND 0.03807f
C13633 XThC.Tn[2].n14 VGND 0.02371f
C13634 XThC.Tn[2].n15 VGND 0.07704f
C13635 XThC.Tn[2].n16 VGND 0.12863f
C13636 XThC.Tn[2].t22 VGND 0.01455f
C13637 XThC.Tn[2].t28 VGND 0.01533f
C13638 XThC.Tn[2].n17 VGND 0.03807f
C13639 XThC.Tn[2].n18 VGND 0.02371f
C13640 XThC.Tn[2].n19 VGND 0.07704f
C13641 XThC.Tn[2].n20 VGND 0.12863f
C13642 XThC.Tn[2].t24 VGND 0.01455f
C13643 XThC.Tn[2].t30 VGND 0.01533f
C13644 XThC.Tn[2].n21 VGND 0.03807f
C13645 XThC.Tn[2].n22 VGND 0.02371f
C13646 XThC.Tn[2].n23 VGND 0.07704f
C13647 XThC.Tn[2].n24 VGND 0.12863f
C13648 XThC.Tn[2].t35 VGND 0.01455f
C13649 XThC.Tn[2].t39 VGND 0.01533f
C13650 XThC.Tn[2].n25 VGND 0.03807f
C13651 XThC.Tn[2].n26 VGND 0.02371f
C13652 XThC.Tn[2].n27 VGND 0.07704f
C13653 XThC.Tn[2].n28 VGND 0.12863f
C13654 XThC.Tn[2].t13 VGND 0.01455f
C13655 XThC.Tn[2].t18 VGND 0.01533f
C13656 XThC.Tn[2].n29 VGND 0.03807f
C13657 XThC.Tn[2].n30 VGND 0.02371f
C13658 XThC.Tn[2].n31 VGND 0.07704f
C13659 XThC.Tn[2].n32 VGND 0.12863f
C13660 XThC.Tn[2].t25 VGND 0.01455f
C13661 XThC.Tn[2].t31 VGND 0.01533f
C13662 XThC.Tn[2].n33 VGND 0.03807f
C13663 XThC.Tn[2].n34 VGND 0.02371f
C13664 XThC.Tn[2].n35 VGND 0.07704f
C13665 XThC.Tn[2].n36 VGND 0.12863f
C13666 XThC.Tn[2].t36 VGND 0.01455f
C13667 XThC.Tn[2].t41 VGND 0.01533f
C13668 XThC.Tn[2].n37 VGND 0.03807f
C13669 XThC.Tn[2].n38 VGND 0.02371f
C13670 XThC.Tn[2].n39 VGND 0.07704f
C13671 XThC.Tn[2].n40 VGND 0.12863f
C13672 XThC.Tn[2].t37 VGND 0.01455f
C13673 XThC.Tn[2].t43 VGND 0.01533f
C13674 XThC.Tn[2].n41 VGND 0.03807f
C13675 XThC.Tn[2].n42 VGND 0.02371f
C13676 XThC.Tn[2].n43 VGND 0.07704f
C13677 XThC.Tn[2].n44 VGND 0.12863f
C13678 XThC.Tn[2].t14 VGND 0.01455f
C13679 XThC.Tn[2].t20 VGND 0.01533f
C13680 XThC.Tn[2].n45 VGND 0.03807f
C13681 XThC.Tn[2].n46 VGND 0.02371f
C13682 XThC.Tn[2].n47 VGND 0.07704f
C13683 XThC.Tn[2].n48 VGND 0.12863f
C13684 XThC.Tn[2].t27 VGND 0.01455f
C13685 XThC.Tn[2].t32 VGND 0.01533f
C13686 XThC.Tn[2].n49 VGND 0.03807f
C13687 XThC.Tn[2].n50 VGND 0.02371f
C13688 XThC.Tn[2].n51 VGND 0.07704f
C13689 XThC.Tn[2].n52 VGND 0.12863f
C13690 XThC.Tn[2].t29 VGND 0.01455f
C13691 XThC.Tn[2].t34 VGND 0.01533f
C13692 XThC.Tn[2].n53 VGND 0.03807f
C13693 XThC.Tn[2].n54 VGND 0.02371f
C13694 XThC.Tn[2].n55 VGND 0.07704f
C13695 XThC.Tn[2].n56 VGND 0.12863f
C13696 XThC.Tn[2].t16 VGND 0.01455f
C13697 XThC.Tn[2].t21 VGND 0.01533f
C13698 XThC.Tn[2].n57 VGND 0.03807f
C13699 XThC.Tn[2].n58 VGND 0.02371f
C13700 XThC.Tn[2].n59 VGND 0.07704f
C13701 XThC.Tn[2].n60 VGND 0.12863f
C13702 XThC.Tn[2].t17 VGND 0.01455f
C13703 XThC.Tn[2].t23 VGND 0.01533f
C13704 XThC.Tn[2].n61 VGND 0.03807f
C13705 XThC.Tn[2].n62 VGND 0.02371f
C13706 XThC.Tn[2].n63 VGND 0.07704f
C13707 XThC.Tn[2].n64 VGND 0.12863f
C13708 XThC.Tn[2].t19 VGND 0.01455f
C13709 XThC.Tn[2].t26 VGND 0.01533f
C13710 XThC.Tn[2].n65 VGND 0.03807f
C13711 XThC.Tn[2].n66 VGND 0.02371f
C13712 XThC.Tn[2].n67 VGND 0.07704f
C13713 XThC.Tn[2].n68 VGND 0.12863f
C13714 XThC.Tn[2].t40 VGND 0.01455f
C13715 XThC.Tn[2].t12 VGND 0.01533f
C13716 XThC.Tn[2].n69 VGND 0.03807f
C13717 XThC.Tn[2].n70 VGND 0.02371f
C13718 XThC.Tn[2].n71 VGND 0.07704f
C13719 XThC.Tn[2].n72 VGND 0.12863f
C13720 XThC.Tn[2].n73 VGND 0.49783f
C13721 XThC.Tn[2].n74 VGND 0.10557f
C13722 XThC.Tn[2].n75 VGND 0.03748f
C13723 XThR.Tn[5].t8 VGND 0.01523f
C13724 XThR.Tn[5].t9 VGND 0.01523f
C13725 XThR.Tn[5].n0 VGND 0.05778f
C13726 XThR.Tn[5].t11 VGND 0.01523f
C13727 XThR.Tn[5].t10 VGND 0.01523f
C13728 XThR.Tn[5].n1 VGND 0.03468f
C13729 XThR.Tn[5].n2 VGND 0.16515f
C13730 XThR.Tn[5].t6 VGND 0.01523f
C13731 XThR.Tn[5].t5 VGND 0.01523f
C13732 XThR.Tn[5].n3 VGND 0.03468f
C13733 XThR.Tn[5].n4 VGND 0.10209f
C13734 XThR.Tn[5].t7 VGND 0.01523f
C13735 XThR.Tn[5].t4 VGND 0.01523f
C13736 XThR.Tn[5].n5 VGND 0.03468f
C13737 XThR.Tn[5].n6 VGND 0.11522f
C13738 XThR.Tn[5].t42 VGND 0.01904f
C13739 XThR.Tn[5].t70 VGND 0.02005f
C13740 XThR.Tn[5].n7 VGND 0.04979f
C13741 XThR.Tn[5].n8 VGND 0.09257f
C13742 XThR.Tn[5].t20 VGND 0.01904f
C13743 XThR.Tn[5].t24 VGND 0.02005f
C13744 XThR.Tn[5].n9 VGND 0.04979f
C13745 XThR.Tn[5].t59 VGND 0.01904f
C13746 XThR.Tn[5].t66 VGND 0.02005f
C13747 XThR.Tn[5].n10 VGND 0.04978f
C13748 XThR.Tn[5].n11 VGND 0.03828f
C13749 XThR.Tn[5].n12 VGND 0.0073f
C13750 XThR.Tn[5].n13 VGND 0.11426f
C13751 XThR.Tn[5].t34 VGND 0.01904f
C13752 XThR.Tn[5].t64 VGND 0.02005f
C13753 XThR.Tn[5].n14 VGND 0.04979f
C13754 XThR.Tn[5].t13 VGND 0.01904f
C13755 XThR.Tn[5].t41 VGND 0.02005f
C13756 XThR.Tn[5].n15 VGND 0.04978f
C13757 XThR.Tn[5].n16 VGND 0.03828f
C13758 XThR.Tn[5].n17 VGND 0.0073f
C13759 XThR.Tn[5].n18 VGND 0.11426f
C13760 XThR.Tn[5].t72 VGND 0.01904f
C13761 XThR.Tn[5].t19 VGND 0.02005f
C13762 XThR.Tn[5].n19 VGND 0.04979f
C13763 XThR.Tn[5].t52 VGND 0.01904f
C13764 XThR.Tn[5].t58 VGND 0.02005f
C13765 XThR.Tn[5].n20 VGND 0.04978f
C13766 XThR.Tn[5].n21 VGND 0.03828f
C13767 XThR.Tn[5].n22 VGND 0.0073f
C13768 XThR.Tn[5].n23 VGND 0.11426f
C13769 XThR.Tn[5].t36 VGND 0.01904f
C13770 XThR.Tn[5].t49 VGND 0.02005f
C13771 XThR.Tn[5].n24 VGND 0.04979f
C13772 XThR.Tn[5].t15 VGND 0.01904f
C13773 XThR.Tn[5].t27 VGND 0.02005f
C13774 XThR.Tn[5].n25 VGND 0.04978f
C13775 XThR.Tn[5].n26 VGND 0.03828f
C13776 XThR.Tn[5].n27 VGND 0.0073f
C13777 XThR.Tn[5].n28 VGND 0.11426f
C13778 XThR.Tn[5].t53 VGND 0.01904f
C13779 XThR.Tn[5].t21 VGND 0.02005f
C13780 XThR.Tn[5].n29 VGND 0.04979f
C13781 XThR.Tn[5].t32 VGND 0.01904f
C13782 XThR.Tn[5].t61 VGND 0.02005f
C13783 XThR.Tn[5].n30 VGND 0.04978f
C13784 XThR.Tn[5].n31 VGND 0.03828f
C13785 XThR.Tn[5].n32 VGND 0.0073f
C13786 XThR.Tn[5].n33 VGND 0.11426f
C13787 XThR.Tn[5].t48 VGND 0.01904f
C13788 XThR.Tn[5].t35 VGND 0.02005f
C13789 XThR.Tn[5].n34 VGND 0.04979f
C13790 XThR.Tn[5].t26 VGND 0.01904f
C13791 XThR.Tn[5].t14 VGND 0.02005f
C13792 XThR.Tn[5].n35 VGND 0.04978f
C13793 XThR.Tn[5].n36 VGND 0.03828f
C13794 XThR.Tn[5].n37 VGND 0.0073f
C13795 XThR.Tn[5].n38 VGND 0.11426f
C13796 XThR.Tn[5].t67 VGND 0.01904f
C13797 XThR.Tn[5].t30 VGND 0.02005f
C13798 XThR.Tn[5].n39 VGND 0.04979f
C13799 XThR.Tn[5].t44 VGND 0.01904f
C13800 XThR.Tn[5].t71 VGND 0.02005f
C13801 XThR.Tn[5].n40 VGND 0.04978f
C13802 XThR.Tn[5].n41 VGND 0.03828f
C13803 XThR.Tn[5].n42 VGND 0.0073f
C13804 XThR.Tn[5].n43 VGND 0.11426f
C13805 XThR.Tn[5].t23 VGND 0.01904f
C13806 XThR.Tn[5].t47 VGND 0.02005f
C13807 XThR.Tn[5].n44 VGND 0.04979f
C13808 XThR.Tn[5].t63 VGND 0.01904f
C13809 XThR.Tn[5].t25 VGND 0.02005f
C13810 XThR.Tn[5].n45 VGND 0.04978f
C13811 XThR.Tn[5].n46 VGND 0.03828f
C13812 XThR.Tn[5].n47 VGND 0.0073f
C13813 XThR.Tn[5].n48 VGND 0.11426f
C13814 XThR.Tn[5].t40 VGND 0.01904f
C13815 XThR.Tn[5].t65 VGND 0.02005f
C13816 XThR.Tn[5].n49 VGND 0.04979f
C13817 XThR.Tn[5].t18 VGND 0.01904f
C13818 XThR.Tn[5].t43 VGND 0.02005f
C13819 XThR.Tn[5].n50 VGND 0.04978f
C13820 XThR.Tn[5].n51 VGND 0.03828f
C13821 XThR.Tn[5].n52 VGND 0.0073f
C13822 XThR.Tn[5].n53 VGND 0.11426f
C13823 XThR.Tn[5].t12 VGND 0.01904f
C13824 XThR.Tn[5].t22 VGND 0.02005f
C13825 XThR.Tn[5].n54 VGND 0.04979f
C13826 XThR.Tn[5].t55 VGND 0.01904f
C13827 XThR.Tn[5].t62 VGND 0.02005f
C13828 XThR.Tn[5].n55 VGND 0.04978f
C13829 XThR.Tn[5].n56 VGND 0.03828f
C13830 XThR.Tn[5].n57 VGND 0.0073f
C13831 XThR.Tn[5].n58 VGND 0.11426f
C13832 XThR.Tn[5].t51 VGND 0.01904f
C13833 XThR.Tn[5].t57 VGND 0.02005f
C13834 XThR.Tn[5].n59 VGND 0.04979f
C13835 XThR.Tn[5].t29 VGND 0.01904f
C13836 XThR.Tn[5].t37 VGND 0.02005f
C13837 XThR.Tn[5].n60 VGND 0.04978f
C13838 XThR.Tn[5].n61 VGND 0.03828f
C13839 XThR.Tn[5].n62 VGND 0.0073f
C13840 XThR.Tn[5].n63 VGND 0.11426f
C13841 XThR.Tn[5].t69 VGND 0.01904f
C13842 XThR.Tn[5].t31 VGND 0.02005f
C13843 XThR.Tn[5].n64 VGND 0.04979f
C13844 XThR.Tn[5].t46 VGND 0.01904f
C13845 XThR.Tn[5].t73 VGND 0.02005f
C13846 XThR.Tn[5].n65 VGND 0.04978f
C13847 XThR.Tn[5].n66 VGND 0.03828f
C13848 XThR.Tn[5].n67 VGND 0.0073f
C13849 XThR.Tn[5].n68 VGND 0.11426f
C13850 XThR.Tn[5].t38 VGND 0.01904f
C13851 XThR.Tn[5].t50 VGND 0.02005f
C13852 XThR.Tn[5].n69 VGND 0.04979f
C13853 XThR.Tn[5].t17 VGND 0.01904f
C13854 XThR.Tn[5].t28 VGND 0.02005f
C13855 XThR.Tn[5].n70 VGND 0.04978f
C13856 XThR.Tn[5].n71 VGND 0.03828f
C13857 XThR.Tn[5].n72 VGND 0.0073f
C13858 XThR.Tn[5].n73 VGND 0.11426f
C13859 XThR.Tn[5].t54 VGND 0.01904f
C13860 XThR.Tn[5].t68 VGND 0.02005f
C13861 XThR.Tn[5].n74 VGND 0.04979f
C13862 XThR.Tn[5].t33 VGND 0.01904f
C13863 XThR.Tn[5].t45 VGND 0.02005f
C13864 XThR.Tn[5].n75 VGND 0.04978f
C13865 XThR.Tn[5].n76 VGND 0.03828f
C13866 XThR.Tn[5].n77 VGND 0.0073f
C13867 XThR.Tn[5].n78 VGND 0.11426f
C13868 XThR.Tn[5].t16 VGND 0.01904f
C13869 XThR.Tn[5].t60 VGND 0.02005f
C13870 XThR.Tn[5].n79 VGND 0.04979f
C13871 XThR.Tn[5].t56 VGND 0.01904f
C13872 XThR.Tn[5].t39 VGND 0.02005f
C13873 XThR.Tn[5].n80 VGND 0.04978f
C13874 XThR.Tn[5].n81 VGND 0.03828f
C13875 XThR.Tn[5].n82 VGND 0.0073f
C13876 XThR.Tn[5].n83 VGND 0.11426f
C13877 XThR.Tn[5].n84 VGND 0.10437f
C13878 XThR.Tn[5].n85 VGND 0.20213f
C13879 XThR.Tn[5].t2 VGND 0.02343f
C13880 XThR.Tn[5].t3 VGND 0.02343f
C13881 XThR.Tn[5].n86 VGND 0.04729f
C13882 XThR.Tn[5].t1 VGND 0.02343f
C13883 XThR.Tn[5].t0 VGND 0.02343f
C13884 XThR.Tn[5].n87 VGND 0.05533f
C13885 XThR.Tn[5].n88 VGND 0.1549f
C13886 XThR.Tn[5].n89 VGND 0.04903f
C13887 XThC.XTB4.Y.t4 VGND 0.02956f
C13888 XThC.XTB4.Y.t13 VGND 0.05016f
C13889 XThC.XTB4.Y.n0 VGND 0.05972f
C13890 XThC.XTB4.Y.t7 VGND 0.02956f
C13891 XThC.XTB4.Y.t17 VGND 0.05016f
C13892 XThC.XTB4.Y.n1 VGND 0.03074f
C13893 XThC.XTB4.Y.t10 VGND 0.02956f
C13894 XThC.XTB4.Y.t2 VGND 0.05016f
C13895 XThC.XTB4.Y.n2 VGND 0.06603f
C13896 XThC.XTB4.Y.t14 VGND 0.02956f
C13897 XThC.XTB4.Y.t3 VGND 0.05016f
C13898 XThC.XTB4.Y.n3 VGND 0.0613f
C13899 XThC.XTB4.Y.n4 VGND 0.03729f
C13900 XThC.XTB4.Y.n5 VGND 0.06174f
C13901 XThC.XTB4.Y.n6 VGND 0.02389f
C13902 XThC.XTB4.Y.n7 VGND 0.02916f
C13903 XThC.XTB4.Y.n8 VGND 0.06603f
C13904 XThC.XTB4.Y.n9 VGND 0.0331f
C13905 XThC.XTB4.Y.n10 VGND 0.06459f
C13906 XThC.XTB4.Y.t5 VGND 0.02956f
C13907 XThC.XTB4.Y.t16 VGND 0.05016f
C13908 XThC.XTB4.Y.n11 VGND 0.06761f
C13909 XThC.XTB4.Y.t9 VGND 0.02956f
C13910 XThC.XTB4.Y.t6 VGND 0.05016f
C13911 XThC.XTB4.Y.t15 VGND 0.02956f
C13912 XThC.XTB4.Y.t12 VGND 0.05016f
C13913 XThC.XTB4.Y.t11 VGND 0.02956f
C13914 XThC.XTB4.Y.t8 VGND 0.05016f
C13915 XThC.XTB4.Y.n12 VGND 0.08416f
C13916 XThC.XTB4.Y.n13 VGND 0.08889f
C13917 XThC.XTB4.Y.n14 VGND 0.03426f
C13918 XThC.XTB4.Y.n15 VGND 0.07234f
C13919 XThC.XTB4.Y.n16 VGND 0.0331f
C13920 XThC.XTB4.Y.n17 VGND 0.02701f
C13921 XThC.XTB4.Y.n18 VGND 0.63971f
C13922 XThC.XTB4.Y.n19 VGND 1.30917f
C13923 XThC.XTB4.Y.t1 VGND 0.06491f
C13924 XThC.XTB4.Y.n20 VGND 0.11223f
C13925 XThC.XTB4.Y.t0 VGND 0.12238f
C13926 XThC.XTB4.Y.n21 VGND 0.16166f
C13927 XThC.Tn[0].t8 VGND 0.01203f
C13928 XThC.Tn[0].t7 VGND 0.01203f
C13929 XThC.Tn[0].n0 VGND 0.02429f
C13930 XThC.Tn[0].t10 VGND 0.01203f
C13931 XThC.Tn[0].t9 VGND 0.01203f
C13932 XThC.Tn[0].n1 VGND 0.02842f
C13933 XThC.Tn[0].n2 VGND 0.07955f
C13934 XThC.Tn[0].t4 VGND 0.00782f
C13935 XThC.Tn[0].t3 VGND 0.00782f
C13936 XThC.Tn[0].n3 VGND 0.01781f
C13937 XThC.Tn[0].t6 VGND 0.00782f
C13938 XThC.Tn[0].t5 VGND 0.00782f
C13939 XThC.Tn[0].n4 VGND 0.01781f
C13940 XThC.Tn[0].t1 VGND 0.00782f
C13941 XThC.Tn[0].t2 VGND 0.00782f
C13942 XThC.Tn[0].n5 VGND 0.01781f
C13943 XThC.Tn[0].t11 VGND 0.00782f
C13944 XThC.Tn[0].t0 VGND 0.00782f
C13945 XThC.Tn[0].n6 VGND 0.02968f
C13946 XThC.Tn[0].n7 VGND 0.08482f
C13947 XThC.Tn[0].n8 VGND 0.05243f
C13948 XThC.Tn[0].n9 VGND 0.05917f
C13949 XThC.Tn[0].t22 VGND 0.00978f
C13950 XThC.Tn[0].t12 VGND 0.0103f
C13951 XThC.Tn[0].n10 VGND 0.02557f
C13952 XThC.Tn[0].n11 VGND 0.01593f
C13953 XThC.Tn[0].n12 VGND 0.05162f
C13954 XThC.Tn[0].t31 VGND 0.00978f
C13955 XThC.Tn[0].t21 VGND 0.0103f
C13956 XThC.Tn[0].n13 VGND 0.02557f
C13957 XThC.Tn[0].n14 VGND 0.01593f
C13958 XThC.Tn[0].n15 VGND 0.05176f
C13959 XThC.Tn[0].n16 VGND 0.08642f
C13960 XThC.Tn[0].t43 VGND 0.00978f
C13961 XThC.Tn[0].t33 VGND 0.0103f
C13962 XThC.Tn[0].n17 VGND 0.02557f
C13963 XThC.Tn[0].n18 VGND 0.01593f
C13964 XThC.Tn[0].n19 VGND 0.05176f
C13965 XThC.Tn[0].n20 VGND 0.08642f
C13966 XThC.Tn[0].t13 VGND 0.00978f
C13967 XThC.Tn[0].t35 VGND 0.0103f
C13968 XThC.Tn[0].n21 VGND 0.02557f
C13969 XThC.Tn[0].n22 VGND 0.01593f
C13970 XThC.Tn[0].n23 VGND 0.05176f
C13971 XThC.Tn[0].n24 VGND 0.08642f
C13972 XThC.Tn[0].t23 VGND 0.00978f
C13973 XThC.Tn[0].t15 VGND 0.0103f
C13974 XThC.Tn[0].n25 VGND 0.02557f
C13975 XThC.Tn[0].n26 VGND 0.01593f
C13976 XThC.Tn[0].n27 VGND 0.05176f
C13977 XThC.Tn[0].n28 VGND 0.08642f
C13978 XThC.Tn[0].t34 VGND 0.00978f
C13979 XThC.Tn[0].t25 VGND 0.0103f
C13980 XThC.Tn[0].n29 VGND 0.02557f
C13981 XThC.Tn[0].n30 VGND 0.01593f
C13982 XThC.Tn[0].n31 VGND 0.05176f
C13983 XThC.Tn[0].n32 VGND 0.08642f
C13984 XThC.Tn[0].t14 VGND 0.00978f
C13985 XThC.Tn[0].t36 VGND 0.0103f
C13986 XThC.Tn[0].n33 VGND 0.02557f
C13987 XThC.Tn[0].n34 VGND 0.01593f
C13988 XThC.Tn[0].n35 VGND 0.05176f
C13989 XThC.Tn[0].n36 VGND 0.08642f
C13990 XThC.Tn[0].t24 VGND 0.00978f
C13991 XThC.Tn[0].t16 VGND 0.0103f
C13992 XThC.Tn[0].n37 VGND 0.02557f
C13993 XThC.Tn[0].n38 VGND 0.01593f
C13994 XThC.Tn[0].n39 VGND 0.05176f
C13995 XThC.Tn[0].n40 VGND 0.08642f
C13996 XThC.Tn[0].t27 VGND 0.00978f
C13997 XThC.Tn[0].t18 VGND 0.0103f
C13998 XThC.Tn[0].n41 VGND 0.02557f
C13999 XThC.Tn[0].n42 VGND 0.01593f
C14000 XThC.Tn[0].n43 VGND 0.05176f
C14001 XThC.Tn[0].n44 VGND 0.08642f
C14002 XThC.Tn[0].t37 VGND 0.00978f
C14003 XThC.Tn[0].t26 VGND 0.0103f
C14004 XThC.Tn[0].n45 VGND 0.02557f
C14005 XThC.Tn[0].n46 VGND 0.01593f
C14006 XThC.Tn[0].n47 VGND 0.05176f
C14007 XThC.Tn[0].n48 VGND 0.08642f
C14008 XThC.Tn[0].t17 VGND 0.00978f
C14009 XThC.Tn[0].t39 VGND 0.0103f
C14010 XThC.Tn[0].n49 VGND 0.02557f
C14011 XThC.Tn[0].n50 VGND 0.01593f
C14012 XThC.Tn[0].n51 VGND 0.05176f
C14013 XThC.Tn[0].n52 VGND 0.08642f
C14014 XThC.Tn[0].t19 VGND 0.00978f
C14015 XThC.Tn[0].t41 VGND 0.0103f
C14016 XThC.Tn[0].n53 VGND 0.02557f
C14017 XThC.Tn[0].n54 VGND 0.01593f
C14018 XThC.Tn[0].n55 VGND 0.05176f
C14019 XThC.Tn[0].n56 VGND 0.08642f
C14020 XThC.Tn[0].t38 VGND 0.00978f
C14021 XThC.Tn[0].t28 VGND 0.0103f
C14022 XThC.Tn[0].n57 VGND 0.02557f
C14023 XThC.Tn[0].n58 VGND 0.01593f
C14024 XThC.Tn[0].n59 VGND 0.05176f
C14025 XThC.Tn[0].n60 VGND 0.08642f
C14026 XThC.Tn[0].t40 VGND 0.00978f
C14027 XThC.Tn[0].t30 VGND 0.0103f
C14028 XThC.Tn[0].n61 VGND 0.02557f
C14029 XThC.Tn[0].n62 VGND 0.01593f
C14030 XThC.Tn[0].n63 VGND 0.05176f
C14031 XThC.Tn[0].n64 VGND 0.08642f
C14032 XThC.Tn[0].t42 VGND 0.00978f
C14033 XThC.Tn[0].t32 VGND 0.0103f
C14034 XThC.Tn[0].n65 VGND 0.02557f
C14035 XThC.Tn[0].n66 VGND 0.01593f
C14036 XThC.Tn[0].n67 VGND 0.05176f
C14037 XThC.Tn[0].n68 VGND 0.08642f
C14038 XThC.Tn[0].t29 VGND 0.00978f
C14039 XThC.Tn[0].t20 VGND 0.0103f
C14040 XThC.Tn[0].n69 VGND 0.02557f
C14041 XThC.Tn[0].n70 VGND 0.01593f
C14042 XThC.Tn[0].n71 VGND 0.05176f
C14043 XThC.Tn[0].n72 VGND 0.08642f
C14044 XThC.Tn[0].n73 VGND 0.53416f
C14045 XThC.Tn[0].n74 VGND 0.06476f
C14046 XThC.Tn[0].n75 VGND 0.02518f
C14047 XThC.Tn[1].t7 VGND 0.01728f
C14048 XThC.Tn[1].t6 VGND 0.01728f
C14049 XThC.Tn[1].n0 VGND 0.03487f
C14050 XThC.Tn[1].t5 VGND 0.01728f
C14051 XThC.Tn[1].t4 VGND 0.01728f
C14052 XThC.Tn[1].n1 VGND 0.0408f
C14053 XThC.Tn[1].n2 VGND 0.12239f
C14054 XThC.Tn[1].t9 VGND 0.01123f
C14055 XThC.Tn[1].t8 VGND 0.01123f
C14056 XThC.Tn[1].n3 VGND 0.02557f
C14057 XThC.Tn[1].t11 VGND 0.01123f
C14058 XThC.Tn[1].t10 VGND 0.01123f
C14059 XThC.Tn[1].n4 VGND 0.02557f
C14060 XThC.Tn[1].t1 VGND 0.01123f
C14061 XThC.Tn[1].t0 VGND 0.01123f
C14062 XThC.Tn[1].n5 VGND 0.02557f
C14063 XThC.Tn[1].t3 VGND 0.01123f
C14064 XThC.Tn[1].t2 VGND 0.01123f
C14065 XThC.Tn[1].n6 VGND 0.04261f
C14066 XThC.Tn[1].n7 VGND 0.12178f
C14067 XThC.Tn[1].n8 VGND 0.07528f
C14068 XThC.Tn[1].n9 VGND 0.08496f
C14069 XThC.Tn[1].t41 VGND 0.01404f
C14070 XThC.Tn[1].t14 VGND 0.01478f
C14071 XThC.Tn[1].n10 VGND 0.03672f
C14072 XThC.Tn[1].n11 VGND 0.02288f
C14073 XThC.Tn[1].n12 VGND 0.07411f
C14074 XThC.Tn[1].t18 VGND 0.01404f
C14075 XThC.Tn[1].t23 VGND 0.01478f
C14076 XThC.Tn[1].n13 VGND 0.03672f
C14077 XThC.Tn[1].n14 VGND 0.02288f
C14078 XThC.Tn[1].n15 VGND 0.07432f
C14079 XThC.Tn[1].n16 VGND 0.12408f
C14080 XThC.Tn[1].t30 VGND 0.01404f
C14081 XThC.Tn[1].t36 VGND 0.01478f
C14082 XThC.Tn[1].n17 VGND 0.03672f
C14083 XThC.Tn[1].n18 VGND 0.02288f
C14084 XThC.Tn[1].n19 VGND 0.07432f
C14085 XThC.Tn[1].n20 VGND 0.12408f
C14086 XThC.Tn[1].t32 VGND 0.01404f
C14087 XThC.Tn[1].t38 VGND 0.01478f
C14088 XThC.Tn[1].n21 VGND 0.03672f
C14089 XThC.Tn[1].n22 VGND 0.02288f
C14090 XThC.Tn[1].n23 VGND 0.07432f
C14091 XThC.Tn[1].n24 VGND 0.12408f
C14092 XThC.Tn[1].t43 VGND 0.01404f
C14093 XThC.Tn[1].t15 VGND 0.01478f
C14094 XThC.Tn[1].n25 VGND 0.03672f
C14095 XThC.Tn[1].n26 VGND 0.02288f
C14096 XThC.Tn[1].n27 VGND 0.07432f
C14097 XThC.Tn[1].n28 VGND 0.12408f
C14098 XThC.Tn[1].t21 VGND 0.01404f
C14099 XThC.Tn[1].t26 VGND 0.01478f
C14100 XThC.Tn[1].n29 VGND 0.03672f
C14101 XThC.Tn[1].n30 VGND 0.02288f
C14102 XThC.Tn[1].n31 VGND 0.07432f
C14103 XThC.Tn[1].n32 VGND 0.12408f
C14104 XThC.Tn[1].t33 VGND 0.01404f
C14105 XThC.Tn[1].t39 VGND 0.01478f
C14106 XThC.Tn[1].n33 VGND 0.03672f
C14107 XThC.Tn[1].n34 VGND 0.02288f
C14108 XThC.Tn[1].n35 VGND 0.07432f
C14109 XThC.Tn[1].n36 VGND 0.12408f
C14110 XThC.Tn[1].t12 VGND 0.01404f
C14111 XThC.Tn[1].t17 VGND 0.01478f
C14112 XThC.Tn[1].n37 VGND 0.03672f
C14113 XThC.Tn[1].n38 VGND 0.02288f
C14114 XThC.Tn[1].n39 VGND 0.07432f
C14115 XThC.Tn[1].n40 VGND 0.12408f
C14116 XThC.Tn[1].t13 VGND 0.01404f
C14117 XThC.Tn[1].t19 VGND 0.01478f
C14118 XThC.Tn[1].n41 VGND 0.03672f
C14119 XThC.Tn[1].n42 VGND 0.02288f
C14120 XThC.Tn[1].n43 VGND 0.07432f
C14121 XThC.Tn[1].n44 VGND 0.12408f
C14122 XThC.Tn[1].t22 VGND 0.01404f
C14123 XThC.Tn[1].t28 VGND 0.01478f
C14124 XThC.Tn[1].n45 VGND 0.03672f
C14125 XThC.Tn[1].n46 VGND 0.02288f
C14126 XThC.Tn[1].n47 VGND 0.07432f
C14127 XThC.Tn[1].n48 VGND 0.12408f
C14128 XThC.Tn[1].t35 VGND 0.01404f
C14129 XThC.Tn[1].t40 VGND 0.01478f
C14130 XThC.Tn[1].n49 VGND 0.03672f
C14131 XThC.Tn[1].n50 VGND 0.02288f
C14132 XThC.Tn[1].n51 VGND 0.07432f
C14133 XThC.Tn[1].n52 VGND 0.12408f
C14134 XThC.Tn[1].t37 VGND 0.01404f
C14135 XThC.Tn[1].t42 VGND 0.01478f
C14136 XThC.Tn[1].n53 VGND 0.03672f
C14137 XThC.Tn[1].n54 VGND 0.02288f
C14138 XThC.Tn[1].n55 VGND 0.07432f
C14139 XThC.Tn[1].n56 VGND 0.12408f
C14140 XThC.Tn[1].t24 VGND 0.01404f
C14141 XThC.Tn[1].t29 VGND 0.01478f
C14142 XThC.Tn[1].n57 VGND 0.03672f
C14143 XThC.Tn[1].n58 VGND 0.02288f
C14144 XThC.Tn[1].n59 VGND 0.07432f
C14145 XThC.Tn[1].n60 VGND 0.12408f
C14146 XThC.Tn[1].t25 VGND 0.01404f
C14147 XThC.Tn[1].t31 VGND 0.01478f
C14148 XThC.Tn[1].n61 VGND 0.03672f
C14149 XThC.Tn[1].n62 VGND 0.02288f
C14150 XThC.Tn[1].n63 VGND 0.07432f
C14151 XThC.Tn[1].n64 VGND 0.12408f
C14152 XThC.Tn[1].t27 VGND 0.01404f
C14153 XThC.Tn[1].t34 VGND 0.01478f
C14154 XThC.Tn[1].n65 VGND 0.03672f
C14155 XThC.Tn[1].n66 VGND 0.02288f
C14156 XThC.Tn[1].n67 VGND 0.07432f
C14157 XThC.Tn[1].n68 VGND 0.12408f
C14158 XThC.Tn[1].t16 VGND 0.01404f
C14159 XThC.Tn[1].t20 VGND 0.01478f
C14160 XThC.Tn[1].n69 VGND 0.03672f
C14161 XThC.Tn[1].n70 VGND 0.02288f
C14162 XThC.Tn[1].n71 VGND 0.07432f
C14163 XThC.Tn[1].n72 VGND 0.12408f
C14164 XThC.Tn[1].n73 VGND 0.63052f
C14165 XThC.Tn[1].n74 VGND 0.11981f
C14166 XThC.Tn[12].t7 VGND 0.01277f
C14167 XThC.Tn[12].t6 VGND 0.01277f
C14168 XThC.Tn[12].n0 VGND 0.03186f
C14169 XThC.Tn[12].t5 VGND 0.01277f
C14170 XThC.Tn[12].t4 VGND 0.01277f
C14171 XThC.Tn[12].n1 VGND 0.02555f
C14172 XThC.Tn[12].n2 VGND 0.06427f
C14173 XThC.Tn[12].t17 VGND 0.01597f
C14174 XThC.Tn[12].t22 VGND 0.01682f
C14175 XThC.Tn[12].n3 VGND 0.04177f
C14176 XThC.Tn[12].n4 VGND 0.02602f
C14177 XThC.Tn[12].n5 VGND 0.08431f
C14178 XThC.Tn[12].t26 VGND 0.01597f
C14179 XThC.Tn[12].t31 VGND 0.01682f
C14180 XThC.Tn[12].n6 VGND 0.04177f
C14181 XThC.Tn[12].n7 VGND 0.02602f
C14182 XThC.Tn[12].n8 VGND 0.08455f
C14183 XThC.Tn[12].n9 VGND 0.14116f
C14184 XThC.Tn[12].t38 VGND 0.01597f
C14185 XThC.Tn[12].t12 VGND 0.01682f
C14186 XThC.Tn[12].n10 VGND 0.04177f
C14187 XThC.Tn[12].n11 VGND 0.02602f
C14188 XThC.Tn[12].n12 VGND 0.08455f
C14189 XThC.Tn[12].n13 VGND 0.14116f
C14190 XThC.Tn[12].t40 VGND 0.01597f
C14191 XThC.Tn[12].t14 VGND 0.01682f
C14192 XThC.Tn[12].n14 VGND 0.04177f
C14193 XThC.Tn[12].n15 VGND 0.02602f
C14194 XThC.Tn[12].n16 VGND 0.08455f
C14195 XThC.Tn[12].n17 VGND 0.14116f
C14196 XThC.Tn[12].t19 VGND 0.01597f
C14197 XThC.Tn[12].t23 VGND 0.01682f
C14198 XThC.Tn[12].n18 VGND 0.04177f
C14199 XThC.Tn[12].n19 VGND 0.02602f
C14200 XThC.Tn[12].n20 VGND 0.08455f
C14201 XThC.Tn[12].n21 VGND 0.14116f
C14202 XThC.Tn[12].t29 VGND 0.01597f
C14203 XThC.Tn[12].t34 VGND 0.01682f
C14204 XThC.Tn[12].n22 VGND 0.04177f
C14205 XThC.Tn[12].n23 VGND 0.02602f
C14206 XThC.Tn[12].n24 VGND 0.08455f
C14207 XThC.Tn[12].n25 VGND 0.14116f
C14208 XThC.Tn[12].t41 VGND 0.01597f
C14209 XThC.Tn[12].t15 VGND 0.01682f
C14210 XThC.Tn[12].n26 VGND 0.04177f
C14211 XThC.Tn[12].n27 VGND 0.02602f
C14212 XThC.Tn[12].n28 VGND 0.08455f
C14213 XThC.Tn[12].n29 VGND 0.14116f
C14214 XThC.Tn[12].t20 VGND 0.01597f
C14215 XThC.Tn[12].t25 VGND 0.01682f
C14216 XThC.Tn[12].n30 VGND 0.04177f
C14217 XThC.Tn[12].n31 VGND 0.02602f
C14218 XThC.Tn[12].n32 VGND 0.08455f
C14219 XThC.Tn[12].n33 VGND 0.14116f
C14220 XThC.Tn[12].t21 VGND 0.01597f
C14221 XThC.Tn[12].t27 VGND 0.01682f
C14222 XThC.Tn[12].n34 VGND 0.04177f
C14223 XThC.Tn[12].n35 VGND 0.02602f
C14224 XThC.Tn[12].n36 VGND 0.08455f
C14225 XThC.Tn[12].n37 VGND 0.14116f
C14226 XThC.Tn[12].t30 VGND 0.01597f
C14227 XThC.Tn[12].t36 VGND 0.01682f
C14228 XThC.Tn[12].n38 VGND 0.04177f
C14229 XThC.Tn[12].n39 VGND 0.02602f
C14230 XThC.Tn[12].n40 VGND 0.08455f
C14231 XThC.Tn[12].n41 VGND 0.14116f
C14232 XThC.Tn[12].t43 VGND 0.01597f
C14233 XThC.Tn[12].t16 VGND 0.01682f
C14234 XThC.Tn[12].n42 VGND 0.04177f
C14235 XThC.Tn[12].n43 VGND 0.02602f
C14236 XThC.Tn[12].n44 VGND 0.08455f
C14237 XThC.Tn[12].n45 VGND 0.14116f
C14238 XThC.Tn[12].t13 VGND 0.01597f
C14239 XThC.Tn[12].t18 VGND 0.01682f
C14240 XThC.Tn[12].n46 VGND 0.04177f
C14241 XThC.Tn[12].n47 VGND 0.02602f
C14242 XThC.Tn[12].n48 VGND 0.08455f
C14243 XThC.Tn[12].n49 VGND 0.14116f
C14244 XThC.Tn[12].t32 VGND 0.01597f
C14245 XThC.Tn[12].t37 VGND 0.01682f
C14246 XThC.Tn[12].n50 VGND 0.04177f
C14247 XThC.Tn[12].n51 VGND 0.02602f
C14248 XThC.Tn[12].n52 VGND 0.08455f
C14249 XThC.Tn[12].n53 VGND 0.14116f
C14250 XThC.Tn[12].t33 VGND 0.01597f
C14251 XThC.Tn[12].t39 VGND 0.01682f
C14252 XThC.Tn[12].n54 VGND 0.04177f
C14253 XThC.Tn[12].n55 VGND 0.02602f
C14254 XThC.Tn[12].n56 VGND 0.08455f
C14255 XThC.Tn[12].n57 VGND 0.14116f
C14256 XThC.Tn[12].t35 VGND 0.01597f
C14257 XThC.Tn[12].t42 VGND 0.01682f
C14258 XThC.Tn[12].n58 VGND 0.04177f
C14259 XThC.Tn[12].n59 VGND 0.02602f
C14260 XThC.Tn[12].n60 VGND 0.08455f
C14261 XThC.Tn[12].n61 VGND 0.14116f
C14262 XThC.Tn[12].t24 VGND 0.01597f
C14263 XThC.Tn[12].t28 VGND 0.01682f
C14264 XThC.Tn[12].n62 VGND 0.04177f
C14265 XThC.Tn[12].n63 VGND 0.02602f
C14266 XThC.Tn[12].n64 VGND 0.08455f
C14267 XThC.Tn[12].n65 VGND 0.14116f
C14268 XThC.Tn[12].n66 VGND 0.67125f
C14269 XThC.Tn[12].n67 VGND 0.23845f
C14270 XThC.Tn[12].t1 VGND 0.01965f
C14271 XThC.Tn[12].t2 VGND 0.01965f
C14272 XThC.Tn[12].n68 VGND 0.04246f
C14273 XThC.Tn[12].t0 VGND 0.01965f
C14274 XThC.Tn[12].t3 VGND 0.01965f
C14275 XThC.Tn[12].n69 VGND 0.06463f
C14276 XThC.Tn[12].n70 VGND 0.17958f
C14277 XThC.Tn[12].n71 VGND 0.02824f
C14278 XThC.Tn[12].t9 VGND 0.01965f
C14279 XThC.Tn[12].t8 VGND 0.01965f
C14280 XThC.Tn[12].n72 VGND 0.05967f
C14281 XThC.Tn[12].t11 VGND 0.01965f
C14282 XThC.Tn[12].t10 VGND 0.01965f
C14283 XThC.Tn[12].n73 VGND 0.04369f
C14284 XThC.Tn[12].n74 VGND 0.19444f
C14285 XThR.Tn[7].t7 VGND 0.01512f
C14286 XThR.Tn[7].t4 VGND 0.01512f
C14287 XThR.Tn[7].n0 VGND 0.04668f
C14288 XThR.Tn[7].t6 VGND 0.01512f
C14289 XThR.Tn[7].t5 VGND 0.01512f
C14290 XThR.Tn[7].n1 VGND 0.0334f
C14291 XThR.Tn[7].n2 VGND 0.1713f
C14292 XThR.Tn[7].t2 VGND 0.02327f
C14293 XThR.Tn[7].t3 VGND 0.02327f
C14294 XThR.Tn[7].n3 VGND 0.07085f
C14295 XThR.Tn[7].t1 VGND 0.02327f
C14296 XThR.Tn[7].t0 VGND 0.02327f
C14297 XThR.Tn[7].n4 VGND 0.05154f
C14298 XThR.Tn[7].n5 VGND 0.22682f
C14299 XThR.Tn[7].n6 VGND 0.02826f
C14300 XThR.Tn[7].t58 VGND 0.01891f
C14301 XThR.Tn[7].t26 VGND 0.01991f
C14302 XThR.Tn[7].n7 VGND 0.04945f
C14303 XThR.Tn[7].n8 VGND 0.09194f
C14304 XThR.Tn[7].t38 VGND 0.01891f
C14305 XThR.Tn[7].t43 VGND 0.01991f
C14306 XThR.Tn[7].n9 VGND 0.04945f
C14307 XThR.Tn[7].t32 VGND 0.01891f
C14308 XThR.Tn[7].t42 VGND 0.01991f
C14309 XThR.Tn[7].n10 VGND 0.04943f
C14310 XThR.Tn[7].n11 VGND 0.03801f
C14311 XThR.Tn[7].n12 VGND 0.00725f
C14312 XThR.Tn[7].n13 VGND 0.11348f
C14313 XThR.Tn[7].t53 VGND 0.01891f
C14314 XThR.Tn[7].t19 VGND 0.01991f
C14315 XThR.Tn[7].n14 VGND 0.04945f
C14316 XThR.Tn[7].t48 VGND 0.01891f
C14317 XThR.Tn[7].t15 VGND 0.01991f
C14318 XThR.Tn[7].n15 VGND 0.04943f
C14319 XThR.Tn[7].n16 VGND 0.03801f
C14320 XThR.Tn[7].n17 VGND 0.00725f
C14321 XThR.Tn[7].n18 VGND 0.11348f
C14322 XThR.Tn[7].t27 VGND 0.01891f
C14323 XThR.Tn[7].t37 VGND 0.01991f
C14324 XThR.Tn[7].n19 VGND 0.04945f
C14325 XThR.Tn[7].t25 VGND 0.01891f
C14326 XThR.Tn[7].t31 VGND 0.01991f
C14327 XThR.Tn[7].n20 VGND 0.04943f
C14328 XThR.Tn[7].n21 VGND 0.03801f
C14329 XThR.Tn[7].n22 VGND 0.00725f
C14330 XThR.Tn[7].n23 VGND 0.11348f
C14331 XThR.Tn[7].t55 VGND 0.01891f
C14332 XThR.Tn[7].t66 VGND 0.01991f
C14333 XThR.Tn[7].n24 VGND 0.04945f
C14334 XThR.Tn[7].t50 VGND 0.01891f
C14335 XThR.Tn[7].t61 VGND 0.01991f
C14336 XThR.Tn[7].n25 VGND 0.04943f
C14337 XThR.Tn[7].n26 VGND 0.03801f
C14338 XThR.Tn[7].n27 VGND 0.00725f
C14339 XThR.Tn[7].n28 VGND 0.11348f
C14340 XThR.Tn[7].t9 VGND 0.01891f
C14341 XThR.Tn[7].t39 VGND 0.01991f
C14342 XThR.Tn[7].n29 VGND 0.04945f
C14343 XThR.Tn[7].t69 VGND 0.01891f
C14344 XThR.Tn[7].t34 VGND 0.01991f
C14345 XThR.Tn[7].n30 VGND 0.04943f
C14346 XThR.Tn[7].n31 VGND 0.03801f
C14347 XThR.Tn[7].n32 VGND 0.00725f
C14348 XThR.Tn[7].n33 VGND 0.11348f
C14349 XThR.Tn[7].t65 VGND 0.01891f
C14350 XThR.Tn[7].t54 VGND 0.01991f
C14351 XThR.Tn[7].n34 VGND 0.04945f
C14352 XThR.Tn[7].t60 VGND 0.01891f
C14353 XThR.Tn[7].t49 VGND 0.01991f
C14354 XThR.Tn[7].n35 VGND 0.04943f
C14355 XThR.Tn[7].n36 VGND 0.03801f
C14356 XThR.Tn[7].n37 VGND 0.00725f
C14357 XThR.Tn[7].n38 VGND 0.11348f
C14358 XThR.Tn[7].t22 VGND 0.01891f
C14359 XThR.Tn[7].t46 VGND 0.01991f
C14360 XThR.Tn[7].n39 VGND 0.04945f
C14361 XThR.Tn[7].t17 VGND 0.01891f
C14362 XThR.Tn[7].t44 VGND 0.01991f
C14363 XThR.Tn[7].n40 VGND 0.04943f
C14364 XThR.Tn[7].n41 VGND 0.03801f
C14365 XThR.Tn[7].n42 VGND 0.00725f
C14366 XThR.Tn[7].n43 VGND 0.11348f
C14367 XThR.Tn[7].t41 VGND 0.01891f
C14368 XThR.Tn[7].t64 VGND 0.01991f
C14369 XThR.Tn[7].n44 VGND 0.04945f
C14370 XThR.Tn[7].t36 VGND 0.01891f
C14371 XThR.Tn[7].t59 VGND 0.01991f
C14372 XThR.Tn[7].n45 VGND 0.04943f
C14373 XThR.Tn[7].n46 VGND 0.03801f
C14374 XThR.Tn[7].n47 VGND 0.00725f
C14375 XThR.Tn[7].n48 VGND 0.11348f
C14376 XThR.Tn[7].t57 VGND 0.01891f
C14377 XThR.Tn[7].t21 VGND 0.01991f
C14378 XThR.Tn[7].n49 VGND 0.04945f
C14379 XThR.Tn[7].t52 VGND 0.01891f
C14380 XThR.Tn[7].t16 VGND 0.01991f
C14381 XThR.Tn[7].n50 VGND 0.04943f
C14382 XThR.Tn[7].n51 VGND 0.03801f
C14383 XThR.Tn[7].n52 VGND 0.00725f
C14384 XThR.Tn[7].n53 VGND 0.11348f
C14385 XThR.Tn[7].t30 VGND 0.01891f
C14386 XThR.Tn[7].t40 VGND 0.01991f
C14387 XThR.Tn[7].n54 VGND 0.04945f
C14388 XThR.Tn[7].t28 VGND 0.01891f
C14389 XThR.Tn[7].t35 VGND 0.01991f
C14390 XThR.Tn[7].n55 VGND 0.04943f
C14391 XThR.Tn[7].n56 VGND 0.03801f
C14392 XThR.Tn[7].n57 VGND 0.00725f
C14393 XThR.Tn[7].n58 VGND 0.11348f
C14394 XThR.Tn[7].t68 VGND 0.01891f
C14395 XThR.Tn[7].t13 VGND 0.01991f
C14396 XThR.Tn[7].n59 VGND 0.04945f
C14397 XThR.Tn[7].t63 VGND 0.01891f
C14398 XThR.Tn[7].t11 VGND 0.01991f
C14399 XThR.Tn[7].n60 VGND 0.04943f
C14400 XThR.Tn[7].n61 VGND 0.03801f
C14401 XThR.Tn[7].n62 VGND 0.00725f
C14402 XThR.Tn[7].n63 VGND 0.11348f
C14403 XThR.Tn[7].t24 VGND 0.01891f
C14404 XThR.Tn[7].t47 VGND 0.01991f
C14405 XThR.Tn[7].n64 VGND 0.04945f
C14406 XThR.Tn[7].t20 VGND 0.01891f
C14407 XThR.Tn[7].t45 VGND 0.01991f
C14408 XThR.Tn[7].n65 VGND 0.04943f
C14409 XThR.Tn[7].n66 VGND 0.03801f
C14410 XThR.Tn[7].n67 VGND 0.00725f
C14411 XThR.Tn[7].n68 VGND 0.11348f
C14412 XThR.Tn[7].t56 VGND 0.01891f
C14413 XThR.Tn[7].t67 VGND 0.01991f
C14414 XThR.Tn[7].n69 VGND 0.04945f
C14415 XThR.Tn[7].t51 VGND 0.01891f
C14416 XThR.Tn[7].t62 VGND 0.01991f
C14417 XThR.Tn[7].n70 VGND 0.04943f
C14418 XThR.Tn[7].n71 VGND 0.03801f
C14419 XThR.Tn[7].n72 VGND 0.00725f
C14420 XThR.Tn[7].n73 VGND 0.11348f
C14421 XThR.Tn[7].t10 VGND 0.01891f
C14422 XThR.Tn[7].t23 VGND 0.01991f
C14423 XThR.Tn[7].n74 VGND 0.04945f
C14424 XThR.Tn[7].t8 VGND 0.01891f
C14425 XThR.Tn[7].t18 VGND 0.01991f
C14426 XThR.Tn[7].n75 VGND 0.04943f
C14427 XThR.Tn[7].n76 VGND 0.03801f
C14428 XThR.Tn[7].n77 VGND 0.00725f
C14429 XThR.Tn[7].n78 VGND 0.11348f
C14430 XThR.Tn[7].t33 VGND 0.01891f
C14431 XThR.Tn[7].t14 VGND 0.01991f
C14432 XThR.Tn[7].n79 VGND 0.04945f
C14433 XThR.Tn[7].t29 VGND 0.01891f
C14434 XThR.Tn[7].t12 VGND 0.01991f
C14435 XThR.Tn[7].n80 VGND 0.04943f
C14436 XThR.Tn[7].n81 VGND 0.03801f
C14437 XThR.Tn[7].n82 VGND 0.00725f
C14438 XThR.Tn[7].n83 VGND 0.11348f
C14439 XThR.Tn[7].n84 VGND 0.10365f
C14440 XThR.Tn[7].n85 VGND 0.42078f
C14441 XThC.Tn[5].t11 VGND 0.01819f
C14442 XThC.Tn[5].t10 VGND 0.01819f
C14443 XThC.Tn[5].n0 VGND 0.03672f
C14444 XThC.Tn[5].t9 VGND 0.01819f
C14445 XThC.Tn[5].t8 VGND 0.01819f
C14446 XThC.Tn[5].n1 VGND 0.04297f
C14447 XThC.Tn[5].n2 VGND 0.12888f
C14448 XThC.Tn[5].t5 VGND 0.01183f
C14449 XThC.Tn[5].t4 VGND 0.01183f
C14450 XThC.Tn[5].n3 VGND 0.02693f
C14451 XThC.Tn[5].t7 VGND 0.01183f
C14452 XThC.Tn[5].t6 VGND 0.01183f
C14453 XThC.Tn[5].n4 VGND 0.02693f
C14454 XThC.Tn[5].t2 VGND 0.01183f
C14455 XThC.Tn[5].t1 VGND 0.01183f
C14456 XThC.Tn[5].n5 VGND 0.02693f
C14457 XThC.Tn[5].t0 VGND 0.01183f
C14458 XThC.Tn[5].t3 VGND 0.01183f
C14459 XThC.Tn[5].n6 VGND 0.04487f
C14460 XThC.Tn[5].n7 VGND 0.12824f
C14461 XThC.Tn[5].n8 VGND 0.07928f
C14462 XThC.Tn[5].n9 VGND 0.08947f
C14463 XThC.Tn[5].t21 VGND 0.01478f
C14464 XThC.Tn[5].t24 VGND 0.01557f
C14465 XThC.Tn[5].n10 VGND 0.03867f
C14466 XThC.Tn[5].n11 VGND 0.02409f
C14467 XThC.Tn[5].n12 VGND 0.07804f
C14468 XThC.Tn[5].t30 VGND 0.01478f
C14469 XThC.Tn[5].t32 VGND 0.01557f
C14470 XThC.Tn[5].n13 VGND 0.03867f
C14471 XThC.Tn[5].n14 VGND 0.02409f
C14472 XThC.Tn[5].n15 VGND 0.07826f
C14473 XThC.Tn[5].n16 VGND 0.13067f
C14474 XThC.Tn[5].t42 VGND 0.01478f
C14475 XThC.Tn[5].t14 VGND 0.01557f
C14476 XThC.Tn[5].n17 VGND 0.03867f
C14477 XThC.Tn[5].n18 VGND 0.02409f
C14478 XThC.Tn[5].n19 VGND 0.07826f
C14479 XThC.Tn[5].n20 VGND 0.13067f
C14480 XThC.Tn[5].t12 VGND 0.01478f
C14481 XThC.Tn[5].t16 VGND 0.01557f
C14482 XThC.Tn[5].n21 VGND 0.03867f
C14483 XThC.Tn[5].n22 VGND 0.02409f
C14484 XThC.Tn[5].n23 VGND 0.07826f
C14485 XThC.Tn[5].n24 VGND 0.13067f
C14486 XThC.Tn[5].t22 VGND 0.01478f
C14487 XThC.Tn[5].t25 VGND 0.01557f
C14488 XThC.Tn[5].n25 VGND 0.03867f
C14489 XThC.Tn[5].n26 VGND 0.02409f
C14490 XThC.Tn[5].n27 VGND 0.07826f
C14491 XThC.Tn[5].n28 VGND 0.13067f
C14492 XThC.Tn[5].t33 VGND 0.01478f
C14493 XThC.Tn[5].t36 VGND 0.01557f
C14494 XThC.Tn[5].n29 VGND 0.03867f
C14495 XThC.Tn[5].n30 VGND 0.02409f
C14496 XThC.Tn[5].n31 VGND 0.07826f
C14497 XThC.Tn[5].n32 VGND 0.13067f
C14498 XThC.Tn[5].t13 VGND 0.01478f
C14499 XThC.Tn[5].t17 VGND 0.01557f
C14500 XThC.Tn[5].n33 VGND 0.03867f
C14501 XThC.Tn[5].n34 VGND 0.02409f
C14502 XThC.Tn[5].n35 VGND 0.07826f
C14503 XThC.Tn[5].n36 VGND 0.13067f
C14504 XThC.Tn[5].t23 VGND 0.01478f
C14505 XThC.Tn[5].t26 VGND 0.01557f
C14506 XThC.Tn[5].n37 VGND 0.03867f
C14507 XThC.Tn[5].n38 VGND 0.02409f
C14508 XThC.Tn[5].n39 VGND 0.07826f
C14509 XThC.Tn[5].n40 VGND 0.13067f
C14510 XThC.Tn[5].t27 VGND 0.01478f
C14511 XThC.Tn[5].t29 VGND 0.01557f
C14512 XThC.Tn[5].n41 VGND 0.03867f
C14513 XThC.Tn[5].n42 VGND 0.02409f
C14514 XThC.Tn[5].n43 VGND 0.07826f
C14515 XThC.Tn[5].n44 VGND 0.13067f
C14516 XThC.Tn[5].t34 VGND 0.01478f
C14517 XThC.Tn[5].t37 VGND 0.01557f
C14518 XThC.Tn[5].n45 VGND 0.03867f
C14519 XThC.Tn[5].n46 VGND 0.02409f
C14520 XThC.Tn[5].n47 VGND 0.07826f
C14521 XThC.Tn[5].n48 VGND 0.13067f
C14522 XThC.Tn[5].t15 VGND 0.01478f
C14523 XThC.Tn[5].t18 VGND 0.01557f
C14524 XThC.Tn[5].n49 VGND 0.03867f
C14525 XThC.Tn[5].n50 VGND 0.02409f
C14526 XThC.Tn[5].n51 VGND 0.07826f
C14527 XThC.Tn[5].n52 VGND 0.13067f
C14528 XThC.Tn[5].t19 VGND 0.01478f
C14529 XThC.Tn[5].t20 VGND 0.01557f
C14530 XThC.Tn[5].n53 VGND 0.03867f
C14531 XThC.Tn[5].n54 VGND 0.02409f
C14532 XThC.Tn[5].n55 VGND 0.07826f
C14533 XThC.Tn[5].n56 VGND 0.13067f
C14534 XThC.Tn[5].t35 VGND 0.01478f
C14535 XThC.Tn[5].t38 VGND 0.01557f
C14536 XThC.Tn[5].n57 VGND 0.03867f
C14537 XThC.Tn[5].n58 VGND 0.02409f
C14538 XThC.Tn[5].n59 VGND 0.07826f
C14539 XThC.Tn[5].n60 VGND 0.13067f
C14540 XThC.Tn[5].t39 VGND 0.01478f
C14541 XThC.Tn[5].t41 VGND 0.01557f
C14542 XThC.Tn[5].n61 VGND 0.03867f
C14543 XThC.Tn[5].n62 VGND 0.02409f
C14544 XThC.Tn[5].n63 VGND 0.07826f
C14545 XThC.Tn[5].n64 VGND 0.13067f
C14546 XThC.Tn[5].t40 VGND 0.01478f
C14547 XThC.Tn[5].t43 VGND 0.01557f
C14548 XThC.Tn[5].n65 VGND 0.03867f
C14549 XThC.Tn[5].n66 VGND 0.02409f
C14550 XThC.Tn[5].n67 VGND 0.07826f
C14551 XThC.Tn[5].n68 VGND 0.13067f
C14552 XThC.Tn[5].t28 VGND 0.01478f
C14553 XThC.Tn[5].t31 VGND 0.01557f
C14554 XThC.Tn[5].n69 VGND 0.03867f
C14555 XThC.Tn[5].n70 VGND 0.02409f
C14556 XThC.Tn[5].n71 VGND 0.07826f
C14557 XThC.Tn[5].n72 VGND 0.13067f
C14558 XThC.Tn[5].n73 VGND 0.1487f
C14559 XThC.Tn[4].t5 VGND 0.0179f
C14560 XThC.Tn[4].t4 VGND 0.0179f
C14561 XThC.Tn[4].n0 VGND 0.03613f
C14562 XThC.Tn[4].t7 VGND 0.0179f
C14563 XThC.Tn[4].t6 VGND 0.0179f
C14564 XThC.Tn[4].n1 VGND 0.04227f
C14565 XThC.Tn[4].n2 VGND 0.11834f
C14566 XThC.Tn[4].t9 VGND 0.01163f
C14567 XThC.Tn[4].t8 VGND 0.01163f
C14568 XThC.Tn[4].n3 VGND 0.02649f
C14569 XThC.Tn[4].t11 VGND 0.01163f
C14570 XThC.Tn[4].t10 VGND 0.01163f
C14571 XThC.Tn[4].n4 VGND 0.02649f
C14572 XThC.Tn[4].t2 VGND 0.01163f
C14573 XThC.Tn[4].t1 VGND 0.01163f
C14574 XThC.Tn[4].n5 VGND 0.02649f
C14575 XThC.Tn[4].t0 VGND 0.01163f
C14576 XThC.Tn[4].t3 VGND 0.01163f
C14577 XThC.Tn[4].n6 VGND 0.04415f
C14578 XThC.Tn[4].n7 VGND 0.12617f
C14579 XThC.Tn[4].n8 VGND 0.078f
C14580 XThC.Tn[4].n9 VGND 0.08802f
C14581 XThC.Tn[4].t39 VGND 0.01455f
C14582 XThC.Tn[4].t12 VGND 0.01532f
C14583 XThC.Tn[4].n10 VGND 0.03804f
C14584 XThC.Tn[4].n11 VGND 0.0237f
C14585 XThC.Tn[4].n12 VGND 0.07678f
C14586 XThC.Tn[4].t16 VGND 0.01455f
C14587 XThC.Tn[4].t21 VGND 0.01532f
C14588 XThC.Tn[4].n13 VGND 0.03804f
C14589 XThC.Tn[4].n14 VGND 0.0237f
C14590 XThC.Tn[4].n15 VGND 0.077f
C14591 XThC.Tn[4].n16 VGND 0.12856f
C14592 XThC.Tn[4].t28 VGND 0.01455f
C14593 XThC.Tn[4].t34 VGND 0.01532f
C14594 XThC.Tn[4].n17 VGND 0.03804f
C14595 XThC.Tn[4].n18 VGND 0.0237f
C14596 XThC.Tn[4].n19 VGND 0.077f
C14597 XThC.Tn[4].n20 VGND 0.12856f
C14598 XThC.Tn[4].t30 VGND 0.01455f
C14599 XThC.Tn[4].t36 VGND 0.01532f
C14600 XThC.Tn[4].n21 VGND 0.03804f
C14601 XThC.Tn[4].n22 VGND 0.0237f
C14602 XThC.Tn[4].n23 VGND 0.077f
C14603 XThC.Tn[4].n24 VGND 0.12856f
C14604 XThC.Tn[4].t41 VGND 0.01455f
C14605 XThC.Tn[4].t13 VGND 0.01532f
C14606 XThC.Tn[4].n25 VGND 0.03804f
C14607 XThC.Tn[4].n26 VGND 0.0237f
C14608 XThC.Tn[4].n27 VGND 0.077f
C14609 XThC.Tn[4].n28 VGND 0.12856f
C14610 XThC.Tn[4].t19 VGND 0.01455f
C14611 XThC.Tn[4].t24 VGND 0.01532f
C14612 XThC.Tn[4].n29 VGND 0.03804f
C14613 XThC.Tn[4].n30 VGND 0.0237f
C14614 XThC.Tn[4].n31 VGND 0.077f
C14615 XThC.Tn[4].n32 VGND 0.12856f
C14616 XThC.Tn[4].t31 VGND 0.01455f
C14617 XThC.Tn[4].t37 VGND 0.01532f
C14618 XThC.Tn[4].n33 VGND 0.03804f
C14619 XThC.Tn[4].n34 VGND 0.0237f
C14620 XThC.Tn[4].n35 VGND 0.077f
C14621 XThC.Tn[4].n36 VGND 0.12856f
C14622 XThC.Tn[4].t42 VGND 0.01455f
C14623 XThC.Tn[4].t15 VGND 0.01532f
C14624 XThC.Tn[4].n37 VGND 0.03804f
C14625 XThC.Tn[4].n38 VGND 0.0237f
C14626 XThC.Tn[4].n39 VGND 0.077f
C14627 XThC.Tn[4].n40 VGND 0.12856f
C14628 XThC.Tn[4].t43 VGND 0.01455f
C14629 XThC.Tn[4].t17 VGND 0.01532f
C14630 XThC.Tn[4].n41 VGND 0.03804f
C14631 XThC.Tn[4].n42 VGND 0.0237f
C14632 XThC.Tn[4].n43 VGND 0.077f
C14633 XThC.Tn[4].n44 VGND 0.12856f
C14634 XThC.Tn[4].t20 VGND 0.01455f
C14635 XThC.Tn[4].t26 VGND 0.01532f
C14636 XThC.Tn[4].n45 VGND 0.03804f
C14637 XThC.Tn[4].n46 VGND 0.0237f
C14638 XThC.Tn[4].n47 VGND 0.077f
C14639 XThC.Tn[4].n48 VGND 0.12856f
C14640 XThC.Tn[4].t33 VGND 0.01455f
C14641 XThC.Tn[4].t38 VGND 0.01532f
C14642 XThC.Tn[4].n49 VGND 0.03804f
C14643 XThC.Tn[4].n50 VGND 0.0237f
C14644 XThC.Tn[4].n51 VGND 0.077f
C14645 XThC.Tn[4].n52 VGND 0.12856f
C14646 XThC.Tn[4].t35 VGND 0.01455f
C14647 XThC.Tn[4].t40 VGND 0.01532f
C14648 XThC.Tn[4].n53 VGND 0.03804f
C14649 XThC.Tn[4].n54 VGND 0.0237f
C14650 XThC.Tn[4].n55 VGND 0.077f
C14651 XThC.Tn[4].n56 VGND 0.12856f
C14652 XThC.Tn[4].t22 VGND 0.01455f
C14653 XThC.Tn[4].t27 VGND 0.01532f
C14654 XThC.Tn[4].n57 VGND 0.03804f
C14655 XThC.Tn[4].n58 VGND 0.0237f
C14656 XThC.Tn[4].n59 VGND 0.077f
C14657 XThC.Tn[4].n60 VGND 0.12856f
C14658 XThC.Tn[4].t23 VGND 0.01455f
C14659 XThC.Tn[4].t29 VGND 0.01532f
C14660 XThC.Tn[4].n61 VGND 0.03804f
C14661 XThC.Tn[4].n62 VGND 0.0237f
C14662 XThC.Tn[4].n63 VGND 0.077f
C14663 XThC.Tn[4].n64 VGND 0.12856f
C14664 XThC.Tn[4].t25 VGND 0.01455f
C14665 XThC.Tn[4].t32 VGND 0.01532f
C14666 XThC.Tn[4].n65 VGND 0.03804f
C14667 XThC.Tn[4].n66 VGND 0.0237f
C14668 XThC.Tn[4].n67 VGND 0.077f
C14669 XThC.Tn[4].n68 VGND 0.12856f
C14670 XThC.Tn[4].t14 VGND 0.01455f
C14671 XThC.Tn[4].t18 VGND 0.01532f
C14672 XThC.Tn[4].n69 VGND 0.03804f
C14673 XThC.Tn[4].n70 VGND 0.0237f
C14674 XThC.Tn[4].n71 VGND 0.077f
C14675 XThC.Tn[4].n72 VGND 0.12856f
C14676 XThC.Tn[4].n73 VGND 0.15757f
C14677 XThC.Tn[4].n74 VGND 0.03746f
C14678 XThC.Tn[6].t7 VGND 0.01833f
C14679 XThC.Tn[6].t6 VGND 0.01833f
C14680 XThC.Tn[6].n0 VGND 0.03699f
C14681 XThC.Tn[6].t5 VGND 0.01833f
C14682 XThC.Tn[6].t4 VGND 0.01833f
C14683 XThC.Tn[6].n1 VGND 0.04329f
C14684 XThC.Tn[6].n2 VGND 0.12118f
C14685 XThC.Tn[6].t8 VGND 0.01191f
C14686 XThC.Tn[6].t11 VGND 0.01191f
C14687 XThC.Tn[6].n3 VGND 0.02713f
C14688 XThC.Tn[6].t10 VGND 0.01191f
C14689 XThC.Tn[6].t9 VGND 0.01191f
C14690 XThC.Tn[6].n4 VGND 0.02713f
C14691 XThC.Tn[6].t1 VGND 0.01191f
C14692 XThC.Tn[6].t0 VGND 0.01191f
C14693 XThC.Tn[6].n5 VGND 0.02713f
C14694 XThC.Tn[6].t3 VGND 0.01191f
C14695 XThC.Tn[6].t2 VGND 0.01191f
C14696 XThC.Tn[6].n6 VGND 0.0452f
C14697 XThC.Tn[6].n7 VGND 0.12919f
C14698 XThC.Tn[6].n8 VGND 0.07987f
C14699 XThC.Tn[6].n9 VGND 0.09013f
C14700 XThC.Tn[6].t32 VGND 0.01489f
C14701 XThC.Tn[6].t13 VGND 0.01568f
C14702 XThC.Tn[6].n10 VGND 0.03895f
C14703 XThC.Tn[6].n11 VGND 0.02427f
C14704 XThC.Tn[6].n12 VGND 0.07862f
C14705 XThC.Tn[6].t42 VGND 0.01489f
C14706 XThC.Tn[6].t23 VGND 0.01568f
C14707 XThC.Tn[6].n13 VGND 0.03895f
C14708 XThC.Tn[6].n14 VGND 0.02427f
C14709 XThC.Tn[6].n15 VGND 0.07884f
C14710 XThC.Tn[6].n16 VGND 0.13164f
C14711 XThC.Tn[6].t22 VGND 0.01489f
C14712 XThC.Tn[6].t36 VGND 0.01568f
C14713 XThC.Tn[6].n17 VGND 0.03895f
C14714 XThC.Tn[6].n18 VGND 0.02427f
C14715 XThC.Tn[6].n19 VGND 0.07884f
C14716 XThC.Tn[6].n20 VGND 0.13164f
C14717 XThC.Tn[6].t24 VGND 0.01489f
C14718 XThC.Tn[6].t37 VGND 0.01568f
C14719 XThC.Tn[6].n21 VGND 0.03895f
C14720 XThC.Tn[6].n22 VGND 0.02427f
C14721 XThC.Tn[6].n23 VGND 0.07884f
C14722 XThC.Tn[6].n24 VGND 0.13164f
C14723 XThC.Tn[6].t34 VGND 0.01489f
C14724 XThC.Tn[6].t16 VGND 0.01568f
C14725 XThC.Tn[6].n25 VGND 0.03895f
C14726 XThC.Tn[6].n26 VGND 0.02427f
C14727 XThC.Tn[6].n27 VGND 0.07884f
C14728 XThC.Tn[6].n28 VGND 0.13164f
C14729 XThC.Tn[6].t12 VGND 0.01489f
C14730 XThC.Tn[6].t27 VGND 0.01568f
C14731 XThC.Tn[6].n29 VGND 0.03895f
C14732 XThC.Tn[6].n30 VGND 0.02427f
C14733 XThC.Tn[6].n31 VGND 0.07884f
C14734 XThC.Tn[6].n32 VGND 0.13164f
C14735 XThC.Tn[6].t25 VGND 0.01489f
C14736 XThC.Tn[6].t38 VGND 0.01568f
C14737 XThC.Tn[6].n33 VGND 0.03895f
C14738 XThC.Tn[6].n34 VGND 0.02427f
C14739 XThC.Tn[6].n35 VGND 0.07884f
C14740 XThC.Tn[6].n36 VGND 0.13164f
C14741 XThC.Tn[6].t35 VGND 0.01489f
C14742 XThC.Tn[6].t17 VGND 0.01568f
C14743 XThC.Tn[6].n37 VGND 0.03895f
C14744 XThC.Tn[6].n38 VGND 0.02427f
C14745 XThC.Tn[6].n39 VGND 0.07884f
C14746 XThC.Tn[6].n40 VGND 0.13164f
C14747 XThC.Tn[6].t39 VGND 0.01489f
C14748 XThC.Tn[6].t19 VGND 0.01568f
C14749 XThC.Tn[6].n41 VGND 0.03895f
C14750 XThC.Tn[6].n42 VGND 0.02427f
C14751 XThC.Tn[6].n43 VGND 0.07884f
C14752 XThC.Tn[6].n44 VGND 0.13164f
C14753 XThC.Tn[6].t14 VGND 0.01489f
C14754 XThC.Tn[6].t28 VGND 0.01568f
C14755 XThC.Tn[6].n45 VGND 0.03895f
C14756 XThC.Tn[6].n46 VGND 0.02427f
C14757 XThC.Tn[6].n47 VGND 0.07884f
C14758 XThC.Tn[6].n48 VGND 0.13164f
C14759 XThC.Tn[6].t26 VGND 0.01489f
C14760 XThC.Tn[6].t40 VGND 0.01568f
C14761 XThC.Tn[6].n49 VGND 0.03895f
C14762 XThC.Tn[6].n50 VGND 0.02427f
C14763 XThC.Tn[6].n51 VGND 0.07884f
C14764 XThC.Tn[6].n52 VGND 0.13164f
C14765 XThC.Tn[6].t30 VGND 0.01489f
C14766 XThC.Tn[6].t43 VGND 0.01568f
C14767 XThC.Tn[6].n53 VGND 0.03895f
C14768 XThC.Tn[6].n54 VGND 0.02427f
C14769 XThC.Tn[6].n55 VGND 0.07884f
C14770 XThC.Tn[6].n56 VGND 0.13164f
C14771 XThC.Tn[6].t15 VGND 0.01489f
C14772 XThC.Tn[6].t29 VGND 0.01568f
C14773 XThC.Tn[6].n57 VGND 0.03895f
C14774 XThC.Tn[6].n58 VGND 0.02427f
C14775 XThC.Tn[6].n59 VGND 0.07884f
C14776 XThC.Tn[6].n60 VGND 0.13164f
C14777 XThC.Tn[6].t18 VGND 0.01489f
C14778 XThC.Tn[6].t31 VGND 0.01568f
C14779 XThC.Tn[6].n61 VGND 0.03895f
C14780 XThC.Tn[6].n62 VGND 0.02427f
C14781 XThC.Tn[6].n63 VGND 0.07884f
C14782 XThC.Tn[6].n64 VGND 0.13164f
C14783 XThC.Tn[6].t20 VGND 0.01489f
C14784 XThC.Tn[6].t33 VGND 0.01568f
C14785 XThC.Tn[6].n65 VGND 0.03895f
C14786 XThC.Tn[6].n66 VGND 0.02427f
C14787 XThC.Tn[6].n67 VGND 0.07884f
C14788 XThC.Tn[6].n68 VGND 0.13164f
C14789 XThC.Tn[6].t41 VGND 0.01489f
C14790 XThC.Tn[6].t21 VGND 0.01568f
C14791 XThC.Tn[6].n69 VGND 0.03895f
C14792 XThC.Tn[6].n70 VGND 0.02427f
C14793 XThC.Tn[6].n71 VGND 0.07884f
C14794 XThC.Tn[6].n72 VGND 0.13164f
C14795 XThC.Tn[6].n73 VGND 0.1464f
C14796 XThC.Tn[6].n74 VGND 0.03835f
C14797 XThC.XTBN.Y.n0 VGND 0.01531f
C14798 XThC.XTBN.Y.t50 VGND 0.01024f
C14799 XThC.XTBN.Y.t118 VGND 0.00603f
C14800 XThC.XTBN.Y.t18 VGND 0.01024f
C14801 XThC.XTBN.Y.t83 VGND 0.00603f
C14802 XThC.XTBN.Y.n1 VGND 0.01477f
C14803 XThC.XTBN.Y.n2 VGND 0.00524f
C14804 XThC.XTBN.Y.t120 VGND 0.01024f
C14805 XThC.XTBN.Y.t71 VGND 0.00603f
C14806 XThC.XTBN.Y.t114 VGND 0.01024f
C14807 XThC.XTBN.Y.t62 VGND 0.00603f
C14808 XThC.XTBN.Y.n3 VGND 0.0138f
C14809 XThC.XTBN.Y.n4 VGND 0.00676f
C14810 XThC.XTBN.Y.n5 VGND 0.01477f
C14811 XThC.XTBN.Y.n6 VGND 0.00676f
C14812 XThC.XTBN.Y.n7 VGND 0.00548f
C14813 XThC.XTBN.Y.n8 VGND 0.00561f
C14814 XThC.XTBN.Y.n9 VGND 0.00676f
C14815 XThC.XTBN.Y.n10 VGND 0.02164f
C14816 XThC.XTBN.Y.n11 VGND 0.00584f
C14817 XThC.XTBN.Y.n12 VGND 0.00877f
C14818 XThC.XTBN.Y.t121 VGND 0.00603f
C14819 XThC.XTBN.Y.t79 VGND 0.01024f
C14820 XThC.XTBN.Y.t84 VGND 0.00603f
C14821 XThC.XTBN.Y.t36 VGND 0.01024f
C14822 XThC.XTBN.Y.n13 VGND 0.01477f
C14823 XThC.XTBN.Y.n14 VGND 0.00524f
C14824 XThC.XTBN.Y.t73 VGND 0.00603f
C14825 XThC.XTBN.Y.t26 VGND 0.01024f
C14826 XThC.XTBN.Y.t64 VGND 0.00603f
C14827 XThC.XTBN.Y.t21 VGND 0.01024f
C14828 XThC.XTBN.Y.n15 VGND 0.0138f
C14829 XThC.XTBN.Y.n16 VGND 0.00676f
C14830 XThC.XTBN.Y.n17 VGND 0.01477f
C14831 XThC.XTBN.Y.n18 VGND 0.00676f
C14832 XThC.XTBN.Y.n19 VGND 0.00548f
C14833 XThC.XTBN.Y.n20 VGND 0.00561f
C14834 XThC.XTBN.Y.n21 VGND 0.00676f
C14835 XThC.XTBN.Y.n22 VGND 0.02164f
C14836 XThC.XTBN.Y.n23 VGND 0.00584f
C14837 XThC.XTBN.Y.n24 VGND 0.00417f
C14838 XThC.XTBN.Y.n25 VGND 0.11789f
C14839 XThC.XTBN.Y.t106 VGND 0.01024f
C14840 XThC.XTBN.Y.t89 VGND 0.00603f
C14841 XThC.XTBN.Y.t70 VGND 0.01024f
C14842 XThC.XTBN.Y.t41 VGND 0.00603f
C14843 XThC.XTBN.Y.n26 VGND 0.01477f
C14844 XThC.XTBN.Y.n27 VGND 0.00524f
C14845 XThC.XTBN.Y.t56 VGND 0.01024f
C14846 XThC.XTBN.Y.t35 VGND 0.00603f
C14847 XThC.XTBN.Y.t48 VGND 0.01024f
C14848 XThC.XTBN.Y.t32 VGND 0.00603f
C14849 XThC.XTBN.Y.n28 VGND 0.0138f
C14850 XThC.XTBN.Y.n29 VGND 0.00676f
C14851 XThC.XTBN.Y.n30 VGND 0.01477f
C14852 XThC.XTBN.Y.n31 VGND 0.00676f
C14853 XThC.XTBN.Y.n32 VGND 0.00548f
C14854 XThC.XTBN.Y.n33 VGND 0.00561f
C14855 XThC.XTBN.Y.n34 VGND 0.00676f
C14856 XThC.XTBN.Y.n35 VGND 0.02164f
C14857 XThC.XTBN.Y.n36 VGND 0.00584f
C14858 XThC.XTBN.Y.n37 VGND 0.00417f
C14859 XThC.XTBN.Y.n38 VGND 0.07443f
C14860 XThC.XTBN.Y.t43 VGND 0.00603f
C14861 XThC.XTBN.Y.t39 VGND 0.01024f
C14862 XThC.XTBN.Y.t10 VGND 0.00603f
C14863 XThC.XTBN.Y.t122 VGND 0.01024f
C14864 XThC.XTBN.Y.n39 VGND 0.01477f
C14865 XThC.XTBN.Y.n40 VGND 0.00524f
C14866 XThC.XTBN.Y.t112 VGND 0.00603f
C14867 XThC.XTBN.Y.t109 VGND 0.01024f
C14868 XThC.XTBN.Y.t108 VGND 0.00603f
C14869 XThC.XTBN.Y.t102 VGND 0.01024f
C14870 XThC.XTBN.Y.n41 VGND 0.0138f
C14871 XThC.XTBN.Y.n42 VGND 0.00676f
C14872 XThC.XTBN.Y.n43 VGND 0.01477f
C14873 XThC.XTBN.Y.n44 VGND 0.00676f
C14874 XThC.XTBN.Y.n45 VGND 0.00548f
C14875 XThC.XTBN.Y.n46 VGND 0.00561f
C14876 XThC.XTBN.Y.n47 VGND 0.00676f
C14877 XThC.XTBN.Y.n48 VGND 0.02164f
C14878 XThC.XTBN.Y.n49 VGND 0.00584f
C14879 XThC.XTBN.Y.n50 VGND 0.00417f
C14880 XThC.XTBN.Y.n51 VGND 0.07443f
C14881 XThC.XTBN.Y.t47 VGND 0.01024f
C14882 XThC.XTBN.Y.t31 VGND 0.00603f
C14883 XThC.XTBN.Y.t17 VGND 0.01024f
C14884 XThC.XTBN.Y.t104 VGND 0.00603f
C14885 XThC.XTBN.Y.n52 VGND 0.01477f
C14886 XThC.XTBN.Y.n53 VGND 0.00524f
C14887 XThC.XTBN.Y.t116 VGND 0.01024f
C14888 XThC.XTBN.Y.t94 VGND 0.00603f
C14889 XThC.XTBN.Y.t111 VGND 0.01024f
C14890 XThC.XTBN.Y.t92 VGND 0.00603f
C14891 XThC.XTBN.Y.n54 VGND 0.0138f
C14892 XThC.XTBN.Y.n55 VGND 0.00676f
C14893 XThC.XTBN.Y.n56 VGND 0.01477f
C14894 XThC.XTBN.Y.n57 VGND 0.00676f
C14895 XThC.XTBN.Y.n58 VGND 0.00548f
C14896 XThC.XTBN.Y.n59 VGND 0.00561f
C14897 XThC.XTBN.Y.n60 VGND 0.00676f
C14898 XThC.XTBN.Y.n61 VGND 0.02164f
C14899 XThC.XTBN.Y.n62 VGND 0.00584f
C14900 XThC.XTBN.Y.n63 VGND 0.00417f
C14901 XThC.XTBN.Y.n64 VGND 0.07443f
C14902 XThC.XTBN.Y.t107 VGND 0.00603f
C14903 XThC.XTBN.Y.t101 VGND 0.01024f
C14904 XThC.XTBN.Y.t72 VGND 0.00603f
C14905 XThC.XTBN.Y.t63 VGND 0.01024f
C14906 XThC.XTBN.Y.n65 VGND 0.01477f
C14907 XThC.XTBN.Y.n66 VGND 0.00524f
C14908 XThC.XTBN.Y.t57 VGND 0.00603f
C14909 XThC.XTBN.Y.t52 VGND 0.01024f
C14910 XThC.XTBN.Y.t49 VGND 0.00603f
C14911 XThC.XTBN.Y.t44 VGND 0.01024f
C14912 XThC.XTBN.Y.n67 VGND 0.0138f
C14913 XThC.XTBN.Y.n68 VGND 0.00676f
C14914 XThC.XTBN.Y.n69 VGND 0.01477f
C14915 XThC.XTBN.Y.n70 VGND 0.00676f
C14916 XThC.XTBN.Y.n71 VGND 0.00548f
C14917 XThC.XTBN.Y.n72 VGND 0.00561f
C14918 XThC.XTBN.Y.n73 VGND 0.00676f
C14919 XThC.XTBN.Y.n74 VGND 0.02164f
C14920 XThC.XTBN.Y.n75 VGND 0.00584f
C14921 XThC.XTBN.Y.n76 VGND 0.00417f
C14922 XThC.XTBN.Y.n77 VGND 0.07443f
C14923 XThC.XTBN.Y.t25 VGND 0.01024f
C14924 XThC.XTBN.Y.t123 VGND 0.00603f
C14925 XThC.XTBN.Y.t100 VGND 0.01024f
C14926 XThC.XTBN.Y.t85 VGND 0.00603f
C14927 XThC.XTBN.Y.n78 VGND 0.01477f
C14928 XThC.XTBN.Y.n79 VGND 0.00524f
C14929 XThC.XTBN.Y.t93 VGND 0.01024f
C14930 XThC.XTBN.Y.t74 VGND 0.00603f
C14931 XThC.XTBN.Y.t90 VGND 0.01024f
C14932 XThC.XTBN.Y.t65 VGND 0.00603f
C14933 XThC.XTBN.Y.n80 VGND 0.0138f
C14934 XThC.XTBN.Y.n81 VGND 0.00676f
C14935 XThC.XTBN.Y.n82 VGND 0.01477f
C14936 XThC.XTBN.Y.n83 VGND 0.00676f
C14937 XThC.XTBN.Y.n84 VGND 0.00548f
C14938 XThC.XTBN.Y.n85 VGND 0.00561f
C14939 XThC.XTBN.Y.n86 VGND 0.00676f
C14940 XThC.XTBN.Y.n87 VGND 0.02164f
C14941 XThC.XTBN.Y.n88 VGND 0.00584f
C14942 XThC.XTBN.Y.n89 VGND 0.00417f
C14943 XThC.XTBN.Y.n90 VGND 0.06646f
C14944 XThC.XTBN.Y.t46 VGND 0.01024f
C14945 XThC.XTBN.Y.t67 VGND 0.00603f
C14946 XThC.XTBN.Y.n91 VGND 0.00619f
C14947 XThC.XTBN.Y.t6 VGND 0.01024f
C14948 XThC.XTBN.Y.t24 VGND 0.00603f
C14949 XThC.XTBN.Y.n92 VGND 0.01243f
C14950 XThC.XTBN.Y.t12 VGND 0.01024f
C14951 XThC.XTBN.Y.t29 VGND 0.00603f
C14952 XThC.XTBN.Y.n93 VGND 0.01348f
C14953 XThC.XTBN.Y.n94 VGND 0.0076f
C14954 XThC.XTBN.Y.n95 VGND 0.01252f
C14955 XThC.XTBN.Y.n96 VGND 0.00434f
C14956 XThC.XTBN.Y.n97 VGND 0.00603f
C14957 XThC.XTBN.Y.n98 VGND 0.01348f
C14958 XThC.XTBN.Y.t54 VGND 0.01024f
C14959 XThC.XTBN.Y.t76 VGND 0.00603f
C14960 XThC.XTBN.Y.n99 VGND 0.01227f
C14961 XThC.XTBN.Y.n100 VGND 0.00676f
C14962 XThC.XTBN.Y.n101 VGND 0.01009f
C14963 XThC.XTBN.Y.t55 VGND 0.00603f
C14964 XThC.XTBN.Y.t38 VGND 0.01024f
C14965 XThC.XTBN.Y.n102 VGND 0.00619f
C14966 XThC.XTBN.Y.t16 VGND 0.00603f
C14967 XThC.XTBN.Y.t113 VGND 0.01024f
C14968 XThC.XTBN.Y.n103 VGND 0.01243f
C14969 XThC.XTBN.Y.t19 VGND 0.00603f
C14970 XThC.XTBN.Y.t119 VGND 0.01024f
C14971 XThC.XTBN.Y.n104 VGND 0.01348f
C14972 XThC.XTBN.Y.n105 VGND 0.0076f
C14973 XThC.XTBN.Y.n106 VGND 0.01252f
C14974 XThC.XTBN.Y.n107 VGND 0.00434f
C14975 XThC.XTBN.Y.n108 VGND 0.00603f
C14976 XThC.XTBN.Y.n109 VGND 0.01348f
C14977 XThC.XTBN.Y.t59 VGND 0.00603f
C14978 XThC.XTBN.Y.t42 VGND 0.01024f
C14979 XThC.XTBN.Y.n110 VGND 0.01227f
C14980 XThC.XTBN.Y.n111 VGND 0.00676f
C14981 XThC.XTBN.Y.n112 VGND 0.00747f
C14982 XThC.XTBN.Y.n113 VGND 0.11256f
C14983 XThC.XTBN.Y.t30 VGND 0.01024f
C14984 XThC.XTBN.Y.t8 VGND 0.00603f
C14985 XThC.XTBN.Y.n114 VGND 0.00619f
C14986 XThC.XTBN.Y.t98 VGND 0.01024f
C14987 XThC.XTBN.Y.t82 VGND 0.00603f
C14988 XThC.XTBN.Y.n115 VGND 0.01243f
C14989 XThC.XTBN.Y.t103 VGND 0.01024f
C14990 XThC.XTBN.Y.t87 VGND 0.00603f
C14991 XThC.XTBN.Y.n116 VGND 0.01348f
C14992 XThC.XTBN.Y.n117 VGND 0.0076f
C14993 XThC.XTBN.Y.n118 VGND 0.01252f
C14994 XThC.XTBN.Y.n119 VGND 0.00434f
C14995 XThC.XTBN.Y.n120 VGND 0.00603f
C14996 XThC.XTBN.Y.n121 VGND 0.01348f
C14997 XThC.XTBN.Y.t34 VGND 0.01024f
C14998 XThC.XTBN.Y.t15 VGND 0.00603f
C14999 XThC.XTBN.Y.n122 VGND 0.01227f
C15000 XThC.XTBN.Y.n123 VGND 0.00676f
C15001 XThC.XTBN.Y.n124 VGND 0.00747f
C15002 XThC.XTBN.Y.n125 VGND 0.07521f
C15003 XThC.XTBN.Y.t110 VGND 0.00603f
C15004 XThC.XTBN.Y.t96 VGND 0.01024f
C15005 XThC.XTBN.Y.n126 VGND 0.00619f
C15006 XThC.XTBN.Y.t68 VGND 0.00603f
C15007 XThC.XTBN.Y.t51 VGND 0.01024f
C15008 XThC.XTBN.Y.n127 VGND 0.01243f
C15009 XThC.XTBN.Y.t77 VGND 0.00603f
C15010 XThC.XTBN.Y.t58 VGND 0.01024f
C15011 XThC.XTBN.Y.n128 VGND 0.01348f
C15012 XThC.XTBN.Y.n129 VGND 0.0076f
C15013 XThC.XTBN.Y.n130 VGND 0.01252f
C15014 XThC.XTBN.Y.n131 VGND 0.00434f
C15015 XThC.XTBN.Y.n132 VGND 0.00603f
C15016 XThC.XTBN.Y.n133 VGND 0.01348f
C15017 XThC.XTBN.Y.t115 VGND 0.00603f
C15018 XThC.XTBN.Y.t99 VGND 0.01024f
C15019 XThC.XTBN.Y.n134 VGND 0.01227f
C15020 XThC.XTBN.Y.n135 VGND 0.00676f
C15021 XThC.XTBN.Y.n136 VGND 0.00747f
C15022 XThC.XTBN.Y.n137 VGND 0.07521f
C15023 XThC.XTBN.Y.t88 VGND 0.01024f
C15024 XThC.XTBN.Y.t60 VGND 0.00603f
C15025 XThC.XTBN.Y.n138 VGND 0.00619f
C15026 XThC.XTBN.Y.t37 VGND 0.01024f
C15027 XThC.XTBN.Y.t20 VGND 0.00603f
C15028 XThC.XTBN.Y.n139 VGND 0.01243f
C15029 XThC.XTBN.Y.t40 VGND 0.01024f
C15030 XThC.XTBN.Y.t22 VGND 0.00603f
C15031 XThC.XTBN.Y.n140 VGND 0.01348f
C15032 XThC.XTBN.Y.n141 VGND 0.0076f
C15033 XThC.XTBN.Y.n142 VGND 0.01252f
C15034 XThC.XTBN.Y.n143 VGND 0.00434f
C15035 XThC.XTBN.Y.n144 VGND 0.00603f
C15036 XThC.XTBN.Y.n145 VGND 0.01348f
C15037 XThC.XTBN.Y.t91 VGND 0.01024f
C15038 XThC.XTBN.Y.t66 VGND 0.00603f
C15039 XThC.XTBN.Y.n146 VGND 0.01227f
C15040 XThC.XTBN.Y.n147 VGND 0.00676f
C15041 XThC.XTBN.Y.n148 VGND 0.00747f
C15042 XThC.XTBN.Y.n149 VGND 0.07534f
C15043 XThC.XTBN.Y.t45 VGND 0.00603f
C15044 XThC.XTBN.Y.t7 VGND 0.01024f
C15045 XThC.XTBN.Y.n150 VGND 0.00619f
C15046 XThC.XTBN.Y.t5 VGND 0.00603f
C15047 XThC.XTBN.Y.t81 VGND 0.01024f
C15048 XThC.XTBN.Y.n151 VGND 0.01243f
C15049 XThC.XTBN.Y.t11 VGND 0.00603f
C15050 XThC.XTBN.Y.t86 VGND 0.01024f
C15051 XThC.XTBN.Y.n152 VGND 0.01348f
C15052 XThC.XTBN.Y.n153 VGND 0.0076f
C15053 XThC.XTBN.Y.n154 VGND 0.01252f
C15054 XThC.XTBN.Y.n155 VGND 0.00434f
C15055 XThC.XTBN.Y.n156 VGND 0.00603f
C15056 XThC.XTBN.Y.n157 VGND 0.01348f
C15057 XThC.XTBN.Y.t53 VGND 0.00603f
C15058 XThC.XTBN.Y.t13 VGND 0.01024f
C15059 XThC.XTBN.Y.n158 VGND 0.01227f
C15060 XThC.XTBN.Y.n159 VGND 0.00676f
C15061 XThC.XTBN.Y.n160 VGND 0.00747f
C15062 XThC.XTBN.Y.n161 VGND 0.07521f
C15063 XThC.XTBN.Y.t23 VGND 0.01024f
C15064 XThC.XTBN.Y.t117 VGND 0.00603f
C15065 XThC.XTBN.Y.n162 VGND 0.00619f
C15066 XThC.XTBN.Y.t95 VGND 0.01024f
C15067 XThC.XTBN.Y.t78 VGND 0.00603f
C15068 XThC.XTBN.Y.n163 VGND 0.01243f
C15069 XThC.XTBN.Y.t97 VGND 0.01024f
C15070 XThC.XTBN.Y.t80 VGND 0.00603f
C15071 XThC.XTBN.Y.n164 VGND 0.01348f
C15072 XThC.XTBN.Y.n165 VGND 0.0076f
C15073 XThC.XTBN.Y.n166 VGND 0.01252f
C15074 XThC.XTBN.Y.n167 VGND 0.00434f
C15075 XThC.XTBN.Y.n168 VGND 0.00603f
C15076 XThC.XTBN.Y.n169 VGND 0.01348f
C15077 XThC.XTBN.Y.t28 VGND 0.01024f
C15078 XThC.XTBN.Y.t4 VGND 0.00603f
C15079 XThC.XTBN.Y.n170 VGND 0.01227f
C15080 XThC.XTBN.Y.n171 VGND 0.00676f
C15081 XThC.XTBN.Y.n172 VGND 0.00747f
C15082 XThC.XTBN.Y.n173 VGND 0.08751f
C15083 XThC.XTBN.Y.n174 VGND 0.11019f
C15084 XThC.XTBN.Y.t105 VGND 0.00603f
C15085 XThC.XTBN.Y.t75 VGND 0.01024f
C15086 XThC.XTBN.Y.t69 VGND 0.00603f
C15087 XThC.XTBN.Y.t33 VGND 0.01024f
C15088 XThC.XTBN.Y.n175 VGND 0.01477f
C15089 XThC.XTBN.Y.t61 VGND 0.00603f
C15090 XThC.XTBN.Y.t27 VGND 0.01024f
C15091 XThC.XTBN.Y.n176 VGND 0.02293f
C15092 XThC.XTBN.Y.n177 VGND 0.00676f
C15093 XThC.XTBN.Y.n178 VGND 0.00561f
C15094 XThC.XTBN.Y.n179 VGND 0.00561f
C15095 XThC.XTBN.Y.n180 VGND 0.00676f
C15096 XThC.XTBN.Y.n181 VGND 0.01477f
C15097 XThC.XTBN.Y.t14 VGND 0.00603f
C15098 XThC.XTBN.Y.t9 VGND 0.01024f
C15099 XThC.XTBN.Y.n182 VGND 0.0138f
C15100 XThC.XTBN.Y.n183 VGND 0.00676f
C15101 XThC.XTBN.Y.n184 VGND 0.00372f
C15102 XThC.XTBN.Y.n185 VGND 0.00408f
C15103 XThC.XTBN.Y.n186 VGND 0.11129f
C15104 XThC.XTBN.Y.n187 VGND 0.02169f
C15105 XThC.XTBN.Y.t3 VGND 0.00428f
C15106 XThC.XTBN.Y.t2 VGND 0.00428f
C15107 XThC.XTBN.Y.n188 VGND 0.0094f
C15108 XThC.XTBN.Y.n189 VGND 0.00607f
C15109 XThC.XTBN.Y.n190 VGND 0.00526f
C15110 XThC.XTBN.Y.t0 VGND 0.00658f
C15111 XThC.XTBN.Y.t1 VGND 0.00658f
C15112 XThC.XTBN.Y.n191 VGND 0.01513f
C15113 XThC.XTBN.Y.n192 VGND 0.0307f
C15114 XThR.Tn[8].t10 VGND 0.0243f
C15115 XThR.Tn[8].t8 VGND 0.0243f
C15116 XThR.Tn[8].n0 VGND 0.07378f
C15117 XThR.Tn[8].t11 VGND 0.0243f
C15118 XThR.Tn[8].t9 VGND 0.0243f
C15119 XThR.Tn[8].n1 VGND 0.05401f
C15120 XThR.Tn[8].n2 VGND 0.2456f
C15121 XThR.Tn[8].t3 VGND 0.01579f
C15122 XThR.Tn[8].t5 VGND 0.01579f
C15123 XThR.Tn[8].n3 VGND 0.03939f
C15124 XThR.Tn[8].t4 VGND 0.01579f
C15125 XThR.Tn[8].t6 VGND 0.01579f
C15126 XThR.Tn[8].n4 VGND 0.03159f
C15127 XThR.Tn[8].n5 VGND 0.07284f
C15128 XThR.Tn[8].t63 VGND 0.01975f
C15129 XThR.Tn[8].t29 VGND 0.02079f
C15130 XThR.Tn[8].n6 VGND 0.05164f
C15131 XThR.Tn[8].n7 VGND 0.09601f
C15132 XThR.Tn[8].t41 VGND 0.01975f
C15133 XThR.Tn[8].t45 VGND 0.02079f
C15134 XThR.Tn[8].n8 VGND 0.05164f
C15135 XThR.Tn[8].t18 VGND 0.01975f
C15136 XThR.Tn[8].t25 VGND 0.02079f
C15137 XThR.Tn[8].n9 VGND 0.05162f
C15138 XThR.Tn[8].n10 VGND 0.0397f
C15139 XThR.Tn[8].n11 VGND 0.00757f
C15140 XThR.Tn[8].n12 VGND 0.11851f
C15141 XThR.Tn[8].t55 VGND 0.01975f
C15142 XThR.Tn[8].t23 VGND 0.02079f
C15143 XThR.Tn[8].n13 VGND 0.05164f
C15144 XThR.Tn[8].t34 VGND 0.01975f
C15145 XThR.Tn[8].t62 VGND 0.02079f
C15146 XThR.Tn[8].n14 VGND 0.05162f
C15147 XThR.Tn[8].n15 VGND 0.0397f
C15148 XThR.Tn[8].n16 VGND 0.00757f
C15149 XThR.Tn[8].n17 VGND 0.11851f
C15150 XThR.Tn[8].t31 VGND 0.01975f
C15151 XThR.Tn[8].t40 VGND 0.02079f
C15152 XThR.Tn[8].n18 VGND 0.05164f
C15153 XThR.Tn[8].t73 VGND 0.01975f
C15154 XThR.Tn[8].t17 VGND 0.02079f
C15155 XThR.Tn[8].n19 VGND 0.05162f
C15156 XThR.Tn[8].n20 VGND 0.0397f
C15157 XThR.Tn[8].n21 VGND 0.00757f
C15158 XThR.Tn[8].n22 VGND 0.11851f
C15159 XThR.Tn[8].t57 VGND 0.01975f
C15160 XThR.Tn[8].t70 VGND 0.02079f
C15161 XThR.Tn[8].n23 VGND 0.05164f
C15162 XThR.Tn[8].t36 VGND 0.01975f
C15163 XThR.Tn[8].t48 VGND 0.02079f
C15164 XThR.Tn[8].n24 VGND 0.05162f
C15165 XThR.Tn[8].n25 VGND 0.0397f
C15166 XThR.Tn[8].n26 VGND 0.00757f
C15167 XThR.Tn[8].n27 VGND 0.11851f
C15168 XThR.Tn[8].t12 VGND 0.01975f
C15169 XThR.Tn[8].t42 VGND 0.02079f
C15170 XThR.Tn[8].n28 VGND 0.05164f
C15171 XThR.Tn[8].t53 VGND 0.01975f
C15172 XThR.Tn[8].t20 VGND 0.02079f
C15173 XThR.Tn[8].n29 VGND 0.05162f
C15174 XThR.Tn[8].n30 VGND 0.0397f
C15175 XThR.Tn[8].n31 VGND 0.00757f
C15176 XThR.Tn[8].n32 VGND 0.11851f
C15177 XThR.Tn[8].t69 VGND 0.01975f
C15178 XThR.Tn[8].t56 VGND 0.02079f
C15179 XThR.Tn[8].n33 VGND 0.05164f
C15180 XThR.Tn[8].t47 VGND 0.01975f
C15181 XThR.Tn[8].t35 VGND 0.02079f
C15182 XThR.Tn[8].n34 VGND 0.05162f
C15183 XThR.Tn[8].n35 VGND 0.0397f
C15184 XThR.Tn[8].n36 VGND 0.00757f
C15185 XThR.Tn[8].n37 VGND 0.11851f
C15186 XThR.Tn[8].t26 VGND 0.01975f
C15187 XThR.Tn[8].t51 VGND 0.02079f
C15188 XThR.Tn[8].n38 VGND 0.05164f
C15189 XThR.Tn[8].t65 VGND 0.01975f
C15190 XThR.Tn[8].t30 VGND 0.02079f
C15191 XThR.Tn[8].n39 VGND 0.05162f
C15192 XThR.Tn[8].n40 VGND 0.0397f
C15193 XThR.Tn[8].n41 VGND 0.00757f
C15194 XThR.Tn[8].n42 VGND 0.11851f
C15195 XThR.Tn[8].t44 VGND 0.01975f
C15196 XThR.Tn[8].t68 VGND 0.02079f
C15197 XThR.Tn[8].n43 VGND 0.05164f
C15198 XThR.Tn[8].t22 VGND 0.01975f
C15199 XThR.Tn[8].t46 VGND 0.02079f
C15200 XThR.Tn[8].n44 VGND 0.05162f
C15201 XThR.Tn[8].n45 VGND 0.0397f
C15202 XThR.Tn[8].n46 VGND 0.00757f
C15203 XThR.Tn[8].n47 VGND 0.11851f
C15204 XThR.Tn[8].t61 VGND 0.01975f
C15205 XThR.Tn[8].t24 VGND 0.02079f
C15206 XThR.Tn[8].n48 VGND 0.05164f
C15207 XThR.Tn[8].t39 VGND 0.01975f
C15208 XThR.Tn[8].t64 VGND 0.02079f
C15209 XThR.Tn[8].n49 VGND 0.05162f
C15210 XThR.Tn[8].n50 VGND 0.0397f
C15211 XThR.Tn[8].n51 VGND 0.00757f
C15212 XThR.Tn[8].n52 VGND 0.11851f
C15213 XThR.Tn[8].t33 VGND 0.01975f
C15214 XThR.Tn[8].t43 VGND 0.02079f
C15215 XThR.Tn[8].n53 VGND 0.05164f
C15216 XThR.Tn[8].t14 VGND 0.01975f
C15217 XThR.Tn[8].t21 VGND 0.02079f
C15218 XThR.Tn[8].n54 VGND 0.05162f
C15219 XThR.Tn[8].n55 VGND 0.0397f
C15220 XThR.Tn[8].n56 VGND 0.00757f
C15221 XThR.Tn[8].n57 VGND 0.11851f
C15222 XThR.Tn[8].t72 VGND 0.01975f
C15223 XThR.Tn[8].t16 VGND 0.02079f
C15224 XThR.Tn[8].n58 VGND 0.05164f
C15225 XThR.Tn[8].t50 VGND 0.01975f
C15226 XThR.Tn[8].t58 VGND 0.02079f
C15227 XThR.Tn[8].n59 VGND 0.05162f
C15228 XThR.Tn[8].n60 VGND 0.0397f
C15229 XThR.Tn[8].n61 VGND 0.00757f
C15230 XThR.Tn[8].n62 VGND 0.11851f
C15231 XThR.Tn[8].t28 VGND 0.01975f
C15232 XThR.Tn[8].t52 VGND 0.02079f
C15233 XThR.Tn[8].n63 VGND 0.05164f
C15234 XThR.Tn[8].t67 VGND 0.01975f
C15235 XThR.Tn[8].t32 VGND 0.02079f
C15236 XThR.Tn[8].n64 VGND 0.05162f
C15237 XThR.Tn[8].n65 VGND 0.0397f
C15238 XThR.Tn[8].n66 VGND 0.00757f
C15239 XThR.Tn[8].n67 VGND 0.11851f
C15240 XThR.Tn[8].t59 VGND 0.01975f
C15241 XThR.Tn[8].t71 VGND 0.02079f
C15242 XThR.Tn[8].n68 VGND 0.05164f
C15243 XThR.Tn[8].t38 VGND 0.01975f
C15244 XThR.Tn[8].t49 VGND 0.02079f
C15245 XThR.Tn[8].n69 VGND 0.05162f
C15246 XThR.Tn[8].n70 VGND 0.0397f
C15247 XThR.Tn[8].n71 VGND 0.00757f
C15248 XThR.Tn[8].n72 VGND 0.11851f
C15249 XThR.Tn[8].t13 VGND 0.01975f
C15250 XThR.Tn[8].t27 VGND 0.02079f
C15251 XThR.Tn[8].n73 VGND 0.05164f
C15252 XThR.Tn[8].t54 VGND 0.01975f
C15253 XThR.Tn[8].t66 VGND 0.02079f
C15254 XThR.Tn[8].n74 VGND 0.05162f
C15255 XThR.Tn[8].n75 VGND 0.0397f
C15256 XThR.Tn[8].n76 VGND 0.00757f
C15257 XThR.Tn[8].n77 VGND 0.11851f
C15258 XThR.Tn[8].t37 VGND 0.01975f
C15259 XThR.Tn[8].t19 VGND 0.02079f
C15260 XThR.Tn[8].n78 VGND 0.05164f
C15261 XThR.Tn[8].t15 VGND 0.01975f
C15262 XThR.Tn[8].t60 VGND 0.02079f
C15263 XThR.Tn[8].n79 VGND 0.05162f
C15264 XThR.Tn[8].n80 VGND 0.0397f
C15265 XThR.Tn[8].n81 VGND 0.00757f
C15266 XThR.Tn[8].n82 VGND 0.11851f
C15267 XThR.Tn[8].n83 VGND 0.10825f
C15268 XThR.Tn[8].n84 VGND 0.33168f
C15269 XThR.Tn[8].t0 VGND 0.0243f
C15270 XThR.Tn[8].t2 VGND 0.0243f
C15271 XThR.Tn[8].n85 VGND 0.0525f
C15272 XThR.Tn[8].t7 VGND 0.0243f
C15273 XThR.Tn[8].t1 VGND 0.0243f
C15274 XThR.Tn[8].n86 VGND 0.07991f
C15275 XThR.Tn[8].n87 VGND 0.22187f
C15276 XThR.Tn[8].n88 VGND 0.01093f
C15277 XThR.Tn[14].t8 VGND 0.0245f
C15278 XThR.Tn[14].t9 VGND 0.0245f
C15279 XThR.Tn[14].n0 VGND 0.07438f
C15280 XThR.Tn[14].t10 VGND 0.0245f
C15281 XThR.Tn[14].t11 VGND 0.0245f
C15282 XThR.Tn[14].n1 VGND 0.05445f
C15283 XThR.Tn[14].n2 VGND 0.2476f
C15284 XThR.Tn[14].t6 VGND 0.01592f
C15285 XThR.Tn[14].t7 VGND 0.01592f
C15286 XThR.Tn[14].n3 VGND 0.03971f
C15287 XThR.Tn[14].t4 VGND 0.01592f
C15288 XThR.Tn[14].t5 VGND 0.01592f
C15289 XThR.Tn[14].n4 VGND 0.03185f
C15290 XThR.Tn[14].n5 VGND 0.07343f
C15291 XThR.Tn[14].t13 VGND 0.01991f
C15292 XThR.Tn[14].t43 VGND 0.02096f
C15293 XThR.Tn[14].n6 VGND 0.05206f
C15294 XThR.Tn[14].n7 VGND 0.09679f
C15295 XThR.Tn[14].t52 VGND 0.01991f
C15296 XThR.Tn[14].t59 VGND 0.02096f
C15297 XThR.Tn[14].n8 VGND 0.05206f
C15298 XThR.Tn[14].t34 VGND 0.01991f
C15299 XThR.Tn[14].t42 VGND 0.02096f
C15300 XThR.Tn[14].n9 VGND 0.05204f
C15301 XThR.Tn[14].n10 VGND 0.04002f
C15302 XThR.Tn[14].n11 VGND 0.00763f
C15303 XThR.Tn[14].n12 VGND 0.11947f
C15304 XThR.Tn[14].t67 VGND 0.01991f
C15305 XThR.Tn[14].t33 VGND 0.02096f
C15306 XThR.Tn[14].n13 VGND 0.05206f
C15307 XThR.Tn[14].t50 VGND 0.01991f
C15308 XThR.Tn[14].t15 VGND 0.02096f
C15309 XThR.Tn[14].n14 VGND 0.05204f
C15310 XThR.Tn[14].n15 VGND 0.04002f
C15311 XThR.Tn[14].n16 VGND 0.00763f
C15312 XThR.Tn[14].n17 VGND 0.11947f
C15313 XThR.Tn[14].t44 VGND 0.01991f
C15314 XThR.Tn[14].t49 VGND 0.02096f
C15315 XThR.Tn[14].n18 VGND 0.05206f
C15316 XThR.Tn[14].t25 VGND 0.01991f
C15317 XThR.Tn[14].t32 VGND 0.02096f
C15318 XThR.Tn[14].n19 VGND 0.05204f
C15319 XThR.Tn[14].n20 VGND 0.04002f
C15320 XThR.Tn[14].n21 VGND 0.00763f
C15321 XThR.Tn[14].n22 VGND 0.11947f
C15322 XThR.Tn[14].t70 VGND 0.01991f
C15323 XThR.Tn[14].t20 VGND 0.02096f
C15324 XThR.Tn[14].n23 VGND 0.05206f
C15325 XThR.Tn[14].t54 VGND 0.01991f
C15326 XThR.Tn[14].t63 VGND 0.02096f
C15327 XThR.Tn[14].n24 VGND 0.05204f
C15328 XThR.Tn[14].n25 VGND 0.04002f
C15329 XThR.Tn[14].n26 VGND 0.00763f
C15330 XThR.Tn[14].n27 VGND 0.11947f
C15331 XThR.Tn[14].t26 VGND 0.01991f
C15332 XThR.Tn[14].t53 VGND 0.02096f
C15333 XThR.Tn[14].n28 VGND 0.05206f
C15334 XThR.Tn[14].t69 VGND 0.01991f
C15335 XThR.Tn[14].t35 VGND 0.02096f
C15336 XThR.Tn[14].n29 VGND 0.05204f
C15337 XThR.Tn[14].n30 VGND 0.04002f
C15338 XThR.Tn[14].n31 VGND 0.00763f
C15339 XThR.Tn[14].n32 VGND 0.11947f
C15340 XThR.Tn[14].t19 VGND 0.01991f
C15341 XThR.Tn[14].t68 VGND 0.02096f
C15342 XThR.Tn[14].n33 VGND 0.05206f
C15343 XThR.Tn[14].t62 VGND 0.01991f
C15344 XThR.Tn[14].t51 VGND 0.02096f
C15345 XThR.Tn[14].n34 VGND 0.05204f
C15346 XThR.Tn[14].n35 VGND 0.04002f
C15347 XThR.Tn[14].n36 VGND 0.00763f
C15348 XThR.Tn[14].n37 VGND 0.11947f
C15349 XThR.Tn[14].t38 VGND 0.01991f
C15350 XThR.Tn[14].t61 VGND 0.02096f
C15351 XThR.Tn[14].n38 VGND 0.05206f
C15352 XThR.Tn[14].t18 VGND 0.01991f
C15353 XThR.Tn[14].t45 VGND 0.02096f
C15354 XThR.Tn[14].n39 VGND 0.05204f
C15355 XThR.Tn[14].n40 VGND 0.04002f
C15356 XThR.Tn[14].n41 VGND 0.00763f
C15357 XThR.Tn[14].n42 VGND 0.11947f
C15358 XThR.Tn[14].t58 VGND 0.01991f
C15359 XThR.Tn[14].t17 VGND 0.02096f
C15360 XThR.Tn[14].n43 VGND 0.05206f
C15361 XThR.Tn[14].t39 VGND 0.01991f
C15362 XThR.Tn[14].t60 VGND 0.02096f
C15363 XThR.Tn[14].n44 VGND 0.05204f
C15364 XThR.Tn[14].n45 VGND 0.04002f
C15365 XThR.Tn[14].n46 VGND 0.00763f
C15366 XThR.Tn[14].n47 VGND 0.11947f
C15367 XThR.Tn[14].t73 VGND 0.01991f
C15368 XThR.Tn[14].t36 VGND 0.02096f
C15369 XThR.Tn[14].n48 VGND 0.05206f
C15370 XThR.Tn[14].t57 VGND 0.01991f
C15371 XThR.Tn[14].t16 VGND 0.02096f
C15372 XThR.Tn[14].n49 VGND 0.05204f
C15373 XThR.Tn[14].n50 VGND 0.04002f
C15374 XThR.Tn[14].n51 VGND 0.00763f
C15375 XThR.Tn[14].n52 VGND 0.11947f
C15376 XThR.Tn[14].t47 VGND 0.01991f
C15377 XThR.Tn[14].t56 VGND 0.02096f
C15378 XThR.Tn[14].n53 VGND 0.05206f
C15379 XThR.Tn[14].t29 VGND 0.01991f
C15380 XThR.Tn[14].t37 VGND 0.02096f
C15381 XThR.Tn[14].n54 VGND 0.05204f
C15382 XThR.Tn[14].n55 VGND 0.04002f
C15383 XThR.Tn[14].n56 VGND 0.00763f
C15384 XThR.Tn[14].n57 VGND 0.11947f
C15385 XThR.Tn[14].t24 VGND 0.01991f
C15386 XThR.Tn[14].t28 VGND 0.02096f
C15387 XThR.Tn[14].n58 VGND 0.05206f
C15388 XThR.Tn[14].t66 VGND 0.01991f
C15389 XThR.Tn[14].t12 VGND 0.02096f
C15390 XThR.Tn[14].n59 VGND 0.05204f
C15391 XThR.Tn[14].n60 VGND 0.04002f
C15392 XThR.Tn[14].n61 VGND 0.00763f
C15393 XThR.Tn[14].n62 VGND 0.11947f
C15394 XThR.Tn[14].t41 VGND 0.01991f
C15395 XThR.Tn[14].t65 VGND 0.02096f
C15396 XThR.Tn[14].n63 VGND 0.05206f
C15397 XThR.Tn[14].t23 VGND 0.01991f
C15398 XThR.Tn[14].t46 VGND 0.02096f
C15399 XThR.Tn[14].n64 VGND 0.05204f
C15400 XThR.Tn[14].n65 VGND 0.04002f
C15401 XThR.Tn[14].n66 VGND 0.00763f
C15402 XThR.Tn[14].n67 VGND 0.11947f
C15403 XThR.Tn[14].t72 VGND 0.01991f
C15404 XThR.Tn[14].t22 VGND 0.02096f
C15405 XThR.Tn[14].n68 VGND 0.05206f
C15406 XThR.Tn[14].t55 VGND 0.01991f
C15407 XThR.Tn[14].t64 VGND 0.02096f
C15408 XThR.Tn[14].n69 VGND 0.05204f
C15409 XThR.Tn[14].n70 VGND 0.04002f
C15410 XThR.Tn[14].n71 VGND 0.00763f
C15411 XThR.Tn[14].n72 VGND 0.11947f
C15412 XThR.Tn[14].t27 VGND 0.01991f
C15413 XThR.Tn[14].t40 VGND 0.02096f
C15414 XThR.Tn[14].n73 VGND 0.05206f
C15415 XThR.Tn[14].t71 VGND 0.01991f
C15416 XThR.Tn[14].t21 VGND 0.02096f
C15417 XThR.Tn[14].n74 VGND 0.05204f
C15418 XThR.Tn[14].n75 VGND 0.04002f
C15419 XThR.Tn[14].n76 VGND 0.00763f
C15420 XThR.Tn[14].n77 VGND 0.11947f
C15421 XThR.Tn[14].t48 VGND 0.01991f
C15422 XThR.Tn[14].t30 VGND 0.02096f
C15423 XThR.Tn[14].n78 VGND 0.05206f
C15424 XThR.Tn[14].t31 VGND 0.01991f
C15425 XThR.Tn[14].t14 VGND 0.02096f
C15426 XThR.Tn[14].n79 VGND 0.05204f
C15427 XThR.Tn[14].n80 VGND 0.04002f
C15428 XThR.Tn[14].n81 VGND 0.00763f
C15429 XThR.Tn[14].n82 VGND 0.11947f
C15430 XThR.Tn[14].n83 VGND 0.10913f
C15431 XThR.Tn[14].n84 VGND 0.43837f
C15432 XThR.Tn[14].t2 VGND 0.0245f
C15433 XThR.Tn[14].t3 VGND 0.0245f
C15434 XThR.Tn[14].n85 VGND 0.05293f
C15435 XThR.Tn[14].t0 VGND 0.0245f
C15436 XThR.Tn[14].t1 VGND 0.0245f
C15437 XThR.Tn[14].n86 VGND 0.08056f
C15438 XThR.Tn[14].n87 VGND 0.22368f
C15439 XThR.Tn[14].n88 VGND 0.01102f
C15440 XThC.Tn[10].t1 VGND 0.013f
C15441 XThC.Tn[10].t5 VGND 0.013f
C15442 XThC.Tn[10].n0 VGND 0.03241f
C15443 XThC.Tn[10].t7 VGND 0.013f
C15444 XThC.Tn[10].t2 VGND 0.013f
C15445 XThC.Tn[10].n1 VGND 0.02599f
C15446 XThC.Tn[10].n2 VGND 0.06539f
C15447 XThC.Tn[10].n3 VGND 0.02837f
C15448 XThC.Tn[10].t41 VGND 0.01625f
C15449 XThC.Tn[10].t22 VGND 0.01711f
C15450 XThC.Tn[10].n4 VGND 0.0425f
C15451 XThC.Tn[10].n5 VGND 0.02647f
C15452 XThC.Tn[10].n6 VGND 0.08577f
C15453 XThC.Tn[10].t19 VGND 0.01625f
C15454 XThC.Tn[10].t32 VGND 0.01711f
C15455 XThC.Tn[10].n7 VGND 0.0425f
C15456 XThC.Tn[10].n8 VGND 0.02647f
C15457 XThC.Tn[10].n9 VGND 0.08601f
C15458 XThC.Tn[10].n10 VGND 0.14361f
C15459 XThC.Tn[10].t31 VGND 0.01625f
C15460 XThC.Tn[10].t13 VGND 0.01711f
C15461 XThC.Tn[10].n11 VGND 0.0425f
C15462 XThC.Tn[10].n12 VGND 0.02647f
C15463 XThC.Tn[10].n13 VGND 0.08601f
C15464 XThC.Tn[10].n14 VGND 0.14361f
C15465 XThC.Tn[10].t33 VGND 0.01625f
C15466 XThC.Tn[10].t14 VGND 0.01711f
C15467 XThC.Tn[10].n15 VGND 0.0425f
C15468 XThC.Tn[10].n16 VGND 0.02647f
C15469 XThC.Tn[10].n17 VGND 0.08601f
C15470 XThC.Tn[10].n18 VGND 0.14361f
C15471 XThC.Tn[10].t43 VGND 0.01625f
C15472 XThC.Tn[10].t25 VGND 0.01711f
C15473 XThC.Tn[10].n19 VGND 0.0425f
C15474 XThC.Tn[10].n20 VGND 0.02647f
C15475 XThC.Tn[10].n21 VGND 0.08601f
C15476 XThC.Tn[10].n22 VGND 0.14361f
C15477 XThC.Tn[10].t21 VGND 0.01625f
C15478 XThC.Tn[10].t36 VGND 0.01711f
C15479 XThC.Tn[10].n23 VGND 0.0425f
C15480 XThC.Tn[10].n24 VGND 0.02647f
C15481 XThC.Tn[10].n25 VGND 0.08601f
C15482 XThC.Tn[10].n26 VGND 0.14361f
C15483 XThC.Tn[10].t34 VGND 0.01625f
C15484 XThC.Tn[10].t15 VGND 0.01711f
C15485 XThC.Tn[10].n27 VGND 0.0425f
C15486 XThC.Tn[10].n28 VGND 0.02647f
C15487 XThC.Tn[10].n29 VGND 0.08601f
C15488 XThC.Tn[10].n30 VGND 0.14361f
C15489 XThC.Tn[10].t12 VGND 0.01625f
C15490 XThC.Tn[10].t26 VGND 0.01711f
C15491 XThC.Tn[10].n31 VGND 0.0425f
C15492 XThC.Tn[10].n32 VGND 0.02647f
C15493 XThC.Tn[10].n33 VGND 0.08601f
C15494 XThC.Tn[10].n34 VGND 0.14361f
C15495 XThC.Tn[10].t16 VGND 0.01625f
C15496 XThC.Tn[10].t28 VGND 0.01711f
C15497 XThC.Tn[10].n35 VGND 0.0425f
C15498 XThC.Tn[10].n36 VGND 0.02647f
C15499 XThC.Tn[10].n37 VGND 0.08601f
C15500 XThC.Tn[10].n38 VGND 0.14361f
C15501 XThC.Tn[10].t23 VGND 0.01625f
C15502 XThC.Tn[10].t37 VGND 0.01711f
C15503 XThC.Tn[10].n39 VGND 0.0425f
C15504 XThC.Tn[10].n40 VGND 0.02647f
C15505 XThC.Tn[10].n41 VGND 0.08601f
C15506 XThC.Tn[10].n42 VGND 0.14361f
C15507 XThC.Tn[10].t35 VGND 0.01625f
C15508 XThC.Tn[10].t17 VGND 0.01711f
C15509 XThC.Tn[10].n43 VGND 0.0425f
C15510 XThC.Tn[10].n44 VGND 0.02647f
C15511 XThC.Tn[10].n45 VGND 0.08601f
C15512 XThC.Tn[10].n46 VGND 0.14361f
C15513 XThC.Tn[10].t38 VGND 0.01625f
C15514 XThC.Tn[10].t20 VGND 0.01711f
C15515 XThC.Tn[10].n47 VGND 0.0425f
C15516 XThC.Tn[10].n48 VGND 0.02647f
C15517 XThC.Tn[10].n49 VGND 0.08601f
C15518 XThC.Tn[10].n50 VGND 0.14361f
C15519 XThC.Tn[10].t24 VGND 0.01625f
C15520 XThC.Tn[10].t39 VGND 0.01711f
C15521 XThC.Tn[10].n51 VGND 0.0425f
C15522 XThC.Tn[10].n52 VGND 0.02647f
C15523 XThC.Tn[10].n53 VGND 0.08601f
C15524 XThC.Tn[10].n54 VGND 0.14361f
C15525 XThC.Tn[10].t27 VGND 0.01625f
C15526 XThC.Tn[10].t40 VGND 0.01711f
C15527 XThC.Tn[10].n55 VGND 0.0425f
C15528 XThC.Tn[10].n56 VGND 0.02647f
C15529 XThC.Tn[10].n57 VGND 0.08601f
C15530 XThC.Tn[10].n58 VGND 0.14361f
C15531 XThC.Tn[10].t29 VGND 0.01625f
C15532 XThC.Tn[10].t42 VGND 0.01711f
C15533 XThC.Tn[10].n59 VGND 0.0425f
C15534 XThC.Tn[10].n60 VGND 0.02647f
C15535 XThC.Tn[10].n61 VGND 0.08601f
C15536 XThC.Tn[10].n62 VGND 0.14361f
C15537 XThC.Tn[10].t18 VGND 0.01625f
C15538 XThC.Tn[10].t30 VGND 0.01711f
C15539 XThC.Tn[10].n63 VGND 0.0425f
C15540 XThC.Tn[10].n64 VGND 0.02647f
C15541 XThC.Tn[10].n65 VGND 0.08601f
C15542 XThC.Tn[10].n66 VGND 0.14361f
C15543 XThC.Tn[10].n67 VGND 0.61605f
C15544 XThC.Tn[10].n68 VGND 0.23449f
C15545 XThC.Tn[10].t4 VGND 0.01999f
C15546 XThC.Tn[10].t3 VGND 0.01999f
C15547 XThC.Tn[10].n69 VGND 0.0432f
C15548 XThC.Tn[10].t6 VGND 0.01999f
C15549 XThC.Tn[10].t9 VGND 0.01999f
C15550 XThC.Tn[10].n70 VGND 0.06575f
C15551 XThC.Tn[10].n71 VGND 0.1827f
C15552 XThC.Tn[10].n72 VGND 0.02873f
C15553 XThC.Tn[10].t11 VGND 0.01999f
C15554 XThC.Tn[10].t10 VGND 0.01999f
C15555 XThC.Tn[10].n73 VGND 0.04445f
C15556 XThC.Tn[10].t0 VGND 0.01999f
C15557 XThC.Tn[10].t8 VGND 0.01999f
C15558 XThC.Tn[10].n74 VGND 0.06071f
C15559 XThC.Tn[10].n75 VGND 0.19782f
C15560 VPWR.n0 VGND 0.04733f
C15561 VPWR.t181 VGND 0.29931f
C15562 VPWR.t1348 VGND 0.13245f
C15563 VPWR.t1007 VGND 0.38188f
C15564 VPWR.t1001 VGND 0.14449f
C15565 VPWR.t0 VGND 0.14449f
C15566 VPWR.t346 VGND 0.14449f
C15567 VPWR.t403 VGND 0.14449f
C15568 VPWR.t1856 VGND 0.14449f
C15569 VPWR.t1852 VGND 0.14449f
C15570 VPWR.t407 VGND 0.10149f
C15571 VPWR.n1 VGND 0.1844f
C15572 VPWR.n2 VGND 0.09757f
C15573 VPWR.t1349 VGND 0.05772f
C15574 VPWR.n3 VGND 0.00929f
C15575 VPWR.t408 VGND 0.01447f
C15576 VPWR.t1853 VGND 0.01447f
C15577 VPWR.n4 VGND 0.03177f
C15578 VPWR.t1857 VGND 0.01447f
C15579 VPWR.t404 VGND 0.01447f
C15580 VPWR.n5 VGND 0.03172f
C15581 VPWR.n6 VGND 0.06514f
C15582 VPWR.n7 VGND 0.18361f
C15583 VPWR.n8 VGND 0.05813f
C15584 VPWR.n9 VGND 0.0427f
C15585 VPWR.n10 VGND 0.07653f
C15586 VPWR.n11 VGND 0.0113f
C15587 VPWR.n12 VGND 0.01646f
C15588 VPWR.n13 VGND 0.01929f
C15589 VPWR.n14 VGND 0.02829f
C15590 VPWR.n15 VGND 0.08565f
C15591 VPWR.n16 VGND 0.01221f
C15592 VPWR.t182 VGND 0.05771f
C15593 VPWR.n17 VGND 0.07422f
C15594 VPWR.n18 VGND 0.33894f
C15595 VPWR.n19 VGND 0.98833f
C15596 VPWR.n20 VGND 0.32171f
C15597 VPWR.n21 VGND 1.02579f
C15598 VPWR.n22 VGND 0.14024f
C15599 VPWR.t2031 VGND 0.01176f
C15600 VPWR.t914 VGND 0.01238f
C15601 VPWR.n23 VGND 0.03075f
C15602 VPWR.n24 VGND 0.07933f
C15603 VPWR.t1976 VGND 0.01176f
C15604 VPWR.t803 VGND 0.01238f
C15605 VPWR.n25 VGND 0.03075f
C15606 VPWR.n26 VGND 0.16128f
C15607 VPWR.t2012 VGND 0.01176f
C15608 VPWR.t945 VGND 0.01238f
C15609 VPWR.n27 VGND 0.03075f
C15610 VPWR.n28 VGND 0.12856f
C15611 VPWR.t1953 VGND 0.01176f
C15612 VPWR.t844 VGND 0.01238f
C15613 VPWR.n29 VGND 0.03075f
C15614 VPWR.n30 VGND 0.12856f
C15615 VPWR.t2013 VGND 0.01176f
C15616 VPWR.t669 VGND 0.01238f
C15617 VPWR.n31 VGND 0.03075f
C15618 VPWR.n32 VGND 0.12856f
C15619 VPWR.t2060 VGND 0.01176f
C15620 VPWR.t835 VGND 0.01238f
C15621 VPWR.n33 VGND 0.03075f
C15622 VPWR.n34 VGND 0.12856f
C15623 VPWR.t2042 VGND 0.01176f
C15624 VPWR.t733 VGND 0.01238f
C15625 VPWR.n35 VGND 0.03075f
C15626 VPWR.n36 VGND 0.12856f
C15627 VPWR.t1937 VGND 0.01176f
C15628 VPWR.t773 VGND 0.01238f
C15629 VPWR.n37 VGND 0.03075f
C15630 VPWR.n38 VGND 0.12856f
C15631 VPWR.t1979 VGND 0.01176f
C15632 VPWR.t672 VGND 0.01238f
C15633 VPWR.n39 VGND 0.03075f
C15634 VPWR.n40 VGND 0.12856f
C15635 VPWR.t2024 VGND 0.01176f
C15636 VPWR.t937 VGND 0.01238f
C15637 VPWR.n41 VGND 0.03075f
C15638 VPWR.n42 VGND 0.12856f
C15639 VPWR.t1969 VGND 0.01176f
C15640 VPWR.t819 VGND 0.01238f
C15641 VPWR.n43 VGND 0.03075f
C15642 VPWR.n44 VGND 0.12856f
C15643 VPWR.t2045 VGND 0.01176f
C15644 VPWR.t985 VGND 0.01238f
C15645 VPWR.n45 VGND 0.03075f
C15646 VPWR.n46 VGND 0.12856f
C15647 VPWR.t1941 VGND 0.01176f
C15648 VPWR.t765 VGND 0.01238f
C15649 VPWR.n47 VGND 0.03075f
C15650 VPWR.n48 VGND 0.12856f
C15651 VPWR.t2017 VGND 0.01176f
C15652 VPWR.t663 VGND 0.01238f
C15653 VPWR.n49 VGND 0.03075f
C15654 VPWR.n50 VGND 0.12856f
C15655 VPWR.t2064 VGND 0.01176f
C15656 VPWR.t931 VGND 0.01238f
C15657 VPWR.n51 VGND 0.03075f
C15658 VPWR.n52 VGND 0.12856f
C15659 VPWR.t1970 VGND 0.01176f
C15660 VPWR.t977 VGND 0.01238f
C15661 VPWR.n53 VGND 0.03075f
C15662 VPWR.n54 VGND 0.1393f
C15663 VPWR.n55 VGND 0.11657f
C15664 VPWR.t871 VGND 0.03709f
C15665 VPWR.t840 VGND 0.0299f
C15666 VPWR.n56 VGND 0.09693f
C15667 VPWR.t755 VGND 0.09401f
C15668 VPWR.t761 VGND 0.03709f
C15669 VPWR.t756 VGND 0.0299f
C15670 VPWR.n57 VGND 0.09693f
C15671 VPWR.n58 VGND 0.0313f
C15672 VPWR.n59 VGND 0.14051f
C15673 VPWR.n60 VGND 0.14051f
C15674 VPWR.n61 VGND 0.0313f
C15675 VPWR.t622 VGND 0.03709f
C15676 VPWR.t617 VGND 0.0299f
C15677 VPWR.n62 VGND 0.09693f
C15678 VPWR.t975 VGND 0.09401f
C15679 VPWR.t882 VGND 0.03709f
C15680 VPWR.t976 VGND 0.0299f
C15681 VPWR.n63 VGND 0.09693f
C15682 VPWR.n64 VGND 0.0313f
C15683 VPWR.n65 VGND 0.14051f
C15684 VPWR.n66 VGND 0.14051f
C15685 VPWR.n67 VGND 0.0313f
C15686 VPWR.t851 VGND 0.03709f
C15687 VPWR.t843 VGND 0.0299f
C15688 VPWR.n68 VGND 0.09693f
C15689 VPWR.t710 VGND 0.09401f
C15690 VPWR.t716 VGND 0.03709f
C15691 VPWR.t711 VGND 0.0299f
C15692 VPWR.n69 VGND 0.09693f
C15693 VPWR.n70 VGND 0.0313f
C15694 VPWR.n71 VGND 0.14051f
C15695 VPWR.n72 VGND 0.14051f
C15696 VPWR.n73 VGND 0.0313f
C15697 VPWR.t973 VGND 0.03709f
C15698 VPWR.t677 VGND 0.0299f
C15699 VPWR.n74 VGND 0.09693f
C15700 VPWR.t828 VGND 0.09401f
C15701 VPWR.t832 VGND 0.03709f
C15702 VPWR.t829 VGND 0.0299f
C15703 VPWR.n75 VGND 0.09693f
C15704 VPWR.n76 VGND 0.0313f
C15705 VPWR.n77 VGND 0.14051f
C15706 VPWR.n78 VGND 0.14051f
C15707 VPWR.n79 VGND 0.0313f
C15708 VPWR.t796 VGND 0.03709f
C15709 VPWR.t813 VGND 0.0299f
C15710 VPWR.n80 VGND 0.09693f
C15711 VPWR.t694 VGND 0.09401f
C15712 VPWR.t700 VGND 0.03709f
C15713 VPWR.t695 VGND 0.0299f
C15714 VPWR.n81 VGND 0.09693f
C15715 VPWR.n82 VGND 0.0313f
C15716 VPWR.n83 VGND 0.14051f
C15717 VPWR.n84 VGND 0.14051f
C15718 VPWR.n85 VGND 0.0313f
C15719 VPWR.t927 VGND 0.03709f
C15720 VPWR.t942 VGND 0.0299f
C15721 VPWR.n86 VGND 0.09693f
C15722 VPWR.t902 VGND 0.09401f
C15723 VPWR.t908 VGND 0.03709f
C15724 VPWR.t903 VGND 0.0299f
C15725 VPWR.n87 VGND 0.09693f
C15726 VPWR.n88 VGND 0.0313f
C15727 VPWR.n89 VGND 0.14051f
C15728 VPWR.n90 VGND 0.14051f
C15729 VPWR.n91 VGND 0.0313f
C15730 VPWR.t690 VGND 0.03709f
C15731 VPWR.t685 VGND 0.0299f
C15732 VPWR.n92 VGND 0.09693f
C15733 VPWR.t646 VGND 0.09401f
C15734 VPWR.t652 VGND 0.03709f
C15735 VPWR.t647 VGND 0.0299f
C15736 VPWR.n93 VGND 0.09693f
C15737 VPWR.n94 VGND 0.0313f
C15738 VPWR.n95 VGND 0.14051f
C15739 VPWR.n96 VGND 0.14051f
C15740 VPWR.n97 VGND 0.0313f
C15741 VPWR.t930 VGND 0.03709f
C15742 VPWR.t635 VGND 0.0299f
C15743 VPWR.n98 VGND 0.09693f
C15744 VPWR.t782 VGND 0.14747f
C15745 VPWR.t780 VGND 0.08295f
C15746 VPWR.t777 VGND 0.09401f
C15747 VPWR.t783 VGND 0.03709f
C15748 VPWR.t778 VGND 0.0299f
C15749 VPWR.n99 VGND 0.09693f
C15750 VPWR.t2041 VGND 0.01176f
C15751 VPWR.t633 VGND 0.01238f
C15752 VPWR.n100 VGND 0.03074f
C15753 VPWR.n101 VGND 0.02885f
C15754 VPWR.n102 VGND 0.01916f
C15755 VPWR.t1983 VGND 0.01176f
C15756 VPWR.t781 VGND 0.01238f
C15757 VPWR.n103 VGND 0.03075f
C15758 VPWR.t1985 VGND 0.01176f
C15759 VPWR.t776 VGND 0.01238f
C15760 VPWR.n104 VGND 0.03074f
C15761 VPWR.n105 VGND 0.02885f
C15762 VPWR.n106 VGND 0.02485f
C15763 VPWR.t1984 VGND 0.01176f
C15764 VPWR.t779 VGND 0.01238f
C15765 VPWR.n107 VGND 0.03074f
C15766 VPWR.n108 VGND 0.02256f
C15767 VPWR.n109 VGND 0.01916f
C15768 VPWR.n110 VGND 0.03605f
C15769 VPWR.t1956 VGND 0.01176f
C15770 VPWR.t838 VGND 0.01238f
C15771 VPWR.n111 VGND 0.03074f
C15772 VPWR.n112 VGND 0.02885f
C15773 VPWR.t1954 VGND 0.01176f
C15774 VPWR.t869 VGND 0.01238f
C15775 VPWR.n113 VGND 0.03074f
C15776 VPWR.n114 VGND 0.04185f
C15777 VPWR.n115 VGND 0.02485f
C15778 VPWR.t1955 VGND 0.01176f
C15779 VPWR.t867 VGND 0.01238f
C15780 VPWR.n116 VGND 0.03074f
C15781 VPWR.n117 VGND 0.02256f
C15782 VPWR.n118 VGND 0.01916f
C15783 VPWR.n119 VGND 0.03491f
C15784 VPWR.t1997 VGND 0.01176f
C15785 VPWR.t754 VGND 0.01238f
C15786 VPWR.n120 VGND 0.03074f
C15787 VPWR.n121 VGND 0.02885f
C15788 VPWR.t1995 VGND 0.01176f
C15789 VPWR.t759 VGND 0.01238f
C15790 VPWR.n122 VGND 0.03074f
C15791 VPWR.n123 VGND 0.04185f
C15792 VPWR.n124 VGND 0.02485f
C15793 VPWR.t1996 VGND 0.01176f
C15794 VPWR.t757 VGND 0.01238f
C15795 VPWR.n125 VGND 0.03074f
C15796 VPWR.n126 VGND 0.02256f
C15797 VPWR.n127 VGND 0.01916f
C15798 VPWR.n128 VGND 0.03332f
C15799 VPWR.n129 VGND 0.21371f
C15800 VPWR.t2054 VGND 0.01176f
C15801 VPWR.t615 VGND 0.01238f
C15802 VPWR.n130 VGND 0.03074f
C15803 VPWR.n131 VGND 0.02885f
C15804 VPWR.t2052 VGND 0.01176f
C15805 VPWR.t620 VGND 0.01238f
C15806 VPWR.n132 VGND 0.03074f
C15807 VPWR.n133 VGND 0.04185f
C15808 VPWR.n134 VGND 0.02485f
C15809 VPWR.t2053 VGND 0.01176f
C15810 VPWR.t618 VGND 0.01238f
C15811 VPWR.n135 VGND 0.03074f
C15812 VPWR.n136 VGND 0.02256f
C15813 VPWR.n137 VGND 0.01916f
C15814 VPWR.n138 VGND 0.03332f
C15815 VPWR.n139 VGND 0.17759f
C15816 VPWR.t2061 VGND 0.01176f
C15817 VPWR.t974 VGND 0.01238f
C15818 VPWR.n140 VGND 0.03074f
C15819 VPWR.n141 VGND 0.02885f
C15820 VPWR.t1950 VGND 0.01176f
C15821 VPWR.t880 VGND 0.01238f
C15822 VPWR.n142 VGND 0.03074f
C15823 VPWR.n143 VGND 0.04185f
C15824 VPWR.n144 VGND 0.02485f
C15825 VPWR.t2059 VGND 0.01176f
C15826 VPWR.t980 VGND 0.01238f
C15827 VPWR.n145 VGND 0.03074f
C15828 VPWR.n146 VGND 0.02256f
C15829 VPWR.n147 VGND 0.01916f
C15830 VPWR.n148 VGND 0.03332f
C15831 VPWR.n149 VGND 0.17759f
C15832 VPWR.t1961 VGND 0.01176f
C15833 VPWR.t841 VGND 0.01238f
C15834 VPWR.n150 VGND 0.03074f
C15835 VPWR.n151 VGND 0.02885f
C15836 VPWR.t1959 VGND 0.01176f
C15837 VPWR.t849 VGND 0.01238f
C15838 VPWR.n152 VGND 0.03074f
C15839 VPWR.n153 VGND 0.04185f
C15840 VPWR.n154 VGND 0.02485f
C15841 VPWR.t1960 VGND 0.01176f
C15842 VPWR.t847 VGND 0.01238f
C15843 VPWR.n155 VGND 0.03074f
C15844 VPWR.n156 VGND 0.02256f
C15845 VPWR.n157 VGND 0.01916f
C15846 VPWR.n158 VGND 0.03332f
C15847 VPWR.n159 VGND 0.17759f
C15848 VPWR.t2011 VGND 0.01176f
C15849 VPWR.t709 VGND 0.01238f
C15850 VPWR.n160 VGND 0.03074f
C15851 VPWR.n161 VGND 0.02885f
C15852 VPWR.t2009 VGND 0.01176f
C15853 VPWR.t714 VGND 0.01238f
C15854 VPWR.n162 VGND 0.03074f
C15855 VPWR.n163 VGND 0.04185f
C15856 VPWR.n164 VGND 0.02485f
C15857 VPWR.t2010 VGND 0.01176f
C15858 VPWR.t712 VGND 0.01238f
C15859 VPWR.n165 VGND 0.03074f
C15860 VPWR.n166 VGND 0.02256f
C15861 VPWR.n167 VGND 0.01916f
C15862 VPWR.n168 VGND 0.03332f
C15863 VPWR.n169 VGND 0.17759f
C15864 VPWR.t2026 VGND 0.01176f
C15865 VPWR.t675 VGND 0.01238f
C15866 VPWR.n170 VGND 0.03074f
C15867 VPWR.n171 VGND 0.02885f
C15868 VPWR.t2062 VGND 0.01176f
C15869 VPWR.t971 VGND 0.01238f
C15870 VPWR.n172 VGND 0.03074f
C15871 VPWR.n173 VGND 0.04185f
C15872 VPWR.n174 VGND 0.02485f
C15873 VPWR.t2063 VGND 0.01176f
C15874 VPWR.t969 VGND 0.01238f
C15875 VPWR.n175 VGND 0.03074f
C15876 VPWR.n176 VGND 0.02256f
C15877 VPWR.n177 VGND 0.01916f
C15878 VPWR.n178 VGND 0.03332f
C15879 VPWR.n179 VGND 0.17759f
C15880 VPWR.t1968 VGND 0.01176f
C15881 VPWR.t827 VGND 0.01238f
C15882 VPWR.n180 VGND 0.03074f
C15883 VPWR.n181 VGND 0.02885f
C15884 VPWR.t1966 VGND 0.01176f
C15885 VPWR.t830 VGND 0.01238f
C15886 VPWR.n182 VGND 0.03074f
C15887 VPWR.n183 VGND 0.04185f
C15888 VPWR.n184 VGND 0.02485f
C15889 VPWR.t1967 VGND 0.01176f
C15890 VPWR.t833 VGND 0.01238f
C15891 VPWR.n185 VGND 0.03074f
C15892 VPWR.n186 VGND 0.02256f
C15893 VPWR.n187 VGND 0.01916f
C15894 VPWR.n188 VGND 0.03332f
C15895 VPWR.n189 VGND 0.17759f
C15896 VPWR.t1975 VGND 0.01176f
C15897 VPWR.t811 VGND 0.01238f
C15898 VPWR.n190 VGND 0.03074f
C15899 VPWR.n191 VGND 0.02885f
C15900 VPWR.t1977 VGND 0.01176f
C15901 VPWR.t794 VGND 0.01238f
C15902 VPWR.n192 VGND 0.03074f
C15903 VPWR.n193 VGND 0.04185f
C15904 VPWR.n194 VGND 0.02485f
C15905 VPWR.t1978 VGND 0.01176f
C15906 VPWR.t792 VGND 0.01238f
C15907 VPWR.n195 VGND 0.03074f
C15908 VPWR.n196 VGND 0.02256f
C15909 VPWR.n197 VGND 0.01916f
C15910 VPWR.n198 VGND 0.03332f
C15911 VPWR.n199 VGND 0.17759f
C15912 VPWR.t2016 VGND 0.01176f
C15913 VPWR.t693 VGND 0.01238f
C15914 VPWR.n200 VGND 0.03074f
C15915 VPWR.n201 VGND 0.02885f
C15916 VPWR.t2014 VGND 0.01176f
C15917 VPWR.t698 VGND 0.01238f
C15918 VPWR.n202 VGND 0.03074f
C15919 VPWR.n203 VGND 0.04185f
C15920 VPWR.n204 VGND 0.02485f
C15921 VPWR.t2015 VGND 0.01176f
C15922 VPWR.t696 VGND 0.01238f
C15923 VPWR.n205 VGND 0.03074f
C15924 VPWR.n206 VGND 0.02256f
C15925 VPWR.n207 VGND 0.01916f
C15926 VPWR.n208 VGND 0.03332f
C15927 VPWR.n209 VGND 0.17759f
C15928 VPWR.t1927 VGND 0.01176f
C15929 VPWR.t940 VGND 0.01238f
C15930 VPWR.n210 VGND 0.03074f
C15931 VPWR.n211 VGND 0.02885f
C15932 VPWR.t1933 VGND 0.01176f
C15933 VPWR.t925 VGND 0.01238f
C15934 VPWR.n212 VGND 0.03074f
C15935 VPWR.n213 VGND 0.04185f
C15936 VPWR.n214 VGND 0.02485f
C15937 VPWR.t1926 VGND 0.01176f
C15938 VPWR.t943 VGND 0.01238f
C15939 VPWR.n215 VGND 0.03074f
C15940 VPWR.n216 VGND 0.02256f
C15941 VPWR.n217 VGND 0.01916f
C15942 VPWR.n218 VGND 0.03332f
C15943 VPWR.n219 VGND 0.17759f
C15944 VPWR.t1936 VGND 0.01176f
C15945 VPWR.t901 VGND 0.01238f
C15946 VPWR.n220 VGND 0.03074f
C15947 VPWR.n221 VGND 0.02885f
C15948 VPWR.t1934 VGND 0.01176f
C15949 VPWR.t906 VGND 0.01238f
C15950 VPWR.n222 VGND 0.03074f
C15951 VPWR.n223 VGND 0.04185f
C15952 VPWR.n224 VGND 0.02485f
C15953 VPWR.t1935 VGND 0.01176f
C15954 VPWR.t904 VGND 0.01238f
C15955 VPWR.n225 VGND 0.03074f
C15956 VPWR.n226 VGND 0.02256f
C15957 VPWR.n227 VGND 0.01916f
C15958 VPWR.n228 VGND 0.03332f
C15959 VPWR.n229 VGND 0.17759f
C15960 VPWR.t2023 VGND 0.01176f
C15961 VPWR.t683 VGND 0.01238f
C15962 VPWR.n230 VGND 0.03074f
C15963 VPWR.n231 VGND 0.02885f
C15964 VPWR.t2021 VGND 0.01176f
C15965 VPWR.t688 VGND 0.01238f
C15966 VPWR.n232 VGND 0.03074f
C15967 VPWR.n233 VGND 0.04185f
C15968 VPWR.n234 VGND 0.02485f
C15969 VPWR.t2022 VGND 0.01176f
C15970 VPWR.t686 VGND 0.01238f
C15971 VPWR.n235 VGND 0.03074f
C15972 VPWR.n236 VGND 0.02256f
C15973 VPWR.n237 VGND 0.01916f
C15974 VPWR.n238 VGND 0.03332f
C15975 VPWR.n239 VGND 0.17759f
C15976 VPWR.t2035 VGND 0.01176f
C15977 VPWR.t645 VGND 0.01238f
C15978 VPWR.n240 VGND 0.03074f
C15979 VPWR.n241 VGND 0.02885f
C15980 VPWR.t2033 VGND 0.01176f
C15981 VPWR.t650 VGND 0.01238f
C15982 VPWR.n242 VGND 0.03074f
C15983 VPWR.n243 VGND 0.04185f
C15984 VPWR.n244 VGND 0.02485f
C15985 VPWR.t2034 VGND 0.01176f
C15986 VPWR.t648 VGND 0.01238f
C15987 VPWR.n245 VGND 0.03074f
C15988 VPWR.n246 VGND 0.02256f
C15989 VPWR.n247 VGND 0.01916f
C15990 VPWR.n248 VGND 0.03332f
C15991 VPWR.n249 VGND 0.17759f
C15992 VPWR.n250 VGND 0.23958f
C15993 VPWR.n251 VGND 0.03332f
C15994 VPWR.t2040 VGND 0.01176f
C15995 VPWR.t636 VGND 0.01238f
C15996 VPWR.n252 VGND 0.03074f
C15997 VPWR.n253 VGND 0.02256f
C15998 VPWR.n254 VGND 0.02485f
C15999 VPWR.t1932 VGND 0.01176f
C16000 VPWR.t928 VGND 0.01238f
C16001 VPWR.n255 VGND 0.03074f
C16002 VPWR.n256 VGND 0.04185f
C16003 VPWR.n257 VGND 0.0313f
C16004 VPWR.t1221 VGND 0.03709f
C16005 VPWR.t1024 VGND 0.0299f
C16006 VPWR.n258 VGND 0.09693f
C16007 VPWR.t1220 VGND 0.14747f
C16008 VPWR.t1664 VGND 0.08295f
C16009 VPWR.t1023 VGND 0.09401f
C16010 VPWR.t474 VGND 0.03709f
C16011 VPWR.t979 VGND 0.0299f
C16012 VPWR.n259 VGND 0.09693f
C16013 VPWR.n260 VGND 0.01815f
C16014 VPWR.n261 VGND 0.08265f
C16015 VPWR.t978 VGND 0.14528f
C16016 VPWR.t1311 VGND 0.08295f
C16017 VPWR.t473 VGND 0.11982f
C16018 VPWR.t1087 VGND 0.03709f
C16019 VPWR.t470 VGND 0.0299f
C16020 VPWR.n262 VGND 0.09693f
C16021 VPWR.n263 VGND 0.01815f
C16022 VPWR.n264 VGND -0.00319f
C16023 VPWR.n265 VGND 0.09471f
C16024 VPWR.t469 VGND 0.09401f
C16025 VPWR.t1665 VGND 0.08295f
C16026 VPWR.t1086 VGND 0.11982f
C16027 VPWR.t1115 VGND 0.03709f
C16028 VPWR.t1651 VGND 0.0299f
C16029 VPWR.n266 VGND 0.09693f
C16030 VPWR.n267 VGND 0.01815f
C16031 VPWR.n268 VGND -0.00319f
C16032 VPWR.n269 VGND 0.09471f
C16033 VPWR.t1650 VGND 0.09401f
C16034 VPWR.t1013 VGND 0.08295f
C16035 VPWR.t1114 VGND 0.11982f
C16036 VPWR.t568 VGND 0.03709f
C16037 VPWR.t1119 VGND 0.0299f
C16038 VPWR.n270 VGND 0.09693f
C16039 VPWR.n271 VGND 0.01815f
C16040 VPWR.n272 VGND -0.00319f
C16041 VPWR.n273 VGND 0.09471f
C16042 VPWR.t1118 VGND 0.09401f
C16043 VPWR.t1014 VGND 0.08295f
C16044 VPWR.t567 VGND 0.11982f
C16045 VPWR.t119 VGND 0.03709f
C16046 VPWR.t263 VGND 0.0299f
C16047 VPWR.n274 VGND 0.09693f
C16048 VPWR.n275 VGND 0.01815f
C16049 VPWR.n276 VGND -0.00319f
C16050 VPWR.n277 VGND 0.09471f
C16051 VPWR.t262 VGND 0.09401f
C16052 VPWR.t1312 VGND 0.08295f
C16053 VPWR.t118 VGND 0.11982f
C16054 VPWR.t317 VGND 0.03709f
C16055 VPWR.t99 VGND 0.0299f
C16056 VPWR.n278 VGND 0.09693f
C16057 VPWR.n279 VGND 0.01815f
C16058 VPWR.n280 VGND -0.00319f
C16059 VPWR.n281 VGND 0.09471f
C16060 VPWR.t98 VGND 0.09401f
C16061 VPWR.t1666 VGND 0.08295f
C16062 VPWR.t316 VGND 0.11982f
C16063 VPWR.t239 VGND 0.03709f
C16064 VPWR.t188 VGND 0.0299f
C16065 VPWR.n282 VGND 0.09693f
C16066 VPWR.n283 VGND 0.01815f
C16067 VPWR.n284 VGND -0.00319f
C16068 VPWR.n285 VGND 0.09471f
C16069 VPWR.t187 VGND 0.09401f
C16070 VPWR.t1015 VGND 0.08295f
C16071 VPWR.t238 VGND 0.11982f
C16072 VPWR.t1864 VGND 0.03709f
C16073 VPWR.t1892 VGND 0.0299f
C16074 VPWR.n286 VGND 0.09693f
C16075 VPWR.n287 VGND 0.01815f
C16076 VPWR.n288 VGND -0.00319f
C16077 VPWR.n289 VGND 0.09471f
C16078 VPWR.t1891 VGND 0.09401f
C16079 VPWR.t1313 VGND 0.08295f
C16080 VPWR.t1863 VGND 0.11982f
C16081 VPWR.t428 VGND 0.03709f
C16082 VPWR.t1868 VGND 0.0299f
C16083 VPWR.n290 VGND 0.09693f
C16084 VPWR.n291 VGND 0.01815f
C16085 VPWR.n292 VGND -0.00319f
C16086 VPWR.n293 VGND 0.09471f
C16087 VPWR.t1867 VGND 0.09401f
C16088 VPWR.t1663 VGND 0.08295f
C16089 VPWR.t427 VGND 0.11982f
C16090 VPWR.t1561 VGND 0.03709f
C16091 VPWR.t1457 VGND 0.0299f
C16092 VPWR.n294 VGND 0.09693f
C16093 VPWR.n295 VGND 0.01815f
C16094 VPWR.n296 VGND -0.00319f
C16095 VPWR.n297 VGND 0.09471f
C16096 VPWR.t1456 VGND 0.09401f
C16097 VPWR.t1667 VGND 0.08295f
C16098 VPWR.t1560 VGND 0.11982f
C16099 VPWR.t1529 VGND 0.03709f
C16100 VPWR.t1517 VGND 0.0299f
C16101 VPWR.n298 VGND 0.09693f
C16102 VPWR.n299 VGND 0.01815f
C16103 VPWR.n300 VGND -0.00319f
C16104 VPWR.n301 VGND 0.09471f
C16105 VPWR.t1516 VGND 0.09401f
C16106 VPWR.t1016 VGND 0.08295f
C16107 VPWR.t1528 VGND 0.11982f
C16108 VPWR.t1288 VGND 0.03709f
C16109 VPWR.t1581 VGND 0.0299f
C16110 VPWR.n302 VGND 0.09693f
C16111 VPWR.n303 VGND 0.01815f
C16112 VPWR.n304 VGND -0.00319f
C16113 VPWR.n305 VGND 0.09471f
C16114 VPWR.t1580 VGND 0.09401f
C16115 VPWR.t1043 VGND 0.08295f
C16116 VPWR.t1287 VGND 0.11982f
C16117 VPWR.t13 VGND 0.03709f
C16118 VPWR.t1469 VGND 0.0299f
C16119 VPWR.n306 VGND 0.09693f
C16120 VPWR.n307 VGND 0.01815f
C16121 VPWR.n308 VGND -0.00319f
C16122 VPWR.n309 VGND 0.09471f
C16123 VPWR.t1468 VGND 0.09401f
C16124 VPWR.t1668 VGND 0.08295f
C16125 VPWR.t12 VGND 0.11982f
C16126 VPWR.t1403 VGND 0.03709f
C16127 VPWR.t23 VGND 0.0299f
C16128 VPWR.n310 VGND 0.09693f
C16129 VPWR.n311 VGND 0.01815f
C16130 VPWR.n312 VGND -0.00319f
C16131 VPWR.n313 VGND 0.09471f
C16132 VPWR.t22 VGND 0.09401f
C16133 VPWR.t1011 VGND 0.08295f
C16134 VPWR.t1402 VGND 0.11982f
C16135 VPWR.t1245 VGND 0.03709f
C16136 VPWR.t1795 VGND 0.0299f
C16137 VPWR.n314 VGND 0.09693f
C16138 VPWR.n315 VGND 0.01815f
C16139 VPWR.n316 VGND -0.00319f
C16140 VPWR.n317 VGND 0.09471f
C16141 VPWR.t1794 VGND 0.09401f
C16142 VPWR.t1012 VGND 0.08295f
C16143 VPWR.t1244 VGND 0.11982f
C16144 VPWR.n318 VGND 0.09471f
C16145 VPWR.n319 VGND -0.00319f
C16146 VPWR.n320 VGND 0.01815f
C16147 VPWR.n321 VGND 0.14051f
C16148 VPWR.n322 VGND 1.01936f
C16149 VPWR.n323 VGND 0.14051f
C16150 VPWR.t1215 VGND 0.03709f
C16151 VPWR.t1032 VGND 0.0299f
C16152 VPWR.n324 VGND 0.09693f
C16153 VPWR.t1214 VGND 0.14747f
C16154 VPWR.t590 VGND 0.08295f
C16155 VPWR.t1031 VGND 0.09401f
C16156 VPWR.t1800 VGND 0.11982f
C16157 VPWR.t1040 VGND 0.03709f
C16158 VPWR.t1537 VGND 0.0299f
C16159 VPWR.n325 VGND 0.09693f
C16160 VPWR.n326 VGND 0.14051f
C16161 VPWR.n327 VGND 0.14051f
C16162 VPWR.t1801 VGND 0.03709f
C16163 VPWR.t43 VGND 0.0299f
C16164 VPWR.n328 VGND 0.09693f
C16165 VPWR.t492 VGND 0.08295f
C16166 VPWR.t42 VGND 0.09401f
C16167 VPWR.t1920 VGND 0.11982f
C16168 VPWR.t21 VGND 0.03709f
C16169 VPWR.t137 VGND 0.0299f
C16170 VPWR.n329 VGND 0.09693f
C16171 VPWR.n330 VGND 0.14051f
C16172 VPWR.n331 VGND 0.14051f
C16173 VPWR.t1921 VGND 0.03709f
C16174 VPWR.t1337 VGND 0.0299f
C16175 VPWR.n332 VGND 0.09693f
C16176 VPWR.t1829 VGND 0.08295f
C16177 VPWR.t1336 VGND 0.09401f
C16178 VPWR.t1810 VGND 0.11982f
C16179 VPWR.t1587 VGND 0.03709f
C16180 VPWR.t215 VGND 0.0299f
C16181 VPWR.n333 VGND 0.09693f
C16182 VPWR.n334 VGND 0.14051f
C16183 VPWR.n335 VGND 0.14051f
C16184 VPWR.t1811 VGND 0.03709f
C16185 VPWR.t273 VGND 0.0299f
C16186 VPWR.n336 VGND 0.09693f
C16187 VPWR.t490 VGND 0.08295f
C16188 VPWR.t272 VGND 0.09401f
C16189 VPWR.t499 VGND 0.11982f
C16190 VPWR.t1105 VGND 0.03709f
C16191 VPWR.t506 VGND 0.0299f
C16192 VPWR.n337 VGND 0.09693f
C16193 VPWR.n338 VGND 0.14051f
C16194 VPWR.n339 VGND 0.14051f
C16195 VPWR.t500 VGND 0.03709f
C16196 VPWR.t1904 VGND 0.0299f
C16197 VPWR.n340 VGND 0.09693f
C16198 VPWR.t588 VGND 0.08295f
C16199 VPWR.t1903 VGND 0.09401f
C16200 VPWR.t185 VGND 0.11982f
C16201 VPWR.t245 VGND 0.03709f
C16202 VPWR.t194 VGND 0.0299f
C16203 VPWR.n341 VGND 0.09693f
C16204 VPWR.n342 VGND 0.14051f
C16205 VPWR.n343 VGND 0.14051f
C16206 VPWR.t186 VGND 0.03709f
C16207 VPWR.t93 VGND 0.0299f
C16208 VPWR.n344 VGND 0.09693f
C16209 VPWR.t489 VGND 0.08295f
C16210 VPWR.t92 VGND 0.09401f
C16211 VPWR.t260 VGND 0.11982f
C16212 VPWR.t111 VGND 0.03709f
C16213 VPWR.t1509 VGND 0.0299f
C16214 VPWR.n345 VGND 0.09693f
C16215 VPWR.n346 VGND 0.14051f
C16216 VPWR.n347 VGND 0.14051f
C16217 VPWR.t261 VGND 0.03709f
C16218 VPWR.t173 VGND 0.0299f
C16219 VPWR.n348 VGND 0.09693f
C16220 VPWR.t1826 VGND 0.08295f
C16221 VPWR.t172 VGND 0.09401f
C16222 VPWR.t1140 VGND 0.11982f
C16223 VPWR.t1125 VGND 0.03709f
C16224 VPWR.t1475 VGND 0.0299f
C16225 VPWR.n349 VGND 0.09693f
C16226 VPWR.n350 VGND 0.14051f
C16227 VPWR.n351 VGND 0.14051f
C16228 VPWR.t1141 VGND 0.03709f
C16229 VPWR.t444 VGND 0.0299f
C16230 VPWR.n352 VGND 0.09693f
C16231 VPWR.t488 VGND 0.08295f
C16232 VPWR.t443 VGND 0.09401f
C16233 VPWR.t464 VGND 0.03709f
C16234 VPWR.t933 VGND 0.0299f
C16235 VPWR.n353 VGND 0.09693f
C16236 VPWR.t1382 VGND 0.03709f
C16237 VPWR.t665 VGND 0.0299f
C16238 VPWR.n354 VGND 0.09693f
C16239 VPWR.t1224 VGND 0.14747f
C16240 VPWR.t151 VGND 0.08295f
C16241 VPWR.t593 VGND 0.09401f
C16242 VPWR.t1225 VGND 0.03709f
C16243 VPWR.t594 VGND 0.0299f
C16244 VPWR.n355 VGND 0.09693f
C16245 VPWR.n356 VGND 0.01815f
C16246 VPWR.n357 VGND -0.00319f
C16247 VPWR.n358 VGND 0.09471f
C16248 VPWR.t1234 VGND 0.11982f
C16249 VPWR.t1047 VGND 0.08295f
C16250 VPWR.t1548 VGND 0.09401f
C16251 VPWR.t1235 VGND 0.03709f
C16252 VPWR.t1549 VGND 0.0299f
C16253 VPWR.n359 VGND 0.09693f
C16254 VPWR.n360 VGND 0.01815f
C16255 VPWR.n361 VGND -0.00319f
C16256 VPWR.n362 VGND 0.09471f
C16257 VPWR.t1542 VGND 0.11982f
C16258 VPWR.t1046 VGND 0.08295f
C16259 VPWR.t28 VGND 0.09401f
C16260 VPWR.t1543 VGND 0.03709f
C16261 VPWR.t29 VGND 0.0299f
C16262 VPWR.n363 VGND 0.09693f
C16263 VPWR.n364 VGND 0.01815f
C16264 VPWR.n365 VGND -0.00319f
C16265 VPWR.n366 VGND 0.09471f
C16266 VPWR.t1273 VGND 0.11982f
C16267 VPWR.t1045 VGND 0.08295f
C16268 VPWR.t551 VGND 0.09401f
C16269 VPWR.t1274 VGND 0.03709f
C16270 VPWR.t552 VGND 0.0299f
C16271 VPWR.n367 VGND 0.09693f
C16272 VPWR.n368 VGND 0.01815f
C16273 VPWR.n369 VGND -0.00319f
C16274 VPWR.n370 VGND 0.09471f
C16275 VPWR.t576 VGND 0.11982f
C16276 VPWR.t1160 VGND 0.08295f
C16277 VPWR.t1524 VGND 0.09401f
C16278 VPWR.t577 VGND 0.03709f
C16279 VPWR.t1525 VGND 0.0299f
C16280 VPWR.n371 VGND 0.09693f
C16281 VPWR.n372 VGND 0.01815f
C16282 VPWR.n373 VGND -0.00319f
C16283 VPWR.n374 VGND 0.09471f
C16284 VPWR.t1596 VGND 0.11982f
C16285 VPWR.t1159 VGND 0.08295f
C16286 VPWR.t1816 VGND 0.09401f
C16287 VPWR.t1597 VGND 0.03709f
C16288 VPWR.t1817 VGND 0.0299f
C16289 VPWR.n375 VGND 0.09693f
C16290 VPWR.n376 VGND 0.01815f
C16291 VPWR.n377 VGND -0.00319f
C16292 VPWR.n378 VGND 0.09471f
C16293 VPWR.t1550 VGND 0.11982f
C16294 VPWR.t1044 VGND 0.08295f
C16295 VPWR.t1106 VGND 0.09401f
C16296 VPWR.t1551 VGND 0.03709f
C16297 VPWR.t1107 VGND 0.0299f
C16298 VPWR.n379 VGND 0.09693f
C16299 VPWR.n380 VGND 0.01815f
C16300 VPWR.n381 VGND -0.00319f
C16301 VPWR.n382 VGND 0.09471f
C16302 VPWR.t545 VGND 0.11982f
C16303 VPWR.t999 VGND 0.08295f
C16304 VPWR.t1395 VGND 0.09401f
C16305 VPWR.t546 VGND 0.03709f
C16306 VPWR.t1396 VGND 0.0299f
C16307 VPWR.n383 VGND 0.09693f
C16308 VPWR.n384 VGND 0.01815f
C16309 VPWR.n385 VGND -0.00319f
C16310 VPWR.n386 VGND 0.09471f
C16311 VPWR.t1389 VGND 0.11982f
C16312 VPWR.t1163 VGND 0.08295f
C16313 VPWR.t374 VGND 0.09401f
C16314 VPWR.t1390 VGND 0.03709f
C16315 VPWR.t375 VGND 0.0299f
C16316 VPWR.n387 VGND 0.09693f
C16317 VPWR.n388 VGND 0.01815f
C16318 VPWR.n389 VGND -0.00319f
C16319 VPWR.n390 VGND 0.09471f
C16320 VPWR.t1182 VGND 0.11982f
C16321 VPWR.t1158 VGND 0.08295f
C16322 VPWR.t359 VGND 0.09401f
C16323 VPWR.t1183 VGND 0.03709f
C16324 VPWR.t360 VGND 0.0299f
C16325 VPWR.n391 VGND 0.09693f
C16326 VPWR.n392 VGND 0.01815f
C16327 VPWR.n393 VGND -0.00319f
C16328 VPWR.n394 VGND 0.09471f
C16329 VPWR.t353 VGND 0.11982f
C16330 VPWR.t153 VGND 0.08295f
C16331 VPWR.t104 VGND 0.09401f
C16332 VPWR.t354 VGND 0.03709f
C16333 VPWR.t105 VGND 0.0299f
C16334 VPWR.n395 VGND 0.09693f
C16335 VPWR.n396 VGND 0.01815f
C16336 VPWR.n397 VGND -0.00319f
C16337 VPWR.n398 VGND 0.09471f
C16338 VPWR.t58 VGND 0.11982f
C16339 VPWR.t1162 VGND 0.08295f
C16340 VPWR.t252 VGND 0.09401f
C16341 VPWR.t59 VGND 0.03709f
C16342 VPWR.t253 VGND 0.0299f
C16343 VPWR.n399 VGND 0.09693f
C16344 VPWR.n400 VGND 0.01815f
C16345 VPWR.n401 VGND -0.00319f
C16346 VPWR.n402 VGND 0.09471f
C16347 VPWR.t246 VGND 0.11982f
C16348 VPWR.t1049 VGND 0.08295f
C16349 VPWR.t1346 VGND 0.09401f
C16350 VPWR.t247 VGND 0.03709f
C16351 VPWR.t1347 VGND 0.0299f
C16352 VPWR.n403 VGND 0.09693f
C16353 VPWR.n404 VGND 0.01815f
C16354 VPWR.n405 VGND -0.00319f
C16355 VPWR.n406 VGND 0.09471f
C16356 VPWR.t1415 VGND 0.11982f
C16357 VPWR.t1048 VGND 0.08295f
C16358 VPWR.t1230 VGND 0.09401f
C16359 VPWR.t1416 VGND 0.03709f
C16360 VPWR.t1231 VGND 0.0299f
C16361 VPWR.n407 VGND 0.09693f
C16362 VPWR.n408 VGND 0.01815f
C16363 VPWR.n409 VGND -0.00319f
C16364 VPWR.n410 VGND 0.09471f
C16365 VPWR.t1484 VGND 0.11982f
C16366 VPWR.t152 VGND 0.08295f
C16367 VPWR.t465 VGND 0.09401f
C16368 VPWR.t1485 VGND 0.03709f
C16369 VPWR.t466 VGND 0.0299f
C16370 VPWR.n411 VGND 0.09693f
C16371 VPWR.n412 VGND 0.01815f
C16372 VPWR.n413 VGND -0.00319f
C16373 VPWR.n414 VGND 0.09471f
C16374 VPWR.t1381 VGND 0.11982f
C16375 VPWR.t1161 VGND 0.08295f
C16376 VPWR.t664 VGND 0.14528f
C16377 VPWR.n415 VGND 0.08265f
C16378 VPWR.n416 VGND 0.01815f
C16379 VPWR.n417 VGND 0.14051f
C16380 VPWR.n418 VGND 1.02579f
C16381 VPWR.n419 VGND 0.14051f
C16382 VPWR.t452 VGND 0.03709f
C16383 VPWR.t767 VGND 0.0299f
C16384 VPWR.n420 VGND 0.09693f
C16385 VPWR.t1383 VGND 0.09401f
C16386 VPWR.t1479 VGND 0.03709f
C16387 VPWR.t1384 VGND 0.0299f
C16388 VPWR.n421 VGND 0.09693f
C16389 VPWR.n422 VGND 0.14051f
C16390 VPWR.n423 VGND 0.14051f
C16391 VPWR.t1601 VGND 0.03709f
C16392 VPWR.t1083 VGND 0.0299f
C16393 VPWR.n424 VGND 0.09693f
C16394 VPWR.t1604 VGND 0.09401f
C16395 VPWR.t1495 VGND 0.03709f
C16396 VPWR.t1605 VGND 0.0299f
C16397 VPWR.n425 VGND 0.09693f
C16398 VPWR.n426 VGND 0.14051f
C16399 VPWR.n427 VGND 0.14051f
C16400 VPWR.t83 VGND 0.03709f
C16401 VPWR.t1499 VGND 0.0299f
C16402 VPWR.n428 VGND 0.09693f
C16403 VPWR.t62 VGND 0.09401f
C16404 VPWR.t1071 VGND 0.03709f
C16405 VPWR.t63 VGND 0.0299f
C16406 VPWR.n429 VGND 0.09693f
C16407 VPWR.n430 VGND 0.14051f
C16408 VPWR.n431 VGND 0.14051f
C16409 VPWR.t1910 VGND 0.03709f
C16410 VPWR.t291 VGND 0.0299f
C16411 VPWR.n432 VGND 0.09693f
C16412 VPWR.t232 VGND 0.09401f
C16413 VPWR.t510 VGND 0.03709f
C16414 VPWR.t233 VGND 0.0299f
C16415 VPWR.n433 VGND 0.09693f
C16416 VPWR.n434 VGND 0.14051f
C16417 VPWR.n435 VGND 0.14051f
C16418 VPWR.t1629 VGND 0.03709f
C16419 VPWR.t514 VGND 0.0299f
C16420 VPWR.n436 VGND 0.09693f
C16421 VPWR.t1385 VGND 0.09401f
C16422 VPWR.t221 VGND 0.03709f
C16423 VPWR.t1386 VGND 0.0299f
C16424 VPWR.n437 VGND 0.09693f
C16425 VPWR.n438 VGND 0.14051f
C16426 VPWR.n439 VGND 0.14051f
C16427 VPWR.t1711 VGND 0.03709f
C16428 VPWR.t1555 VGND 0.0299f
C16429 VPWR.n440 VGND 0.09693f
C16430 VPWR.t1714 VGND 0.09401f
C16431 VPWR.t1465 VGND 0.03709f
C16432 VPWR.t1715 VGND 0.0299f
C16433 VPWR.n441 VGND 0.09693f
C16434 VPWR.n442 VGND 0.14051f
C16435 VPWR.n443 VGND 0.14051f
C16436 VPWR.t1888 VGND 0.03709f
C16437 VPWR.t1925 VGND 0.0299f
C16438 VPWR.n444 VGND 0.09693f
C16439 VPWR.t38 VGND 0.09401f
C16440 VPWR.t1443 VGND 0.03709f
C16441 VPWR.t39 VGND 0.0299f
C16442 VPWR.n445 VGND 0.09693f
C16443 VPWR.n446 VGND 0.14051f
C16444 VPWR.n447 VGND 0.14051f
C16445 VPWR.t1847 VGND 0.03709f
C16446 VPWR.t177 VGND 0.0299f
C16447 VPWR.n448 VGND 0.09693f
C16448 VPWR.t1200 VGND 0.14747f
C16449 VPWR.t1818 VGND 0.08295f
C16450 VPWR.t1240 VGND 0.09401f
C16451 VPWR.t1201 VGND 0.03709f
C16452 VPWR.t1241 VGND 0.0299f
C16453 VPWR.n449 VGND 0.09693f
C16454 VPWR.t1223 VGND 0.03709f
C16455 VPWR.t1022 VGND 0.0299f
C16456 VPWR.n450 VGND 0.09693f
C16457 VPWR.t1222 VGND 0.14747f
C16458 VPWR.t328 VGND 0.08295f
C16459 VPWR.t1021 VGND 0.09401f
C16460 VPWR.t472 VGND 0.03709f
C16461 VPWR.t987 VGND 0.0299f
C16462 VPWR.n451 VGND 0.09693f
C16463 VPWR.n452 VGND 0.01815f
C16464 VPWR.n453 VGND 0.08265f
C16465 VPWR.t986 VGND 0.14528f
C16466 VPWR.t324 VGND 0.08295f
C16467 VPWR.t471 VGND 0.11982f
C16468 VPWR.t1085 VGND 0.03709f
C16469 VPWR.t468 VGND 0.0299f
C16470 VPWR.n454 VGND 0.09693f
C16471 VPWR.n455 VGND 0.01815f
C16472 VPWR.n456 VGND -0.00319f
C16473 VPWR.n457 VGND 0.09471f
C16474 VPWR.t467 VGND 0.09401f
C16475 VPWR.t329 VGND 0.08295f
C16476 VPWR.t1084 VGND 0.11982f
C16477 VPWR.t1113 VGND 0.03709f
C16478 VPWR.t1649 VGND 0.0299f
C16479 VPWR.n458 VGND 0.09693f
C16480 VPWR.n459 VGND 0.01815f
C16481 VPWR.n460 VGND -0.00319f
C16482 VPWR.n461 VGND 0.09471f
C16483 VPWR.t1648 VGND 0.09401f
C16484 VPWR.t366 VGND 0.08295f
C16485 VPWR.t1112 VGND 0.11982f
C16486 VPWR.t566 VGND 0.03709f
C16487 VPWR.t1117 VGND 0.0299f
C16488 VPWR.n462 VGND 0.09693f
C16489 VPWR.n463 VGND 0.01815f
C16490 VPWR.n464 VGND -0.00319f
C16491 VPWR.n465 VGND 0.09471f
C16492 VPWR.t1116 VGND 0.09401f
C16493 VPWR.t367 VGND 0.08295f
C16494 VPWR.t565 VGND 0.11982f
C16495 VPWR.t117 VGND 0.03709f
C16496 VPWR.t259 VGND 0.0299f
C16497 VPWR.n466 VGND 0.09693f
C16498 VPWR.n467 VGND 0.01815f
C16499 VPWR.n468 VGND -0.00319f
C16500 VPWR.n469 VGND 0.09471f
C16501 VPWR.t258 VGND 0.09401f
C16502 VPWR.t325 VGND 0.08295f
C16503 VPWR.t116 VGND 0.11982f
C16504 VPWR.t315 VGND 0.03709f
C16505 VPWR.t95 VGND 0.0299f
C16506 VPWR.n470 VGND 0.09693f
C16507 VPWR.n471 VGND 0.01815f
C16508 VPWR.n472 VGND -0.00319f
C16509 VPWR.n473 VGND 0.09471f
C16510 VPWR.t94 VGND 0.09401f
C16511 VPWR.t361 VGND 0.08295f
C16512 VPWR.t314 VGND 0.11982f
C16513 VPWR.t237 VGND 0.03709f
C16514 VPWR.t323 VGND 0.0299f
C16515 VPWR.n474 VGND 0.09693f
C16516 VPWR.n475 VGND 0.01815f
C16517 VPWR.n476 VGND -0.00319f
C16518 VPWR.n477 VGND 0.09471f
C16519 VPWR.t322 VGND 0.09401f
C16520 VPWR.t368 VGND 0.08295f
C16521 VPWR.t236 VGND 0.11982f
C16522 VPWR.t1862 VGND 0.03709f
C16523 VPWR.t1843 VGND 0.0299f
C16524 VPWR.n478 VGND 0.09693f
C16525 VPWR.n479 VGND 0.01815f
C16526 VPWR.n480 VGND -0.00319f
C16527 VPWR.n481 VGND 0.09471f
C16528 VPWR.t1842 VGND 0.09401f
C16529 VPWR.t326 VGND 0.08295f
C16530 VPWR.t1861 VGND 0.11982f
C16531 VPWR.t426 VGND 0.03709f
C16532 VPWR.t1866 VGND 0.0299f
C16533 VPWR.n482 VGND 0.09693f
C16534 VPWR.n483 VGND 0.01815f
C16535 VPWR.n484 VGND -0.00319f
C16536 VPWR.n485 VGND 0.09471f
C16537 VPWR.t1865 VGND 0.09401f
C16538 VPWR.t327 VGND 0.08295f
C16539 VPWR.t425 VGND 0.11982f
C16540 VPWR.t1559 VGND 0.03709f
C16541 VPWR.t1455 VGND 0.0299f
C16542 VPWR.n486 VGND 0.09693f
C16543 VPWR.n487 VGND 0.01815f
C16544 VPWR.n488 VGND -0.00319f
C16545 VPWR.n489 VGND 0.09471f
C16546 VPWR.t1454 VGND 0.09401f
C16547 VPWR.t362 VGND 0.08295f
C16548 VPWR.t1558 VGND 0.11982f
C16549 VPWR.t1527 VGND 0.03709f
C16550 VPWR.t1513 VGND 0.0299f
C16551 VPWR.n490 VGND 0.09693f
C16552 VPWR.n491 VGND 0.01815f
C16553 VPWR.n492 VGND -0.00319f
C16554 VPWR.n493 VGND 0.09471f
C16555 VPWR.t1512 VGND 0.09401f
C16556 VPWR.t369 VGND 0.08295f
C16557 VPWR.t1526 VGND 0.11982f
C16558 VPWR.t1286 VGND 0.03709f
C16559 VPWR.t1579 VGND 0.0299f
C16560 VPWR.n494 VGND 0.09693f
C16561 VPWR.n495 VGND 0.01815f
C16562 VPWR.n496 VGND -0.00319f
C16563 VPWR.n497 VGND 0.09471f
C16564 VPWR.t1578 VGND 0.09401f
C16565 VPWR.t341 VGND 0.08295f
C16566 VPWR.t1285 VGND 0.11982f
C16567 VPWR.t31 VGND 0.03709f
C16568 VPWR.t1467 VGND 0.0299f
C16569 VPWR.n498 VGND 0.09693f
C16570 VPWR.n499 VGND 0.01815f
C16571 VPWR.n500 VGND -0.00319f
C16572 VPWR.n501 VGND 0.09471f
C16573 VPWR.t1466 VGND 0.09401f
C16574 VPWR.t363 VGND 0.08295f
C16575 VPWR.t30 VGND 0.11982f
C16576 VPWR.t1401 VGND 0.03709f
C16577 VPWR.t19 VGND 0.0299f
C16578 VPWR.n502 VGND 0.09693f
C16579 VPWR.n503 VGND 0.01815f
C16580 VPWR.n504 VGND -0.00319f
C16581 VPWR.n505 VGND 0.09471f
C16582 VPWR.t18 VGND 0.09401f
C16583 VPWR.t364 VGND 0.08295f
C16584 VPWR.t1400 VGND 0.11982f
C16585 VPWR.t1243 VGND 0.03709f
C16586 VPWR.t1793 VGND 0.0299f
C16587 VPWR.n506 VGND 0.09693f
C16588 VPWR.n507 VGND 0.01815f
C16589 VPWR.n508 VGND -0.00319f
C16590 VPWR.n509 VGND 0.09471f
C16591 VPWR.t1792 VGND 0.09401f
C16592 VPWR.t365 VGND 0.08295f
C16593 VPWR.t1242 VGND 0.11982f
C16594 VPWR.n510 VGND 0.09471f
C16595 VPWR.n511 VGND -0.00319f
C16596 VPWR.n512 VGND 0.01815f
C16597 VPWR.n513 VGND 0.14051f
C16598 VPWR.n514 VGND 1.01936f
C16599 VPWR.n515 VGND 0.14051f
C16600 VPWR.t1207 VGND 0.03709f
C16601 VPWR.t335 VGND 0.0299f
C16602 VPWR.n516 VGND 0.09693f
C16603 VPWR.t1206 VGND 0.14747f
C16604 VPWR.t1334 VGND 0.08295f
C16605 VPWR.t334 VGND 0.09401f
C16606 VPWR.t1683 VGND 0.11982f
C16607 VPWR.t1020 VGND 0.03709f
C16608 VPWR.t1690 VGND 0.0299f
C16609 VPWR.n517 VGND 0.09693f
C16610 VPWR.n518 VGND 0.14051f
C16611 VPWR.n519 VGND 0.14051f
C16612 VPWR.t1684 VGND 0.03709f
C16613 VPWR.t1882 VGND 0.0299f
C16614 VPWR.n520 VGND 0.09693f
C16615 VPWR.t379 VGND 0.08295f
C16616 VPWR.t1881 VGND 0.09401f
C16617 VPWR.t584 VGND 0.11982f
C16618 VPWR.t998 VGND 0.03709f
C16619 VPWR.t1284 VGND 0.0299f
C16620 VPWR.n521 VGND 0.09693f
C16621 VPWR.n522 VGND 0.14051f
C16622 VPWR.n523 VGND 0.14051f
C16623 VPWR.t585 VGND 0.03709f
C16624 VPWR.t1703 VGND 0.0299f
C16625 VPWR.n524 VGND 0.09693f
C16626 VPWR.t1329 VGND 0.08295f
C16627 VPWR.t1702 VGND 0.09401f
C16628 VPWR.t1520 VGND 0.11982f
C16629 VPWR.t1255 VGND 0.03709f
C16630 VPWR.t281 VGND 0.0299f
C16631 VPWR.n525 VGND 0.09693f
C16632 VPWR.n526 VGND 0.14051f
C16633 VPWR.n527 VGND 0.14051f
C16634 VPWR.t1521 VGND 0.03709f
C16635 VPWR.t1095 VGND 0.0299f
C16636 VPWR.n528 VGND 0.09693f
C16637 VPWR.t377 VGND 0.08295f
C16638 VPWR.t1094 VGND 0.09401f
C16639 VPWR.t1424 VGND 0.11982f
C16640 VPWR.t271 VGND 0.03709f
C16641 VPWR.t1431 VGND 0.0299f
C16642 VPWR.n529 VGND 0.09693f
C16643 VPWR.n530 VGND 0.14051f
C16644 VPWR.n531 VGND 0.14051f
C16645 VPWR.t1425 VGND 0.03709f
C16646 VPWR.t1175 VGND 0.0299f
C16647 VPWR.n532 VGND 0.09693f
C16648 VPWR.t1332 VGND 0.08295f
C16649 VPWR.t1174 VGND 0.09401f
C16650 VPWR.t304 VGND 0.11982f
C16651 VPWR.t1896 VGND 0.03709f
C16652 VPWR.t1065 VGND 0.0299f
C16653 VPWR.n533 VGND 0.09693f
C16654 VPWR.n534 VGND 0.14051f
C16655 VPWR.n535 VGND 0.14051f
C16656 VPWR.t305 VGND 0.03709f
C16657 VPWR.t67 VGND 0.0299f
C16658 VPWR.n536 VGND 0.09693f
C16659 VPWR.t376 VGND 0.08295f
C16660 VPWR.t66 VGND 0.09401f
C16661 VPWR.t423 VGND 0.11982f
C16662 VPWR.t85 VGND 0.03709f
C16663 VPWR.t1489 VGND 0.0299f
C16664 VPWR.n537 VGND 0.09693f
C16665 VPWR.n538 VGND 0.14051f
C16666 VPWR.n539 VGND 0.14051f
C16667 VPWR.t424 VGND 0.03709f
C16668 VPWR.t1358 VGND 0.0299f
C16669 VPWR.n540 VGND 0.09693f
C16670 VPWR.t1323 VGND 0.08295f
C16671 VPWR.t1357 VGND 0.09401f
C16672 VPWR.t1646 VGND 0.11982f
C16673 VPWR.t1613 VGND 0.03709f
C16674 VPWR.t1659 VGND 0.0299f
C16675 VPWR.n541 VGND 0.09693f
C16676 VPWR.n542 VGND 0.14051f
C16677 VPWR.n543 VGND 0.14051f
C16678 VPWR.t1647 VGND 0.03709f
C16679 VPWR.t1372 VGND 0.0299f
C16680 VPWR.n544 VGND 0.09693f
C16681 VPWR.t1335 VGND 0.08295f
C16682 VPWR.t1371 VGND 0.09401f
C16683 VPWR.t442 VGND 0.03709f
C16684 VPWR.t821 VGND 0.0299f
C16685 VPWR.n545 VGND 0.09693f
C16686 VPWR.t458 VGND 0.03709f
C16687 VPWR.t939 VGND 0.0299f
C16688 VPWR.n546 VGND 0.09693f
C16689 VPWR.t1216 VGND 0.14747f
C16690 VPWR.t296 VGND 0.08295f
C16691 VPWR.t1029 VGND 0.09401f
C16692 VPWR.t1217 VGND 0.03709f
C16693 VPWR.t1030 VGND 0.0299f
C16694 VPWR.n547 VGND 0.09693f
C16695 VPWR.n548 VGND 0.01815f
C16696 VPWR.n549 VGND -0.00319f
C16697 VPWR.n550 VGND 0.09471f
C16698 VPWR.t1037 VGND 0.11982f
C16699 VPWR.t1262 VGND 0.08295f
C16700 VPWR.t1534 VGND 0.09401f
C16701 VPWR.t1038 VGND 0.03709f
C16702 VPWR.t1535 VGND 0.0299f
C16703 VPWR.n551 VGND 0.09693f
C16704 VPWR.n552 VGND 0.01815f
C16705 VPWR.n553 VGND -0.00319f
C16706 VPWR.n554 VGND 0.09471f
C16707 VPWR.t1798 VGND 0.11982f
C16708 VPWR.t1261 VGND 0.08295f
C16709 VPWR.t40 VGND 0.09401f
C16710 VPWR.t1799 VGND 0.03709f
C16711 VPWR.t41 VGND 0.0299f
C16712 VPWR.n555 VGND 0.09693f
C16713 VPWR.n556 VGND 0.01815f
C16714 VPWR.n557 VGND -0.00319f
C16715 VPWR.n558 VGND 0.09471f
C16716 VPWR.t16 VGND 0.11982f
C16717 VPWR.t1260 VGND 0.08295f
C16718 VPWR.t1295 VGND 0.09401f
C16719 VPWR.t17 VGND 0.03709f
C16720 VPWR.t1296 VGND 0.0299f
C16721 VPWR.n559 VGND 0.09693f
C16722 VPWR.n560 VGND 0.01815f
C16723 VPWR.n561 VGND -0.00319f
C16724 VPWR.n562 VGND 0.09471f
C16725 VPWR.t1918 VGND 0.11982f
C16726 VPWR.t340 VGND 0.08295f
C16727 VPWR.t1590 VGND 0.09401f
C16728 VPWR.t1919 VGND 0.03709f
C16729 VPWR.t1591 VGND 0.0299f
C16730 VPWR.n563 VGND 0.09693f
C16731 VPWR.n564 VGND 0.01815f
C16732 VPWR.n565 VGND -0.00319f
C16733 VPWR.n566 VGND 0.09471f
C16734 VPWR.t1584 VGND 0.11982f
C16735 VPWR.t1266 VGND 0.08295f
C16736 VPWR.t210 VGND 0.09401f
C16737 VPWR.t1585 VGND 0.03709f
C16738 VPWR.t211 VGND 0.0299f
C16739 VPWR.n567 VGND 0.09693f
C16740 VPWR.n568 VGND 0.01815f
C16741 VPWR.n569 VGND -0.00319f
C16742 VPWR.n570 VGND 0.09471f
C16743 VPWR.t1808 VGND 0.11982f
C16744 VPWR.t1259 VGND 0.08295f
C16745 VPWR.t268 VGND 0.09401f
C16746 VPWR.t1809 VGND 0.03709f
C16747 VPWR.t269 VGND 0.0299f
C16748 VPWR.n571 VGND 0.09693f
C16749 VPWR.n572 VGND 0.01815f
C16750 VPWR.n573 VGND -0.00319f
C16751 VPWR.n574 VGND 0.09471f
C16752 VPWR.t431 VGND 0.11982f
C16753 VPWR.t295 VGND 0.08295f
C16754 VPWR.t503 VGND 0.09401f
C16755 VPWR.t432 VGND 0.03709f
C16756 VPWR.t504 VGND 0.0299f
C16757 VPWR.n575 VGND 0.09693f
C16758 VPWR.n576 VGND 0.01815f
C16759 VPWR.n577 VGND -0.00319f
C16760 VPWR.n578 VGND 0.09471f
C16761 VPWR.t497 VGND 0.11982f
C16762 VPWR.t294 VGND 0.08295f
C16763 VPWR.t1899 VGND 0.09401f
C16764 VPWR.t498 VGND 0.03709f
C16765 VPWR.t1900 VGND 0.0299f
C16766 VPWR.n579 VGND 0.09693f
C16767 VPWR.n580 VGND 0.01815f
C16768 VPWR.n581 VGND -0.00319f
C16769 VPWR.n582 VGND 0.09471f
C16770 VPWR.t242 VGND 0.11982f
C16771 VPWR.t1265 VGND 0.08295f
C16772 VPWR.t191 VGND 0.09401f
C16773 VPWR.t243 VGND 0.03709f
C16774 VPWR.t192 VGND 0.0299f
C16775 VPWR.n583 VGND 0.09693f
C16776 VPWR.n584 VGND 0.01815f
C16777 VPWR.n585 VGND -0.00319f
C16778 VPWR.n586 VGND 0.09471f
C16779 VPWR.t320 VGND 0.11982f
C16780 VPWR.t1258 VGND 0.08295f
C16781 VPWR.t88 VGND 0.09401f
C16782 VPWR.t321 VGND 0.03709f
C16783 VPWR.t89 VGND 0.0299f
C16784 VPWR.n587 VGND 0.09693f
C16785 VPWR.n588 VGND 0.01815f
C16786 VPWR.n589 VGND -0.00319f
C16787 VPWR.n590 VGND 0.09471f
C16788 VPWR.t108 VGND 0.11982f
C16789 VPWR.t293 VGND 0.08295f
C16790 VPWR.t1506 VGND 0.09401f
C16791 VPWR.t109 VGND 0.03709f
C16792 VPWR.t1507 VGND 0.0299f
C16793 VPWR.n591 VGND 0.09693f
C16794 VPWR.n592 VGND 0.01815f
C16795 VPWR.n593 VGND -0.00319f
C16796 VPWR.n594 VGND 0.09471f
C16797 VPWR.t256 VGND 0.11982f
C16798 VPWR.t1264 VGND 0.08295f
C16799 VPWR.t170 VGND 0.09401f
C16800 VPWR.t257 VGND 0.03709f
C16801 VPWR.t171 VGND 0.0299f
C16802 VPWR.n595 VGND 0.09693f
C16803 VPWR.n596 VGND 0.01815f
C16804 VPWR.n597 VGND -0.00319f
C16805 VPWR.n598 VGND 0.09471f
C16806 VPWR.t1122 VGND 0.11982f
C16807 VPWR.t1263 VGND 0.08295f
C16808 VPWR.t1472 VGND 0.09401f
C16809 VPWR.t1123 VGND 0.03709f
C16810 VPWR.t1473 VGND 0.0299f
C16811 VPWR.n599 VGND 0.09693f
C16812 VPWR.n600 VGND 0.01815f
C16813 VPWR.n601 VGND -0.00319f
C16814 VPWR.n602 VGND 0.09471f
C16815 VPWR.t601 VGND 0.11982f
C16816 VPWR.t297 VGND 0.08295f
C16817 VPWR.t439 VGND 0.09401f
C16818 VPWR.t602 VGND 0.03709f
C16819 VPWR.t440 VGND 0.0299f
C16820 VPWR.n603 VGND 0.09693f
C16821 VPWR.n604 VGND 0.01815f
C16822 VPWR.n605 VGND -0.00319f
C16823 VPWR.n606 VGND 0.09471f
C16824 VPWR.t457 VGND 0.11982f
C16825 VPWR.t292 VGND 0.08295f
C16826 VPWR.t938 VGND 0.14528f
C16827 VPWR.n607 VGND 0.08265f
C16828 VPWR.n608 VGND 0.01815f
C16829 VPWR.n609 VGND 0.14051f
C16830 VPWR.n610 VGND 1.02579f
C16831 VPWR.n611 VGND 0.14051f
C16832 VPWR.t1376 VGND 0.03709f
C16833 VPWR.t674 VGND 0.0299f
C16834 VPWR.n612 VGND 0.09693f
C16835 VPWR.t459 VGND 0.09401f
C16836 VPWR.t1481 VGND 0.03709f
C16837 VPWR.t460 VGND 0.0299f
C16838 VPWR.n613 VGND 0.09693f
C16839 VPWR.n614 VGND 0.14051f
C16840 VPWR.n615 VGND 0.14051f
C16841 VPWR.t1412 VGND 0.03709f
C16842 VPWR.t1143 VGND 0.0299f
C16843 VPWR.n616 VGND 0.09693f
C16844 VPWR.t1342 VGND 0.09401f
C16845 VPWR.t1109 VGND 0.03709f
C16846 VPWR.t1343 VGND 0.0299f
C16847 VPWR.n617 VGND 0.09693f
C16848 VPWR.n618 VGND 0.14051f
C16849 VPWR.n619 VGND 0.14051f
C16850 VPWR.t71 VGND 0.03709f
C16851 VPWR.t249 VGND 0.0299f
C16852 VPWR.n620 VGND 0.09693f
C16853 VPWR.t112 VGND 0.09401f
C16854 VPWR.t350 VGND 0.03709f
C16855 VPWR.t113 VGND 0.0299f
C16856 VPWR.n621 VGND 0.09693f
C16857 VPWR.n622 VGND 0.14051f
C16858 VPWR.n623 VGND 0.14051f
C16859 VPWR.t1179 VGND 0.03709f
C16860 VPWR.t356 VGND 0.0299f
C16861 VPWR.n624 VGND 0.09693f
C16862 VPWR.t370 VGND 0.09401f
C16863 VPWR.t520 VGND 0.03709f
C16864 VPWR.t371 VGND 0.0299f
C16865 VPWR.n625 VGND 0.09693f
C16866 VPWR.n626 VGND 0.14051f
C16867 VPWR.n627 VGND 0.14051f
C16868 VPWR.t540 VGND 0.03709f
C16869 VPWR.t1392 VGND 0.0299f
C16870 VPWR.n628 VGND 0.09693f
C16871 VPWR.t1100 VGND 0.09401f
C16872 VPWR.t285 VGND 0.03709f
C16873 VPWR.t1101 VGND 0.0299f
C16874 VPWR.n629 VGND 0.09693f
C16875 VPWR.n630 VGND 0.14051f
C16876 VPWR.n631 VGND 0.14051f
C16877 VPWR.t1593 VGND 0.03709f
C16878 VPWR.t1813 VGND 0.0299f
C16879 VPWR.n632 VGND 0.09693f
C16880 VPWR.t1598 VGND 0.09401f
C16881 VPWR.t141 VGND 0.03709f
C16882 VPWR.t1599 VGND 0.0299f
C16883 VPWR.n633 VGND 0.09693f
C16884 VPWR.n634 VGND 0.14051f
C16885 VPWR.n635 VGND 0.14051f
C16886 VPWR.t1270 VGND 0.03709f
C16887 VPWR.t548 VGND 0.0299f
C16888 VPWR.n636 VGND 0.09693f
C16889 VPWR.t1275 VGND 0.09401f
C16890 VPWR.t1694 VGND 0.03709f
C16891 VPWR.t1276 VGND 0.0299f
C16892 VPWR.n637 VGND 0.09693f
C16893 VPWR.n638 VGND 0.14051f
C16894 VPWR.n639 VGND 0.14051f
C16895 VPWR.t337 VGND 0.03709f
C16896 VPWR.t1545 VGND 0.0299f
C16897 VPWR.n640 VGND 0.09693f
C16898 VPWR.t1228 VGND 0.14747f
C16899 VPWR.t183 VGND 0.08295f
C16900 VPWR.t479 VGND 0.09401f
C16901 VPWR.t1229 VGND 0.03709f
C16902 VPWR.t480 VGND 0.0299f
C16903 VPWR.n641 VGND 0.09693f
C16904 VPWR.t1203 VGND 0.03709f
C16905 VPWR.t1239 VGND 0.0299f
C16906 VPWR.n642 VGND 0.09693f
C16907 VPWR.t1202 VGND 0.14747f
C16908 VPWR.t1661 VGND 0.08295f
C16909 VPWR.t1238 VGND 0.09401f
C16910 VPWR.t450 VGND 0.03709f
C16911 VPWR.t775 VGND 0.0299f
C16912 VPWR.n643 VGND 0.09693f
C16913 VPWR.n644 VGND 0.01815f
C16914 VPWR.n645 VGND 0.08265f
C16915 VPWR.t774 VGND 0.14528f
C16916 VPWR.t1839 VGND 0.08295f
C16917 VPWR.t449 VGND 0.11982f
C16918 VPWR.t1477 VGND 0.03709f
C16919 VPWR.t1378 VGND 0.0299f
C16920 VPWR.n646 VGND 0.09693f
C16921 VPWR.n647 VGND 0.01815f
C16922 VPWR.n648 VGND -0.00319f
C16923 VPWR.n649 VGND 0.09471f
C16924 VPWR.t1377 VGND 0.09401f
C16925 VPWR.t1662 VGND 0.08295f
C16926 VPWR.t1476 VGND 0.11982f
C16927 VPWR.t1364 VGND 0.03709f
C16928 VPWR.t1081 VGND 0.0299f
C16929 VPWR.n650 VGND 0.09693f
C16930 VPWR.n651 VGND 0.01815f
C16931 VPWR.n652 VGND -0.00319f
C16932 VPWR.n653 VGND 0.09471f
C16933 VPWR.t1080 VGND 0.09401f
C16934 VPWR.t523 VGND 0.08295f
C16935 VPWR.t1363 VGND 0.11982f
C16936 VPWR.t1491 VGND 0.03709f
C16937 VPWR.t1603 VGND 0.0299f
C16938 VPWR.n654 VGND 0.09693f
C16939 VPWR.n655 VGND 0.01815f
C16940 VPWR.n656 VGND -0.00319f
C16941 VPWR.n657 VGND 0.09471f
C16942 VPWR.t1602 VGND 0.09401f
C16943 VPWR.t524 VGND 0.08295f
C16944 VPWR.t1490 VGND 0.11982f
C16945 VPWR.t81 VGND 0.03709f
C16946 VPWR.t1497 VGND 0.0299f
C16947 VPWR.n658 VGND 0.09693f
C16948 VPWR.n659 VGND 0.01815f
C16949 VPWR.n660 VGND -0.00319f
C16950 VPWR.n661 VGND 0.09471f
C16951 VPWR.t1496 VGND 0.09401f
C16952 VPWR.t1840 VGND 0.08295f
C16953 VPWR.t80 VGND 0.11982f
C16954 VPWR.t1067 VGND 0.03709f
C16955 VPWR.t61 VGND 0.0299f
C16956 VPWR.n662 VGND 0.09693f
C16957 VPWR.n663 VGND 0.01815f
C16958 VPWR.n664 VGND -0.00319f
C16959 VPWR.n665 VGND 0.09471f
C16960 VPWR.t60 VGND 0.09401f
C16961 VPWR.t1326 VGND 0.08295f
C16962 VPWR.t1066 VGND 0.11982f
C16963 VPWR.t1908 VGND 0.03709f
C16964 VPWR.t289 VGND 0.0299f
C16965 VPWR.n666 VGND 0.09693f
C16966 VPWR.n667 VGND 0.01815f
C16967 VPWR.n668 VGND -0.00319f
C16968 VPWR.n669 VGND 0.09471f
C16969 VPWR.t288 VGND 0.09401f
C16970 VPWR.t525 VGND 0.08295f
C16971 VPWR.t1907 VGND 0.11982f
C16972 VPWR.t1437 VGND 0.03709f
C16973 VPWR.t231 VGND 0.0299f
C16974 VPWR.n670 VGND 0.09693f
C16975 VPWR.n671 VGND 0.01815f
C16976 VPWR.n672 VGND -0.00319f
C16977 VPWR.n673 VGND 0.09471f
C16978 VPWR.t230 VGND 0.09401f
C16979 VPWR.t1841 VGND 0.08295f
C16980 VPWR.t1436 VGND 0.11982f
C16981 VPWR.t1627 VGND 0.03709f
C16982 VPWR.t512 VGND 0.0299f
C16983 VPWR.n674 VGND 0.09693f
C16984 VPWR.n675 VGND 0.01815f
C16985 VPWR.n676 VGND -0.00319f
C16986 VPWR.n677 VGND 0.09471f
C16987 VPWR.t511 VGND 0.09401f
C16988 VPWR.t1660 VGND 0.08295f
C16989 VPWR.t1626 VGND 0.11982f
C16990 VPWR.t219 VGND 0.03709f
C16991 VPWR.t542 VGND 0.0299f
C16992 VPWR.n678 VGND 0.09693f
C16993 VPWR.n679 VGND 0.01815f
C16994 VPWR.n680 VGND -0.00319f
C16995 VPWR.n681 VGND 0.09471f
C16996 VPWR.t541 VGND 0.09401f
C16997 VPWR.t1327 VGND 0.08295f
C16998 VPWR.t218 VGND 0.11982f
C16999 VPWR.t1709 VGND 0.03709f
C17000 VPWR.t1553 VGND 0.0299f
C17001 VPWR.n682 VGND 0.09693f
C17002 VPWR.n683 VGND 0.01815f
C17003 VPWR.n684 VGND -0.00319f
C17004 VPWR.n685 VGND 0.09471f
C17005 VPWR.t1552 VGND 0.09401f
C17006 VPWR.t526 VGND 0.08295f
C17007 VPWR.t1708 VGND 0.11982f
C17008 VPWR.t1463 VGND 0.03709f
C17009 VPWR.t1713 VGND 0.0299f
C17010 VPWR.n686 VGND 0.09693f
C17011 VPWR.n687 VGND 0.01815f
C17012 VPWR.n688 VGND -0.00319f
C17013 VPWR.n689 VGND 0.09471f
C17014 VPWR.t1712 VGND 0.09401f
C17015 VPWR.t1838 VGND 0.08295f
C17016 VPWR.t1462 VGND 0.11982f
C17017 VPWR.t1884 VGND 0.03709f
C17018 VPWR.t1923 VGND 0.0299f
C17019 VPWR.n690 VGND 0.09693f
C17020 VPWR.n691 VGND 0.01815f
C17021 VPWR.n692 VGND -0.00319f
C17022 VPWR.n693 VGND 0.09471f
C17023 VPWR.t1922 VGND 0.09401f
C17024 VPWR.t1328 VGND 0.08295f
C17025 VPWR.t1883 VGND 0.11982f
C17026 VPWR.t1441 VGND 0.03709f
C17027 VPWR.t37 VGND 0.0299f
C17028 VPWR.n694 VGND 0.09693f
C17029 VPWR.n695 VGND 0.01815f
C17030 VPWR.n696 VGND -0.00319f
C17031 VPWR.n697 VGND 0.09471f
C17032 VPWR.t36 VGND 0.09401f
C17033 VPWR.t521 VGND 0.08295f
C17034 VPWR.t1440 VGND 0.11982f
C17035 VPWR.t1845 VGND 0.03709f
C17036 VPWR.t1445 VGND 0.0299f
C17037 VPWR.n698 VGND 0.09693f
C17038 VPWR.n699 VGND 0.01815f
C17039 VPWR.n700 VGND -0.00319f
C17040 VPWR.n701 VGND 0.09471f
C17041 VPWR.t1444 VGND 0.09401f
C17042 VPWR.t522 VGND 0.08295f
C17043 VPWR.t1844 VGND 0.11982f
C17044 VPWR.n702 VGND 0.09471f
C17045 VPWR.n703 VGND -0.00319f
C17046 VPWR.n704 VGND 0.01815f
C17047 VPWR.n705 VGND 0.14051f
C17048 VPWR.n706 VGND 1.01936f
C17049 VPWR.n707 VGND 0.14051f
C17050 VPWR.t1199 VGND 0.03709f
C17051 VPWR.t1034 VGND 0.0299f
C17052 VPWR.n708 VGND 0.09693f
C17053 VPWR.t1198 VGND 0.14747f
C17054 VPWR.t313 VGND 0.08295f
C17055 VPWR.t1033 VGND 0.09401f
C17056 VPWR.t178 VGND 0.11982f
C17057 VPWR.t1851 VGND 0.03709f
C17058 VPWR.t1692 VGND 0.0299f
C17059 VPWR.n709 VGND 0.09693f
C17060 VPWR.n710 VGND 0.14051f
C17061 VPWR.n711 VGND 0.14051f
C17062 VPWR.t179 VGND 0.03709f
C17063 VPWR.t1268 VGND 0.0299f
C17064 VPWR.n712 VGND 0.09693f
C17065 VPWR.t1790 VGND 0.08295f
C17066 VPWR.t1267 VGND 0.09401f
C17067 VPWR.t1291 VGND 0.11982f
C17068 VPWR.t57 VGND 0.03709f
C17069 VPWR.t1057 VGND 0.0299f
C17070 VPWR.n713 VGND 0.09693f
C17071 VPWR.n714 VGND 0.14051f
C17072 VPWR.n715 VGND 0.14051f
C17073 VPWR.t1292 VGND 0.03709f
C17074 VPWR.t1698 VGND 0.0299f
C17075 VPWR.n716 VGND 0.09693f
C17076 VPWR.t1397 VGND 0.08295f
C17077 VPWR.t1697 VGND 0.09401f
C17078 VPWR.t46 VGND 0.11982f
C17079 VPWR.t1696 VGND 0.03709f
C17080 VPWR.t1557 VGND 0.0299f
C17081 VPWR.n717 VGND 0.09693f
C17082 VPWR.n718 VGND 0.14051f
C17083 VPWR.n719 VGND 0.14051f
C17084 VPWR.t47 VGND 0.03709f
C17085 VPWR.t165 VGND 0.0299f
C17086 VPWR.n720 VGND 0.09693f
C17087 VPWR.t1788 VGND 0.08295f
C17088 VPWR.t164 VGND 0.09401f
C17089 VPWR.t515 VGND 0.11982f
C17090 VPWR.t1091 VGND 0.03709f
C17091 VPWR.t518 VGND 0.0299f
C17092 VPWR.n721 VGND 0.09693f
C17093 VPWR.n722 VGND 0.14051f
C17094 VPWR.n723 VGND 0.14051f
C17095 VPWR.t516 VGND 0.03709f
C17096 VPWR.t235 VGND 0.0299f
C17097 VPWR.n724 VGND 0.09693f
C17098 VPWR.t311 VGND 0.08295f
C17099 VPWR.t234 VGND 0.09401f
C17100 VPWR.t342 VGND 0.11982f
C17101 VPWR.t1169 VGND 0.03709f
C17102 VPWR.t345 VGND 0.0299f
C17103 VPWR.n725 VGND 0.09693f
C17104 VPWR.n726 VGND 0.14051f
C17105 VPWR.n727 VGND 0.14051f
C17106 VPWR.t343 VGND 0.03709f
C17107 VPWR.t115 VGND 0.0299f
C17108 VPWR.n728 VGND 0.09693f
C17109 VPWR.t575 VGND 0.08295f
C17110 VPWR.t114 VGND 0.09401f
C17111 VPWR.t1614 VGND 0.11982f
C17112 VPWR.t75 VGND 0.03709f
C17113 VPWR.t1617 VGND 0.0299f
C17114 VPWR.n729 VGND 0.09693f
C17115 VPWR.n730 VGND 0.14051f
C17116 VPWR.n731 VGND 0.14051f
C17117 VPWR.t1615 VGND 0.03709f
C17118 VPWR.t1410 VGND 0.0299f
C17119 VPWR.n732 VGND 0.09693f
C17120 VPWR.t307 VGND 0.08295f
C17121 VPWR.t1409 VGND 0.09401f
C17122 VPWR.t1074 VGND 0.11982f
C17123 VPWR.t1607 VGND 0.03709f
C17124 VPWR.t598 VGND 0.0299f
C17125 VPWR.n733 VGND 0.09693f
C17126 VPWR.n734 VGND 0.14051f
C17127 VPWR.n735 VGND 0.14051f
C17128 VPWR.t1075 VGND 0.03709f
C17129 VPWR.t494 VGND 0.0299f
C17130 VPWR.n736 VGND 0.09693f
C17131 VPWR.t1399 VGND 0.08295f
C17132 VPWR.t493 VGND 0.09401f
C17133 VPWR.t1368 VGND 0.03709f
C17134 VPWR.t735 VGND 0.0299f
C17135 VPWR.n737 VGND 0.09693f
C17136 VPWR.t438 VGND 0.03709f
C17137 VPWR.t837 VGND 0.0299f
C17138 VPWR.n738 VGND 0.09693f
C17139 VPWR.t1208 VGND 0.14747f
C17140 VPWR.t1306 VGND 0.08295f
C17141 VPWR.t332 VGND 0.09401f
C17142 VPWR.t1209 VGND 0.03709f
C17143 VPWR.t333 VGND 0.0299f
C17144 VPWR.n739 VGND 0.09693f
C17145 VPWR.n740 VGND 0.01815f
C17146 VPWR.n741 VGND -0.00319f
C17147 VPWR.n742 VGND 0.09471f
C17148 VPWR.t1017 VGND 0.11982f
C17149 VPWR.t150 VGND 0.08295f
C17150 VPWR.t1687 VGND 0.09401f
C17151 VPWR.t1018 VGND 0.03709f
C17152 VPWR.t1688 VGND 0.0299f
C17153 VPWR.n743 VGND 0.09693f
C17154 VPWR.n744 VGND 0.01815f
C17155 VPWR.n745 VGND -0.00319f
C17156 VPWR.n746 VGND 0.09471f
C17157 VPWR.t1681 VGND 0.11982f
C17158 VPWR.t149 VGND 0.08295f
C17159 VPWR.t1879 VGND 0.09401f
C17160 VPWR.t1682 VGND 0.03709f
C17161 VPWR.t1880 VGND 0.0299f
C17162 VPWR.n747 VGND 0.09693f
C17163 VPWR.n748 VGND 0.01815f
C17164 VPWR.n749 VGND -0.00319f
C17165 VPWR.n750 VGND 0.09471f
C17166 VPWR.t995 VGND 0.11982f
C17167 VPWR.t1310 VGND 0.08295f
C17168 VPWR.t1281 VGND 0.09401f
C17169 VPWR.t996 VGND 0.03709f
C17170 VPWR.t1282 VGND 0.0299f
C17171 VPWR.n751 VGND 0.09693f
C17172 VPWR.n752 VGND 0.01815f
C17173 VPWR.n753 VGND -0.00319f
C17174 VPWR.n754 VGND 0.09471f
C17175 VPWR.t582 VGND 0.11982f
C17176 VPWR.t148 VGND 0.08295f
C17177 VPWR.t1700 VGND 0.09401f
C17178 VPWR.t583 VGND 0.03709f
C17179 VPWR.t1701 VGND 0.0299f
C17180 VPWR.n755 VGND 0.09693f
C17181 VPWR.n756 VGND 0.01815f
C17182 VPWR.n757 VGND -0.00319f
C17183 VPWR.n758 VGND 0.09471f
C17184 VPWR.t1252 VGND 0.11982f
C17185 VPWR.t147 VGND 0.08295f
C17186 VPWR.t278 VGND 0.09401f
C17187 VPWR.t1253 VGND 0.03709f
C17188 VPWR.t279 VGND 0.0299f
C17189 VPWR.n759 VGND 0.09693f
C17190 VPWR.n760 VGND 0.01815f
C17191 VPWR.n761 VGND -0.00319f
C17192 VPWR.n762 VGND 0.09471f
C17193 VPWR.t1518 VGND 0.11982f
C17194 VPWR.t1309 VGND 0.08295f
C17195 VPWR.t1092 VGND 0.09401f
C17196 VPWR.t1519 VGND 0.03709f
C17197 VPWR.t1093 VGND 0.0299f
C17198 VPWR.n763 VGND 0.09693f
C17199 VPWR.n764 VGND 0.01815f
C17200 VPWR.n765 VGND -0.00319f
C17201 VPWR.n766 VGND 0.09471f
C17202 VPWR.t266 VGND 0.11982f
C17203 VPWR.t1305 VGND 0.08295f
C17204 VPWR.t1428 VGND 0.09401f
C17205 VPWR.t267 VGND 0.03709f
C17206 VPWR.t1429 VGND 0.0299f
C17207 VPWR.n767 VGND 0.09693f
C17208 VPWR.n768 VGND 0.01815f
C17209 VPWR.n769 VGND -0.00319f
C17210 VPWR.n770 VGND 0.09471f
C17211 VPWR.t1422 VGND 0.11982f
C17212 VPWR.t1304 VGND 0.08295f
C17213 VPWR.t1172 VGND 0.09401f
C17214 VPWR.t1423 VGND 0.03709f
C17215 VPWR.t1173 VGND 0.0299f
C17216 VPWR.n771 VGND 0.09693f
C17217 VPWR.n772 VGND 0.01815f
C17218 VPWR.n773 VGND -0.00319f
C17219 VPWR.n774 VGND 0.09471f
C17220 VPWR.t1893 VGND 0.11982f
C17221 VPWR.t146 VGND 0.08295f
C17222 VPWR.t1062 VGND 0.09401f
C17223 VPWR.t1894 VGND 0.03709f
C17224 VPWR.t1063 VGND 0.0299f
C17225 VPWR.n775 VGND 0.09693f
C17226 VPWR.n776 VGND 0.01815f
C17227 VPWR.n777 VGND -0.00319f
C17228 VPWR.n778 VGND 0.09471f
C17229 VPWR.t302 VGND 0.11982f
C17230 VPWR.t1308 VGND 0.08295f
C17231 VPWR.t64 VGND 0.09401f
C17232 VPWR.t303 VGND 0.03709f
C17233 VPWR.t65 VGND 0.0299f
C17234 VPWR.n779 VGND 0.09693f
C17235 VPWR.n780 VGND 0.01815f
C17236 VPWR.n781 VGND -0.00319f
C17237 VPWR.n782 VGND 0.09471f
C17238 VPWR.t100 VGND 0.11982f
C17239 VPWR.t1303 VGND 0.08295f
C17240 VPWR.t563 VGND 0.09401f
C17241 VPWR.t101 VGND 0.03709f
C17242 VPWR.t564 VGND 0.0299f
C17243 VPWR.n783 VGND 0.09693f
C17244 VPWR.n784 VGND 0.01815f
C17245 VPWR.n785 VGND -0.00319f
C17246 VPWR.n786 VGND 0.09471f
C17247 VPWR.t421 VGND 0.11982f
C17248 VPWR.t145 VGND 0.08295f
C17249 VPWR.t1355 VGND 0.09401f
C17250 VPWR.t422 VGND 0.03709f
C17251 VPWR.t1356 VGND 0.0299f
C17252 VPWR.n787 VGND 0.09693f
C17253 VPWR.n788 VGND 0.01815f
C17254 VPWR.n789 VGND -0.00319f
C17255 VPWR.n790 VGND 0.09471f
C17256 VPWR.t1610 VGND 0.11982f
C17257 VPWR.t144 VGND 0.08295f
C17258 VPWR.t1656 VGND 0.09401f
C17259 VPWR.t1611 VGND 0.03709f
C17260 VPWR.t1657 VGND 0.0299f
C17261 VPWR.n791 VGND 0.09693f
C17262 VPWR.n792 VGND 0.01815f
C17263 VPWR.n793 VGND -0.00319f
C17264 VPWR.n794 VGND 0.09471f
C17265 VPWR.t1644 VGND 0.11982f
C17266 VPWR.t1307 VGND 0.08295f
C17267 VPWR.t1369 VGND 0.09401f
C17268 VPWR.t1645 VGND 0.03709f
C17269 VPWR.t1370 VGND 0.0299f
C17270 VPWR.n795 VGND 0.09693f
C17271 VPWR.n796 VGND 0.01815f
C17272 VPWR.n797 VGND -0.00319f
C17273 VPWR.n798 VGND 0.09471f
C17274 VPWR.t437 VGND 0.11982f
C17275 VPWR.t1302 VGND 0.08295f
C17276 VPWR.t836 VGND 0.14528f
C17277 VPWR.n799 VGND 0.08265f
C17278 VPWR.n800 VGND 0.01815f
C17279 VPWR.n801 VGND 0.14051f
C17280 VPWR.n802 VGND 1.02579f
C17281 VPWR.n803 VGND 0.14051f
C17282 VPWR.t1380 VGND 0.03709f
C17283 VPWR.t671 VGND 0.0299f
C17284 VPWR.n804 VGND 0.09693f
C17285 VPWR.t461 VGND 0.09401f
C17286 VPWR.t1483 VGND 0.03709f
C17287 VPWR.t462 VGND 0.0299f
C17288 VPWR.n805 VGND 0.09693f
C17289 VPWR.n806 VGND 0.14051f
C17290 VPWR.n807 VGND 0.14051f
C17291 VPWR.t1414 VGND 0.03709f
C17292 VPWR.t1145 VGND 0.0299f
C17293 VPWR.n808 VGND 0.09693f
C17294 VPWR.t1344 VGND 0.09401f
C17295 VPWR.t1111 VGND 0.03709f
C17296 VPWR.t1345 VGND 0.0299f
C17297 VPWR.n809 VGND 0.09693f
C17298 VPWR.n810 VGND 0.14051f
C17299 VPWR.n811 VGND 0.14051f
C17300 VPWR.t73 VGND 0.03709f
C17301 VPWR.t251 VGND 0.0299f
C17302 VPWR.n812 VGND 0.09693f
C17303 VPWR.t102 VGND 0.09401f
C17304 VPWR.t352 VGND 0.03709f
C17305 VPWR.t103 VGND 0.0299f
C17306 VPWR.n813 VGND 0.09693f
C17307 VPWR.n814 VGND 0.14051f
C17308 VPWR.n815 VGND 0.14051f
C17309 VPWR.t1181 VGND 0.03709f
C17310 VPWR.t358 VGND 0.0299f
C17311 VPWR.n816 VGND 0.09693f
C17312 VPWR.t372 VGND 0.09401f
C17313 VPWR.t1388 VGND 0.03709f
C17314 VPWR.t373 VGND 0.0299f
C17315 VPWR.n817 VGND 0.09693f
C17316 VPWR.n818 VGND 0.14051f
C17317 VPWR.n819 VGND 0.14051f
C17318 VPWR.t544 VGND 0.03709f
C17319 VPWR.t1394 VGND 0.0299f
C17320 VPWR.n820 VGND 0.09693f
C17321 VPWR.t1102 VGND 0.09401f
C17322 VPWR.t287 VGND 0.03709f
C17323 VPWR.t1103 VGND 0.0299f
C17324 VPWR.n821 VGND 0.09693f
C17325 VPWR.n822 VGND 0.14051f
C17326 VPWR.n823 VGND 0.14051f
C17327 VPWR.t1595 VGND 0.03709f
C17328 VPWR.t1815 VGND 0.0299f
C17329 VPWR.n824 VGND 0.09693f
C17330 VPWR.t1522 VGND 0.09401f
C17331 VPWR.t143 VGND 0.03709f
C17332 VPWR.t1523 VGND 0.0299f
C17333 VPWR.n825 VGND 0.09693f
C17334 VPWR.n826 VGND 0.14051f
C17335 VPWR.n827 VGND 0.14051f
C17336 VPWR.t1272 VGND 0.03709f
C17337 VPWR.t550 VGND 0.0299f
C17338 VPWR.n828 VGND 0.09693f
C17339 VPWR.t26 VGND 0.09401f
C17340 VPWR.t1541 VGND 0.03709f
C17341 VPWR.t27 VGND 0.0299f
C17342 VPWR.n829 VGND 0.09693f
C17343 VPWR.n830 VGND 0.14051f
C17344 VPWR.n831 VGND 0.14051f
C17345 VPWR.t339 VGND 0.03709f
C17346 VPWR.t1547 VGND 0.0299f
C17347 VPWR.n832 VGND 0.09693f
C17348 VPWR.t1226 VGND 0.14747f
C17349 VPWR.t1098 VGND 0.08295f
C17350 VPWR.t591 VGND 0.09401f
C17351 VPWR.t1227 VGND 0.03709f
C17352 VPWR.t592 VGND 0.0299f
C17353 VPWR.n833 VGND 0.09693f
C17354 VPWR.t1213 VGND 0.03709f
C17355 VPWR.t331 VGND 0.0299f
C17356 VPWR.n834 VGND 0.09693f
C17357 VPWR.t1212 VGND 0.14747f
C17358 VPWR.t1577 VGND 0.08295f
C17359 VPWR.t330 VGND 0.09401f
C17360 VPWR.t434 VGND 0.03709f
C17361 VPWR.t846 VGND 0.0299f
C17362 VPWR.n835 VGND 0.09693f
C17363 VPWR.n836 VGND 0.01815f
C17364 VPWR.n837 VGND 0.08265f
C17365 VPWR.t845 VGND 0.14528f
C17366 VPWR.t1573 VGND 0.08295f
C17367 VPWR.t433 VGND 0.11982f
C17368 VPWR.t1233 VGND 0.03709f
C17369 VPWR.t1366 VGND 0.0299f
C17370 VPWR.n838 VGND 0.09693f
C17371 VPWR.n839 VGND 0.01815f
C17372 VPWR.n840 VGND -0.00319f
C17373 VPWR.n841 VGND 0.09471f
C17374 VPWR.t1365 VGND 0.09401f
C17375 VPWR.t1675 VGND 0.08295f
C17376 VPWR.t1232 VGND 0.11982f
C17377 VPWR.t1609 VGND 0.03709f
C17378 VPWR.t1655 VGND 0.0299f
C17379 VPWR.n842 VGND 0.09693f
C17380 VPWR.n843 VGND 0.01815f
C17381 VPWR.n844 VGND -0.00319f
C17382 VPWR.n845 VGND 0.09471f
C17383 VPWR.t1654 VGND 0.09401f
C17384 VPWR.t1277 VGND 0.08295f
C17385 VPWR.t1608 VGND 0.11982f
C17386 VPWR.t420 VGND 0.03709f
C17387 VPWR.t1354 VGND 0.0299f
C17388 VPWR.n846 VGND 0.09693f
C17389 VPWR.n847 VGND 0.01815f
C17390 VPWR.n848 VGND -0.00319f
C17391 VPWR.n849 VGND 0.09471f
C17392 VPWR.t1353 VGND 0.09401f
C17393 VPWR.t1278 VGND 0.08295f
C17394 VPWR.t419 VGND 0.11982f
C17395 VPWR.t97 VGND 0.03709f
C17396 VPWR.t562 VGND 0.0299f
C17397 VPWR.n850 VGND 0.09693f
C17398 VPWR.n851 VGND 0.01815f
C17399 VPWR.n852 VGND -0.00319f
C17400 VPWR.n853 VGND 0.09471f
C17401 VPWR.t561 VGND 0.09401f
C17402 VPWR.t1574 VGND 0.08295f
C17403 VPWR.t96 VGND 0.11982f
C17404 VPWR.t301 VGND 0.03709f
C17405 VPWR.t77 VGND 0.0299f
C17406 VPWR.n854 VGND 0.09693f
C17407 VPWR.n855 VGND 0.01815f
C17408 VPWR.n856 VGND -0.00319f
C17409 VPWR.n857 VGND 0.09471f
C17410 VPWR.t76 VGND 0.09401f
C17411 VPWR.t1676 VGND 0.08295f
C17412 VPWR.t300 VGND 0.11982f
C17413 VPWR.t1890 VGND 0.03709f
C17414 VPWR.t1061 VGND 0.0299f
C17415 VPWR.n858 VGND 0.09693f
C17416 VPWR.n859 VGND 0.01815f
C17417 VPWR.n860 VGND -0.00319f
C17418 VPWR.n861 VGND 0.09471f
C17419 VPWR.t1060 VGND 0.09401f
C17420 VPWR.t1279 VGND 0.08295f
C17421 VPWR.t1889 VGND 0.11982f
C17422 VPWR.t1421 VGND 0.03709f
C17423 VPWR.t1171 VGND 0.0299f
C17424 VPWR.n862 VGND 0.09693f
C17425 VPWR.n863 VGND 0.01815f
C17426 VPWR.n864 VGND -0.00319f
C17427 VPWR.n865 VGND 0.09471f
C17428 VPWR.t1170 VGND 0.09401f
C17429 VPWR.t1575 VGND 0.08295f
C17430 VPWR.t1420 VGND 0.11982f
C17431 VPWR.t1459 VGND 0.03709f
C17432 VPWR.t1427 VGND 0.0299f
C17433 VPWR.n866 VGND 0.09693f
C17434 VPWR.n867 VGND 0.01815f
C17435 VPWR.n868 VGND -0.00319f
C17436 VPWR.n869 VGND 0.09471f
C17437 VPWR.t1426 VGND 0.09401f
C17438 VPWR.t1576 VGND 0.08295f
C17439 VPWR.t1458 VGND 0.11982f
C17440 VPWR.t1515 VGND 0.03709f
C17441 VPWR.t1089 VGND 0.0299f
C17442 VPWR.n870 VGND 0.09693f
C17443 VPWR.n871 VGND 0.01815f
C17444 VPWR.n872 VGND -0.00319f
C17445 VPWR.n873 VGND 0.09471f
C17446 VPWR.t1088 VGND 0.09401f
C17447 VPWR.t1677 VGND 0.08295f
C17448 VPWR.t1514 VGND 0.11982f
C17449 VPWR.t1251 VGND 0.03709f
C17450 VPWR.t277 VGND 0.0299f
C17451 VPWR.n874 VGND 0.09693f
C17452 VPWR.n875 VGND 0.01815f
C17453 VPWR.n876 VGND -0.00319f
C17454 VPWR.n877 VGND 0.09471f
C17455 VPWR.t276 VGND 0.09401f
C17456 VPWR.t1280 VGND 0.08295f
C17457 VPWR.t1250 VGND 0.11982f
C17458 VPWR.t581 VGND 0.03709f
C17459 VPWR.t1257 VGND 0.0299f
C17460 VPWR.n878 VGND 0.09693f
C17461 VPWR.n879 VGND 0.01815f
C17462 VPWR.n880 VGND -0.00319f
C17463 VPWR.n881 VGND 0.09471f
C17464 VPWR.t1256 VGND 0.09401f
C17465 VPWR.t1572 VGND 0.08295f
C17466 VPWR.t580 VGND 0.11982f
C17467 VPWR.t994 VGND 0.03709f
C17468 VPWR.t579 VGND 0.0299f
C17469 VPWR.n882 VGND 0.09693f
C17470 VPWR.n883 VGND 0.01815f
C17471 VPWR.n884 VGND -0.00319f
C17472 VPWR.n885 VGND 0.09471f
C17473 VPWR.t578 VGND 0.09401f
C17474 VPWR.t1678 VGND 0.08295f
C17475 VPWR.t993 VGND 0.11982f
C17476 VPWR.t1418 VGND 0.03709f
C17477 VPWR.t387 VGND 0.0299f
C17478 VPWR.n886 VGND 0.09693f
C17479 VPWR.n887 VGND 0.01815f
C17480 VPWR.n888 VGND -0.00319f
C17481 VPWR.n889 VGND 0.09471f
C17482 VPWR.t386 VGND 0.09401f
C17483 VPWR.t1679 VGND 0.08295f
C17484 VPWR.t1417 VGND 0.11982f
C17485 VPWR.t596 VGND 0.03709f
C17486 VPWR.t1686 VGND 0.0299f
C17487 VPWR.n890 VGND 0.09693f
C17488 VPWR.n891 VGND 0.01815f
C17489 VPWR.n892 VGND -0.00319f
C17490 VPWR.n893 VGND 0.09471f
C17491 VPWR.t1685 VGND 0.09401f
C17492 VPWR.t1680 VGND 0.08295f
C17493 VPWR.t595 VGND 0.11982f
C17494 VPWR.n894 VGND 0.09471f
C17495 VPWR.n895 VGND -0.00319f
C17496 VPWR.n896 VGND 0.01815f
C17497 VPWR.n897 VGND 0.14051f
C17498 VPWR.n898 VGND 1.01936f
C17499 VPWR.n899 VGND 0.14051f
C17500 VPWR.t1219 VGND 0.03709f
C17501 VPWR.t1028 VGND 0.0299f
C17502 VPWR.n900 VGND 0.09693f
C17503 VPWR.t1218 VGND 0.14747f
C17504 VPWR.t1248 VGND 0.08295f
C17505 VPWR.t1027 VGND 0.09401f
C17506 VPWR.t1796 VGND 0.11982f
C17507 VPWR.t1036 VGND 0.03709f
C17508 VPWR.t1803 VGND 0.0299f
C17509 VPWR.n901 VGND 0.09693f
C17510 VPWR.n902 VGND 0.14051f
C17511 VPWR.n903 VGND 0.14051f
C17512 VPWR.t1797 VGND 0.03709f
C17513 VPWR.t25 VGND 0.0299f
C17514 VPWR.n904 VGND 0.09693f
C17515 VPWR.t1565 VGND 0.08295f
C17516 VPWR.t24 VGND 0.09401f
C17517 VPWR.t1916 VGND 0.11982f
C17518 VPWR.t15 VGND 0.03709f
C17519 VPWR.t1294 VGND 0.0299f
C17520 VPWR.n905 VGND 0.09693f
C17521 VPWR.n906 VGND 0.14051f
C17522 VPWR.n907 VGND 0.14051f
C17523 VPWR.t1917 VGND 0.03709f
C17524 VPWR.t1589 VGND 0.0299f
C17525 VPWR.n908 VGND 0.09693f
C17526 VPWR.t1571 VGND 0.08295f
C17527 VPWR.t1588 VGND 0.09401f
C17528 VPWR.t1806 VGND 0.11982f
C17529 VPWR.t1583 VGND 0.03709f
C17530 VPWR.t209 VGND 0.0299f
C17531 VPWR.n909 VGND 0.09693f
C17532 VPWR.n910 VGND 0.14051f
C17533 VPWR.n911 VGND 0.14051f
C17534 VPWR.t1807 VGND 0.03709f
C17535 VPWR.t265 VGND 0.0299f
C17536 VPWR.n912 VGND 0.09693f
C17537 VPWR.t1563 VGND 0.08295f
C17538 VPWR.t264 VGND 0.09401f
C17539 VPWR.t495 VGND 0.11982f
C17540 VPWR.t430 VGND 0.03709f
C17541 VPWR.t502 VGND 0.0299f
C17542 VPWR.n913 VGND 0.09693f
C17543 VPWR.n914 VGND 0.14051f
C17544 VPWR.n915 VGND 0.14051f
C17545 VPWR.t496 VGND 0.03709f
C17546 VPWR.t1898 VGND 0.0299f
C17547 VPWR.n916 VGND 0.09693f
C17548 VPWR.t1246 VGND 0.08295f
C17549 VPWR.t1897 VGND 0.09401f
C17550 VPWR.t318 VGND 0.11982f
C17551 VPWR.t241 VGND 0.03709f
C17552 VPWR.t190 VGND 0.0299f
C17553 VPWR.n917 VGND 0.09693f
C17554 VPWR.n918 VGND 0.14051f
C17555 VPWR.n919 VGND 0.14051f
C17556 VPWR.t319 VGND 0.03709f
C17557 VPWR.t87 VGND 0.0299f
C17558 VPWR.n920 VGND 0.09693f
C17559 VPWR.t1562 VGND 0.08295f
C17560 VPWR.t86 VGND 0.09401f
C17561 VPWR.t254 VGND 0.11982f
C17562 VPWR.t107 VGND 0.03709f
C17563 VPWR.t1505 VGND 0.0299f
C17564 VPWR.n921 VGND 0.09693f
C17565 VPWR.n922 VGND 0.14051f
C17566 VPWR.n923 VGND 0.14051f
C17567 VPWR.t255 VGND 0.03709f
C17568 VPWR.t169 VGND 0.0299f
C17569 VPWR.n924 VGND 0.09693f
C17570 VPWR.t1568 VGND 0.08295f
C17571 VPWR.t168 VGND 0.09401f
C17572 VPWR.t599 VGND 0.11982f
C17573 VPWR.t1121 VGND 0.03709f
C17574 VPWR.t1471 VGND 0.0299f
C17575 VPWR.n925 VGND 0.09693f
C17576 VPWR.n926 VGND 0.14051f
C17577 VPWR.n927 VGND 0.14051f
C17578 VPWR.t600 VGND 0.03709f
C17579 VPWR.t436 VGND 0.0299f
C17580 VPWR.n928 VGND 0.09693f
C17581 VPWR.t1249 VGND 0.08295f
C17582 VPWR.t435 VGND 0.09401f
C17583 VPWR.t456 VGND 0.03709f
C17584 VPWR.t947 VGND 0.0299f
C17585 VPWR.n929 VGND 0.09693f
C17586 VPWR.t446 VGND 0.03709f
C17587 VPWR.t805 VGND 0.0299f
C17588 VPWR.n930 VGND 0.09693f
C17589 VPWR.t1204 VGND 0.14747f
C17590 VPWR.t1531 VGND 0.08295f
C17591 VPWR.t1236 VGND 0.09401f
C17592 VPWR.t1205 VGND 0.03709f
C17593 VPWR.t1237 VGND 0.0299f
C17594 VPWR.n931 VGND 0.09693f
C17595 VPWR.n932 VGND 0.01815f
C17596 VPWR.n933 VGND -0.00319f
C17597 VPWR.n934 VGND 0.09471f
C17598 VPWR.t1025 VGND 0.11982f
C17599 VPWR.t1533 VGND 0.08295f
C17600 VPWR.t1438 VGND 0.09401f
C17601 VPWR.t1026 VGND 0.03709f
C17602 VPWR.t1439 VGND 0.0299f
C17603 VPWR.n935 VGND 0.09693f
C17604 VPWR.n936 VGND 0.01815f
C17605 VPWR.n937 VGND -0.00319f
C17606 VPWR.n938 VGND 0.09471f
C17607 VPWR.t1407 VGND 0.11982f
C17608 VPWR.t527 VGND 0.08295f
C17609 VPWR.t1885 VGND 0.09401f
C17610 VPWR.t1408 VGND 0.03709f
C17611 VPWR.t1886 VGND 0.0299f
C17612 VPWR.n939 VGND 0.09693f
C17613 VPWR.n940 VGND 0.01815f
C17614 VPWR.n941 VGND -0.00319f
C17615 VPWR.n942 VGND 0.09471f
C17616 VPWR.t384 VGND 0.11982f
C17617 VPWR.t1674 VGND 0.08295f
C17618 VPWR.t1289 VGND 0.09401f
C17619 VPWR.t385 VGND 0.03709f
C17620 VPWR.t1290 VGND 0.0299f
C17621 VPWR.n943 VGND 0.09693f
C17622 VPWR.n944 VGND 0.01815f
C17623 VPWR.n945 VGND -0.00319f
C17624 VPWR.n946 VGND 0.09471f
C17625 VPWR.t553 VGND 0.11982f
C17626 VPWR.t1500 VGND 0.08295f
C17627 VPWR.t1706 VGND 0.09401f
C17628 VPWR.t554 VGND 0.03709f
C17629 VPWR.t1707 VGND 0.0299f
C17630 VPWR.n947 VGND 0.09693f
C17631 VPWR.n948 VGND 0.01815f
C17632 VPWR.n949 VGND -0.00319f
C17633 VPWR.n950 VGND 0.09471f
C17634 VPWR.t1704 VGND 0.11982f
C17635 VPWR.t1341 VGND 0.08295f
C17636 VPWR.t282 VGND 0.09401f
C17637 VPWR.t1705 VGND 0.03709f
C17638 VPWR.t283 VGND 0.0299f
C17639 VPWR.n951 VGND 0.09693f
C17640 VPWR.n952 VGND 0.01815f
C17641 VPWR.n953 VGND -0.00319f
C17642 VPWR.n954 VGND 0.09471f
C17643 VPWR.t212 VGND 0.11982f
C17644 VPWR.t1673 VGND 0.08295f
C17645 VPWR.t537 VGND 0.09401f
C17646 VPWR.t213 VGND 0.03709f
C17647 VPWR.t538 VGND 0.0299f
C17648 VPWR.n955 VGND 0.09693f
C17649 VPWR.n956 VGND 0.01815f
C17650 VPWR.n957 VGND -0.00319f
C17651 VPWR.n958 VGND 0.09471f
C17652 VPWR.t1622 VGND 0.11982f
C17653 VPWR.t1530 VGND 0.08295f
C17654 VPWR.t1434 VGND 0.09401f
C17655 VPWR.t1623 VGND 0.03709f
C17656 VPWR.t1435 VGND 0.0299f
C17657 VPWR.n959 VGND 0.09693f
C17658 VPWR.n960 VGND 0.01815f
C17659 VPWR.n961 VGND -0.00319f
C17660 VPWR.n962 VGND 0.09471f
C17661 VPWR.t1432 VGND 0.11982f
C17662 VPWR.t1503 VGND 0.08295f
C17663 VPWR.t1176 VGND 0.09401f
C17664 VPWR.t1433 VGND 0.03709f
C17665 VPWR.t1177 VGND 0.0299f
C17666 VPWR.n963 VGND 0.09693f
C17667 VPWR.n964 VGND 0.01815f
C17668 VPWR.n965 VGND -0.00319f
C17669 VPWR.n966 VGND 0.09471f
C17670 VPWR.t1901 VGND 0.11982f
C17671 VPWR.t1340 VGND 0.08295f
C17672 VPWR.t1068 VGND 0.09401f
C17673 VPWR.t1902 VGND 0.03709f
C17674 VPWR.t1069 VGND 0.0299f
C17675 VPWR.n967 VGND 0.09693f
C17676 VPWR.n968 VGND 0.01815f
C17677 VPWR.n969 VGND -0.00319f
C17678 VPWR.n970 VGND 0.09471f
C17679 VPWR.t1058 VGND 0.11982f
C17680 VPWR.t1672 VGND 0.08295f
C17681 VPWR.t68 VGND 0.09401f
C17682 VPWR.t1059 VGND 0.03709f
C17683 VPWR.t69 VGND 0.0299f
C17684 VPWR.n971 VGND 0.09693f
C17685 VPWR.n972 VGND 0.01815f
C17686 VPWR.n973 VGND -0.00319f
C17687 VPWR.n974 VGND 0.09471f
C17688 VPWR.t90 VGND 0.11982f
C17689 VPWR.t1502 VGND 0.08295f
C17690 VPWR.t1492 VGND 0.09401f
C17691 VPWR.t91 VGND 0.03709f
C17692 VPWR.t1493 VGND 0.0299f
C17693 VPWR.n975 VGND 0.09693f
C17694 VPWR.n976 VGND 0.01815f
C17695 VPWR.n977 VGND -0.00319f
C17696 VPWR.n978 VGND 0.09471f
C17697 VPWR.t559 VGND 0.11982f
C17698 VPWR.t1339 VGND 0.08295f
C17699 VPWR.t1361 VGND 0.09401f
C17700 VPWR.t560 VGND 0.03709f
C17701 VPWR.t1362 VGND 0.0299f
C17702 VPWR.n979 VGND 0.09693f
C17703 VPWR.n980 VGND 0.01815f
C17704 VPWR.n981 VGND -0.00319f
C17705 VPWR.n982 VGND 0.09471f
C17706 VPWR.t1359 VGND 0.11982f
C17707 VPWR.t1338 VGND 0.08295f
C17708 VPWR.t1486 VGND 0.09401f
C17709 VPWR.t1360 VGND 0.03709f
C17710 VPWR.t1487 VGND 0.0299f
C17711 VPWR.n983 VGND 0.09693f
C17712 VPWR.n984 VGND 0.01815f
C17713 VPWR.n985 VGND -0.00319f
C17714 VPWR.n986 VGND 0.09471f
C17715 VPWR.t1652 VGND 0.11982f
C17716 VPWR.t1532 VGND 0.08295f
C17717 VPWR.t1373 VGND 0.09401f
C17718 VPWR.t1653 VGND 0.03709f
C17719 VPWR.t1374 VGND 0.0299f
C17720 VPWR.n987 VGND 0.09693f
C17721 VPWR.n988 VGND 0.01815f
C17722 VPWR.n989 VGND -0.00319f
C17723 VPWR.n990 VGND 0.09471f
C17724 VPWR.t445 VGND 0.11982f
C17725 VPWR.t1501 VGND 0.08295f
C17726 VPWR.t804 VGND 0.14528f
C17727 VPWR.n991 VGND 0.08265f
C17728 VPWR.n992 VGND 0.01815f
C17729 VPWR.n993 VGND 0.14051f
C17730 VPWR.n994 VGND 6.08253f
C17731 VPWR.n995 VGND 0.06632f
C17732 VPWR.n996 VGND -0.01884f
C17733 VPWR.t2027 VGND 0.01176f
C17734 VPWR.t922 VGND 0.01238f
C17735 VPWR.n997 VGND 0.03f
C17736 VPWR.n998 VGND 0.01873f
C17737 VPWR.t924 VGND 0.02986f
C17738 VPWR.n999 VGND 0.0649f
C17739 VPWR.t916 VGND 0.0299f
C17740 VPWR.n1000 VGND 0.04757f
C17741 VPWR.t447 VGND 0.09401f
C17742 VPWR.t1928 VGND 0.01176f
C17743 VPWR.t808 VGND 0.01238f
C17744 VPWR.n1001 VGND 0.03f
C17745 VPWR.n1002 VGND 0.01873f
C17746 VPWR.t810 VGND 0.02986f
C17747 VPWR.n1003 VGND 0.0649f
C17748 VPWR.t448 VGND 0.0299f
C17749 VPWR.n1004 VGND 0.04757f
C17750 VPWR.n1005 VGND -0.01884f
C17751 VPWR.n1006 VGND 0.06632f
C17752 VPWR.t2037 VGND 0.01176f
C17753 VPWR.t891 VGND 0.01238f
C17754 VPWR.n1007 VGND 0.03075f
C17755 VPWR.n1008 VGND 0.01916f
C17756 VPWR.n1009 VGND 0.06224f
C17757 VPWR.n1010 VGND 0.09842f
C17758 VPWR.n1011 VGND 0.05494f
C17759 VPWR.n1012 VGND 0.06632f
C17760 VPWR.n1013 VGND -0.01884f
C17761 VPWR.t2036 VGND 0.01176f
C17762 VPWR.t896 VGND 0.01238f
C17763 VPWR.n1014 VGND 0.03f
C17764 VPWR.n1015 VGND 0.01873f
C17765 VPWR.t898 VGND 0.02986f
C17766 VPWR.n1016 VGND 0.0649f
C17767 VPWR.t1511 VGND 0.0299f
C17768 VPWR.n1017 VGND 0.04757f
C17769 VPWR.t1510 VGND 0.09401f
C17770 VPWR.t667 VGND 0.11982f
C17771 VPWR.t2025 VGND 0.01176f
C17772 VPWR.t888 VGND 0.01238f
C17773 VPWR.n1018 VGND 0.03f
C17774 VPWR.n1019 VGND 0.01873f
C17775 VPWR.t890 VGND 0.02986f
C17776 VPWR.n1020 VGND 0.0649f
C17777 VPWR.t175 VGND 0.0299f
C17778 VPWR.n1021 VGND 0.04757f
C17779 VPWR.n1022 VGND 0.02426f
C17780 VPWR.n1023 VGND 0.19562f
C17781 VPWR.n1024 VGND 0.08433f
C17782 VPWR.n1025 VGND 0.0313f
C17783 VPWR.t879 VGND 0.03709f
C17784 VPWR.t874 VGND 0.0299f
C17785 VPWR.n1026 VGND 0.09693f
C17786 VPWR.t873 VGND 0.09401f
C17787 VPWR.t742 VGND 0.11982f
C17788 VPWR.t632 VGND 0.03709f
C17789 VPWR.t627 VGND 0.0299f
C17790 VPWR.n1027 VGND 0.09693f
C17791 VPWR.t743 VGND 0.03709f
C17792 VPWR.t738 VGND 0.0299f
C17793 VPWR.n1028 VGND 0.09693f
C17794 VPWR.t740 VGND 0.08295f
C17795 VPWR.t737 VGND 0.14528f
C17796 VPWR.n1029 VGND 0.08262f
C17797 VPWR.n1030 VGND 0.00608f
C17798 VPWR.n1031 VGND 0.02407f
C17799 VPWR.t1989 VGND 0.01176f
C17800 VPWR.t736 VGND 0.01238f
C17801 VPWR.n1032 VGND 0.03074f
C17802 VPWR.n1033 VGND 0.02885f
C17803 VPWR.n1034 VGND 0.01916f
C17804 VPWR.n1035 VGND 0.17759f
C17805 VPWR.t1943 VGND 0.01176f
C17806 VPWR.t872 VGND 0.01238f
C17807 VPWR.n1036 VGND 0.03074f
C17808 VPWR.n1037 VGND 0.02885f
C17809 VPWR.n1038 VGND 0.01916f
C17810 VPWR.n1039 VGND 0.03332f
C17811 VPWR.t1944 VGND 0.01176f
C17812 VPWR.t860 VGND 0.01238f
C17813 VPWR.n1040 VGND 0.03074f
C17814 VPWR.n1041 VGND 0.02256f
C17815 VPWR.n1042 VGND 0.02426f
C17816 VPWR.t1993 VGND 0.01176f
C17817 VPWR.t728 VGND 0.01238f
C17818 VPWR.n1043 VGND 0.03074f
C17819 VPWR.n1044 VGND 0.02256f
C17820 VPWR.n1045 VGND 0.02426f
C17821 VPWR.t2044 VGND 0.01176f
C17822 VPWR.t988 VGND 0.01238f
C17823 VPWR.n1046 VGND 0.03074f
C17824 VPWR.n1047 VGND 0.02256f
C17825 VPWR.n1048 VGND 0.02426f
C17826 VPWR.t1949 VGND 0.01176f
C17827 VPWR.t852 VGND 0.01238f
C17828 VPWR.n1049 VGND 0.03074f
C17829 VPWR.n1050 VGND 0.02256f
C17830 VPWR.n1051 VGND 0.02426f
C17831 VPWR.t2000 VGND 0.01176f
C17832 VPWR.t720 VGND 0.01238f
C17833 VPWR.n1052 VGND 0.03074f
C17834 VPWR.n1053 VGND 0.02256f
C17835 VPWR.n1054 VGND 0.02426f
C17836 VPWR.t2008 VGND 0.01176f
C17837 VPWR.t678 VGND 0.01238f
C17838 VPWR.n1055 VGND 0.03074f
C17839 VPWR.n1056 VGND 0.02256f
C17840 VPWR.n1057 VGND 0.02426f
C17841 VPWR.t2050 VGND 0.01176f
C17842 VPWR.t959 VGND 0.01238f
C17843 VPWR.n1058 VGND 0.03074f
C17844 VPWR.n1059 VGND 0.02256f
C17845 VPWR.n1060 VGND 0.02426f
C17846 VPWR.t1957 VGND 0.01176f
C17847 VPWR.t817 VGND 0.01238f
C17848 VPWR.n1061 VGND 0.03074f
C17849 VPWR.n1062 VGND 0.02256f
C17850 VPWR.n1063 VGND 0.02426f
C17851 VPWR.t1973 VGND 0.01176f
C17852 VPWR.t787 VGND 0.01238f
C17853 VPWR.n1064 VGND 0.03074f
C17854 VPWR.n1065 VGND 0.02256f
C17855 VPWR.n1066 VGND 0.02426f
C17856 VPWR.t2056 VGND 0.01176f
C17857 VPWR.t951 VGND 0.01238f
C17858 VPWR.n1067 VGND 0.03074f
C17859 VPWR.n1068 VGND 0.02256f
C17860 VPWR.n1069 VGND 0.02426f
C17861 VPWR.t2068 VGND 0.01176f
C17862 VPWR.t912 VGND 0.01238f
C17863 VPWR.n1070 VGND 0.03074f
C17864 VPWR.n1071 VGND 0.02256f
C17865 VPWR.n1072 VGND 0.02426f
C17866 VPWR.t1930 VGND 0.01176f
C17867 VPWR.t899 VGND 0.01238f
C17868 VPWR.n1073 VGND 0.03074f
C17869 VPWR.n1074 VGND 0.02256f
C17870 VPWR.t2018 VGND 0.01176f
C17871 VPWR.t658 VGND 0.01238f
C17872 VPWR.n1075 VGND 0.03075f
C17873 VPWR.n1076 VGND 0.01916f
C17874 VPWR.n1077 VGND 0.01916f
C17875 VPWR.n1078 VGND 0.03332f
C17876 VPWR.n1079 VGND 0.17759f
C17877 VPWR.n1080 VGND 0.01916f
C17878 VPWR.n1081 VGND 0.03332f
C17879 VPWR.n1082 VGND 0.17759f
C17880 VPWR.n1083 VGND 0.01916f
C17881 VPWR.n1084 VGND 0.03332f
C17882 VPWR.n1085 VGND 0.17759f
C17883 VPWR.n1086 VGND 0.01916f
C17884 VPWR.n1087 VGND 0.03332f
C17885 VPWR.n1088 VGND 0.17759f
C17886 VPWR.n1089 VGND 0.01916f
C17887 VPWR.n1090 VGND 0.03332f
C17888 VPWR.n1091 VGND 0.17759f
C17889 VPWR.n1092 VGND 0.01916f
C17890 VPWR.n1093 VGND 0.03332f
C17891 VPWR.n1094 VGND 0.17759f
C17892 VPWR.n1095 VGND 0.01916f
C17893 VPWR.n1096 VGND 0.03332f
C17894 VPWR.n1097 VGND 0.17759f
C17895 VPWR.n1098 VGND 0.01916f
C17896 VPWR.n1099 VGND 0.03332f
C17897 VPWR.n1100 VGND 0.17759f
C17898 VPWR.n1101 VGND 0.01916f
C17899 VPWR.n1102 VGND 0.03332f
C17900 VPWR.n1103 VGND 0.17759f
C17901 VPWR.n1104 VGND 0.01916f
C17902 VPWR.n1105 VGND 0.03332f
C17903 VPWR.n1106 VGND 0.17759f
C17904 VPWR.n1107 VGND 0.01916f
C17905 VPWR.n1108 VGND 0.03332f
C17906 VPWR.n1109 VGND 0.23958f
C17907 VPWR.n1110 VGND 0.03605f
C17908 VPWR.t2019 VGND 0.01176f
C17909 VPWR.t656 VGND 0.01238f
C17910 VPWR.n1111 VGND 0.03074f
C17911 VPWR.n1112 VGND 0.02256f
C17912 VPWR.n1113 VGND 0.02485f
C17913 VPWR.t2020 VGND 0.01176f
C17914 VPWR.t653 VGND 0.01238f
C17915 VPWR.n1114 VGND 0.03074f
C17916 VPWR.n1115 VGND 0.02885f
C17917 VPWR.t660 VGND 0.03709f
C17918 VPWR.t655 VGND 0.0299f
C17919 VPWR.n1116 VGND 0.09693f
C17920 VPWR.t659 VGND 0.14747f
C17921 VPWR.t657 VGND 0.08295f
C17922 VPWR.t654 VGND 0.09401f
C17923 VPWR.t876 VGND 0.08295f
C17924 VPWR.t878 VGND 0.11982f
C17925 VPWR.t764 VGND 0.03709f
C17926 VPWR.t859 VGND 0.0299f
C17927 VPWR.n1117 VGND 0.09693f
C17928 VPWR.n1118 VGND 0.00608f
C17929 VPWR.n1119 VGND -0.00323f
C17930 VPWR.n1120 VGND 0.09471f
C17931 VPWR.t858 VGND 0.09401f
C17932 VPWR.t861 VGND 0.08295f
C17933 VPWR.t763 VGND 0.11982f
C17934 VPWR.t732 VGND 0.03709f
C17935 VPWR.t727 VGND 0.0299f
C17936 VPWR.n1121 VGND 0.09693f
C17937 VPWR.n1122 VGND 0.00608f
C17938 VPWR.n1123 VGND -0.00323f
C17939 VPWR.n1124 VGND 0.09471f
C17940 VPWR.t726 VGND 0.09401f
C17941 VPWR.t729 VGND 0.08295f
C17942 VPWR.t731 VGND 0.11982f
C17943 VPWR.t992 VGND 0.03709f
C17944 VPWR.t984 VGND 0.0299f
C17945 VPWR.n1125 VGND 0.09693f
C17946 VPWR.n1126 VGND 0.00608f
C17947 VPWR.n1127 VGND -0.00323f
C17948 VPWR.n1128 VGND 0.09471f
C17949 VPWR.t983 VGND 0.09401f
C17950 VPWR.t989 VGND 0.08295f
C17951 VPWR.t991 VGND 0.11982f
C17952 VPWR.t856 VGND 0.03709f
C17953 VPWR.t936 VGND 0.0299f
C17954 VPWR.n1129 VGND 0.09693f
C17955 VPWR.n1130 VGND 0.00608f
C17956 VPWR.n1131 VGND -0.00323f
C17957 VPWR.n1132 VGND 0.09471f
C17958 VPWR.t935 VGND 0.09401f
C17959 VPWR.t853 VGND 0.08295f
C17960 VPWR.t855 VGND 0.11982f
C17961 VPWR.t724 VGND 0.03709f
C17962 VPWR.t719 VGND 0.0299f
C17963 VPWR.n1133 VGND 0.09693f
C17964 VPWR.n1134 VGND 0.00608f
C17965 VPWR.n1135 VGND -0.00323f
C17966 VPWR.n1136 VGND 0.09471f
C17967 VPWR.t718 VGND 0.09401f
C17968 VPWR.t721 VGND 0.08295f
C17969 VPWR.t723 VGND 0.11982f
C17970 VPWR.t682 VGND 0.03709f
C17971 VPWR.t703 VGND 0.0299f
C17972 VPWR.n1137 VGND 0.09693f
C17973 VPWR.n1138 VGND 0.00608f
C17974 VPWR.n1139 VGND -0.00323f
C17975 VPWR.n1140 VGND 0.09471f
C17976 VPWR.t702 VGND 0.09401f
C17977 VPWR.t679 VGND 0.08295f
C17978 VPWR.t681 VGND 0.11982f
C17979 VPWR.t963 VGND 0.03709f
C17980 VPWR.t958 VGND 0.0299f
C17981 VPWR.n1141 VGND 0.09693f
C17982 VPWR.n1142 VGND 0.00608f
C17983 VPWR.n1143 VGND -0.00323f
C17984 VPWR.n1144 VGND 0.09471f
C17985 VPWR.t957 VGND 0.09401f
C17986 VPWR.t960 VGND 0.08295f
C17987 VPWR.t962 VGND 0.11982f
C17988 VPWR.t799 VGND 0.03709f
C17989 VPWR.t816 VGND 0.0299f
C17990 VPWR.n1145 VGND 0.09693f
C17991 VPWR.n1146 VGND 0.00608f
C17992 VPWR.n1147 VGND -0.00323f
C17993 VPWR.n1148 VGND 0.09471f
C17994 VPWR.t815 VGND 0.09401f
C17995 VPWR.t818 VGND 0.08295f
C17996 VPWR.t798 VGND 0.11982f
C17997 VPWR.t791 VGND 0.03709f
C17998 VPWR.t786 VGND 0.0299f
C17999 VPWR.n1149 VGND 0.09693f
C18000 VPWR.n1150 VGND 0.00608f
C18001 VPWR.n1151 VGND -0.00323f
C18002 VPWR.n1152 VGND 0.09471f
C18003 VPWR.t785 VGND 0.09401f
C18004 VPWR.t788 VGND 0.08295f
C18005 VPWR.t790 VGND 0.11982f
C18006 VPWR.t955 VGND 0.03709f
C18007 VPWR.t950 VGND 0.0299f
C18008 VPWR.n1153 VGND 0.09693f
C18009 VPWR.n1154 VGND 0.00608f
C18010 VPWR.n1155 VGND -0.00323f
C18011 VPWR.n1156 VGND 0.09471f
C18012 VPWR.t949 VGND 0.09401f
C18013 VPWR.t952 VGND 0.08295f
C18014 VPWR.t954 VGND 0.11982f
C18015 VPWR.t919 VGND 0.03709f
C18016 VPWR.t911 VGND 0.0299f
C18017 VPWR.n1157 VGND 0.09693f
C18018 VPWR.n1158 VGND 0.00608f
C18019 VPWR.n1159 VGND -0.00323f
C18020 VPWR.n1160 VGND 0.09471f
C18021 VPWR.t910 VGND 0.09401f
C18022 VPWR.t913 VGND 0.08295f
C18023 VPWR.t918 VGND 0.11982f
C18024 VPWR.t802 VGND 0.03709f
C18025 VPWR.t895 VGND 0.0299f
C18026 VPWR.n1161 VGND 0.09693f
C18027 VPWR.n1162 VGND 0.00608f
C18028 VPWR.n1163 VGND -0.00323f
C18029 VPWR.n1164 VGND 0.09471f
C18030 VPWR.t894 VGND 0.09401f
C18031 VPWR.t900 VGND 0.08295f
C18032 VPWR.t801 VGND 0.11982f
C18033 VPWR.n1165 VGND 0.09471f
C18034 VPWR.n1166 VGND -0.00323f
C18035 VPWR.n1167 VGND 0.00608f
C18036 VPWR.n1168 VGND 0.14051f
C18037 VPWR.n1169 VGND 0.01815f
C18038 VPWR.n1170 VGND 0.06632f
C18039 VPWR.n1171 VGND 0.05494f
C18040 VPWR.n1172 VGND 0.04733f
C18041 VPWR.t156 VGND 0.98528f
C18042 VPWR.n1173 VGND 0.53738f
C18043 VPWR.t161 VGND 0.98528f
C18044 VPWR.n1174 VGND 0.41792f
C18045 VPWR.n1175 VGND 0.29367f
C18046 VPWR.t1351 VGND 0.05772f
C18047 VPWR.n1176 VGND 0.00929f
C18048 VPWR.t166 VGND 0.01447f
C18049 VPWR.t604 VGND 0.01447f
C18050 VPWR.n1177 VGND 0.03177f
C18051 VPWR.t605 VGND 0.01447f
C18052 VPWR.t1041 VGND 0.01447f
C18053 VPWR.n1178 VGND 0.03172f
C18054 VPWR.t204 VGND 0.01447f
C18055 VPWR.t203 VGND 0.01447f
C18056 VPWR.n1179 VGND 0.03172f
C18057 VPWR.n1180 VGND 0.10523f
C18058 VPWR.n1181 VGND 0.18361f
C18059 VPWR.n1182 VGND 0.05813f
C18060 VPWR.n1183 VGND 0.0427f
C18061 VPWR.t199 VGND 0.01447f
C18062 VPWR.t205 VGND 0.01447f
C18063 VPWR.n1184 VGND 0.03177f
C18064 VPWR.n1185 VGND 0.13029f
C18065 VPWR.n1186 VGND 0.0113f
C18066 VPWR.n1187 VGND 0.01646f
C18067 VPWR.n1188 VGND 0.01929f
C18068 VPWR.n1189 VGND 0.02829f
C18069 VPWR.t1350 VGND 0.05772f
C18070 VPWR.n1190 VGND 0.15208f
C18071 VPWR.n1191 VGND 0.01221f
C18072 VPWR.t1804 VGND 0.05771f
C18073 VPWR.t453 VGND 0.05771f
C18074 VPWR.n1192 VGND 0.13578f
C18075 VPWR.n1193 VGND 0.33894f
C18076 VPWR.n1194 VGND 1.65711f
C18077 VPWR.n1195 VGND 0.04733f
C18078 VPWR.t160 VGND 0.98528f
C18079 VPWR.n1196 VGND 0.53738f
C18080 VPWR.t1005 VGND 0.98528f
C18081 VPWR.n1197 VGND 0.41792f
C18082 VPWR.n1198 VGND 0.29631f
C18083 VPWR.n1199 VGND 0.00929f
C18084 VPWR.t416 VGND 0.01447f
C18085 VPWR.t414 VGND 0.01447f
C18086 VPWR.n1200 VGND 0.03177f
C18087 VPWR.t413 VGND 0.01447f
C18088 VPWR.t411 VGND 0.01447f
C18089 VPWR.n1201 VGND 0.03172f
C18090 VPWR.t1449 VGND 0.01447f
C18091 VPWR.t1450 VGND 0.01447f
C18092 VPWR.n1202 VGND 0.03172f
C18093 VPWR.n1203 VGND 0.10523f
C18094 VPWR.n1204 VGND 0.18361f
C18095 VPWR.n1205 VGND 0.05813f
C18096 VPWR.n1206 VGND 0.0427f
C18097 VPWR.t1821 VGND 0.01447f
C18098 VPWR.t1823 VGND 0.01447f
C18099 VPWR.n1207 VGND 0.03177f
C18100 VPWR.n1208 VGND 0.13029f
C18101 VPWR.n1209 VGND 0.0113f
C18102 VPWR.n1210 VGND 0.01646f
C18103 VPWR.n1211 VGND 0.01929f
C18104 VPWR.n1212 VGND 0.02778f
C18105 VPWR.n1213 VGND 0.00774f
C18106 VPWR.t1352 VGND 0.05764f
C18107 VPWR.n1214 VGND 0.06161f
C18108 VPWR.n1215 VGND 0.00738f
C18109 VPWR.t180 VGND 0.05776f
C18110 VPWR.n1216 VGND 0.092f
C18111 VPWR.n1217 VGND 0.33894f
C18112 VPWR.n1218 VGND 1.65711f
C18113 VPWR.n1219 VGND 0.04733f
C18114 VPWR.t8 VGND 0.98528f
C18115 VPWR.n1220 VGND 0.53738f
C18116 VPWR.t1 VGND 0.98528f
C18117 VPWR.n1221 VGND 0.41792f
C18118 VPWR.n1222 VGND 0.29631f
C18119 VPWR.n1223 VGND 0.00929f
C18120 VPWR.t55 VGND 0.01447f
C18121 VPWR.t53 VGND 0.01447f
C18122 VPWR.n1224 VGND 0.03177f
C18123 VPWR.t52 VGND 0.01447f
C18124 VPWR.t51 VGND 0.01447f
C18125 VPWR.n1225 VGND 0.03172f
C18126 VPWR.t1314 VGND 0.01447f
C18127 VPWR.t1321 VGND 0.01447f
C18128 VPWR.n1226 VGND 0.03172f
C18129 VPWR.n1227 VGND 0.10523f
C18130 VPWR.n1228 VGND 0.18361f
C18131 VPWR.n1229 VGND 0.05813f
C18132 VPWR.n1230 VGND 0.0427f
C18133 VPWR.t1318 VGND 0.01447f
C18134 VPWR.t1315 VGND 0.01447f
C18135 VPWR.n1231 VGND 0.03177f
C18136 VPWR.n1232 VGND 0.13029f
C18137 VPWR.n1233 VGND 0.0113f
C18138 VPWR.n1234 VGND 0.01646f
C18139 VPWR.n1235 VGND 0.01929f
C18140 VPWR.n1236 VGND 0.02778f
C18141 VPWR.n1237 VGND 0.01412f
C18142 VPWR.n1238 VGND 0.01321f
C18143 VPWR.t1805 VGND 0.05776f
C18144 VPWR.t454 VGND 0.05776f
C18145 VPWR.n1239 VGND 0.1706f
C18146 VPWR.n1240 VGND 0.33894f
C18147 VPWR.n1241 VGND 1.65711f
C18148 VPWR.t196 VGND 0.05767f
C18149 VPWR.t487 VGND 0.05776f
C18150 VPWR.t198 VGND 0.05728f
C18151 VPWR.n1242 VGND 0.14851f
C18152 VPWR.t155 VGND 0.05662f
C18153 VPWR.n1243 VGND 0.06842f
C18154 VPWR.n1244 VGND 0.04733f
C18155 VPWR.t1448 VGND 0.0545f
C18156 VPWR.n1245 VGND 0.05184f
C18157 VPWR.t402 VGND 0.01447f
C18158 VPWR.t1831 VGND 0.01447f
C18159 VPWR.n1246 VGND 0.03162f
C18160 VPWR.t348 VGND 0.05064f
C18161 VPWR.n1247 VGND 0.07595f
C18162 VPWR.n1248 VGND 0.04733f
C18163 VPWR.t10 VGND 0.0577f
C18164 VPWR.n1249 VGND 0.07264f
C18165 VPWR.n1250 VGND 0.02778f
C18166 VPWR.n1251 VGND 0.04733f
C18167 VPWR.n1252 VGND 0.01221f
C18168 VPWR.t1833 VGND 0.01447f
C18169 VPWR.t1835 VGND 0.01447f
C18170 VPWR.n1253 VGND 0.03162f
C18171 VPWR.n1254 VGND 0.04633f
C18172 VPWR.n1255 VGND 0.01221f
C18173 VPWR.n1256 VGND 0.0355f
C18174 VPWR.n1257 VGND 0.0355f
C18175 VPWR.n1258 VGND 0.04733f
C18176 VPWR.n1259 VGND 0.00838f
C18177 VPWR.t1855 VGND 0.01447f
C18178 VPWR.t406 VGND 0.01447f
C18179 VPWR.n1260 VGND 0.03162f
C18180 VPWR.n1261 VGND 0.0364f
C18181 VPWR.t158 VGND 0.01447f
C18182 VPWR.t229 VGND 0.01447f
C18183 VPWR.n1262 VGND 0.03162f
C18184 VPWR.n1263 VGND 0.04023f
C18185 VPWR.n1264 VGND 0.01066f
C18186 VPWR.n1265 VGND 0.04296f
C18187 VPWR.n1266 VGND 0.0162f
C18188 VPWR.n1267 VGND 0.00638f
C18189 VPWR.t1419 VGND 0.04853f
C18190 VPWR.t195 VGND 0.10919f
C18191 VPWR.t486 VGND 0.12739f
C18192 VPWR.t197 VGND 0.23658f
C18193 VPWR.t9 VGND 0.12729f
C18194 VPWR.t1834 VGND 0.14449f
C18195 VPWR.t1832 VGND 0.14048f
C18196 VPWR.t1830 VGND 0.22466f
C18197 VPWR.t401 VGND 0.19108f
C18198 VPWR.t347 VGND 0.12739f
C18199 VPWR.t405 VGND 0.12739f
C18200 VPWR.t228 VGND 0.12739f
C18201 VPWR.t1854 VGND 0.12739f
C18202 VPWR.t157 VGND 0.12739f
C18203 VPWR.t1447 VGND 0.12739f
C18204 VPWR.t154 VGND 0.12587f
C18205 VPWR.n1268 VGND 0.43293f
C18206 VPWR.n1269 VGND 0.17591f
C18207 VPWR.n1270 VGND 0.01929f
C18208 VPWR.n1271 VGND 0.0355f
C18209 VPWR.n1272 VGND 0.0427f
C18210 VPWR.n1273 VGND 0.01093f
C18211 VPWR.n1274 VGND 0.06419f
C18212 VPWR.n1275 VGND 0.31964f
C18213 VPWR.n1276 VGND 1.65711f
C18214 VPWR.t1050 VGND 0.05674f
C18215 VPWR.t1055 VGND 0.05658f
C18216 VPWR.t485 VGND 0.05771f
C18217 VPWR.n1277 VGND 0.08042f
C18218 VPWR.t606 VGND 0.05509f
C18219 VPWR.t206 VGND 0.05509f
C18220 VPWR.n1278 VGND 0.09995f
C18221 VPWR.n1279 VGND 0.04733f
C18222 VPWR.n1280 VGND 0.0092f
C18223 VPWR.n1281 VGND 0.04733f
C18224 VPWR.t167 VGND 0.01447f
C18225 VPWR.t1786 VGND 0.01447f
C18226 VPWR.n1282 VGND 0.03162f
C18227 VPWR.t207 VGND 0.01447f
C18228 VPWR.t1000 VGND 0.01447f
C18229 VPWR.n1283 VGND 0.03162f
C18230 VPWR.n1284 VGND 0.06442f
C18231 VPWR.t1002 VGND 0.0577f
C18232 VPWR.t1836 VGND 0.0577f
C18233 VPWR.n1285 VGND 0.13299f
C18234 VPWR.n1286 VGND 0.02778f
C18235 VPWR.n1287 VGND 0.04733f
C18236 VPWR.n1288 VGND 0.01221f
C18237 VPWR.t1669 VGND 0.01447f
C18238 VPWR.t3 VGND 0.01447f
C18239 VPWR.n1289 VGND 0.03162f
C18240 VPWR.t1006 VGND 0.01447f
C18241 VPWR.t225 VGND 0.01447f
C18242 VPWR.n1290 VGND 0.03162f
C18243 VPWR.n1291 VGND 0.0728f
C18244 VPWR.n1292 VGND 0.01221f
C18245 VPWR.n1293 VGND 0.04733f
C18246 VPWR.n1294 VGND 0.04733f
C18247 VPWR.n1295 VGND 0.04733f
C18248 VPWR.n1296 VGND 0.01139f
C18249 VPWR.t1042 VGND 0.01447f
C18250 VPWR.t603 VGND 0.01447f
C18251 VPWR.n1297 VGND 0.03162f
C18252 VPWR.t202 VGND 0.01447f
C18253 VPWR.t201 VGND 0.01447f
C18254 VPWR.n1298 VGND 0.03162f
C18255 VPWR.n1299 VGND 0.06442f
C18256 VPWR.n1300 VGND 0.01066f
C18257 VPWR.n1301 VGND 0.00993f
C18258 VPWR.n1302 VGND 0.04733f
C18259 VPWR.n1303 VGND 0.0355f
C18260 VPWR.n1304 VGND 0.00802f
C18261 VPWR.t2 VGND 0.98528f
C18262 VPWR.n1305 VGND 0.53738f
C18263 VPWR.t200 VGND 0.98528f
C18264 VPWR.n1306 VGND 0.41792f
C18265 VPWR.n1307 VGND 0.29367f
C18266 VPWR.n1308 VGND 0.01929f
C18267 VPWR.n1309 VGND 0.0355f
C18268 VPWR.n1310 VGND 0.04296f
C18269 VPWR.n1311 VGND 0.01075f
C18270 VPWR.n1312 VGND 0.05885f
C18271 VPWR.n1313 VGND 0.07971f
C18272 VPWR.n1314 VGND 0.31939f
C18273 VPWR.n1315 VGND 1.65711f
C18274 VPWR.t1630 VGND 0.05764f
C18275 VPWR.t1858 VGND 0.05764f
C18276 VPWR.n1316 VGND 0.01412f
C18277 VPWR.t412 VGND 0.05509f
C18278 VPWR.t1822 VGND 0.05509f
C18279 VPWR.n1317 VGND 0.09995f
C18280 VPWR.n1318 VGND 0.04733f
C18281 VPWR.n1319 VGND 0.0092f
C18282 VPWR.n1320 VGND 0.04733f
C18283 VPWR.t417 VGND 0.01447f
C18284 VPWR.t1003 VGND 0.01447f
C18285 VPWR.n1321 VGND 0.03162f
C18286 VPWR.t1010 VGND 0.01447f
C18287 VPWR.t1837 VGND 0.01447f
C18288 VPWR.n1322 VGND 0.03162f
C18289 VPWR.n1323 VGND 0.06442f
C18290 VPWR.t1784 VGND 0.0577f
C18291 VPWR.t163 VGND 0.0577f
C18292 VPWR.n1324 VGND 0.13299f
C18293 VPWR.n1325 VGND 0.02778f
C18294 VPWR.n1326 VGND 0.04733f
C18295 VPWR.n1327 VGND 0.01221f
C18296 VPWR.t1008 VGND 0.01447f
C18297 VPWR.t227 VGND 0.01447f
C18298 VPWR.n1328 VGND 0.03162f
C18299 VPWR.t1785 VGND 0.01447f
C18300 VPWR.t1671 VGND 0.01447f
C18301 VPWR.n1329 VGND 0.03162f
C18302 VPWR.n1330 VGND 0.0728f
C18303 VPWR.n1331 VGND 0.01221f
C18304 VPWR.n1332 VGND 0.04733f
C18305 VPWR.n1333 VGND 0.04733f
C18306 VPWR.n1334 VGND 0.04733f
C18307 VPWR.n1335 VGND 0.01139f
C18308 VPWR.t418 VGND 0.01447f
C18309 VPWR.t415 VGND 0.01447f
C18310 VPWR.n1336 VGND 0.03162f
C18311 VPWR.t1009 VGND 0.01447f
C18312 VPWR.t1820 VGND 0.01447f
C18313 VPWR.n1337 VGND 0.03162f
C18314 VPWR.n1338 VGND 0.06442f
C18315 VPWR.n1339 VGND 0.01066f
C18316 VPWR.n1340 VGND 0.00993f
C18317 VPWR.n1341 VGND 0.04733f
C18318 VPWR.n1342 VGND 0.0355f
C18319 VPWR.n1343 VGND 0.00802f
C18320 VPWR.t226 VGND 0.98528f
C18321 VPWR.n1344 VGND 0.53738f
C18322 VPWR.t162 VGND 0.98528f
C18323 VPWR.n1345 VGND 0.41792f
C18324 VPWR.n1346 VGND 0.29631f
C18325 VPWR.n1347 VGND 0.01929f
C18326 VPWR.n1348 VGND 0.0355f
C18327 VPWR.n1349 VGND 0.04296f
C18328 VPWR.n1350 VGND 0.01093f
C18329 VPWR.n1351 VGND 0.11651f
C18330 VPWR.n1352 VGND 0.32454f
C18331 VPWR.n1353 VGND 1.65711f
C18332 VPWR.t54 VGND 0.05509f
C18333 VPWR.t1316 VGND 0.05509f
C18334 VPWR.n1354 VGND 0.09995f
C18335 VPWR.n1355 VGND 0.04733f
C18336 VPWR.n1356 VGND 0.0092f
C18337 VPWR.n1357 VGND 0.04733f
C18338 VPWR.t49 VGND 0.01447f
C18339 VPWR.t1787 VGND 0.01447f
C18340 VPWR.n1358 VGND 0.03162f
C18341 VPWR.t1317 VGND 0.01447f
C18342 VPWR.t7 VGND 0.01447f
C18343 VPWR.n1359 VGND 0.03162f
C18344 VPWR.n1360 VGND 0.06442f
C18345 VPWR.t1004 VGND 0.0577f
C18346 VPWR.t1699 VGND 0.0577f
C18347 VPWR.n1361 VGND 0.13299f
C18348 VPWR.n1362 VGND 0.02778f
C18349 VPWR.n1363 VGND 0.04733f
C18350 VPWR.n1364 VGND 0.01221f
C18351 VPWR.t1670 VGND 0.01447f
C18352 VPWR.t5 VGND 0.01447f
C18353 VPWR.n1365 VGND 0.03162f
C18354 VPWR.t11 VGND 0.01447f
C18355 VPWR.t159 VGND 0.01447f
C18356 VPWR.n1366 VGND 0.03162f
C18357 VPWR.n1367 VGND 0.0728f
C18358 VPWR.n1368 VGND 0.01221f
C18359 VPWR.n1369 VGND 0.04733f
C18360 VPWR.n1370 VGND 0.04733f
C18361 VPWR.n1371 VGND 0.04733f
C18362 VPWR.n1372 VGND 0.01139f
C18363 VPWR.t50 VGND 0.01447f
C18364 VPWR.t48 VGND 0.01447f
C18365 VPWR.n1373 VGND 0.03162f
C18366 VPWR.t1320 VGND 0.01447f
C18367 VPWR.t1319 VGND 0.01447f
C18368 VPWR.n1374 VGND 0.03162f
C18369 VPWR.n1375 VGND 0.06442f
C18370 VPWR.n1376 VGND 0.01066f
C18371 VPWR.n1377 VGND 0.00993f
C18372 VPWR.n1378 VGND 0.04733f
C18373 VPWR.n1379 VGND 0.0355f
C18374 VPWR.n1380 VGND 0.00802f
C18375 VPWR.t4 VGND 0.75581f
C18376 VPWR.n1381 VGND 0.43242f
C18377 VPWR.t6 VGND 0.75581f
C18378 VPWR.n1382 VGND 0.33884f
C18379 VPWR.n1383 VGND 0.28407f
C18380 VPWR.n1384 VGND 0.43427f
C18381 VPWR.n1385 VGND 6.23731f
C18382 VPWR.n1386 VGND 9.66078f
C18383 VPWR.n1387 VGND 1.11067f
C18384 VPWR.n1388 VGND 1.01936f
C18385 VPWR.n1389 VGND 0.05494f
C18386 VPWR.n1390 VGND 0.06546f
C18387 VPWR.t2066 VGND 0.01176f
C18388 VPWR.t822 VGND 0.01238f
C18389 VPWR.n1391 VGND 0.03075f
C18390 VPWR.n1392 VGND 0.01916f
C18391 VPWR.n1393 VGND 0.06224f
C18392 VPWR.n1394 VGND 0.07839f
C18393 VPWR.n1395 VGND 0.09265f
C18394 VPWR.t1972 VGND 0.01176f
C18395 VPWR.t691 VGND 0.01238f
C18396 VPWR.n1396 VGND 0.03075f
C18397 VPWR.n1397 VGND 0.01916f
C18398 VPWR.n1398 VGND 0.06224f
C18399 VPWR.n1399 VGND 0.09842f
C18400 VPWR.n1400 VGND 0.06632f
C18401 VPWR.n1401 VGND 0.06632f
C18402 VPWR.n1402 VGND 0.06632f
C18403 VPWR.n1403 VGND 0.06632f
C18404 VPWR.n1404 VGND 0.06632f
C18405 VPWR.n1405 VGND 0.06632f
C18406 VPWR.n1406 VGND 0.06632f
C18407 VPWR.n1407 VGND 0.05494f
C18408 VPWR.n1408 VGND -0.01884f
C18409 VPWR.t1990 VGND 0.01176f
C18410 VPWR.t640 VGND 0.01238f
C18411 VPWR.n1409 VGND 0.03f
C18412 VPWR.n1410 VGND 0.01873f
C18413 VPWR.t642 VGND 0.02986f
C18414 VPWR.n1411 VGND 0.0649f
C18415 VPWR.t299 VGND 0.0299f
C18416 VPWR.n1412 VGND 0.04757f
C18417 VPWR.t298 VGND 0.09401f
C18418 VPWR.t892 VGND 0.08295f
C18419 VPWR.t897 VGND 0.11982f
C18420 VPWR.t1938 VGND 0.01176f
C18421 VPWR.t770 VGND 0.01238f
C18422 VPWR.n1413 VGND 0.03f
C18423 VPWR.n1414 VGND 0.01873f
C18424 VPWR.t772 VGND 0.02986f
C18425 VPWR.n1415 VGND 0.0649f
C18426 VPWR.t79 VGND 0.0299f
C18427 VPWR.n1416 VGND 0.04757f
C18428 VPWR.t2038 VGND 0.01176f
C18429 VPWR.t885 VGND 0.01238f
C18430 VPWR.n1417 VGND 0.03f
C18431 VPWR.n1418 VGND 0.01873f
C18432 VPWR.t887 VGND 0.02986f
C18433 VPWR.n1419 VGND 0.0649f
C18434 VPWR.t1906 VGND 0.0299f
C18435 VPWR.n1420 VGND 0.04757f
C18436 VPWR.t507 VGND 0.09401f
C18437 VPWR.t2047 VGND 0.01176f
C18438 VPWR.t864 VGND 0.01238f
C18439 VPWR.n1421 VGND 0.03f
C18440 VPWR.n1422 VGND 0.01873f
C18441 VPWR.t866 VGND 0.02986f
C18442 VPWR.n1423 VGND 0.0649f
C18443 VPWR.t508 VGND 0.0299f
C18444 VPWR.n1424 VGND 0.04757f
C18445 VPWR.t1946 VGND 0.01176f
C18446 VPWR.t751 VGND 0.01238f
C18447 VPWR.n1425 VGND 0.03f
C18448 VPWR.n1426 VGND 0.01873f
C18449 VPWR.t753 VGND 0.02986f
C18450 VPWR.n1427 VGND 0.0649f
C18451 VPWR.t1625 VGND 0.0299f
C18452 VPWR.n1428 VGND 0.04757f
C18453 VPWR.t216 VGND 0.09401f
C18454 VPWR.t2004 VGND 0.01176f
C18455 VPWR.t609 VGND 0.01238f
C18456 VPWR.n1429 VGND 0.03f
C18457 VPWR.n1430 VGND 0.01873f
C18458 VPWR.t611 VGND 0.02986f
C18459 VPWR.n1431 VGND 0.0649f
C18460 VPWR.t217 VGND 0.0299f
C18461 VPWR.n1432 VGND 0.04757f
C18462 VPWR.t2005 VGND 0.01176f
C18463 VPWR.t966 VGND 0.01238f
C18464 VPWR.n1433 VGND 0.03f
C18465 VPWR.n1434 VGND 0.01873f
C18466 VPWR.t968 VGND 0.02986f
C18467 VPWR.n1435 VGND 0.0649f
C18468 VPWR.t608 VGND 0.0299f
C18469 VPWR.n1436 VGND 0.04757f
C18470 VPWR.t138 VGND 0.09401f
C18471 VPWR.t1951 VGND 0.01176f
C18472 VPWR.t746 VGND 0.01238f
C18473 VPWR.n1437 VGND 0.03f
C18474 VPWR.n1438 VGND 0.01873f
C18475 VPWR.t748 VGND 0.02986f
C18476 VPWR.n1439 VGND 0.0649f
C18477 VPWR.t139 VGND 0.0299f
C18478 VPWR.n1440 VGND 0.04757f
C18479 VPWR.t1962 VGND 0.01176f
C18480 VPWR.t706 VGND 0.01238f
C18481 VPWR.n1441 VGND 0.03f
C18482 VPWR.n1442 VGND 0.01873f
C18483 VPWR.t708 VGND 0.02986f
C18484 VPWR.n1443 VGND 0.0649f
C18485 VPWR.t45 VGND 0.0299f
C18486 VPWR.n1444 VGND 0.04757f
C18487 VPWR.t825 VGND 0.14747f
C18488 VPWR.t823 VGND 0.08295f
C18489 VPWR.t1848 VGND 0.09401f
C18490 VPWR.t2065 VGND 0.01176f
C18491 VPWR.t824 VGND 0.01238f
C18492 VPWR.n1445 VGND 0.03f
C18493 VPWR.n1446 VGND 0.01873f
C18494 VPWR.t826 VGND 0.02986f
C18495 VPWR.n1447 VGND 0.0649f
C18496 VPWR.t1849 VGND 0.0299f
C18497 VPWR.n1448 VGND 0.04757f
C18498 VPWR.n1449 VGND 0.01815f
C18499 VPWR.n1450 VGND -0.00319f
C18500 VPWR.n1451 VGND 0.09471f
C18501 VPWR.t613 VGND 0.11982f
C18502 VPWR.t692 VGND 0.08295f
C18503 VPWR.t1538 VGND 0.09401f
C18504 VPWR.t2003 VGND 0.01176f
C18505 VPWR.t612 VGND 0.01238f
C18506 VPWR.n1452 VGND 0.03f
C18507 VPWR.n1453 VGND 0.01873f
C18508 VPWR.t614 VGND 0.02986f
C18509 VPWR.n1454 VGND 0.0649f
C18510 VPWR.t1539 VGND 0.0299f
C18511 VPWR.n1455 VGND 0.04757f
C18512 VPWR.n1456 VGND -0.00319f
C18513 VPWR.n1457 VGND 0.09471f
C18514 VPWR.t707 VGND 0.11982f
C18515 VPWR.t705 VGND 0.08295f
C18516 VPWR.t44 VGND 0.09401f
C18517 VPWR.t745 VGND 0.08295f
C18518 VPWR.t747 VGND 0.11982f
C18519 VPWR.n1458 VGND 0.09471f
C18520 VPWR.n1459 VGND -0.00319f
C18521 VPWR.n1460 VGND 0.01815f
C18522 VPWR.n1461 VGND 0.14051f
C18523 VPWR.n1462 VGND -0.01884f
C18524 VPWR.n1463 VGND 0.08433f
C18525 VPWR.n1464 VGND 0.08433f
C18526 VPWR.n1465 VGND -0.01884f
C18527 VPWR.n1466 VGND 0.05494f
C18528 VPWR.n1467 VGND 0.14051f
C18529 VPWR.n1468 VGND 0.01815f
C18530 VPWR.n1469 VGND -0.00319f
C18531 VPWR.n1470 VGND 0.09471f
C18532 VPWR.t967 VGND 0.11982f
C18533 VPWR.t965 VGND 0.08295f
C18534 VPWR.t607 VGND 0.09401f
C18535 VPWR.t624 VGND 0.08295f
C18536 VPWR.t610 VGND 0.11982f
C18537 VPWR.n1471 VGND 0.09471f
C18538 VPWR.n1472 VGND -0.00319f
C18539 VPWR.n1473 VGND 0.01815f
C18540 VPWR.n1474 VGND 0.05494f
C18541 VPWR.n1475 VGND 0.14051f
C18542 VPWR.n1476 VGND -0.01884f
C18543 VPWR.n1477 VGND 0.08433f
C18544 VPWR.n1478 VGND 0.08433f
C18545 VPWR.n1479 VGND -0.01884f
C18546 VPWR.n1480 VGND 0.05494f
C18547 VPWR.n1481 VGND 0.14051f
C18548 VPWR.n1482 VGND 0.01815f
C18549 VPWR.n1483 VGND -0.00319f
C18550 VPWR.n1484 VGND 0.09471f
C18551 VPWR.t752 VGND 0.11982f
C18552 VPWR.t750 VGND 0.08295f
C18553 VPWR.t1624 VGND 0.09401f
C18554 VPWR.t863 VGND 0.08295f
C18555 VPWR.t865 VGND 0.11982f
C18556 VPWR.n1485 VGND 0.09471f
C18557 VPWR.n1486 VGND -0.00319f
C18558 VPWR.n1487 VGND 0.01815f
C18559 VPWR.n1488 VGND 0.05494f
C18560 VPWR.n1489 VGND 0.14051f
C18561 VPWR.n1490 VGND -0.01884f
C18562 VPWR.n1491 VGND 0.08433f
C18563 VPWR.n1492 VGND 0.08433f
C18564 VPWR.n1493 VGND -0.01884f
C18565 VPWR.n1494 VGND 0.05494f
C18566 VPWR.n1495 VGND 0.14051f
C18567 VPWR.n1496 VGND 0.01815f
C18568 VPWR.n1497 VGND -0.00319f
C18569 VPWR.n1498 VGND 0.09471f
C18570 VPWR.t886 VGND 0.11982f
C18571 VPWR.t884 VGND 0.08295f
C18572 VPWR.t1905 VGND 0.09401f
C18573 VPWR.t639 VGND 0.08295f
C18574 VPWR.t641 VGND 0.11982f
C18575 VPWR.n1499 VGND 0.09471f
C18576 VPWR.n1500 VGND -0.00319f
C18577 VPWR.n1501 VGND 0.01815f
C18578 VPWR.n1502 VGND 0.05494f
C18579 VPWR.n1503 VGND 0.14051f
C18580 VPWR.n1504 VGND -0.01884f
C18581 VPWR.n1505 VGND 0.08433f
C18582 VPWR.n1506 VGND 0.08433f
C18583 VPWR.n1507 VGND 0.08433f
C18584 VPWR.n1508 VGND 0.08433f
C18585 VPWR.n1509 VGND -0.01884f
C18586 VPWR.n1510 VGND 0.14051f
C18587 VPWR.n1511 VGND 0.01815f
C18588 VPWR.n1512 VGND -0.00319f
C18589 VPWR.n1513 VGND 0.09471f
C18590 VPWR.t78 VGND 0.09401f
C18591 VPWR.t769 VGND 0.08295f
C18592 VPWR.t771 VGND 0.11982f
C18593 VPWR.n1514 VGND 0.09471f
C18594 VPWR.n1515 VGND -0.00319f
C18595 VPWR.n1516 VGND 0.01815f
C18596 VPWR.n1517 VGND 0.14051f
C18597 VPWR.n1518 VGND 0.05494f
C18598 VPWR.n1519 VGND 0.06632f
C18599 VPWR.n1520 VGND 0.09265f
C18600 VPWR.t1940 VGND 0.01176f
C18601 VPWR.t768 VGND 0.01238f
C18602 VPWR.n1521 VGND 0.03075f
C18603 VPWR.n1522 VGND 0.01916f
C18604 VPWR.n1523 VGND 0.06224f
C18605 VPWR.n1524 VGND 0.09842f
C18606 VPWR.n1525 VGND 0.09265f
C18607 VPWR.t1991 VGND 0.01176f
C18608 VPWR.t638 VGND 0.01238f
C18609 VPWR.n1526 VGND 0.03075f
C18610 VPWR.n1527 VGND 0.01916f
C18611 VPWR.n1528 VGND 0.06224f
C18612 VPWR.n1529 VGND 0.09842f
C18613 VPWR.n1530 VGND 0.09265f
C18614 VPWR.t2039 VGND 0.01176f
C18615 VPWR.t883 VGND 0.01238f
C18616 VPWR.n1531 VGND 0.03075f
C18617 VPWR.n1532 VGND 0.01916f
C18618 VPWR.n1533 VGND 0.06224f
C18619 VPWR.n1534 VGND 0.09842f
C18620 VPWR.n1535 VGND 0.09265f
C18621 VPWR.t2049 VGND 0.01176f
C18622 VPWR.t862 VGND 0.01238f
C18623 VPWR.n1536 VGND 0.03075f
C18624 VPWR.n1537 VGND 0.01916f
C18625 VPWR.n1538 VGND 0.06224f
C18626 VPWR.n1539 VGND 0.09842f
C18627 VPWR.n1540 VGND 0.09265f
C18628 VPWR.t1948 VGND 0.01176f
C18629 VPWR.t749 VGND 0.01238f
C18630 VPWR.n1541 VGND 0.03075f
C18631 VPWR.n1542 VGND 0.01916f
C18632 VPWR.n1543 VGND 0.06224f
C18633 VPWR.n1544 VGND 0.09842f
C18634 VPWR.n1545 VGND 0.09265f
C18635 VPWR.t1998 VGND 0.01176f
C18636 VPWR.t623 VGND 0.01238f
C18637 VPWR.n1546 VGND 0.03075f
C18638 VPWR.n1547 VGND 0.01916f
C18639 VPWR.n1548 VGND 0.06224f
C18640 VPWR.n1549 VGND 0.09842f
C18641 VPWR.n1550 VGND 0.09265f
C18642 VPWR.t2006 VGND 0.01176f
C18643 VPWR.t964 VGND 0.01238f
C18644 VPWR.n1551 VGND 0.03075f
C18645 VPWR.n1552 VGND 0.01916f
C18646 VPWR.n1553 VGND 0.06224f
C18647 VPWR.n1554 VGND 0.09842f
C18648 VPWR.n1555 VGND 0.09265f
C18649 VPWR.t1952 VGND 0.01176f
C18650 VPWR.t744 VGND 0.01238f
C18651 VPWR.n1556 VGND 0.03075f
C18652 VPWR.n1557 VGND 0.01916f
C18653 VPWR.n1558 VGND 0.06224f
C18654 VPWR.n1559 VGND 0.09842f
C18655 VPWR.n1560 VGND 0.09265f
C18656 VPWR.t1964 VGND 0.01176f
C18657 VPWR.t704 VGND 0.01238f
C18658 VPWR.n1561 VGND 0.03075f
C18659 VPWR.n1562 VGND 0.01916f
C18660 VPWR.n1563 VGND 0.06224f
C18661 VPWR.n1564 VGND 0.09842f
C18662 VPWR.n1565 VGND 0.09265f
C18663 VPWR.n1566 VGND 0.06632f
C18664 VPWR.n1567 VGND 0.05494f
C18665 VPWR.n1568 VGND 0.14051f
C18666 VPWR.n1569 VGND -0.01884f
C18667 VPWR.n1570 VGND 0.08433f
C18668 VPWR.n1571 VGND 0.08433f
C18669 VPWR.n1572 VGND -0.01884f
C18670 VPWR.n1573 VGND 0.02426f
C18671 VPWR.n1574 VGND 0.0313f
C18672 VPWR.t1963 VGND 0.01176f
C18673 VPWR.t800 VGND 0.01238f
C18674 VPWR.n1575 VGND 0.03074f
C18675 VPWR.n1576 VGND 0.04185f
C18676 VPWR.n1577 VGND 0.02485f
C18677 VPWR.t1931 VGND 0.01176f
C18678 VPWR.t893 VGND 0.01238f
C18679 VPWR.n1578 VGND 0.03074f
C18680 VPWR.n1579 VGND 0.02885f
C18681 VPWR.n1580 VGND 0.0313f
C18682 VPWR.t2067 VGND 0.01176f
C18683 VPWR.t917 VGND 0.01238f
C18684 VPWR.n1581 VGND 0.03074f
C18685 VPWR.n1582 VGND 0.04185f
C18686 VPWR.n1583 VGND 0.02485f
C18687 VPWR.t2069 VGND 0.01176f
C18688 VPWR.t909 VGND 0.01238f
C18689 VPWR.n1584 VGND 0.03074f
C18690 VPWR.n1585 VGND 0.02885f
C18691 VPWR.n1586 VGND 0.0313f
C18692 VPWR.t2055 VGND 0.01176f
C18693 VPWR.t953 VGND 0.01238f
C18694 VPWR.n1587 VGND 0.03074f
C18695 VPWR.n1588 VGND 0.04185f
C18696 VPWR.n1589 VGND 0.02485f
C18697 VPWR.t2057 VGND 0.01176f
C18698 VPWR.t948 VGND 0.01238f
C18699 VPWR.n1590 VGND 0.03074f
C18700 VPWR.n1591 VGND 0.02885f
C18701 VPWR.n1592 VGND 0.0313f
C18702 VPWR.t1971 VGND 0.01176f
C18703 VPWR.t789 VGND 0.01238f
C18704 VPWR.n1593 VGND 0.03074f
C18705 VPWR.n1594 VGND 0.04185f
C18706 VPWR.n1595 VGND 0.02485f
C18707 VPWR.t1974 VGND 0.01176f
C18708 VPWR.t784 VGND 0.01238f
C18709 VPWR.n1596 VGND 0.03074f
C18710 VPWR.n1597 VGND 0.02885f
C18711 VPWR.n1598 VGND 0.0313f
C18712 VPWR.t1965 VGND 0.01176f
C18713 VPWR.t797 VGND 0.01238f
C18714 VPWR.n1599 VGND 0.03074f
C18715 VPWR.n1600 VGND 0.04185f
C18716 VPWR.n1601 VGND 0.02485f
C18717 VPWR.t1958 VGND 0.01176f
C18718 VPWR.t814 VGND 0.01238f
C18719 VPWR.n1602 VGND 0.03074f
C18720 VPWR.n1603 VGND 0.02885f
C18721 VPWR.n1604 VGND 0.0313f
C18722 VPWR.t2048 VGND 0.01176f
C18723 VPWR.t961 VGND 0.01238f
C18724 VPWR.n1605 VGND 0.03074f
C18725 VPWR.n1606 VGND 0.04185f
C18726 VPWR.n1607 VGND 0.02485f
C18727 VPWR.t2051 VGND 0.01176f
C18728 VPWR.t956 VGND 0.01238f
C18729 VPWR.n1608 VGND 0.03074f
C18730 VPWR.n1609 VGND 0.02885f
C18731 VPWR.n1610 VGND 0.0313f
C18732 VPWR.t2007 VGND 0.01176f
C18733 VPWR.t680 VGND 0.01238f
C18734 VPWR.n1611 VGND 0.03074f
C18735 VPWR.n1612 VGND 0.04185f
C18736 VPWR.n1613 VGND 0.02485f
C18737 VPWR.t2002 VGND 0.01176f
C18738 VPWR.t701 VGND 0.01238f
C18739 VPWR.n1614 VGND 0.03074f
C18740 VPWR.n1615 VGND 0.02885f
C18741 VPWR.n1616 VGND 0.0313f
C18742 VPWR.t1999 VGND 0.01176f
C18743 VPWR.t722 VGND 0.01238f
C18744 VPWR.n1617 VGND 0.03074f
C18745 VPWR.n1618 VGND 0.04185f
C18746 VPWR.n1619 VGND 0.02485f
C18747 VPWR.t2001 VGND 0.01176f
C18748 VPWR.t717 VGND 0.01238f
C18749 VPWR.n1620 VGND 0.03074f
C18750 VPWR.n1621 VGND 0.02885f
C18751 VPWR.n1622 VGND 0.0313f
C18752 VPWR.t1947 VGND 0.01176f
C18753 VPWR.t854 VGND 0.01238f
C18754 VPWR.n1623 VGND 0.03074f
C18755 VPWR.n1624 VGND 0.04185f
C18756 VPWR.n1625 VGND 0.02485f
C18757 VPWR.t2058 VGND 0.01176f
C18758 VPWR.t934 VGND 0.01238f
C18759 VPWR.n1626 VGND 0.03074f
C18760 VPWR.n1627 VGND 0.02885f
C18761 VPWR.n1628 VGND 0.0313f
C18762 VPWR.t2043 VGND 0.01176f
C18763 VPWR.t990 VGND 0.01238f
C18764 VPWR.n1629 VGND 0.03074f
C18765 VPWR.n1630 VGND 0.04185f
C18766 VPWR.n1631 VGND 0.02485f
C18767 VPWR.t2046 VGND 0.01176f
C18768 VPWR.t982 VGND 0.01238f
C18769 VPWR.n1632 VGND 0.03074f
C18770 VPWR.n1633 VGND 0.02885f
C18771 VPWR.n1634 VGND 0.0313f
C18772 VPWR.t1992 VGND 0.01176f
C18773 VPWR.t730 VGND 0.01238f
C18774 VPWR.n1635 VGND 0.03074f
C18775 VPWR.n1636 VGND 0.04185f
C18776 VPWR.n1637 VGND 0.02485f
C18777 VPWR.t1994 VGND 0.01176f
C18778 VPWR.t725 VGND 0.01238f
C18779 VPWR.n1638 VGND 0.03074f
C18780 VPWR.n1639 VGND 0.02885f
C18781 VPWR.n1640 VGND 0.0313f
C18782 VPWR.t1981 VGND 0.01176f
C18783 VPWR.t762 VGND 0.01238f
C18784 VPWR.n1641 VGND 0.03074f
C18785 VPWR.n1642 VGND 0.04185f
C18786 VPWR.n1643 VGND 0.02485f
C18787 VPWR.t1945 VGND 0.01176f
C18788 VPWR.t857 VGND 0.01238f
C18789 VPWR.n1644 VGND 0.03074f
C18790 VPWR.n1645 VGND 0.02885f
C18791 VPWR.n1646 VGND 0.0313f
C18792 VPWR.t1939 VGND 0.01176f
C18793 VPWR.t877 VGND 0.01238f
C18794 VPWR.n1647 VGND 0.03074f
C18795 VPWR.n1648 VGND 0.04185f
C18796 VPWR.n1649 VGND 0.02485f
C18797 VPWR.t1942 VGND 0.01176f
C18798 VPWR.t875 VGND 0.01238f
C18799 VPWR.n1650 VGND 0.03074f
C18800 VPWR.n1651 VGND 0.02256f
C18801 VPWR.n1652 VGND 0.01916f
C18802 VPWR.n1653 VGND 0.03332f
C18803 VPWR.n1654 VGND 0.17759f
C18804 VPWR.t2032 VGND 0.01176f
C18805 VPWR.t625 VGND 0.01238f
C18806 VPWR.n1655 VGND 0.03074f
C18807 VPWR.n1656 VGND 0.02885f
C18808 VPWR.t2028 VGND 0.01176f
C18809 VPWR.t630 VGND 0.01238f
C18810 VPWR.n1657 VGND 0.03074f
C18811 VPWR.n1658 VGND 0.04185f
C18812 VPWR.n1659 VGND 0.02485f
C18813 VPWR.t2030 VGND 0.01176f
C18814 VPWR.t628 VGND 0.01238f
C18815 VPWR.n1660 VGND 0.03074f
C18816 VPWR.n1661 VGND 0.02256f
C18817 VPWR.n1662 VGND 0.01916f
C18818 VPWR.n1663 VGND 0.03332f
C18819 VPWR.n1664 VGND 0.21371f
C18820 VPWR.n1665 VGND 0.03491f
C18821 VPWR.t1988 VGND 0.01176f
C18822 VPWR.t739 VGND 0.01238f
C18823 VPWR.n1666 VGND 0.03074f
C18824 VPWR.n1667 VGND 0.02256f
C18825 VPWR.n1668 VGND 0.02485f
C18826 VPWR.t1986 VGND 0.01176f
C18827 VPWR.t741 VGND 0.01238f
C18828 VPWR.n1669 VGND 0.03074f
C18829 VPWR.n1670 VGND 0.04185f
C18830 VPWR.n1671 VGND 0.0313f
C18831 VPWR.n1672 VGND 0.02426f
C18832 VPWR.n1673 VGND 0.00608f
C18833 VPWR.n1674 VGND -0.00323f
C18834 VPWR.n1675 VGND 0.09471f
C18835 VPWR.t626 VGND 0.09401f
C18836 VPWR.t629 VGND 0.08295f
C18837 VPWR.t631 VGND 0.11982f
C18838 VPWR.n1676 VGND 0.09471f
C18839 VPWR.n1677 VGND -0.00323f
C18840 VPWR.n1678 VGND 0.00608f
C18841 VPWR.n1679 VGND 0.02426f
C18842 VPWR.n1680 VGND 0.05494f
C18843 VPWR.t1980 VGND 0.01176f
C18844 VPWR.t666 VGND 0.01238f
C18845 VPWR.n1681 VGND 0.03f
C18846 VPWR.n1682 VGND 0.01873f
C18847 VPWR.t668 VGND 0.02986f
C18848 VPWR.n1683 VGND 0.0649f
C18849 VPWR.t1073 VGND 0.0299f
C18850 VPWR.n1684 VGND 0.04757f
C18851 VPWR.t662 VGND 0.08295f
C18852 VPWR.t1072 VGND 0.09401f
C18853 VPWR.t807 VGND 0.08295f
C18854 VPWR.t809 VGND 0.11982f
C18855 VPWR.n1685 VGND 0.09471f
C18856 VPWR.n1686 VGND -0.00319f
C18857 VPWR.n1687 VGND 0.01815f
C18858 VPWR.n1688 VGND 0.14051f
C18859 VPWR.n1689 VGND -0.01884f
C18860 VPWR.n1690 VGND 0.08433f
C18861 VPWR.n1691 VGND 0.08433f
C18862 VPWR.n1692 VGND -0.01884f
C18863 VPWR.n1693 VGND 0.14051f
C18864 VPWR.n1694 VGND 0.01815f
C18865 VPWR.n1695 VGND -0.00319f
C18866 VPWR.n1696 VGND 0.09471f
C18867 VPWR.t174 VGND 0.09401f
C18868 VPWR.t644 VGND 0.08295f
C18869 VPWR.t889 VGND 0.11982f
C18870 VPWR.n1697 VGND 0.09471f
C18871 VPWR.n1698 VGND -0.00319f
C18872 VPWR.n1699 VGND 0.01815f
C18873 VPWR.n1700 VGND 0.14051f
C18874 VPWR.n1701 VGND 0.05494f
C18875 VPWR.n1702 VGND 0.06632f
C18876 VPWR.n1703 VGND 0.09265f
C18877 VPWR.t1987 VGND 0.01176f
C18878 VPWR.t643 VGND 0.01238f
C18879 VPWR.n1704 VGND 0.03075f
C18880 VPWR.n1705 VGND 0.01916f
C18881 VPWR.n1706 VGND 0.06224f
C18882 VPWR.n1707 VGND 0.09842f
C18883 VPWR.n1708 VGND 0.09265f
C18884 VPWR.t1982 VGND 0.01176f
C18885 VPWR.t661 VGND 0.01238f
C18886 VPWR.n1709 VGND 0.03075f
C18887 VPWR.n1710 VGND 0.01916f
C18888 VPWR.n1711 VGND 0.06224f
C18889 VPWR.n1712 VGND 0.09842f
C18890 VPWR.t2029 VGND 0.01176f
C18891 VPWR.t920 VGND 0.01238f
C18892 VPWR.n1713 VGND 0.03075f
C18893 VPWR.n1714 VGND 0.01916f
C18894 VPWR.n1715 VGND 0.06223f
C18895 VPWR.n1716 VGND 0.05189f
C18896 VPWR.t1929 VGND 0.01176f
C18897 VPWR.t806 VGND 0.01238f
C18898 VPWR.n1717 VGND 0.03075f
C18899 VPWR.n1718 VGND 0.01916f
C18900 VPWR.n1719 VGND 0.06224f
C18901 VPWR.n1720 VGND 0.09842f
C18902 VPWR.n1721 VGND 0.09265f
C18903 VPWR.n1722 VGND 0.06632f
C18904 VPWR.n1723 VGND 0.05494f
C18905 VPWR.n1724 VGND 0.14051f
C18906 VPWR.n1725 VGND 0.01815f
C18907 VPWR.n1726 VGND -0.00319f
C18908 VPWR.n1727 VGND 0.09471f
C18909 VPWR.t923 VGND 0.11982f
C18910 VPWR.t921 VGND 0.08295f
C18911 VPWR.t915 VGND 0.14528f
C18912 VPWR.n1728 VGND 0.08265f
C18913 VPWR.n1729 VGND 0.01815f
C18914 VPWR.n1730 VGND 0.14051f
C18915 VPWR.n1731 VGND 0.16623f
C18916 VPWR.n1732 VGND 1.02579f
C18917 VPWR.n1733 VGND 0.08433f
C18918 VPWR.n1734 VGND 0.08433f
C18919 VPWR.n1735 VGND 0.08433f
C18920 VPWR.n1736 VGND 0.08433f
C18921 VPWR.n1737 VGND 0.08433f
C18922 VPWR.n1738 VGND 0.08433f
C18923 VPWR.n1739 VGND 0.08433f
C18924 VPWR.n1740 VGND 0.08433f
C18925 VPWR.n1741 VGND 0.08433f
C18926 VPWR.n1742 VGND 0.08433f
C18927 VPWR.n1743 VGND 0.08433f
C18928 VPWR.n1744 VGND 0.08433f
C18929 VPWR.n1745 VGND 0.08433f
C18930 VPWR.n1746 VGND 0.08433f
C18931 VPWR.n1747 VGND 0.08433f
C18932 VPWR.n1748 VGND 0.19562f
C18933 VPWR.n1749 VGND 1.02579f
C18934 VPWR.n1750 VGND 1.02579f
C18935 VPWR.n1751 VGND 0.19562f
C18936 VPWR.n1752 VGND 0.14051f
C18937 VPWR.n1753 VGND 0.01815f
C18938 VPWR.n1754 VGND 0.08265f
C18939 VPWR.t946 VGND 0.14528f
C18940 VPWR.t409 VGND 0.08295f
C18941 VPWR.t455 VGND 0.11982f
C18942 VPWR.n1755 VGND 0.09471f
C18943 VPWR.n1756 VGND -0.00319f
C18944 VPWR.n1757 VGND 0.01815f
C18945 VPWR.n1758 VGND 0.14051f
C18946 VPWR.n1759 VGND 0.08433f
C18947 VPWR.n1760 VGND 0.08433f
C18948 VPWR.n1761 VGND 0.14051f
C18949 VPWR.n1762 VGND 0.01815f
C18950 VPWR.n1763 VGND -0.00319f
C18951 VPWR.n1764 VGND 0.09471f
C18952 VPWR.t1470 VGND 0.09401f
C18953 VPWR.t1567 VGND 0.08295f
C18954 VPWR.t1120 VGND 0.11982f
C18955 VPWR.n1765 VGND 0.09471f
C18956 VPWR.n1766 VGND -0.00319f
C18957 VPWR.n1767 VGND 0.01815f
C18958 VPWR.n1768 VGND 0.14051f
C18959 VPWR.n1769 VGND 0.08433f
C18960 VPWR.n1770 VGND 0.08433f
C18961 VPWR.n1771 VGND 0.14051f
C18962 VPWR.n1772 VGND 0.01815f
C18963 VPWR.n1773 VGND -0.00319f
C18964 VPWR.n1774 VGND 0.09471f
C18965 VPWR.t1504 VGND 0.09401f
C18966 VPWR.t410 VGND 0.08295f
C18967 VPWR.t106 VGND 0.11982f
C18968 VPWR.n1775 VGND 0.09471f
C18969 VPWR.n1776 VGND -0.00319f
C18970 VPWR.n1777 VGND 0.01815f
C18971 VPWR.n1778 VGND 0.14051f
C18972 VPWR.n1779 VGND 0.08433f
C18973 VPWR.n1780 VGND 0.08433f
C18974 VPWR.n1781 VGND 0.14051f
C18975 VPWR.n1782 VGND 0.01815f
C18976 VPWR.n1783 VGND -0.00319f
C18977 VPWR.n1784 VGND 0.09471f
C18978 VPWR.t189 VGND 0.09401f
C18979 VPWR.t1569 VGND 0.08295f
C18980 VPWR.t240 VGND 0.11982f
C18981 VPWR.n1785 VGND 0.09471f
C18982 VPWR.n1786 VGND -0.00319f
C18983 VPWR.n1787 VGND 0.01815f
C18984 VPWR.n1788 VGND 0.14051f
C18985 VPWR.n1789 VGND 0.08433f
C18986 VPWR.n1790 VGND 0.08433f
C18987 VPWR.n1791 VGND 0.14051f
C18988 VPWR.n1792 VGND 0.01815f
C18989 VPWR.n1793 VGND -0.00319f
C18990 VPWR.n1794 VGND 0.09471f
C18991 VPWR.t501 VGND 0.09401f
C18992 VPWR.t1247 VGND 0.08295f
C18993 VPWR.t429 VGND 0.11982f
C18994 VPWR.n1795 VGND 0.09471f
C18995 VPWR.n1796 VGND -0.00319f
C18996 VPWR.n1797 VGND 0.01815f
C18997 VPWR.n1798 VGND 0.14051f
C18998 VPWR.n1799 VGND 0.08433f
C18999 VPWR.n1800 VGND 0.08433f
C19000 VPWR.n1801 VGND 0.14051f
C19001 VPWR.n1802 VGND 0.01815f
C19002 VPWR.n1803 VGND -0.00319f
C19003 VPWR.n1804 VGND 0.09471f
C19004 VPWR.t208 VGND 0.09401f
C19005 VPWR.t1570 VGND 0.08295f
C19006 VPWR.t1582 VGND 0.11982f
C19007 VPWR.n1805 VGND 0.09471f
C19008 VPWR.n1806 VGND -0.00319f
C19009 VPWR.n1807 VGND 0.01815f
C19010 VPWR.n1808 VGND 0.14051f
C19011 VPWR.n1809 VGND 0.08433f
C19012 VPWR.n1810 VGND 0.08433f
C19013 VPWR.n1811 VGND 0.14051f
C19014 VPWR.n1812 VGND 0.01815f
C19015 VPWR.n1813 VGND -0.00319f
C19016 VPWR.n1814 VGND 0.09471f
C19017 VPWR.t1293 VGND 0.09401f
C19018 VPWR.t1564 VGND 0.08295f
C19019 VPWR.t14 VGND 0.11982f
C19020 VPWR.n1815 VGND 0.09471f
C19021 VPWR.n1816 VGND -0.00319f
C19022 VPWR.n1817 VGND 0.01815f
C19023 VPWR.n1818 VGND 0.14051f
C19024 VPWR.n1819 VGND 0.08433f
C19025 VPWR.n1820 VGND 0.08433f
C19026 VPWR.n1821 VGND 0.14051f
C19027 VPWR.n1822 VGND 0.01815f
C19028 VPWR.n1823 VGND -0.00319f
C19029 VPWR.n1824 VGND 0.09471f
C19030 VPWR.t1802 VGND 0.09401f
C19031 VPWR.t1566 VGND 0.08295f
C19032 VPWR.t1035 VGND 0.11982f
C19033 VPWR.n1825 VGND 0.09471f
C19034 VPWR.n1826 VGND -0.00319f
C19035 VPWR.n1827 VGND 0.01815f
C19036 VPWR.n1828 VGND 0.14051f
C19037 VPWR.n1829 VGND 0.08433f
C19038 VPWR.n1830 VGND 1.01936f
C19039 VPWR.n1831 VGND 0.19562f
C19040 VPWR.n1832 VGND 0.08433f
C19041 VPWR.n1833 VGND 0.08433f
C19042 VPWR.n1834 VGND 0.08433f
C19043 VPWR.n1835 VGND 0.08433f
C19044 VPWR.n1836 VGND 0.08433f
C19045 VPWR.n1837 VGND 0.08433f
C19046 VPWR.n1838 VGND 0.08433f
C19047 VPWR.n1839 VGND 0.08433f
C19048 VPWR.n1840 VGND 0.08433f
C19049 VPWR.n1841 VGND 0.08433f
C19050 VPWR.n1842 VGND 0.08433f
C19051 VPWR.n1843 VGND 0.08433f
C19052 VPWR.n1844 VGND 0.08433f
C19053 VPWR.n1845 VGND 0.08433f
C19054 VPWR.n1846 VGND 0.08433f
C19055 VPWR.n1847 VGND 1.01936f
C19056 VPWR.n1848 VGND 1.01936f
C19057 VPWR.n1849 VGND 0.08433f
C19058 VPWR.n1850 VGND 0.14051f
C19059 VPWR.n1851 VGND 0.01815f
C19060 VPWR.n1852 VGND -0.00319f
C19061 VPWR.n1853 VGND 0.09471f
C19062 VPWR.t338 VGND 0.11982f
C19063 VPWR.t1298 VGND 0.08295f
C19064 VPWR.t1546 VGND 0.09401f
C19065 VPWR.t1297 VGND 0.08295f
C19066 VPWR.t1540 VGND 0.11982f
C19067 VPWR.n1854 VGND 0.09471f
C19068 VPWR.n1855 VGND -0.00319f
C19069 VPWR.n1856 VGND 0.01815f
C19070 VPWR.n1857 VGND 0.14051f
C19071 VPWR.n1858 VGND 0.08433f
C19072 VPWR.n1859 VGND 0.08433f
C19073 VPWR.n1860 VGND 0.14051f
C19074 VPWR.n1861 VGND 0.01815f
C19075 VPWR.n1862 VGND -0.00319f
C19076 VPWR.n1863 VGND 0.09471f
C19077 VPWR.t1271 VGND 0.11982f
C19078 VPWR.t1453 VGND 0.08295f
C19079 VPWR.t549 VGND 0.09401f
C19080 VPWR.t484 VGND 0.08295f
C19081 VPWR.t142 VGND 0.11982f
C19082 VPWR.n1864 VGND 0.09471f
C19083 VPWR.n1865 VGND -0.00319f
C19084 VPWR.n1866 VGND 0.01815f
C19085 VPWR.n1867 VGND 0.14051f
C19086 VPWR.n1868 VGND 0.08433f
C19087 VPWR.n1869 VGND 0.08433f
C19088 VPWR.n1870 VGND 0.14051f
C19089 VPWR.n1871 VGND 0.01815f
C19090 VPWR.n1872 VGND -0.00319f
C19091 VPWR.n1873 VGND 0.09471f
C19092 VPWR.t1594 VGND 0.11982f
C19093 VPWR.t483 VGND 0.08295f
C19094 VPWR.t1814 VGND 0.09401f
C19095 VPWR.t1452 VGND 0.08295f
C19096 VPWR.t286 VGND 0.11982f
C19097 VPWR.n1874 VGND 0.09471f
C19098 VPWR.n1875 VGND -0.00319f
C19099 VPWR.n1876 VGND 0.01815f
C19100 VPWR.n1877 VGND 0.14051f
C19101 VPWR.n1878 VGND 0.08433f
C19102 VPWR.n1879 VGND 0.08433f
C19103 VPWR.n1880 VGND 0.14051f
C19104 VPWR.n1881 VGND 0.01815f
C19105 VPWR.n1882 VGND -0.00319f
C19106 VPWR.n1883 VGND 0.09471f
C19107 VPWR.t543 VGND 0.11982f
C19108 VPWR.t572 VGND 0.08295f
C19109 VPWR.t1393 VGND 0.09401f
C19110 VPWR.t571 VGND 0.08295f
C19111 VPWR.t1387 VGND 0.11982f
C19112 VPWR.n1884 VGND 0.09471f
C19113 VPWR.n1885 VGND -0.00319f
C19114 VPWR.n1886 VGND 0.01815f
C19115 VPWR.n1887 VGND 0.14051f
C19116 VPWR.n1888 VGND 0.08433f
C19117 VPWR.n1889 VGND 0.08433f
C19118 VPWR.n1890 VGND 0.14051f
C19119 VPWR.n1891 VGND 0.01815f
C19120 VPWR.n1892 VGND -0.00319f
C19121 VPWR.n1893 VGND 0.09471f
C19122 VPWR.t1180 VGND 0.11982f
C19123 VPWR.t482 VGND 0.08295f
C19124 VPWR.t357 VGND 0.09401f
C19125 VPWR.t1451 VGND 0.08295f
C19126 VPWR.t351 VGND 0.11982f
C19127 VPWR.n1894 VGND 0.09471f
C19128 VPWR.n1895 VGND -0.00319f
C19129 VPWR.n1896 VGND 0.01815f
C19130 VPWR.n1897 VGND 0.14051f
C19131 VPWR.n1898 VGND 0.08433f
C19132 VPWR.n1899 VGND 0.08433f
C19133 VPWR.n1900 VGND 0.14051f
C19134 VPWR.n1901 VGND 0.01815f
C19135 VPWR.n1902 VGND -0.00319f
C19136 VPWR.n1903 VGND 0.09471f
C19137 VPWR.t72 VGND 0.11982f
C19138 VPWR.t570 VGND 0.08295f
C19139 VPWR.t250 VGND 0.09401f
C19140 VPWR.t481 VGND 0.08295f
C19141 VPWR.t1110 VGND 0.11982f
C19142 VPWR.n1904 VGND 0.09471f
C19143 VPWR.n1905 VGND -0.00319f
C19144 VPWR.n1906 VGND 0.01815f
C19145 VPWR.n1907 VGND 0.14051f
C19146 VPWR.n1908 VGND 0.08433f
C19147 VPWR.n1909 VGND 0.08433f
C19148 VPWR.n1910 VGND 0.14051f
C19149 VPWR.n1911 VGND 0.01815f
C19150 VPWR.n1912 VGND -0.00319f
C19151 VPWR.n1913 VGND 0.09471f
C19152 VPWR.t1413 VGND 0.11982f
C19153 VPWR.t1299 VGND 0.08295f
C19154 VPWR.t1144 VGND 0.09401f
C19155 VPWR.t1099 VGND 0.08295f
C19156 VPWR.t1482 VGND 0.11982f
C19157 VPWR.n1914 VGND 0.09471f
C19158 VPWR.n1915 VGND -0.00319f
C19159 VPWR.n1916 VGND 0.01815f
C19160 VPWR.n1917 VGND 0.14051f
C19161 VPWR.n1918 VGND 0.08433f
C19162 VPWR.n1919 VGND 0.08433f
C19163 VPWR.n1920 VGND 0.14051f
C19164 VPWR.n1921 VGND 0.01815f
C19165 VPWR.n1922 VGND -0.00319f
C19166 VPWR.n1923 VGND 0.09471f
C19167 VPWR.t1379 VGND 0.11982f
C19168 VPWR.t569 VGND 0.08295f
C19169 VPWR.t670 VGND 0.14528f
C19170 VPWR.n1924 VGND 0.08265f
C19171 VPWR.n1925 VGND 0.01815f
C19172 VPWR.n1926 VGND 0.14051f
C19173 VPWR.n1927 VGND 0.19562f
C19174 VPWR.n1928 VGND 1.02579f
C19175 VPWR.n1929 VGND 0.08433f
C19176 VPWR.n1930 VGND 0.08433f
C19177 VPWR.n1931 VGND 0.08433f
C19178 VPWR.n1932 VGND 0.08433f
C19179 VPWR.n1933 VGND 0.08433f
C19180 VPWR.n1934 VGND 0.08433f
C19181 VPWR.n1935 VGND 0.08433f
C19182 VPWR.n1936 VGND 0.08433f
C19183 VPWR.n1937 VGND 0.08433f
C19184 VPWR.n1938 VGND 0.08433f
C19185 VPWR.n1939 VGND 0.08433f
C19186 VPWR.n1940 VGND 0.08433f
C19187 VPWR.n1941 VGND 0.08433f
C19188 VPWR.n1942 VGND 0.08433f
C19189 VPWR.n1943 VGND 0.08433f
C19190 VPWR.n1944 VGND 0.19562f
C19191 VPWR.n1945 VGND 1.02579f
C19192 VPWR.n1946 VGND 1.02579f
C19193 VPWR.n1947 VGND 0.19562f
C19194 VPWR.n1948 VGND 0.14051f
C19195 VPWR.n1949 VGND 0.01815f
C19196 VPWR.n1950 VGND 0.08265f
C19197 VPWR.t734 VGND 0.14528f
C19198 VPWR.t1398 VGND 0.08295f
C19199 VPWR.t1367 VGND 0.11982f
C19200 VPWR.n1951 VGND 0.09471f
C19201 VPWR.n1952 VGND -0.00319f
C19202 VPWR.n1953 VGND 0.01815f
C19203 VPWR.n1954 VGND 0.14051f
C19204 VPWR.n1955 VGND 0.08433f
C19205 VPWR.n1956 VGND 0.08433f
C19206 VPWR.n1957 VGND 0.14051f
C19207 VPWR.n1958 VGND 0.01815f
C19208 VPWR.n1959 VGND -0.00319f
C19209 VPWR.n1960 VGND 0.09471f
C19210 VPWR.t597 VGND 0.09401f
C19211 VPWR.t306 VGND 0.08295f
C19212 VPWR.t1606 VGND 0.11982f
C19213 VPWR.n1961 VGND 0.09471f
C19214 VPWR.n1962 VGND -0.00319f
C19215 VPWR.n1963 VGND 0.01815f
C19216 VPWR.n1964 VGND 0.14051f
C19217 VPWR.n1965 VGND 0.08433f
C19218 VPWR.n1966 VGND 0.08433f
C19219 VPWR.n1967 VGND 0.14051f
C19220 VPWR.n1968 VGND 0.01815f
C19221 VPWR.n1969 VGND -0.00319f
C19222 VPWR.n1970 VGND 0.09471f
C19223 VPWR.t1616 VGND 0.09401f
C19224 VPWR.t310 VGND 0.08295f
C19225 VPWR.t74 VGND 0.11982f
C19226 VPWR.n1971 VGND 0.09471f
C19227 VPWR.n1972 VGND -0.00319f
C19228 VPWR.n1973 VGND 0.01815f
C19229 VPWR.n1974 VGND 0.14051f
C19230 VPWR.n1975 VGND 0.08433f
C19231 VPWR.n1976 VGND 0.08433f
C19232 VPWR.n1977 VGND 0.14051f
C19233 VPWR.n1978 VGND 0.01815f
C19234 VPWR.n1979 VGND -0.00319f
C19235 VPWR.n1980 VGND 0.09471f
C19236 VPWR.t344 VGND 0.09401f
C19237 VPWR.t308 VGND 0.08295f
C19238 VPWR.t1168 VGND 0.11982f
C19239 VPWR.n1981 VGND 0.09471f
C19240 VPWR.n1982 VGND -0.00319f
C19241 VPWR.n1983 VGND 0.01815f
C19242 VPWR.n1984 VGND 0.14051f
C19243 VPWR.n1985 VGND 0.08433f
C19244 VPWR.n1986 VGND 0.08433f
C19245 VPWR.n1987 VGND 0.14051f
C19246 VPWR.n1988 VGND 0.01815f
C19247 VPWR.n1989 VGND -0.00319f
C19248 VPWR.n1990 VGND 0.09471f
C19249 VPWR.t517 VGND 0.09401f
C19250 VPWR.t312 VGND 0.08295f
C19251 VPWR.t1090 VGND 0.11982f
C19252 VPWR.n1991 VGND 0.09471f
C19253 VPWR.n1992 VGND -0.00319f
C19254 VPWR.n1993 VGND 0.01815f
C19255 VPWR.n1994 VGND 0.14051f
C19256 VPWR.n1995 VGND 0.08433f
C19257 VPWR.n1996 VGND 0.08433f
C19258 VPWR.n1997 VGND 0.14051f
C19259 VPWR.n1998 VGND 0.01815f
C19260 VPWR.n1999 VGND -0.00319f
C19261 VPWR.n2000 VGND 0.09471f
C19262 VPWR.t1556 VGND 0.09401f
C19263 VPWR.t309 VGND 0.08295f
C19264 VPWR.t1695 VGND 0.11982f
C19265 VPWR.n2001 VGND 0.09471f
C19266 VPWR.n2002 VGND -0.00319f
C19267 VPWR.n2003 VGND 0.01815f
C19268 VPWR.n2004 VGND 0.14051f
C19269 VPWR.n2005 VGND 0.08433f
C19270 VPWR.n2006 VGND 0.08433f
C19271 VPWR.n2007 VGND 0.14051f
C19272 VPWR.n2008 VGND 0.01815f
C19273 VPWR.n2009 VGND -0.00319f
C19274 VPWR.n2010 VGND 0.09471f
C19275 VPWR.t1056 VGND 0.09401f
C19276 VPWR.t1789 VGND 0.08295f
C19277 VPWR.t56 VGND 0.11982f
C19278 VPWR.n2011 VGND 0.09471f
C19279 VPWR.n2012 VGND -0.00319f
C19280 VPWR.n2013 VGND 0.01815f
C19281 VPWR.n2014 VGND 0.14051f
C19282 VPWR.n2015 VGND 0.08433f
C19283 VPWR.n2016 VGND 0.08433f
C19284 VPWR.n2017 VGND 0.14051f
C19285 VPWR.n2018 VGND 0.01815f
C19286 VPWR.n2019 VGND -0.00319f
C19287 VPWR.n2020 VGND 0.09471f
C19288 VPWR.t1691 VGND 0.09401f
C19289 VPWR.t1791 VGND 0.08295f
C19290 VPWR.t1850 VGND 0.11982f
C19291 VPWR.n2021 VGND 0.09471f
C19292 VPWR.n2022 VGND -0.00319f
C19293 VPWR.n2023 VGND 0.01815f
C19294 VPWR.n2024 VGND 0.14051f
C19295 VPWR.n2025 VGND 0.08433f
C19296 VPWR.n2026 VGND 1.01936f
C19297 VPWR.n2027 VGND 0.19562f
C19298 VPWR.n2028 VGND 0.08433f
C19299 VPWR.n2029 VGND 0.08433f
C19300 VPWR.n2030 VGND 0.08433f
C19301 VPWR.n2031 VGND 0.08433f
C19302 VPWR.n2032 VGND 0.08433f
C19303 VPWR.n2033 VGND 0.08433f
C19304 VPWR.n2034 VGND 0.08433f
C19305 VPWR.n2035 VGND 0.08433f
C19306 VPWR.n2036 VGND 0.08433f
C19307 VPWR.n2037 VGND 0.08433f
C19308 VPWR.n2038 VGND 0.08433f
C19309 VPWR.n2039 VGND 0.08433f
C19310 VPWR.n2040 VGND 0.08433f
C19311 VPWR.n2041 VGND 0.08433f
C19312 VPWR.n2042 VGND 0.08433f
C19313 VPWR.n2043 VGND 1.01936f
C19314 VPWR.n2044 VGND 1.01936f
C19315 VPWR.n2045 VGND 0.08433f
C19316 VPWR.n2046 VGND 0.14051f
C19317 VPWR.n2047 VGND 0.01815f
C19318 VPWR.n2048 VGND -0.00319f
C19319 VPWR.n2049 VGND 0.09471f
C19320 VPWR.t336 VGND 0.11982f
C19321 VPWR.t1076 VGND 0.08295f
C19322 VPWR.t1544 VGND 0.09401f
C19323 VPWR.t478 VGND 0.08295f
C19324 VPWR.t1693 VGND 0.11982f
C19325 VPWR.n2050 VGND 0.09471f
C19326 VPWR.n2051 VGND -0.00319f
C19327 VPWR.n2052 VGND 0.01815f
C19328 VPWR.n2053 VGND 0.14051f
C19329 VPWR.n2054 VGND 0.08433f
C19330 VPWR.n2055 VGND 0.08433f
C19331 VPWR.n2056 VGND 0.14051f
C19332 VPWR.n2057 VGND 0.01815f
C19333 VPWR.n2058 VGND -0.00319f
C19334 VPWR.n2059 VGND 0.09471f
C19335 VPWR.t1269 VGND 0.11982f
C19336 VPWR.t477 VGND 0.08295f
C19337 VPWR.t547 VGND 0.09401f
C19338 VPWR.t1138 VGND 0.08295f
C19339 VPWR.t140 VGND 0.11982f
C19340 VPWR.n2060 VGND 0.09471f
C19341 VPWR.n2061 VGND -0.00319f
C19342 VPWR.n2062 VGND 0.01815f
C19343 VPWR.n2063 VGND 0.14051f
C19344 VPWR.n2064 VGND 0.08433f
C19345 VPWR.n2065 VGND 0.08433f
C19346 VPWR.n2066 VGND 0.14051f
C19347 VPWR.n2067 VGND 0.01815f
C19348 VPWR.n2068 VGND -0.00319f
C19349 VPWR.n2069 VGND 0.09471f
C19350 VPWR.t1592 VGND 0.11982f
C19351 VPWR.t1137 VGND 0.08295f
C19352 VPWR.t1812 VGND 0.09401f
C19353 VPWR.t476 VGND 0.08295f
C19354 VPWR.t284 VGND 0.11982f
C19355 VPWR.n2070 VGND 0.09471f
C19356 VPWR.n2071 VGND -0.00319f
C19357 VPWR.n2072 VGND 0.01815f
C19358 VPWR.n2073 VGND 0.14051f
C19359 VPWR.n2074 VGND 0.08433f
C19360 VPWR.n2075 VGND 0.08433f
C19361 VPWR.n2076 VGND 0.14051f
C19362 VPWR.n2077 VGND 0.01815f
C19363 VPWR.n2078 VGND -0.00319f
C19364 VPWR.n2079 VGND 0.09471f
C19365 VPWR.t539 VGND 0.11982f
C19366 VPWR.t530 VGND 0.08295f
C19367 VPWR.t1391 VGND 0.09401f
C19368 VPWR.t529 VGND 0.08295f
C19369 VPWR.t519 VGND 0.11982f
C19370 VPWR.n2080 VGND 0.09471f
C19371 VPWR.n2081 VGND -0.00319f
C19372 VPWR.n2082 VGND 0.01815f
C19373 VPWR.n2083 VGND 0.14051f
C19374 VPWR.n2084 VGND 0.08433f
C19375 VPWR.n2085 VGND 0.08433f
C19376 VPWR.n2086 VGND 0.14051f
C19377 VPWR.n2087 VGND 0.01815f
C19378 VPWR.n2088 VGND -0.00319f
C19379 VPWR.n2089 VGND 0.09471f
C19380 VPWR.t1178 VGND 0.11982f
C19381 VPWR.t1079 VGND 0.08295f
C19382 VPWR.t355 VGND 0.09401f
C19383 VPWR.t475 VGND 0.08295f
C19384 VPWR.t349 VGND 0.11982f
C19385 VPWR.n2090 VGND 0.09471f
C19386 VPWR.n2091 VGND -0.00319f
C19387 VPWR.n2092 VGND 0.01815f
C19388 VPWR.n2093 VGND 0.14051f
C19389 VPWR.n2094 VGND 0.08433f
C19390 VPWR.n2095 VGND 0.08433f
C19391 VPWR.n2096 VGND 0.14051f
C19392 VPWR.n2097 VGND 0.01815f
C19393 VPWR.n2098 VGND -0.00319f
C19394 VPWR.n2099 VGND 0.09471f
C19395 VPWR.t70 VGND 0.11982f
C19396 VPWR.t528 VGND 0.08295f
C19397 VPWR.t248 VGND 0.09401f
C19398 VPWR.t1078 VGND 0.08295f
C19399 VPWR.t1108 VGND 0.11982f
C19400 VPWR.n2100 VGND 0.09471f
C19401 VPWR.n2101 VGND -0.00319f
C19402 VPWR.n2102 VGND 0.01815f
C19403 VPWR.n2103 VGND 0.14051f
C19404 VPWR.n2104 VGND 0.08433f
C19405 VPWR.n2105 VGND 0.08433f
C19406 VPWR.n2106 VGND 0.14051f
C19407 VPWR.n2107 VGND 0.01815f
C19408 VPWR.n2108 VGND -0.00319f
C19409 VPWR.n2109 VGND 0.09471f
C19410 VPWR.t1411 VGND 0.11982f
C19411 VPWR.t1077 VGND 0.08295f
C19412 VPWR.t1142 VGND 0.09401f
C19413 VPWR.t184 VGND 0.08295f
C19414 VPWR.t1480 VGND 0.11982f
C19415 VPWR.n2110 VGND 0.09471f
C19416 VPWR.n2111 VGND -0.00319f
C19417 VPWR.n2112 VGND 0.01815f
C19418 VPWR.n2113 VGND 0.14051f
C19419 VPWR.n2114 VGND 0.08433f
C19420 VPWR.n2115 VGND 0.08433f
C19421 VPWR.n2116 VGND 0.14051f
C19422 VPWR.n2117 VGND 0.01815f
C19423 VPWR.n2118 VGND -0.00319f
C19424 VPWR.n2119 VGND 0.09471f
C19425 VPWR.t1375 VGND 0.11982f
C19426 VPWR.t1139 VGND 0.08295f
C19427 VPWR.t673 VGND 0.14528f
C19428 VPWR.n2120 VGND 0.08265f
C19429 VPWR.n2121 VGND 0.01815f
C19430 VPWR.n2122 VGND 0.14051f
C19431 VPWR.n2123 VGND 0.19562f
C19432 VPWR.n2124 VGND 1.02579f
C19433 VPWR.n2125 VGND 0.08433f
C19434 VPWR.n2126 VGND 0.08433f
C19435 VPWR.n2127 VGND 0.08433f
C19436 VPWR.n2128 VGND 0.08433f
C19437 VPWR.n2129 VGND 0.08433f
C19438 VPWR.n2130 VGND 0.08433f
C19439 VPWR.n2131 VGND 0.08433f
C19440 VPWR.n2132 VGND 0.08433f
C19441 VPWR.n2133 VGND 0.08433f
C19442 VPWR.n2134 VGND 0.08433f
C19443 VPWR.n2135 VGND 0.08433f
C19444 VPWR.n2136 VGND 0.08433f
C19445 VPWR.n2137 VGND 0.08433f
C19446 VPWR.n2138 VGND 0.08433f
C19447 VPWR.n2139 VGND 0.08433f
C19448 VPWR.n2140 VGND 0.19562f
C19449 VPWR.n2141 VGND 1.02579f
C19450 VPWR.n2142 VGND 1.02579f
C19451 VPWR.n2143 VGND 0.19562f
C19452 VPWR.n2144 VGND 0.14051f
C19453 VPWR.n2145 VGND 0.01815f
C19454 VPWR.n2146 VGND 0.08265f
C19455 VPWR.t820 VGND 0.14528f
C19456 VPWR.t1330 VGND 0.08295f
C19457 VPWR.t441 VGND 0.11982f
C19458 VPWR.n2147 VGND 0.09471f
C19459 VPWR.n2148 VGND -0.00319f
C19460 VPWR.n2149 VGND 0.01815f
C19461 VPWR.n2150 VGND 0.14051f
C19462 VPWR.n2151 VGND 0.08433f
C19463 VPWR.n2152 VGND 0.08433f
C19464 VPWR.n2153 VGND 0.14051f
C19465 VPWR.n2154 VGND 0.01815f
C19466 VPWR.n2155 VGND -0.00319f
C19467 VPWR.n2156 VGND 0.09471f
C19468 VPWR.t1658 VGND 0.09401f
C19469 VPWR.t1322 VGND 0.08295f
C19470 VPWR.t1612 VGND 0.11982f
C19471 VPWR.n2157 VGND 0.09471f
C19472 VPWR.n2158 VGND -0.00319f
C19473 VPWR.n2159 VGND 0.01815f
C19474 VPWR.n2160 VGND 0.14051f
C19475 VPWR.n2161 VGND 0.08433f
C19476 VPWR.n2162 VGND 0.08433f
C19477 VPWR.n2163 VGND 0.14051f
C19478 VPWR.n2164 VGND 0.01815f
C19479 VPWR.n2165 VGND -0.00319f
C19480 VPWR.n2166 VGND 0.09471f
C19481 VPWR.t1488 VGND 0.09401f
C19482 VPWR.t1331 VGND 0.08295f
C19483 VPWR.t84 VGND 0.11982f
C19484 VPWR.n2167 VGND 0.09471f
C19485 VPWR.n2168 VGND -0.00319f
C19486 VPWR.n2169 VGND 0.01815f
C19487 VPWR.n2170 VGND 0.14051f
C19488 VPWR.n2171 VGND 0.08433f
C19489 VPWR.n2172 VGND 0.08433f
C19490 VPWR.n2173 VGND 0.14051f
C19491 VPWR.n2174 VGND 0.01815f
C19492 VPWR.n2175 VGND -0.00319f
C19493 VPWR.n2176 VGND 0.09471f
C19494 VPWR.t1064 VGND 0.09401f
C19495 VPWR.t1324 VGND 0.08295f
C19496 VPWR.t1895 VGND 0.11982f
C19497 VPWR.n2177 VGND 0.09471f
C19498 VPWR.n2178 VGND -0.00319f
C19499 VPWR.n2179 VGND 0.01815f
C19500 VPWR.n2180 VGND 0.14051f
C19501 VPWR.n2181 VGND 0.08433f
C19502 VPWR.n2182 VGND 0.08433f
C19503 VPWR.n2183 VGND 0.14051f
C19504 VPWR.n2184 VGND 0.01815f
C19505 VPWR.n2185 VGND -0.00319f
C19506 VPWR.n2186 VGND 0.09471f
C19507 VPWR.t1430 VGND 0.09401f
C19508 VPWR.t1333 VGND 0.08295f
C19509 VPWR.t270 VGND 0.11982f
C19510 VPWR.n2187 VGND 0.09471f
C19511 VPWR.n2188 VGND -0.00319f
C19512 VPWR.n2189 VGND 0.01815f
C19513 VPWR.n2190 VGND 0.14051f
C19514 VPWR.n2191 VGND 0.08433f
C19515 VPWR.n2192 VGND 0.08433f
C19516 VPWR.n2193 VGND 0.14051f
C19517 VPWR.n2194 VGND 0.01815f
C19518 VPWR.n2195 VGND -0.00319f
C19519 VPWR.n2196 VGND 0.09471f
C19520 VPWR.t280 VGND 0.09401f
C19521 VPWR.t1325 VGND 0.08295f
C19522 VPWR.t1254 VGND 0.11982f
C19523 VPWR.n2197 VGND 0.09471f
C19524 VPWR.n2198 VGND -0.00319f
C19525 VPWR.n2199 VGND 0.01815f
C19526 VPWR.n2200 VGND 0.14051f
C19527 VPWR.n2201 VGND 0.08433f
C19528 VPWR.n2202 VGND 0.08433f
C19529 VPWR.n2203 VGND 0.14051f
C19530 VPWR.n2204 VGND 0.01815f
C19531 VPWR.n2205 VGND -0.00319f
C19532 VPWR.n2206 VGND 0.09471f
C19533 VPWR.t1283 VGND 0.09401f
C19534 VPWR.t378 VGND 0.08295f
C19535 VPWR.t997 VGND 0.11982f
C19536 VPWR.n2207 VGND 0.09471f
C19537 VPWR.n2208 VGND -0.00319f
C19538 VPWR.n2209 VGND 0.01815f
C19539 VPWR.n2210 VGND 0.14051f
C19540 VPWR.n2211 VGND 0.08433f
C19541 VPWR.n2212 VGND 0.08433f
C19542 VPWR.n2213 VGND 0.14051f
C19543 VPWR.n2214 VGND 0.01815f
C19544 VPWR.n2215 VGND -0.00319f
C19545 VPWR.n2216 VGND 0.09471f
C19546 VPWR.t1689 VGND 0.09401f
C19547 VPWR.t380 VGND 0.08295f
C19548 VPWR.t1019 VGND 0.11982f
C19549 VPWR.n2217 VGND 0.09471f
C19550 VPWR.n2218 VGND -0.00319f
C19551 VPWR.n2219 VGND 0.01815f
C19552 VPWR.n2220 VGND 0.14051f
C19553 VPWR.n2221 VGND 0.08433f
C19554 VPWR.n2222 VGND 1.01936f
C19555 VPWR.n2223 VGND 0.19562f
C19556 VPWR.n2224 VGND 0.08433f
C19557 VPWR.n2225 VGND 0.08433f
C19558 VPWR.n2226 VGND 0.08433f
C19559 VPWR.n2227 VGND 0.08433f
C19560 VPWR.n2228 VGND 0.08433f
C19561 VPWR.n2229 VGND 0.08433f
C19562 VPWR.n2230 VGND 0.08433f
C19563 VPWR.n2231 VGND 0.08433f
C19564 VPWR.n2232 VGND 0.08433f
C19565 VPWR.n2233 VGND 0.08433f
C19566 VPWR.n2234 VGND 0.08433f
C19567 VPWR.n2235 VGND 0.08433f
C19568 VPWR.n2236 VGND 0.08433f
C19569 VPWR.n2237 VGND 0.08433f
C19570 VPWR.n2238 VGND 0.08433f
C19571 VPWR.n2239 VGND 1.01936f
C19572 VPWR.n2240 VGND 1.01936f
C19573 VPWR.n2241 VGND 0.08433f
C19574 VPWR.n2242 VGND 0.14051f
C19575 VPWR.n2243 VGND 0.01815f
C19576 VPWR.n2244 VGND -0.00319f
C19577 VPWR.n2245 VGND 0.09471f
C19578 VPWR.t1846 VGND 0.11982f
C19579 VPWR.t1878 VGND 0.08295f
C19580 VPWR.t176 VGND 0.09401f
C19581 VPWR.t1877 VGND 0.08295f
C19582 VPWR.t1442 VGND 0.11982f
C19583 VPWR.n2246 VGND 0.09471f
C19584 VPWR.n2247 VGND -0.00319f
C19585 VPWR.n2248 VGND 0.01815f
C19586 VPWR.n2249 VGND 0.14051f
C19587 VPWR.n2250 VGND 0.08433f
C19588 VPWR.n2251 VGND 0.08433f
C19589 VPWR.n2252 VGND 0.14051f
C19590 VPWR.n2253 VGND 0.01815f
C19591 VPWR.n2254 VGND -0.00319f
C19592 VPWR.n2255 VGND 0.09471f
C19593 VPWR.t1887 VGND 0.11982f
C19594 VPWR.t224 VGND 0.08295f
C19595 VPWR.t1924 VGND 0.09401f
C19596 VPWR.t382 VGND 0.08295f
C19597 VPWR.t1464 VGND 0.11982f
C19598 VPWR.n2256 VGND 0.09471f
C19599 VPWR.n2257 VGND -0.00319f
C19600 VPWR.n2258 VGND 0.01815f
C19601 VPWR.n2259 VGND 0.14051f
C19602 VPWR.n2260 VGND 0.08433f
C19603 VPWR.n2261 VGND 0.08433f
C19604 VPWR.n2262 VGND 0.14051f
C19605 VPWR.n2263 VGND 0.01815f
C19606 VPWR.n2264 VGND -0.00319f
C19607 VPWR.n2265 VGND 0.09471f
C19608 VPWR.t1710 VGND 0.11982f
C19609 VPWR.t381 VGND 0.08295f
C19610 VPWR.t1554 VGND 0.09401f
C19611 VPWR.t223 VGND 0.08295f
C19612 VPWR.t220 VGND 0.11982f
C19613 VPWR.n2266 VGND 0.09471f
C19614 VPWR.n2267 VGND -0.00319f
C19615 VPWR.n2268 VGND 0.01815f
C19616 VPWR.n2269 VGND 0.14051f
C19617 VPWR.n2270 VGND 0.08433f
C19618 VPWR.n2271 VGND 0.08433f
C19619 VPWR.n2272 VGND 0.14051f
C19620 VPWR.n2273 VGND 0.01815f
C19621 VPWR.n2274 VGND -0.00319f
C19622 VPWR.n2275 VGND 0.09471f
C19623 VPWR.t1628 VGND 0.11982f
C19624 VPWR.t1406 VGND 0.08295f
C19625 VPWR.t513 VGND 0.09401f
C19626 VPWR.t1405 VGND 0.08295f
C19627 VPWR.t509 VGND 0.11982f
C19628 VPWR.n2276 VGND 0.09471f
C19629 VPWR.n2277 VGND -0.00319f
C19630 VPWR.n2278 VGND 0.01815f
C19631 VPWR.n2279 VGND 0.14051f
C19632 VPWR.n2280 VGND 0.08433f
C19633 VPWR.n2281 VGND 0.08433f
C19634 VPWR.n2282 VGND 0.14051f
C19635 VPWR.n2283 VGND 0.01815f
C19636 VPWR.n2284 VGND -0.00319f
C19637 VPWR.n2285 VGND 0.09471f
C19638 VPWR.t1909 VGND 0.11982f
C19639 VPWR.t398 VGND 0.08295f
C19640 VPWR.t290 VGND 0.09401f
C19641 VPWR.t222 VGND 0.08295f
C19642 VPWR.t1070 VGND 0.11982f
C19643 VPWR.n2286 VGND 0.09471f
C19644 VPWR.n2287 VGND -0.00319f
C19645 VPWR.n2288 VGND 0.01815f
C19646 VPWR.n2289 VGND 0.14051f
C19647 VPWR.n2290 VGND 0.08433f
C19648 VPWR.n2291 VGND 0.08433f
C19649 VPWR.n2292 VGND 0.14051f
C19650 VPWR.n2293 VGND 0.01815f
C19651 VPWR.n2294 VGND -0.00319f
C19652 VPWR.n2295 VGND 0.09471f
C19653 VPWR.t82 VGND 0.11982f
C19654 VPWR.t1404 VGND 0.08295f
C19655 VPWR.t1498 VGND 0.09401f
C19656 VPWR.t397 VGND 0.08295f
C19657 VPWR.t1494 VGND 0.11982f
C19658 VPWR.n2296 VGND 0.09471f
C19659 VPWR.n2297 VGND -0.00319f
C19660 VPWR.n2298 VGND 0.01815f
C19661 VPWR.n2299 VGND 0.14051f
C19662 VPWR.n2300 VGND 0.08433f
C19663 VPWR.n2301 VGND 0.08433f
C19664 VPWR.n2302 VGND 0.14051f
C19665 VPWR.n2303 VGND 0.01815f
C19666 VPWR.n2304 VGND -0.00319f
C19667 VPWR.n2305 VGND 0.09471f
C19668 VPWR.t1600 VGND 0.11982f
C19669 VPWR.t396 VGND 0.08295f
C19670 VPWR.t1082 VGND 0.09401f
C19671 VPWR.t1819 VGND 0.08295f
C19672 VPWR.t1478 VGND 0.11982f
C19673 VPWR.n2306 VGND 0.09471f
C19674 VPWR.n2307 VGND -0.00319f
C19675 VPWR.n2308 VGND 0.01815f
C19676 VPWR.n2309 VGND 0.14051f
C19677 VPWR.n2310 VGND 0.08433f
C19678 VPWR.n2311 VGND 0.08433f
C19679 VPWR.n2312 VGND 0.14051f
C19680 VPWR.n2313 VGND 0.01815f
C19681 VPWR.n2314 VGND -0.00319f
C19682 VPWR.n2315 VGND 0.09471f
C19683 VPWR.t451 VGND 0.11982f
C19684 VPWR.t383 VGND 0.08295f
C19685 VPWR.t766 VGND 0.14528f
C19686 VPWR.n2316 VGND 0.08265f
C19687 VPWR.n2317 VGND 0.01815f
C19688 VPWR.n2318 VGND 0.14051f
C19689 VPWR.n2319 VGND 0.19562f
C19690 VPWR.n2320 VGND 1.02579f
C19691 VPWR.n2321 VGND 0.08433f
C19692 VPWR.n2322 VGND 0.08433f
C19693 VPWR.n2323 VGND 0.08433f
C19694 VPWR.n2324 VGND 0.08433f
C19695 VPWR.n2325 VGND 0.08433f
C19696 VPWR.n2326 VGND 0.08433f
C19697 VPWR.n2327 VGND 0.08433f
C19698 VPWR.n2328 VGND 0.08433f
C19699 VPWR.n2329 VGND 0.08433f
C19700 VPWR.n2330 VGND 0.08433f
C19701 VPWR.n2331 VGND 0.08433f
C19702 VPWR.n2332 VGND 0.08433f
C19703 VPWR.n2333 VGND 0.08433f
C19704 VPWR.n2334 VGND 0.08433f
C19705 VPWR.n2335 VGND 0.08433f
C19706 VPWR.n2336 VGND 0.19562f
C19707 VPWR.n2337 VGND 1.02579f
C19708 VPWR.n2338 VGND 1.02579f
C19709 VPWR.n2339 VGND 0.19562f
C19710 VPWR.n2340 VGND 0.14051f
C19711 VPWR.n2341 VGND 0.01815f
C19712 VPWR.n2342 VGND 0.08265f
C19713 VPWR.t932 VGND 0.14528f
C19714 VPWR.t586 VGND 0.08295f
C19715 VPWR.t463 VGND 0.11982f
C19716 VPWR.n2343 VGND 0.09471f
C19717 VPWR.n2344 VGND -0.00319f
C19718 VPWR.n2345 VGND 0.01815f
C19719 VPWR.n2346 VGND 0.14051f
C19720 VPWR.n2347 VGND 0.08433f
C19721 VPWR.n2348 VGND 0.08433f
C19722 VPWR.n2349 VGND 0.14051f
C19723 VPWR.n2350 VGND 0.01815f
C19724 VPWR.n2351 VGND -0.00319f
C19725 VPWR.n2352 VGND 0.09471f
C19726 VPWR.t1474 VGND 0.09401f
C19727 VPWR.t1825 VGND 0.08295f
C19728 VPWR.t1124 VGND 0.11982f
C19729 VPWR.n2353 VGND 0.09471f
C19730 VPWR.n2354 VGND -0.00319f
C19731 VPWR.n2355 VGND 0.01815f
C19732 VPWR.n2356 VGND 0.14051f
C19733 VPWR.n2357 VGND 0.08433f
C19734 VPWR.n2358 VGND 0.08433f
C19735 VPWR.n2359 VGND 0.14051f
C19736 VPWR.n2360 VGND 0.01815f
C19737 VPWR.n2361 VGND -0.00319f
C19738 VPWR.n2362 VGND 0.09471f
C19739 VPWR.t1508 VGND 0.09401f
C19740 VPWR.t587 VGND 0.08295f
C19741 VPWR.t110 VGND 0.11982f
C19742 VPWR.n2363 VGND 0.09471f
C19743 VPWR.n2364 VGND -0.00319f
C19744 VPWR.n2365 VGND 0.01815f
C19745 VPWR.n2366 VGND 0.14051f
C19746 VPWR.n2367 VGND 0.08433f
C19747 VPWR.n2368 VGND 0.08433f
C19748 VPWR.n2369 VGND 0.14051f
C19749 VPWR.n2370 VGND 0.01815f
C19750 VPWR.n2371 VGND -0.00319f
C19751 VPWR.n2372 VGND 0.09471f
C19752 VPWR.t193 VGND 0.09401f
C19753 VPWR.t1827 VGND 0.08295f
C19754 VPWR.t244 VGND 0.11982f
C19755 VPWR.n2373 VGND 0.09471f
C19756 VPWR.n2374 VGND -0.00319f
C19757 VPWR.n2375 VGND 0.01815f
C19758 VPWR.n2376 VGND 0.14051f
C19759 VPWR.n2377 VGND 0.08433f
C19760 VPWR.n2378 VGND 0.08433f
C19761 VPWR.n2379 VGND 0.14051f
C19762 VPWR.n2380 VGND 0.01815f
C19763 VPWR.n2381 VGND -0.00319f
C19764 VPWR.n2382 VGND 0.09471f
C19765 VPWR.t505 VGND 0.09401f
C19766 VPWR.t589 VGND 0.08295f
C19767 VPWR.t1104 VGND 0.11982f
C19768 VPWR.n2383 VGND 0.09471f
C19769 VPWR.n2384 VGND -0.00319f
C19770 VPWR.n2385 VGND 0.01815f
C19771 VPWR.n2386 VGND 0.14051f
C19772 VPWR.n2387 VGND 0.08433f
C19773 VPWR.n2388 VGND 0.08433f
C19774 VPWR.n2389 VGND 0.14051f
C19775 VPWR.n2390 VGND 0.01815f
C19776 VPWR.n2391 VGND -0.00319f
C19777 VPWR.n2392 VGND 0.09471f
C19778 VPWR.t214 VGND 0.09401f
C19779 VPWR.t1828 VGND 0.08295f
C19780 VPWR.t1586 VGND 0.11982f
C19781 VPWR.n2393 VGND 0.09471f
C19782 VPWR.n2394 VGND -0.00319f
C19783 VPWR.n2395 VGND 0.01815f
C19784 VPWR.n2396 VGND 0.14051f
C19785 VPWR.n2397 VGND 0.08433f
C19786 VPWR.n2398 VGND 0.08433f
C19787 VPWR.n2399 VGND 0.14051f
C19788 VPWR.n2400 VGND 0.01815f
C19789 VPWR.n2401 VGND -0.00319f
C19790 VPWR.n2402 VGND 0.09471f
C19791 VPWR.t136 VGND 0.09401f
C19792 VPWR.t491 VGND 0.08295f
C19793 VPWR.t20 VGND 0.11982f
C19794 VPWR.n2403 VGND 0.09471f
C19795 VPWR.n2404 VGND -0.00319f
C19796 VPWR.n2405 VGND 0.01815f
C19797 VPWR.n2406 VGND 0.14051f
C19798 VPWR.n2407 VGND 0.08433f
C19799 VPWR.n2408 VGND 0.08433f
C19800 VPWR.n2409 VGND 0.14051f
C19801 VPWR.n2410 VGND 0.01815f
C19802 VPWR.n2411 VGND -0.00319f
C19803 VPWR.n2412 VGND 0.09471f
C19804 VPWR.t1536 VGND 0.09401f
C19805 VPWR.t1824 VGND 0.08295f
C19806 VPWR.t1039 VGND 0.11982f
C19807 VPWR.n2413 VGND 0.09471f
C19808 VPWR.n2414 VGND -0.00319f
C19809 VPWR.n2415 VGND 0.01815f
C19810 VPWR.n2416 VGND 0.14051f
C19811 VPWR.n2417 VGND 0.08433f
C19812 VPWR.n2418 VGND 1.01936f
C19813 VPWR.n2419 VGND 0.19562f
C19814 VPWR.n2420 VGND 0.08433f
C19815 VPWR.n2421 VGND 0.08433f
C19816 VPWR.n2422 VGND 0.08433f
C19817 VPWR.n2423 VGND 0.08433f
C19818 VPWR.n2424 VGND 0.08433f
C19819 VPWR.n2425 VGND 0.08433f
C19820 VPWR.n2426 VGND 0.08433f
C19821 VPWR.n2427 VGND 0.08433f
C19822 VPWR.n2428 VGND 0.08433f
C19823 VPWR.n2429 VGND 0.08433f
C19824 VPWR.n2430 VGND 0.08433f
C19825 VPWR.n2431 VGND 0.08433f
C19826 VPWR.n2432 VGND 0.08433f
C19827 VPWR.n2433 VGND 0.08433f
C19828 VPWR.n2434 VGND 0.08433f
C19829 VPWR.n2435 VGND 1.01936f
C19830 VPWR.n2436 VGND 0.57693f
C19831 VPWR.n2437 VGND 0.08433f
C19832 VPWR.n2438 VGND 0.08739f
C19833 VPWR.n2439 VGND 0.02426f
C19834 VPWR.n2440 VGND 0.00608f
C19835 VPWR.n2441 VGND -0.00323f
C19836 VPWR.n2442 VGND 0.09471f
C19837 VPWR.t929 VGND 0.11982f
C19838 VPWR.t637 VGND 0.08295f
C19839 VPWR.t634 VGND 0.09401f
C19840 VPWR.t649 VGND 0.08295f
C19841 VPWR.t651 VGND 0.11982f
C19842 VPWR.n2443 VGND 0.09471f
C19843 VPWR.n2444 VGND -0.00323f
C19844 VPWR.n2445 VGND 0.00608f
C19845 VPWR.n2446 VGND 0.02426f
C19846 VPWR.n2447 VGND 0.08739f
C19847 VPWR.n2448 VGND 0.08433f
C19848 VPWR.n2449 VGND 0.08433f
C19849 VPWR.n2450 VGND 0.08739f
C19850 VPWR.n2451 VGND 0.02426f
C19851 VPWR.n2452 VGND 0.00608f
C19852 VPWR.n2453 VGND -0.00323f
C19853 VPWR.n2454 VGND 0.09471f
C19854 VPWR.t689 VGND 0.11982f
C19855 VPWR.t687 VGND 0.08295f
C19856 VPWR.t684 VGND 0.09401f
C19857 VPWR.t905 VGND 0.08295f
C19858 VPWR.t907 VGND 0.11982f
C19859 VPWR.n2455 VGND 0.09471f
C19860 VPWR.n2456 VGND -0.00323f
C19861 VPWR.n2457 VGND 0.00608f
C19862 VPWR.n2458 VGND 0.02426f
C19863 VPWR.n2459 VGND 0.08739f
C19864 VPWR.n2460 VGND 0.08433f
C19865 VPWR.n2461 VGND 0.08433f
C19866 VPWR.n2462 VGND 0.08739f
C19867 VPWR.n2463 VGND 0.02426f
C19868 VPWR.n2464 VGND 0.00608f
C19869 VPWR.n2465 VGND -0.00323f
C19870 VPWR.n2466 VGND 0.09471f
C19871 VPWR.t926 VGND 0.11982f
C19872 VPWR.t944 VGND 0.08295f
C19873 VPWR.t941 VGND 0.09401f
C19874 VPWR.t697 VGND 0.08295f
C19875 VPWR.t699 VGND 0.11982f
C19876 VPWR.n2467 VGND 0.09471f
C19877 VPWR.n2468 VGND -0.00323f
C19878 VPWR.n2469 VGND 0.00608f
C19879 VPWR.n2470 VGND 0.02426f
C19880 VPWR.n2471 VGND 0.08739f
C19881 VPWR.n2472 VGND 0.08433f
C19882 VPWR.n2473 VGND 0.08433f
C19883 VPWR.n2474 VGND 0.08739f
C19884 VPWR.n2475 VGND 0.02426f
C19885 VPWR.n2476 VGND 0.00608f
C19886 VPWR.n2477 VGND -0.00323f
C19887 VPWR.n2478 VGND 0.09471f
C19888 VPWR.t795 VGND 0.11982f
C19889 VPWR.t793 VGND 0.08295f
C19890 VPWR.t812 VGND 0.09401f
C19891 VPWR.t834 VGND 0.08295f
C19892 VPWR.t831 VGND 0.11982f
C19893 VPWR.n2479 VGND 0.09471f
C19894 VPWR.n2480 VGND -0.00323f
C19895 VPWR.n2481 VGND 0.00608f
C19896 VPWR.n2482 VGND 0.02426f
C19897 VPWR.n2483 VGND 0.08739f
C19898 VPWR.n2484 VGND 0.08433f
C19899 VPWR.n2485 VGND 0.08433f
C19900 VPWR.n2486 VGND 0.08739f
C19901 VPWR.n2487 VGND 0.02426f
C19902 VPWR.n2488 VGND 0.00608f
C19903 VPWR.n2489 VGND -0.00323f
C19904 VPWR.n2490 VGND 0.09471f
C19905 VPWR.t972 VGND 0.11982f
C19906 VPWR.t970 VGND 0.08295f
C19907 VPWR.t676 VGND 0.09401f
C19908 VPWR.t713 VGND 0.08295f
C19909 VPWR.t715 VGND 0.11982f
C19910 VPWR.n2491 VGND 0.09471f
C19911 VPWR.n2492 VGND -0.00323f
C19912 VPWR.n2493 VGND 0.00608f
C19913 VPWR.n2494 VGND 0.02426f
C19914 VPWR.n2495 VGND 0.08739f
C19915 VPWR.n2496 VGND 0.08433f
C19916 VPWR.n2497 VGND 0.08433f
C19917 VPWR.n2498 VGND 0.08739f
C19918 VPWR.n2499 VGND 0.02426f
C19919 VPWR.n2500 VGND 0.00608f
C19920 VPWR.n2501 VGND -0.00323f
C19921 VPWR.n2502 VGND 0.09471f
C19922 VPWR.t850 VGND 0.11982f
C19923 VPWR.t848 VGND 0.08295f
C19924 VPWR.t842 VGND 0.09401f
C19925 VPWR.t981 VGND 0.08295f
C19926 VPWR.t881 VGND 0.11982f
C19927 VPWR.n2503 VGND 0.09471f
C19928 VPWR.n2504 VGND -0.00323f
C19929 VPWR.n2505 VGND 0.00608f
C19930 VPWR.n2506 VGND 0.02426f
C19931 VPWR.n2507 VGND 0.08739f
C19932 VPWR.n2508 VGND 0.08433f
C19933 VPWR.n2509 VGND 0.08433f
C19934 VPWR.n2510 VGND 0.08739f
C19935 VPWR.n2511 VGND 0.02426f
C19936 VPWR.n2512 VGND 0.00608f
C19937 VPWR.n2513 VGND -0.00323f
C19938 VPWR.n2514 VGND 0.09471f
C19939 VPWR.t621 VGND 0.11982f
C19940 VPWR.t619 VGND 0.08295f
C19941 VPWR.t616 VGND 0.09401f
C19942 VPWR.t758 VGND 0.08295f
C19943 VPWR.t760 VGND 0.11982f
C19944 VPWR.n2515 VGND 0.09471f
C19945 VPWR.n2516 VGND -0.00323f
C19946 VPWR.n2517 VGND 0.00608f
C19947 VPWR.n2518 VGND 0.02426f
C19948 VPWR.n2519 VGND 0.08739f
C19949 VPWR.n2520 VGND 0.08433f
C19950 VPWR.n2521 VGND 0.08433f
C19951 VPWR.n2522 VGND 0.08739f
C19952 VPWR.n2523 VGND 0.02426f
C19953 VPWR.n2524 VGND 0.00608f
C19954 VPWR.n2525 VGND -0.00323f
C19955 VPWR.n2526 VGND 0.09471f
C19956 VPWR.t870 VGND 0.11982f
C19957 VPWR.t868 VGND 0.08295f
C19958 VPWR.t839 VGND 0.14528f
C19959 VPWR.n2527 VGND 0.08262f
C19960 VPWR.n2528 VGND 0.00608f
C19961 VPWR.n2529 VGND 0.02407f
C19962 VPWR.n2530 VGND 0.1096f
C19963 VPWR.n2531 VGND 0.19562f
C19964 VPWR.n2532 VGND 2.68892f
C19965 VPWR.n2533 VGND 1.09505f
C19966 VPWR.n2534 VGND 0.45882f
C19967 VPWR.t1870 VGND 0.05509f
C19968 VPWR.t125 VGND 0.05509f
C19969 VPWR.n2535 VGND 0.09995f
C19970 VPWR.n2536 VGND 0.04733f
C19971 VPWR.t1869 VGND 0.01447f
C19972 VPWR.t1873 VGND 0.01447f
C19973 VPWR.n2537 VGND 0.03106f
C19974 VPWR.t135 VGND 0.01447f
C19975 VPWR.t123 VGND 0.01447f
C19976 VPWR.n2538 VGND 0.03106f
C19977 VPWR.n2539 VGND 0.01075f
C19978 VPWR.n2540 VGND 0.04733f
C19979 VPWR.t1776 VGND 0.01447f
C19980 VPWR.t1757 VGND 0.01447f
C19981 VPWR.n2541 VGND 0.03106f
C19982 VPWR.t1739 VGND 0.01447f
C19983 VPWR.t1746 VGND 0.01447f
C19984 VPWR.n2542 VGND 0.03106f
C19985 VPWR.t1753 VGND 0.0577f
C19986 VPWR.t1732 VGND 0.0577f
C19987 VPWR.n2543 VGND 0.13306f
C19988 VPWR.n2544 VGND 0.0427f
C19989 VPWR.n2545 VGND 0.01376f
C19990 VPWR.n2546 VGND 0.06244f
C19991 VPWR.n2547 VGND 0.00929f
C19992 VPWR.t1734 VGND 0.01447f
C19993 VPWR.t1872 VGND 0.01447f
C19994 VPWR.n2548 VGND 0.03106f
C19995 VPWR.t1752 VGND 0.01447f
C19996 VPWR.t131 VGND 0.01447f
C19997 VPWR.n2549 VGND 0.03106f
C19998 VPWR.n2550 VGND 0.06244f
C19999 VPWR.n2551 VGND 0.01439f
C20000 VPWR.n2552 VGND 0.04733f
C20001 VPWR.n2553 VGND 0.04733f
C20002 VPWR.n2554 VGND 0.04733f
C20003 VPWR.n2555 VGND 0.01294f
C20004 VPWR.n2556 VGND 0.06244f
C20005 VPWR.n2557 VGND 0.01221f
C20006 VPWR.n2558 VGND 0.00993f
C20007 VPWR.n2559 VGND 0.04733f
C20008 VPWR.n2560 VGND 0.0355f
C20009 VPWR.n2561 VGND 0.00802f
C20010 VPWR.t1731 VGND 0.17289f
C20011 VPWR.t1738 VGND 0.25478f
C20012 VPWR.t1745 VGND 0.25478f
C20013 VPWR.t1733 VGND 0.25478f
C20014 VPWR.t130 VGND 0.25478f
C20015 VPWR.t134 VGND 0.25478f
C20016 VPWR.t122 VGND 0.25478f
C20017 VPWR.t124 VGND 0.56722f
C20018 VPWR.n2562 VGND 0.61911f
C20019 VPWR.n2563 VGND 0.01801f
C20020 VPWR.n2564 VGND 1.08592f
C20021 VPWR.n2565 VGND 0.04733f
C20022 VPWR.t1729 VGND 0.17289f
C20023 VPWR.t1742 VGND 0.25478f
C20024 VPWR.t1716 VGND 0.25478f
C20025 VPWR.t1768 VGND 0.25478f
C20026 VPWR.t1148 VGND 0.25478f
C20027 VPWR.t1185 VGND 0.25478f
C20028 VPWR.t1146 VGND 0.25478f
C20029 VPWR.t1189 VGND 0.41857f
C20030 VPWR.t1096 VGND 0.44435f
C20031 VPWR.n2566 VGND 0.62705f
C20032 VPWR.n2567 VGND 0.17837f
C20033 VPWR.n2568 VGND 0.04733f
C20034 VPWR.t1619 VGND 0.01447f
C20035 VPWR.t1147 VGND 0.01447f
C20036 VPWR.n2569 VGND 0.03106f
C20037 VPWR.t1186 VGND 0.01447f
C20038 VPWR.t1195 VGND 0.01447f
C20039 VPWR.n2570 VGND 0.03106f
C20040 VPWR.n2571 VGND 0.06244f
C20041 VPWR.n2572 VGND 0.04733f
C20042 VPWR.t1779 VGND 0.01447f
C20043 VPWR.t1149 VGND 0.01447f
C20044 VPWR.n2573 VGND 0.03106f
C20045 VPWR.t1769 VGND 0.01447f
C20046 VPWR.t1193 VGND 0.01447f
C20047 VPWR.n2574 VGND 0.03106f
C20048 VPWR.n2575 VGND 0.00929f
C20049 VPWR.t1730 VGND 0.0577f
C20050 VPWR.t1778 VGND 0.0577f
C20051 VPWR.n2576 VGND 0.13306f
C20052 VPWR.t1761 VGND 0.01447f
C20053 VPWR.t1736 VGND 0.01447f
C20054 VPWR.n2577 VGND 0.03106f
C20055 VPWR.t1743 VGND 0.01447f
C20056 VPWR.t1717 VGND 0.01447f
C20057 VPWR.n2578 VGND 0.03106f
C20058 VPWR.n2579 VGND 0.06244f
C20059 VPWR.n2580 VGND 0.01376f
C20060 VPWR.n2581 VGND 0.0427f
C20061 VPWR.n2582 VGND 0.04733f
C20062 VPWR.n2583 VGND 0.04733f
C20063 VPWR.n2584 VGND 0.01439f
C20064 VPWR.n2585 VGND 0.06244f
C20065 VPWR.n2586 VGND 0.01075f
C20066 VPWR.n2587 VGND 0.01294f
C20067 VPWR.n2588 VGND 0.04733f
C20068 VPWR.n2589 VGND 0.04733f
C20069 VPWR.n2590 VGND 0.01221f
C20070 VPWR.n2591 VGND 0.00993f
C20071 VPWR.t1618 VGND 0.05509f
C20072 VPWR.t1190 VGND 0.05509f
C20073 VPWR.n2592 VGND 0.09995f
C20074 VPWR.n2593 VGND 0.00802f
C20075 VPWR.n2594 VGND 0.0355f
C20076 VPWR.n2595 VGND 0.01801f
C20077 VPWR.n2596 VGND 0.0355f
C20078 VPWR.n2597 VGND 0.01412f
C20079 VPWR.n2598 VGND 0.01093f
C20080 VPWR.t1631 VGND 0.05764f
C20081 VPWR.t1097 VGND 0.05764f
C20082 VPWR.n2599 VGND 0.11651f
C20083 VPWR.n2600 VGND 0.03293f
C20084 VPWR.n2601 VGND 1.65272f
C20085 VPWR.n2602 VGND 0.04733f
C20086 VPWR.t275 VGND 0.05658f
C20087 VPWR.t1763 VGND 0.17289f
C20088 VPWR.t1720 VGND 0.25478f
C20089 VPWR.t1770 VGND 0.25478f
C20090 VPWR.t1747 VGND 0.25478f
C20091 VPWR.t1640 VGND 0.25478f
C20092 VPWR.t1634 VGND 0.25478f
C20093 VPWR.t1053 VGND 0.25478f
C20094 VPWR.t1636 VGND 0.41857f
C20095 VPWR.t1196 VGND 0.16075f
C20096 VPWR.t274 VGND 0.12739f
C20097 VPWR.t1300 VGND 0.28359f
C20098 VPWR.n2603 VGND 0.55577f
C20099 VPWR.n2604 VGND 0.17573f
C20100 VPWR.n2605 VGND 0.04733f
C20101 VPWR.t1635 VGND 0.01447f
C20102 VPWR.t1642 VGND 0.01447f
C20103 VPWR.n2606 VGND 0.03106f
C20104 VPWR.t1915 VGND 0.01447f
C20105 VPWR.t1054 VGND 0.01447f
C20106 VPWR.n2607 VGND 0.03106f
C20107 VPWR.n2608 VGND 0.06244f
C20108 VPWR.n2609 VGND 0.04733f
C20109 VPWR.t1765 VGND 0.01447f
C20110 VPWR.t1641 VGND 0.01447f
C20111 VPWR.n2610 VGND 0.03106f
C20112 VPWR.t1748 VGND 0.01447f
C20113 VPWR.t1912 VGND 0.01447f
C20114 VPWR.n2611 VGND 0.03106f
C20115 VPWR.n2612 VGND 0.00929f
C20116 VPWR.t1777 VGND 0.0577f
C20117 VPWR.t1764 VGND 0.0577f
C20118 VPWR.n2613 VGND 0.13306f
C20119 VPWR.t1740 VGND 0.01447f
C20120 VPWR.t1783 VGND 0.01447f
C20121 VPWR.n2614 VGND 0.03106f
C20122 VPWR.t1721 VGND 0.01447f
C20123 VPWR.t1771 VGND 0.01447f
C20124 VPWR.n2615 VGND 0.03106f
C20125 VPWR.n2616 VGND 0.06244f
C20126 VPWR.n2617 VGND 0.01376f
C20127 VPWR.n2618 VGND 0.0427f
C20128 VPWR.n2619 VGND 0.04733f
C20129 VPWR.n2620 VGND 0.04733f
C20130 VPWR.n2621 VGND 0.01439f
C20131 VPWR.n2622 VGND 0.06244f
C20132 VPWR.n2623 VGND 0.01075f
C20133 VPWR.n2624 VGND 0.01294f
C20134 VPWR.n2625 VGND 0.04733f
C20135 VPWR.n2626 VGND 0.04733f
C20136 VPWR.n2627 VGND 0.01221f
C20137 VPWR.n2628 VGND 0.00993f
C20138 VPWR.t1637 VGND 0.05509f
C20139 VPWR.t1914 VGND 0.05509f
C20140 VPWR.n2629 VGND 0.09995f
C20141 VPWR.n2630 VGND 0.00802f
C20142 VPWR.n2631 VGND 0.0355f
C20143 VPWR.n2632 VGND 0.01801f
C20144 VPWR.n2633 VGND 0.0355f
C20145 VPWR.t1301 VGND 0.05771f
C20146 VPWR.n2634 VGND 0.08042f
C20147 VPWR.n2635 VGND 0.01075f
C20148 VPWR.n2636 VGND 0.05885f
C20149 VPWR.t1197 VGND 0.05673f
C20150 VPWR.n2637 VGND 0.07353f
C20151 VPWR.n2638 VGND 0.02804f
C20152 VPWR.n2639 VGND 1.65272f
C20153 VPWR.n2640 VGND 0.04733f
C20154 VPWR.t1766 VGND 0.09805f
C20155 VPWR.t1724 VGND 0.14449f
C20156 VPWR.t1772 VGND 0.14048f
C20157 VPWR.t1750 VGND 0.22466f
C20158 VPWR.t388 VGND 0.19108f
C20159 VPWR.t1754 VGND 0.12739f
C20160 VPWR.t394 VGND 0.12739f
C20161 VPWR.t1726 VGND 0.12739f
C20162 VPWR.t1156 VGND 0.12739f
C20163 VPWR.t1758 VGND 0.12739f
C20164 VPWR.t392 VGND 0.12739f
C20165 VPWR.t1781 VGND 0.17743f
C20166 VPWR.t1446 VGND 0.10009f
C20167 VPWR.t531 VGND 0.10919f
C20168 VPWR.t1126 VGND 0.12739f
C20169 VPWR.t533 VGND 0.23658f
C20170 VPWR.n2641 VGND 0.38137f
C20171 VPWR.n2642 VGND 0.17591f
C20172 VPWR.t534 VGND 0.05728f
C20173 VPWR.n2643 VGND 0.04733f
C20174 VPWR.t1782 VGND 0.05662f
C20175 VPWR.t393 VGND 0.0545f
C20176 VPWR.t1727 VGND 0.01447f
C20177 VPWR.t1759 VGND 0.01447f
C20178 VPWR.n2644 VGND 0.03106f
C20179 VPWR.t395 VGND 0.01447f
C20180 VPWR.t1157 VGND 0.01447f
C20181 VPWR.n2645 VGND 0.03106f
C20182 VPWR.n2646 VGND 0.03541f
C20183 VPWR.n2647 VGND 0.04733f
C20184 VPWR.t1751 VGND 0.01447f
C20185 VPWR.t389 VGND 0.01447f
C20186 VPWR.n2648 VGND 0.03106f
C20187 VPWR.n2649 VGND 0.00929f
C20188 VPWR.t1767 VGND 0.0577f
C20189 VPWR.n2650 VGND 0.07271f
C20190 VPWR.t1725 VGND 0.01447f
C20191 VPWR.t1773 VGND 0.01447f
C20192 VPWR.n2651 VGND 0.03106f
C20193 VPWR.n2652 VGND 0.03541f
C20194 VPWR.n2653 VGND 0.01376f
C20195 VPWR.n2654 VGND 0.0427f
C20196 VPWR.n2655 VGND 0.04733f
C20197 VPWR.n2656 VGND 0.04733f
C20198 VPWR.n2657 VGND 0.01439f
C20199 VPWR.n2658 VGND 0.03459f
C20200 VPWR.t1755 VGND 0.05064f
C20201 VPWR.n2659 VGND 0.04037f
C20202 VPWR.n2660 VGND 0.00993f
C20203 VPWR.n2661 VGND 0.04733f
C20204 VPWR.n2662 VGND 0.04733f
C20205 VPWR.n2663 VGND 0.03924f
C20206 VPWR.n2664 VGND 0.01221f
C20207 VPWR.n2665 VGND 0.05193f
C20208 VPWR.n2666 VGND 0.06842f
C20209 VPWR.n2667 VGND 0.00629f
C20210 VPWR.n2668 VGND 0.02804f
C20211 VPWR.n2669 VGND 0.01801f
C20212 VPWR.n2670 VGND 0.0355f
C20213 VPWR.t1127 VGND 0.05776f
C20214 VPWR.n2671 VGND 0.14851f
C20215 VPWR.n2672 VGND 0.01093f
C20216 VPWR.t532 VGND 0.05767f
C20217 VPWR.n2673 VGND 0.06419f
C20218 VPWR.n2674 VGND 0.02778f
C20219 VPWR.n2675 VGND 1.65272f
C20220 VPWR.n2676 VGND 0.0427f
C20221 VPWR.t1760 VGND 0.67334f
C20222 VPWR.t1719 VGND 0.25478f
C20223 VPWR.t1749 VGND 0.25478f
C20224 VPWR.t1723 VGND 0.25478f
C20225 VPWR.t128 VGND 0.25478f
C20226 VPWR.t126 VGND 0.25478f
C20227 VPWR.t132 VGND 0.25478f
C20228 VPWR.t120 VGND 0.23051f
C20229 VPWR.t555 VGND 0.55809f
C20230 VPWR.t1130 VGND 0.15469f
C20231 VPWR.n2677 VGND 0.33436f
C20232 VPWR.n2678 VGND 0.17837f
C20233 VPWR.t1874 VGND 0.01447f
C20234 VPWR.t1871 VGND 0.01447f
C20235 VPWR.n2679 VGND 0.03172f
C20236 VPWR.t129 VGND 0.01447f
C20237 VPWR.t127 VGND 0.01447f
C20238 VPWR.n2680 VGND 0.03172f
C20239 VPWR.n2681 VGND 0.12037f
C20240 VPWR.n2682 VGND 0.09759f
C20241 VPWR.t1875 VGND 0.01447f
C20242 VPWR.t1876 VGND 0.01447f
C20243 VPWR.n2683 VGND 0.03177f
C20244 VPWR.t133 VGND 0.01447f
C20245 VPWR.t121 VGND 0.01447f
C20246 VPWR.n2684 VGND 0.03177f
C20247 VPWR.n2685 VGND 0.13194f
C20248 VPWR.n2686 VGND 0.0113f
C20249 VPWR.n2687 VGND 0.38113f
C20250 VPWR.n2688 VGND 0.01801f
C20251 VPWR.n2689 VGND 0.01646f
C20252 VPWR.n2690 VGND 0.01412f
C20253 VPWR.n2691 VGND 0.01321f
C20254 VPWR.t556 VGND 0.05776f
C20255 VPWR.t1461 VGND 0.05776f
C20256 VPWR.n2692 VGND 0.1706f
C20257 VPWR.n2693 VGND 0.0355f
C20258 VPWR.n2694 VGND 1.65272f
C20259 VPWR.n2695 VGND 0.0427f
C20260 VPWR.t1741 VGND 0.67334f
C20261 VPWR.t1774 VGND 0.25478f
C20262 VPWR.t1728 VGND 0.25478f
C20263 VPWR.t1775 VGND 0.25478f
C20264 VPWR.t535 VGND 0.25478f
C20265 VPWR.t1150 VGND 0.25478f
C20266 VPWR.t1187 VGND 0.25478f
C20267 VPWR.t1191 VGND 0.23051f
C20268 VPWR.t34 VGND 0.49591f
C20269 VPWR.t1132 VGND 0.10919f
C20270 VPWR.t1136 VGND 0.10768f
C20271 VPWR.n2696 VGND 0.33284f
C20272 VPWR.n2697 VGND 0.17837f
C20273 VPWR.t536 VGND 0.01447f
C20274 VPWR.t1151 VGND 0.01447f
C20275 VPWR.n2698 VGND 0.03172f
C20276 VPWR.t1184 VGND 0.01447f
C20277 VPWR.t1194 VGND 0.01447f
C20278 VPWR.n2699 VGND 0.03172f
C20279 VPWR.n2700 VGND 0.12037f
C20280 VPWR.n2701 VGND 0.09759f
C20281 VPWR.t1621 VGND 0.01447f
C20282 VPWR.t1620 VGND 0.01447f
C20283 VPWR.n2702 VGND 0.03177f
C20284 VPWR.t1188 VGND 0.01447f
C20285 VPWR.t1192 VGND 0.01447f
C20286 VPWR.n2703 VGND 0.03177f
C20287 VPWR.n2704 VGND 0.13194f
C20288 VPWR.n2705 VGND 0.0113f
C20289 VPWR.n2706 VGND 0.38113f
C20290 VPWR.n2707 VGND 0.01801f
C20291 VPWR.n2708 VGND 0.0162f
C20292 VPWR.n2709 VGND 0.00774f
C20293 VPWR.t1133 VGND 0.05764f
C20294 VPWR.n2710 VGND 0.06161f
C20295 VPWR.n2711 VGND 0.00738f
C20296 VPWR.t35 VGND 0.05776f
C20297 VPWR.n2712 VGND 0.092f
C20298 VPWR.n2713 VGND 0.0355f
C20299 VPWR.n2714 VGND 1.65272f
C20300 VPWR.n2715 VGND 0.04321f
C20301 VPWR.t1722 VGND 0.67334f
C20302 VPWR.t1735 VGND 0.25478f
C20303 VPWR.t1762 VGND 0.25478f
C20304 VPWR.t1737 VGND 0.25478f
C20305 VPWR.t1051 VGND 0.25478f
C20306 VPWR.t1638 VGND 0.25478f
C20307 VPWR.t1166 VGND 0.25478f
C20308 VPWR.t1164 VGND 0.23051f
C20309 VPWR.t557 VGND 0.52776f
C20310 VPWR.t1128 VGND 0.18199f
C20311 VPWR.n2716 VGND 0.33133f
C20312 VPWR.n2717 VGND 0.17573f
C20313 VPWR.t1131 VGND 0.05772f
C20314 VPWR.t1643 VGND 0.01447f
C20315 VPWR.t1639 VGND 0.01447f
C20316 VPWR.n2718 VGND 0.03172f
C20317 VPWR.t1052 VGND 0.01447f
C20318 VPWR.t1913 VGND 0.01447f
C20319 VPWR.n2719 VGND 0.03172f
C20320 VPWR.n2720 VGND 0.12037f
C20321 VPWR.n2721 VGND 0.09759f
C20322 VPWR.t1632 VGND 0.01447f
C20323 VPWR.t1633 VGND 0.01447f
C20324 VPWR.n2722 VGND 0.03177f
C20325 VPWR.t1167 VGND 0.01447f
C20326 VPWR.t1165 VGND 0.01447f
C20327 VPWR.n2723 VGND 0.03177f
C20328 VPWR.n2724 VGND 0.13194f
C20329 VPWR.n2725 VGND 0.0113f
C20330 VPWR.n2726 VGND 0.38113f
C20331 VPWR.n2727 VGND 0.01801f
C20332 VPWR.n2728 VGND 0.01595f
C20333 VPWR.t1129 VGND 0.05772f
C20334 VPWR.n2729 VGND 0.15208f
C20335 VPWR.n2730 VGND 0.01221f
C20336 VPWR.t558 VGND 0.05771f
C20337 VPWR.t1460 VGND 0.05771f
C20338 VPWR.n2731 VGND 0.13578f
C20339 VPWR.n2732 VGND 0.0355f
C20340 VPWR.n2733 VGND 1.65272f
C20341 VPWR.n2734 VGND 0.04321f
C20342 VPWR.t33 VGND 0.05771f
C20343 VPWR.n2735 VGND 0.01595f
C20344 VPWR.t1135 VGND 0.05772f
C20345 VPWR.n2736 VGND 0.01801f
C20346 VPWR.t1756 VGND 0.38188f
C20347 VPWR.t1780 VGND 0.14449f
C20348 VPWR.t1744 VGND 0.14449f
C20349 VPWR.t1718 VGND 0.14449f
C20350 VPWR.t390 VGND 0.14449f
C20351 VPWR.t573 VGND 0.14449f
C20352 VPWR.t1154 VGND 0.14449f
C20353 VPWR.t1152 VGND 0.13073f
C20354 VPWR.t32 VGND 0.29931f
C20355 VPWR.t1134 VGND 0.10321f
C20356 VPWR.n2737 VGND 0.1844f
C20357 VPWR.t1155 VGND 0.01447f
C20358 VPWR.t1153 VGND 0.01447f
C20359 VPWR.n2738 VGND 0.03177f
C20360 VPWR.n2739 VGND 0.07818f
C20361 VPWR.t391 VGND 0.01447f
C20362 VPWR.t574 VGND 0.01447f
C20363 VPWR.n2740 VGND 0.03306f
C20364 VPWR.n2741 VGND 0.17652f
C20365 VPWR.n2742 VGND 0.38113f
C20366 VPWR.n2743 VGND 0.0113f
C20367 VPWR.n2744 VGND 0.09757f
C20368 VPWR.n2745 VGND 0.08565f
C20369 VPWR.n2746 VGND 0.01221f
C20370 VPWR.n2747 VGND 0.07422f
C20371 VPWR.n2748 VGND 0.0355f
C20372 VPWR.n2749 VGND 2.4051f
C20373 VPWR.n2750 VGND 1.94782f
C20374 VPWR.t400 VGND 0.02934f
C20375 VPWR.n2751 VGND 0.13152f
C20376 VPWR.n2752 VGND 0.28949f
C20377 VPWR.n2753 VGND 0.07634f
C20378 VPWR.n2754 VGND 0.03626f
C20379 VPWR.n2755 VGND 0.04427f
C20380 VPWR.n2756 VGND 0.08973f
C20381 VPWR.n2757 VGND 0.11697f
C20382 VPWR.n2758 VGND 0.08973f
C20383 VPWR.t1210 VGND 2.82254f
C20384 VPWR.t399 VGND 0.89146f
C20385 VPWR.n2759 VGND 0.11789f
C20386 VPWR.n2760 VGND 0.46644f
C20387 VPWR.t1911 VGND 0.02933f
C20388 VPWR.n2761 VGND 0.17958f
C20389 VPWR.n2762 VGND 0.01813f
C20390 VPWR.n2763 VGND 0.09893f
C20391 VPWR.n2764 VGND 0.08882f
C20392 VPWR.n2765 VGND 0.11789f
C20393 VPWR.n2766 VGND 0.07425f
C20394 VPWR.t1211 VGND 0.02933f
C20395 VPWR.n2767 VGND 0.17958f
C20396 VPWR.n2768 VGND 0.01813f
C20397 VPWR.n2769 VGND 0.11789f
C20398 VPWR.n2770 VGND 0.07715f
C20399 VPWR.n2771 VGND 0.08799f
C20400 VPWR.n2772 VGND 1.68677f
C20401 VPWR.n2773 VGND 0.08799f
C20402 VPWR.n2774 VGND 0.07715f
C20403 VPWR.n2775 VGND 0.11789f
C20404 VPWR.n2776 VGND 0.09884f
C20405 VPWR.n2777 VGND 0.08176f
C20406 VPWR.n2778 VGND 1.01392f
C20407 VPWR.n2779 VGND 0.0638f
C20408 VPWR.n2780 VGND 0.08924f
C20409 VPWR.n2781 VGND 0.06203f
C20410 VPWR.n2782 VGND 0.01813f
C20411 VPWR.n2783 VGND 0.0638f
C20412 VPWR.n2784 VGND 0.04898f
C20413 VPWR.n2785 VGND 0.17527f
C20414 VPWR.n2786 VGND 0.06905f
C20415 VPWR.n2787 VGND 0.04427f
C20416 VPWR.t1859 VGND 0.34902f
C20417 VPWR.n2788 VGND 0.08176f
C20418 VPWR.n2789 VGND 0.09884f
C20419 VPWR.n2790 VGND 0.03626f
C20420 VPWR.n2791 VGND 2.04283f
C20421 VPWR.n2792 VGND 0.03626f
C20422 VPWR.n2793 VGND 0.03626f
C20423 VPWR.n2794 VGND 0.0901f
C20424 VPWR.n2795 VGND 0.04947f
C20425 VPWR.n2796 VGND 0.38311f
C20426 VPWR.n2797 VGND 0.31521f
C20427 VPWR.t1860 VGND 0.02932f
C20428 VPWR.n2798 VGND 0.22184f
C20429 VPWR.n2799 VGND 3.38263f
C20430 Iout.n0 VGND 0.23929f
C20431 Iout.n1 VGND 1.25122f
C20432 Iout.n2 VGND 0.23929f
C20433 Iout.n3 VGND 0.23929f
C20434 Iout.t244 VGND 0.02304f
C20435 Iout.n4 VGND 0.05124f
C20436 Iout.n5 VGND 0.20242f
C20437 Iout.n6 VGND 0.23929f
C20438 Iout.n7 VGND 1.25122f
C20439 Iout.n8 VGND 0.23929f
C20440 Iout.t28 VGND 0.02304f
C20441 Iout.n9 VGND 0.05124f
C20442 Iout.n10 VGND 0.20242f
C20443 Iout.n11 VGND 0.23929f
C20444 Iout.n12 VGND 1.25122f
C20445 Iout.n13 VGND 0.23929f
C20446 Iout.t119 VGND 0.02304f
C20447 Iout.n14 VGND 0.05124f
C20448 Iout.n15 VGND 0.20242f
C20449 Iout.n16 VGND 0.23929f
C20450 Iout.n17 VGND 1.25122f
C20451 Iout.n18 VGND 0.23929f
C20452 Iout.t89 VGND 0.02304f
C20453 Iout.n19 VGND 0.05124f
C20454 Iout.n20 VGND 0.20242f
C20455 Iout.n21 VGND 0.49611f
C20456 Iout.t168 VGND 0.02304f
C20457 Iout.n22 VGND 0.05124f
C20458 Iout.n23 VGND 0.29851f
C20459 Iout.n24 VGND 0.23929f
C20460 Iout.n25 VGND 0.23929f
C20461 Iout.n26 VGND 0.23929f
C20462 Iout.n27 VGND 0.23929f
C20463 Iout.n28 VGND 0.23929f
C20464 Iout.n29 VGND 0.23929f
C20465 Iout.n30 VGND 0.23929f
C20466 Iout.n31 VGND 0.23929f
C20467 Iout.n32 VGND 0.23929f
C20468 Iout.n33 VGND 0.23929f
C20469 Iout.n34 VGND 0.23929f
C20470 Iout.n35 VGND 0.23929f
C20471 Iout.n36 VGND 0.23929f
C20472 Iout.n37 VGND 0.23929f
C20473 Iout.t212 VGND 0.02304f
C20474 Iout.n38 VGND 0.05124f
C20475 Iout.n39 VGND 0.02606f
C20476 Iout.n40 VGND 0.23929f
C20477 Iout.n41 VGND 0.04775f
C20478 Iout.t45 VGND 0.02304f
C20479 Iout.n42 VGND 0.05124f
C20480 Iout.n43 VGND 0.02606f
C20481 Iout.t61 VGND 0.02304f
C20482 Iout.n44 VGND 0.05124f
C20483 Iout.n45 VGND 0.02606f
C20484 Iout.n46 VGND 0.23929f
C20485 Iout.t204 VGND 0.02304f
C20486 Iout.n47 VGND 0.05124f
C20487 Iout.n48 VGND 0.02606f
C20488 Iout.n49 VGND 0.23929f
C20489 Iout.t229 VGND 0.02304f
C20490 Iout.n50 VGND 0.05124f
C20491 Iout.n51 VGND 0.02606f
C20492 Iout.n52 VGND 0.23929f
C20493 Iout.t133 VGND 0.02304f
C20494 Iout.n53 VGND 0.05124f
C20495 Iout.n54 VGND 0.02606f
C20496 Iout.n55 VGND 0.23929f
C20497 Iout.t254 VGND 0.02304f
C20498 Iout.n56 VGND 0.05124f
C20499 Iout.n57 VGND 0.02606f
C20500 Iout.n58 VGND 0.23929f
C20501 Iout.t15 VGND 0.02304f
C20502 Iout.n59 VGND 0.05124f
C20503 Iout.n60 VGND 0.02606f
C20504 Iout.n61 VGND 0.23929f
C20505 Iout.t184 VGND 0.02304f
C20506 Iout.n62 VGND 0.05124f
C20507 Iout.n63 VGND 0.02606f
C20508 Iout.n64 VGND 0.23929f
C20509 Iout.t146 VGND 0.02304f
C20510 Iout.n65 VGND 0.05124f
C20511 Iout.n66 VGND 0.02606f
C20512 Iout.n67 VGND 0.23929f
C20513 Iout.t22 VGND 0.02304f
C20514 Iout.n68 VGND 0.05124f
C20515 Iout.n69 VGND 0.02606f
C20516 Iout.n70 VGND 0.23929f
C20517 Iout.t60 VGND 0.02304f
C20518 Iout.n71 VGND 0.05124f
C20519 Iout.n72 VGND 0.02606f
C20520 Iout.n73 VGND 0.23929f
C20521 Iout.t170 VGND 0.02304f
C20522 Iout.n74 VGND 0.05124f
C20523 Iout.n75 VGND 0.02606f
C20524 Iout.n76 VGND 0.23929f
C20525 Iout.t154 VGND 0.02304f
C20526 Iout.n77 VGND 0.05124f
C20527 Iout.n78 VGND 0.02606f
C20528 Iout.n79 VGND 0.23929f
C20529 Iout.n80 VGND 0.23929f
C20530 Iout.t90 VGND 0.02304f
C20531 Iout.n81 VGND 0.05124f
C20532 Iout.n82 VGND 0.02606f
C20533 Iout.n83 VGND 0.23929f
C20534 Iout.n84 VGND 0.04775f
C20535 Iout.t106 VGND 0.02304f
C20536 Iout.n85 VGND 0.05124f
C20537 Iout.n86 VGND 0.02606f
C20538 Iout.t21 VGND 0.02304f
C20539 Iout.n87 VGND 0.05124f
C20540 Iout.n88 VGND 0.02606f
C20541 Iout.n89 VGND 0.23929f
C20542 Iout.t197 VGND 0.02304f
C20543 Iout.n90 VGND 0.05124f
C20544 Iout.n91 VGND 0.02606f
C20545 Iout.n92 VGND 0.23929f
C20546 Iout.t173 VGND 0.02304f
C20547 Iout.n93 VGND 0.05124f
C20548 Iout.n94 VGND 0.02606f
C20549 Iout.n95 VGND 0.23929f
C20550 Iout.t214 VGND 0.02304f
C20551 Iout.n96 VGND 0.05124f
C20552 Iout.n97 VGND 0.02606f
C20553 Iout.n98 VGND 0.23929f
C20554 Iout.t179 VGND 0.02304f
C20555 Iout.n99 VGND 0.05124f
C20556 Iout.n100 VGND 0.02606f
C20557 Iout.n101 VGND 0.23929f
C20558 Iout.t56 VGND 0.02304f
C20559 Iout.n102 VGND 0.05124f
C20560 Iout.n103 VGND 0.02606f
C20561 Iout.n104 VGND 0.23929f
C20562 Iout.t13 VGND 0.02304f
C20563 Iout.n105 VGND 0.05124f
C20564 Iout.n106 VGND 0.02606f
C20565 Iout.n107 VGND 0.23929f
C20566 Iout.t79 VGND 0.02304f
C20567 Iout.n108 VGND 0.05124f
C20568 Iout.n109 VGND 0.02606f
C20569 Iout.n110 VGND 0.23929f
C20570 Iout.t55 VGND 0.02304f
C20571 Iout.n111 VGND 0.05124f
C20572 Iout.n112 VGND 0.02606f
C20573 Iout.n113 VGND 0.23929f
C20574 Iout.t117 VGND 0.02304f
C20575 Iout.n114 VGND 0.05124f
C20576 Iout.n115 VGND 0.02606f
C20577 Iout.n116 VGND 0.23929f
C20578 Iout.t240 VGND 0.02304f
C20579 Iout.n117 VGND 0.05124f
C20580 Iout.n118 VGND 0.02606f
C20581 Iout.n119 VGND 0.23929f
C20582 Iout.t118 VGND 0.02304f
C20583 Iout.n120 VGND 0.05124f
C20584 Iout.n121 VGND 0.02606f
C20585 Iout.n122 VGND 0.04775f
C20586 Iout.t14 VGND 0.02304f
C20587 Iout.n123 VGND 0.05124f
C20588 Iout.n124 VGND 0.02606f
C20589 Iout.n125 VGND 0.23929f
C20590 Iout.n126 VGND 0.23929f
C20591 Iout.t188 VGND 0.02304f
C20592 Iout.n127 VGND 0.05124f
C20593 Iout.n128 VGND 0.02606f
C20594 Iout.n129 VGND 0.04775f
C20595 Iout.t203 VGND 0.02304f
C20596 Iout.n130 VGND 0.05124f
C20597 Iout.n131 VGND 0.02606f
C20598 Iout.n132 VGND 0.23929f
C20599 Iout.t123 VGND 0.02304f
C20600 Iout.n133 VGND 0.05124f
C20601 Iout.n134 VGND 0.02606f
C20602 Iout.n135 VGND 0.04775f
C20603 Iout.t248 VGND 0.02304f
C20604 Iout.n136 VGND 0.05124f
C20605 Iout.n137 VGND 0.02606f
C20606 Iout.n138 VGND 0.23929f
C20607 Iout.n139 VGND 0.23929f
C20608 Iout.t53 VGND 0.02304f
C20609 Iout.n140 VGND 0.05124f
C20610 Iout.n141 VGND 0.02606f
C20611 Iout.n142 VGND 0.04775f
C20612 Iout.t171 VGND 0.02304f
C20613 Iout.n143 VGND 0.05124f
C20614 Iout.n144 VGND 0.02606f
C20615 Iout.n145 VGND 0.14126f
C20616 Iout.t255 VGND 0.02304f
C20617 Iout.n146 VGND 0.05124f
C20618 Iout.n147 VGND 0.02606f
C20619 Iout.n148 VGND 0.04775f
C20620 Iout.t157 VGND 0.02304f
C20621 Iout.n149 VGND 0.05124f
C20622 Iout.n150 VGND 0.02606f
C20623 Iout.n151 VGND 0.23929f
C20624 Iout.n152 VGND 0.14126f
C20625 Iout.n153 VGND 0.23929f
C20626 Iout.n154 VGND 0.23929f
C20627 Iout.n155 VGND 0.23929f
C20628 Iout.t165 VGND 0.02304f
C20629 Iout.n156 VGND 0.05124f
C20630 Iout.n157 VGND 0.02606f
C20631 Iout.n158 VGND 0.23929f
C20632 Iout.n159 VGND 0.23929f
C20633 Iout.n160 VGND 0.23929f
C20634 Iout.n161 VGND 0.23929f
C20635 Iout.n162 VGND 0.23929f
C20636 Iout.n163 VGND 0.23929f
C20637 Iout.n164 VGND 0.23929f
C20638 Iout.n165 VGND 0.23929f
C20639 Iout.n166 VGND 0.23929f
C20640 Iout.n167 VGND 0.23929f
C20641 Iout.t195 VGND 0.02304f
C20642 Iout.n168 VGND 0.05124f
C20643 Iout.n169 VGND 0.02606f
C20644 Iout.n170 VGND 0.23929f
C20645 Iout.n171 VGND 0.04775f
C20646 Iout.t211 VGND 0.02304f
C20647 Iout.n172 VGND 0.05124f
C20648 Iout.n173 VGND 0.02606f
C20649 Iout.t242 VGND 0.02304f
C20650 Iout.n174 VGND 0.05124f
C20651 Iout.n175 VGND 0.02606f
C20652 Iout.n176 VGND 0.23929f
C20653 Iout.t103 VGND 0.02304f
C20654 Iout.n177 VGND 0.05124f
C20655 Iout.n178 VGND 0.02606f
C20656 Iout.n179 VGND 0.23929f
C20657 Iout.t59 VGND 0.02304f
C20658 Iout.n180 VGND 0.05124f
C20659 Iout.n181 VGND 0.02606f
C20660 Iout.n182 VGND 0.23929f
C20661 Iout.t39 VGND 0.02304f
C20662 Iout.n183 VGND 0.05124f
C20663 Iout.n184 VGND 0.02606f
C20664 Iout.n185 VGND 0.23929f
C20665 Iout.t172 VGND 0.02304f
C20666 Iout.n186 VGND 0.05124f
C20667 Iout.n187 VGND 0.02606f
C20668 Iout.n188 VGND 0.23929f
C20669 Iout.t216 VGND 0.02304f
C20670 Iout.n189 VGND 0.05124f
C20671 Iout.n190 VGND 0.02606f
C20672 Iout.n191 VGND 0.14126f
C20673 Iout.t155 VGND 0.02304f
C20674 Iout.n192 VGND 0.05124f
C20675 Iout.n193 VGND 0.02606f
C20676 Iout.n194 VGND 0.04775f
C20677 Iout.t0 VGND 0.02304f
C20678 Iout.n195 VGND 0.05124f
C20679 Iout.n196 VGND 0.02606f
C20680 Iout.n197 VGND 0.14126f
C20681 Iout.n198 VGND 0.04775f
C20682 Iout.t75 VGND 0.02304f
C20683 Iout.n199 VGND 0.05124f
C20684 Iout.n200 VGND 0.02606f
C20685 Iout.n201 VGND 0.04775f
C20686 Iout.t8 VGND 0.02304f
C20687 Iout.n202 VGND 0.05124f
C20688 Iout.n203 VGND 0.02606f
C20689 Iout.n204 VGND 0.14126f
C20690 Iout.n205 VGND 0.04775f
C20691 Iout.t98 VGND 0.02304f
C20692 Iout.n206 VGND 0.05124f
C20693 Iout.n207 VGND 0.02606f
C20694 Iout.n208 VGND 0.14126f
C20695 Iout.n209 VGND 0.04775f
C20696 Iout.t94 VGND 0.02304f
C20697 Iout.n210 VGND 0.05124f
C20698 Iout.n211 VGND 0.02606f
C20699 Iout.n212 VGND 0.14126f
C20700 Iout.n213 VGND 0.04775f
C20701 Iout.t4 VGND 0.02304f
C20702 Iout.n214 VGND 0.05124f
C20703 Iout.n215 VGND 0.02606f
C20704 Iout.n216 VGND 0.14126f
C20705 Iout.n217 VGND 0.04775f
C20706 Iout.t50 VGND 0.02304f
C20707 Iout.n218 VGND 0.05124f
C20708 Iout.n219 VGND 0.02606f
C20709 Iout.n220 VGND 0.14126f
C20710 Iout.n221 VGND 0.04775f
C20711 Iout.t114 VGND 0.02304f
C20712 Iout.n222 VGND 0.05124f
C20713 Iout.n223 VGND 0.02606f
C20714 Iout.n224 VGND 0.14126f
C20715 Iout.n225 VGND 0.04775f
C20716 Iout.t126 VGND 0.02304f
C20717 Iout.n226 VGND 0.05124f
C20718 Iout.n227 VGND 0.02606f
C20719 Iout.n228 VGND 0.04775f
C20720 Iout.n229 VGND 0.14126f
C20721 Iout.n230 VGND 0.23929f
C20722 Iout.n231 VGND 0.04775f
C20723 Iout.t40 VGND 0.02304f
C20724 Iout.n232 VGND 0.05124f
C20725 Iout.n233 VGND 0.02606f
C20726 Iout.n234 VGND 0.04775f
C20727 Iout.t66 VGND 0.02304f
C20728 Iout.n235 VGND 0.05124f
C20729 Iout.n236 VGND 0.02606f
C20730 Iout.n237 VGND 0.04775f
C20731 Iout.t205 VGND 0.02304f
C20732 Iout.n238 VGND 0.05124f
C20733 Iout.n239 VGND 0.02606f
C20734 Iout.n240 VGND 0.04775f
C20735 Iout.t131 VGND 0.02304f
C20736 Iout.n241 VGND 0.05124f
C20737 Iout.n242 VGND 0.02606f
C20738 Iout.n243 VGND 0.04775f
C20739 Iout.t6 VGND 0.02304f
C20740 Iout.n244 VGND 0.05124f
C20741 Iout.n245 VGND 0.02606f
C20742 Iout.n246 VGND 0.04775f
C20743 Iout.t174 VGND 0.02304f
C20744 Iout.n247 VGND 0.05124f
C20745 Iout.n248 VGND 0.02606f
C20746 Iout.n249 VGND 0.04775f
C20747 Iout.t105 VGND 0.02304f
C20748 Iout.n250 VGND 0.05124f
C20749 Iout.n251 VGND 0.02606f
C20750 Iout.t198 VGND 0.02304f
C20751 Iout.n252 VGND 0.05124f
C20752 Iout.n253 VGND 0.02606f
C20753 Iout.n254 VGND 0.04775f
C20754 Iout.t111 VGND 0.02304f
C20755 Iout.n255 VGND 0.05124f
C20756 Iout.n256 VGND 0.02606f
C20757 Iout.n257 VGND 0.04775f
C20758 Iout.n258 VGND 0.23929f
C20759 Iout.t32 VGND 0.02304f
C20760 Iout.n259 VGND 0.05124f
C20761 Iout.n260 VGND 0.02606f
C20762 Iout.n261 VGND 0.04775f
C20763 Iout.n262 VGND 0.23929f
C20764 Iout.n263 VGND 0.23929f
C20765 Iout.n264 VGND 0.04775f
C20766 Iout.t92 VGND 0.02304f
C20767 Iout.n265 VGND 0.05124f
C20768 Iout.n266 VGND 0.02606f
C20769 Iout.n267 VGND 0.04775f
C20770 Iout.n268 VGND 0.23929f
C20771 Iout.n269 VGND 0.23929f
C20772 Iout.n270 VGND 0.04775f
C20773 Iout.t37 VGND 0.02304f
C20774 Iout.n271 VGND 0.05124f
C20775 Iout.n272 VGND 0.02606f
C20776 Iout.n273 VGND 0.04775f
C20777 Iout.n274 VGND 0.23929f
C20778 Iout.n275 VGND 0.23929f
C20779 Iout.n276 VGND 0.04775f
C20780 Iout.t70 VGND 0.02304f
C20781 Iout.n277 VGND 0.05124f
C20782 Iout.n278 VGND 0.02606f
C20783 Iout.n279 VGND 0.04775f
C20784 Iout.n280 VGND 0.23929f
C20785 Iout.n281 VGND 0.23929f
C20786 Iout.n282 VGND 0.04775f
C20787 Iout.t237 VGND 0.02304f
C20788 Iout.n283 VGND 0.05124f
C20789 Iout.n284 VGND 0.02606f
C20790 Iout.n285 VGND 0.04775f
C20791 Iout.n286 VGND 0.23929f
C20792 Iout.n287 VGND 0.23929f
C20793 Iout.n288 VGND 0.04775f
C20794 Iout.t228 VGND 0.02304f
C20795 Iout.n289 VGND 0.05124f
C20796 Iout.n290 VGND 0.02606f
C20797 Iout.n291 VGND 0.04775f
C20798 Iout.n292 VGND 0.23929f
C20799 Iout.n293 VGND 0.23929f
C20800 Iout.n294 VGND 0.04775f
C20801 Iout.t24 VGND 0.02304f
C20802 Iout.n295 VGND 0.05124f
C20803 Iout.n296 VGND 0.02606f
C20804 Iout.n297 VGND 0.04775f
C20805 Iout.n298 VGND 0.23929f
C20806 Iout.n299 VGND 0.23929f
C20807 Iout.n300 VGND 0.04775f
C20808 Iout.t189 VGND 0.02304f
C20809 Iout.n301 VGND 0.05124f
C20810 Iout.n302 VGND 0.02606f
C20811 Iout.n303 VGND 0.04775f
C20812 Iout.n304 VGND 0.23929f
C20813 Iout.t26 VGND 0.02304f
C20814 Iout.n305 VGND 0.05124f
C20815 Iout.n306 VGND 0.02606f
C20816 Iout.n307 VGND 0.04775f
C20817 Iout.t80 VGND 0.02304f
C20818 Iout.n308 VGND 0.05124f
C20819 Iout.n309 VGND 0.02606f
C20820 Iout.n310 VGND 0.04775f
C20821 Iout.t226 VGND 0.02304f
C20822 Iout.n311 VGND 0.05124f
C20823 Iout.n312 VGND 0.02606f
C20824 Iout.n313 VGND 0.04775f
C20825 Iout.t83 VGND 0.02304f
C20826 Iout.n314 VGND 0.05124f
C20827 Iout.n315 VGND 0.02606f
C20828 Iout.n316 VGND 0.04775f
C20829 Iout.t113 VGND 0.02304f
C20830 Iout.n317 VGND 0.05124f
C20831 Iout.n318 VGND 0.02606f
C20832 Iout.n319 VGND 0.04775f
C20833 Iout.t67 VGND 0.02304f
C20834 Iout.n320 VGND 0.05124f
C20835 Iout.n321 VGND 0.02606f
C20836 Iout.n322 VGND 0.04775f
C20837 Iout.t18 VGND 0.02304f
C20838 Iout.n323 VGND 0.05124f
C20839 Iout.n324 VGND 0.02606f
C20840 Iout.n325 VGND 0.04775f
C20841 Iout.t46 VGND 0.02304f
C20842 Iout.n326 VGND 0.05124f
C20843 Iout.n327 VGND 0.02606f
C20844 Iout.n328 VGND 0.04775f
C20845 Iout.t150 VGND 0.02304f
C20846 Iout.n329 VGND 0.05124f
C20847 Iout.n330 VGND 0.02606f
C20848 Iout.n331 VGND 0.04775f
C20849 Iout.n332 VGND 0.23929f
C20850 Iout.t182 VGND 0.02304f
C20851 Iout.n333 VGND 0.05124f
C20852 Iout.n334 VGND 0.02606f
C20853 Iout.n335 VGND 0.04775f
C20854 Iout.t209 VGND 0.02304f
C20855 Iout.n336 VGND 0.05124f
C20856 Iout.n337 VGND 0.02606f
C20857 Iout.n338 VGND 0.04775f
C20858 Iout.t225 VGND 0.02304f
C20859 Iout.n339 VGND 0.05124f
C20860 Iout.n340 VGND 0.02606f
C20861 Iout.n341 VGND 0.04775f
C20862 Iout.t219 VGND 0.02304f
C20863 Iout.n342 VGND 0.05124f
C20864 Iout.n343 VGND 0.02606f
C20865 Iout.n344 VGND 0.04775f
C20866 Iout.t192 VGND 0.02304f
C20867 Iout.n345 VGND 0.05124f
C20868 Iout.n346 VGND 0.02606f
C20869 Iout.n347 VGND 0.04775f
C20870 Iout.t149 VGND 0.02304f
C20871 Iout.n348 VGND 0.05124f
C20872 Iout.n349 VGND 0.02606f
C20873 Iout.n350 VGND 0.04775f
C20874 Iout.t207 VGND 0.02304f
C20875 Iout.n351 VGND 0.05124f
C20876 Iout.n352 VGND 0.02606f
C20877 Iout.n353 VGND 0.04775f
C20878 Iout.t145 VGND 0.02304f
C20879 Iout.n354 VGND 0.05124f
C20880 Iout.n355 VGND 0.02606f
C20881 Iout.n356 VGND 0.04775f
C20882 Iout.t115 VGND 0.02304f
C20883 Iout.n357 VGND 0.05124f
C20884 Iout.n358 VGND 0.02606f
C20885 Iout.n359 VGND 0.04775f
C20886 Iout.t76 VGND 0.02304f
C20887 Iout.n360 VGND 0.05124f
C20888 Iout.n361 VGND 0.02606f
C20889 Iout.n362 VGND 0.04775f
C20890 Iout.t251 VGND 0.02304f
C20891 Iout.n363 VGND 0.05124f
C20892 Iout.n364 VGND 0.02606f
C20893 Iout.n365 VGND 0.04775f
C20894 Iout.t187 VGND 0.02304f
C20895 Iout.n366 VGND 0.05124f
C20896 Iout.n367 VGND 0.02606f
C20897 Iout.n368 VGND 0.04775f
C20898 Iout.n369 VGND 0.23929f
C20899 Iout.t190 VGND 0.02304f
C20900 Iout.n370 VGND 0.05124f
C20901 Iout.n371 VGND 0.02606f
C20902 Iout.n372 VGND 0.04775f
C20903 Iout.n373 VGND 0.23929f
C20904 Iout.n374 VGND 0.23929f
C20905 Iout.n375 VGND 0.04775f
C20906 Iout.t183 VGND 0.02304f
C20907 Iout.n376 VGND 0.05124f
C20908 Iout.n377 VGND 0.02606f
C20909 Iout.t112 VGND 0.02304f
C20910 Iout.n378 VGND 0.05124f
C20911 Iout.n379 VGND 0.02606f
C20912 Iout.n380 VGND 0.04775f
C20913 Iout.n381 VGND 0.23929f
C20914 Iout.n382 VGND 0.23929f
C20915 Iout.n383 VGND 0.04775f
C20916 Iout.t243 VGND 0.02304f
C20917 Iout.n384 VGND 0.05124f
C20918 Iout.n385 VGND 0.02606f
C20919 Iout.t194 VGND 0.02304f
C20920 Iout.n386 VGND 0.05124f
C20921 Iout.n387 VGND 0.02606f
C20922 Iout.n388 VGND 0.04775f
C20923 Iout.n389 VGND 0.23929f
C20924 Iout.n390 VGND 0.23929f
C20925 Iout.n391 VGND 0.04775f
C20926 Iout.t253 VGND 0.02304f
C20927 Iout.n392 VGND 0.05124f
C20928 Iout.n393 VGND 0.02606f
C20929 Iout.t73 VGND 0.02304f
C20930 Iout.n394 VGND 0.05124f
C20931 Iout.n395 VGND 0.02606f
C20932 Iout.n396 VGND 0.04775f
C20933 Iout.n397 VGND 0.23929f
C20934 Iout.n398 VGND 0.23929f
C20935 Iout.n399 VGND 0.04775f
C20936 Iout.t132 VGND 0.02304f
C20937 Iout.n400 VGND 0.05124f
C20938 Iout.n401 VGND 0.02606f
C20939 Iout.t99 VGND 0.02304f
C20940 Iout.n402 VGND 0.05124f
C20941 Iout.n403 VGND 0.02606f
C20942 Iout.n404 VGND 0.04775f
C20943 Iout.n405 VGND 0.23929f
C20944 Iout.n406 VGND 0.23929f
C20945 Iout.n407 VGND 0.04775f
C20946 Iout.t199 VGND 0.02304f
C20947 Iout.n408 VGND 0.05124f
C20948 Iout.n409 VGND 0.02606f
C20949 Iout.t91 VGND 0.02304f
C20950 Iout.n410 VGND 0.05124f
C20951 Iout.n411 VGND 0.02606f
C20952 Iout.n412 VGND 0.04775f
C20953 Iout.n413 VGND 0.23929f
C20954 Iout.n414 VGND 0.23929f
C20955 Iout.n415 VGND 0.04775f
C20956 Iout.t49 VGND 0.02304f
C20957 Iout.n416 VGND 0.05124f
C20958 Iout.n417 VGND 0.02606f
C20959 Iout.t85 VGND 0.02304f
C20960 Iout.n418 VGND 0.05124f
C20961 Iout.n419 VGND 0.02606f
C20962 Iout.n420 VGND 0.04775f
C20963 Iout.n421 VGND 0.23929f
C20964 Iout.n422 VGND 0.23929f
C20965 Iout.n423 VGND 0.04775f
C20966 Iout.t246 VGND 0.02304f
C20967 Iout.n424 VGND 0.05124f
C20968 Iout.n425 VGND 0.02606f
C20969 Iout.t206 VGND 0.02304f
C20970 Iout.n426 VGND 0.05124f
C20971 Iout.n427 VGND 0.02606f
C20972 Iout.n428 VGND 0.04775f
C20973 Iout.n429 VGND 0.23929f
C20974 Iout.n430 VGND 0.23929f
C20975 Iout.n431 VGND 0.04775f
C20976 Iout.t20 VGND 0.02304f
C20977 Iout.n432 VGND 0.05124f
C20978 Iout.n433 VGND 0.02606f
C20979 Iout.t78 VGND 0.02304f
C20980 Iout.n434 VGND 0.05124f
C20981 Iout.n435 VGND 0.02606f
C20982 Iout.n436 VGND 0.23929f
C20983 Iout.n437 VGND 0.04775f
C20984 Iout.t104 VGND 0.02304f
C20985 Iout.n438 VGND 0.05124f
C20986 Iout.n439 VGND 0.02606f
C20987 Iout.n440 VGND 0.04775f
C20988 Iout.t41 VGND 0.02304f
C20989 Iout.n441 VGND 0.05124f
C20990 Iout.n442 VGND 0.02606f
C20991 Iout.n443 VGND 0.04775f
C20992 Iout.n444 VGND 0.23929f
C20993 Iout.n445 VGND 0.23929f
C20994 Iout.n446 VGND 0.04775f
C20995 Iout.t176 VGND 0.02304f
C20996 Iout.n447 VGND 0.05124f
C20997 Iout.n448 VGND 0.02606f
C20998 Iout.t164 VGND 0.02304f
C20999 Iout.n449 VGND 0.05124f
C21000 Iout.n450 VGND 0.02606f
C21001 Iout.n451 VGND 0.04775f
C21002 Iout.t186 VGND 0.02304f
C21003 Iout.n452 VGND 0.05124f
C21004 Iout.n453 VGND 0.02606f
C21005 Iout.n454 VGND 0.04775f
C21006 Iout.n455 VGND 0.23929f
C21007 Iout.n456 VGND 0.23929f
C21008 Iout.n457 VGND 0.04775f
C21009 Iout.t160 VGND 0.02304f
C21010 Iout.n458 VGND 0.05124f
C21011 Iout.n459 VGND 0.02606f
C21012 Iout.t29 VGND 0.02304f
C21013 Iout.n460 VGND 0.05124f
C21014 Iout.n461 VGND 0.02606f
C21015 Iout.n462 VGND 0.04775f
C21016 Iout.t221 VGND 0.02304f
C21017 Iout.n463 VGND 0.05124f
C21018 Iout.n464 VGND 0.02606f
C21019 Iout.n465 VGND 0.04775f
C21020 Iout.n466 VGND 0.23929f
C21021 Iout.n467 VGND 0.23929f
C21022 Iout.n468 VGND 0.04775f
C21023 Iout.t9 VGND 0.02304f
C21024 Iout.n469 VGND 0.05124f
C21025 Iout.n470 VGND 0.02606f
C21026 Iout.n471 VGND 0.04775f
C21027 Iout.t177 VGND 0.02304f
C21028 Iout.n472 VGND 0.05124f
C21029 Iout.n473 VGND 0.02606f
C21030 Iout.n474 VGND 0.04775f
C21031 Iout.n475 VGND 0.23929f
C21032 Iout.n476 VGND 0.23929f
C21033 Iout.n477 VGND 0.04775f
C21034 Iout.t65 VGND 0.02304f
C21035 Iout.n478 VGND 0.05124f
C21036 Iout.n479 VGND 0.02606f
C21037 Iout.t196 VGND 0.02304f
C21038 Iout.n480 VGND 0.05124f
C21039 Iout.n481 VGND 0.02606f
C21040 Iout.n482 VGND 0.04775f
C21041 Iout.t58 VGND 0.02304f
C21042 Iout.n483 VGND 0.05124f
C21043 Iout.n484 VGND 0.02606f
C21044 Iout.n485 VGND 0.04775f
C21045 Iout.n486 VGND 0.23929f
C21046 Iout.n487 VGND 0.23929f
C21047 Iout.n488 VGND 0.04775f
C21048 Iout.t81 VGND 0.02304f
C21049 Iout.n489 VGND 0.05124f
C21050 Iout.n490 VGND 0.02606f
C21051 Iout.t129 VGND 0.02304f
C21052 Iout.n491 VGND 0.05124f
C21053 Iout.n492 VGND 0.02606f
C21054 Iout.n493 VGND 0.04775f
C21055 Iout.t178 VGND 0.02304f
C21056 Iout.n494 VGND 0.05124f
C21057 Iout.n495 VGND 0.02606f
C21058 Iout.n496 VGND 0.04775f
C21059 Iout.n497 VGND 0.23929f
C21060 Iout.n498 VGND 0.14126f
C21061 Iout.n499 VGND 0.04775f
C21062 Iout.t142 VGND 0.02304f
C21063 Iout.n500 VGND 0.05124f
C21064 Iout.n501 VGND 0.02606f
C21065 Iout.n502 VGND 0.14126f
C21066 Iout.n503 VGND 0.04775f
C21067 Iout.t7 VGND 0.02304f
C21068 Iout.n504 VGND 0.05124f
C21069 Iout.n505 VGND 0.02606f
C21070 Iout.n506 VGND 0.04775f
C21071 Iout.t124 VGND 0.02304f
C21072 Iout.n507 VGND 0.05124f
C21073 Iout.n508 VGND 0.02606f
C21074 Iout.t201 VGND 0.02304f
C21075 Iout.n509 VGND 0.05124f
C21076 Iout.n510 VGND 0.02606f
C21077 Iout.n511 VGND 0.14126f
C21078 Iout.n512 VGND 0.04775f
C21079 Iout.t158 VGND 0.02304f
C21080 Iout.n513 VGND 0.05124f
C21081 Iout.n514 VGND 0.02606f
C21082 Iout.n515 VGND 0.04775f
C21083 Iout.n516 VGND 0.14126f
C21084 Iout.n517 VGND 0.23929f
C21085 Iout.n518 VGND 0.04775f
C21086 Iout.t139 VGND 0.02304f
C21087 Iout.n519 VGND 0.05124f
C21088 Iout.n520 VGND 0.02606f
C21089 Iout.n521 VGND 0.04775f
C21090 Iout.n522 VGND 0.23929f
C21091 Iout.n523 VGND 0.23929f
C21092 Iout.n524 VGND 0.04775f
C21093 Iout.t231 VGND 0.02304f
C21094 Iout.n525 VGND 0.05124f
C21095 Iout.n526 VGND 0.02606f
C21096 Iout.n527 VGND 0.04775f
C21097 Iout.n528 VGND 0.23929f
C21098 Iout.n529 VGND 0.23929f
C21099 Iout.n530 VGND 0.04775f
C21100 Iout.t10 VGND 0.02304f
C21101 Iout.n531 VGND 0.05124f
C21102 Iout.n532 VGND 0.02606f
C21103 Iout.n533 VGND 0.04775f
C21104 Iout.t213 VGND 0.02304f
C21105 Iout.n534 VGND 0.05124f
C21106 Iout.n535 VGND 0.02606f
C21107 Iout.t69 VGND 0.02304f
C21108 Iout.n536 VGND 0.05124f
C21109 Iout.n537 VGND 0.02606f
C21110 Iout.n538 VGND 0.04775f
C21111 Iout.n539 VGND 0.23929f
C21112 Iout.n540 VGND 0.23929f
C21113 Iout.n541 VGND 0.04775f
C21114 Iout.t31 VGND 0.02304f
C21115 Iout.n542 VGND 0.05124f
C21116 Iout.n543 VGND 0.02606f
C21117 Iout.n544 VGND 0.04775f
C21118 Iout.n545 VGND 0.23929f
C21119 Iout.n546 VGND 0.23929f
C21120 Iout.n547 VGND 0.04775f
C21121 Iout.t191 VGND 0.02304f
C21122 Iout.n548 VGND 0.05124f
C21123 Iout.n549 VGND 0.02606f
C21124 Iout.n550 VGND 0.04775f
C21125 Iout.n551 VGND 0.23929f
C21126 Iout.n552 VGND 0.23929f
C21127 Iout.n553 VGND 0.04775f
C21128 Iout.t25 VGND 0.02304f
C21129 Iout.n554 VGND 0.05124f
C21130 Iout.n555 VGND 0.02606f
C21131 Iout.n556 VGND 0.04775f
C21132 Iout.t34 VGND 0.02304f
C21133 Iout.n557 VGND 0.05124f
C21134 Iout.n558 VGND 0.02606f
C21135 Iout.t169 VGND 0.02304f
C21136 Iout.n559 VGND 0.05124f
C21137 Iout.n560 VGND 0.02606f
C21138 Iout.n561 VGND 0.04775f
C21139 Iout.n562 VGND 0.23929f
C21140 Iout.t125 VGND 0.02304f
C21141 Iout.n563 VGND 0.05124f
C21142 Iout.n564 VGND 0.02606f
C21143 Iout.n565 VGND 0.04775f
C21144 Iout.n566 VGND 0.23929f
C21145 Iout.n567 VGND 0.23929f
C21146 Iout.n568 VGND 0.04775f
C21147 Iout.t48 VGND 0.02304f
C21148 Iout.n569 VGND 0.05124f
C21149 Iout.n570 VGND 0.02606f
C21150 Iout.n571 VGND 0.04775f
C21151 Iout.n572 VGND 0.23929f
C21152 Iout.t82 VGND 0.02304f
C21153 Iout.n573 VGND 0.05124f
C21154 Iout.n574 VGND 0.02606f
C21155 Iout.n575 VGND 0.04775f
C21156 Iout.t233 VGND 0.02304f
C21157 Iout.n576 VGND 0.05124f
C21158 Iout.n577 VGND 0.02606f
C21159 Iout.n578 VGND 0.04775f
C21160 Iout.n579 VGND 0.23929f
C21161 Iout.n580 VGND 0.23929f
C21162 Iout.n581 VGND 0.04775f
C21163 Iout.t222 VGND 0.02304f
C21164 Iout.n582 VGND 0.05124f
C21165 Iout.n583 VGND 0.02606f
C21166 Iout.n584 VGND 0.04775f
C21167 Iout.n585 VGND 0.23929f
C21168 Iout.n586 VGND 0.23929f
C21169 Iout.n587 VGND 0.04775f
C21170 Iout.t235 VGND 0.02304f
C21171 Iout.n588 VGND 0.05124f
C21172 Iout.n589 VGND 0.02606f
C21173 Iout.n590 VGND 0.04775f
C21174 Iout.n591 VGND 0.23929f
C21175 Iout.n592 VGND 0.23929f
C21176 Iout.n593 VGND 0.04775f
C21177 Iout.t128 VGND 0.02304f
C21178 Iout.n594 VGND 0.05124f
C21179 Iout.n595 VGND 0.02606f
C21180 Iout.n596 VGND 0.04775f
C21181 Iout.n597 VGND 0.23929f
C21182 Iout.n598 VGND 0.23929f
C21183 Iout.n599 VGND 0.04775f
C21184 Iout.t134 VGND 0.02304f
C21185 Iout.n600 VGND 0.05124f
C21186 Iout.n601 VGND 0.02606f
C21187 Iout.n602 VGND 0.04775f
C21188 Iout.n603 VGND 0.23929f
C21189 Iout.n604 VGND 0.23929f
C21190 Iout.n605 VGND 0.04775f
C21191 Iout.t151 VGND 0.02304f
C21192 Iout.n606 VGND 0.05124f
C21193 Iout.n607 VGND 0.02606f
C21194 Iout.n608 VGND 0.04775f
C21195 Iout.n609 VGND 0.23929f
C21196 Iout.n610 VGND 0.23929f
C21197 Iout.n611 VGND 0.04775f
C21198 Iout.t33 VGND 0.02304f
C21199 Iout.n612 VGND 0.05124f
C21200 Iout.n613 VGND 0.02606f
C21201 Iout.n614 VGND 0.04775f
C21202 Iout.n615 VGND 0.23929f
C21203 Iout.n616 VGND 0.23929f
C21204 Iout.n617 VGND 0.04775f
C21205 Iout.t72 VGND 0.02304f
C21206 Iout.n618 VGND 0.05124f
C21207 Iout.n619 VGND 0.02606f
C21208 Iout.n620 VGND 0.04775f
C21209 Iout.n621 VGND 0.23929f
C21210 Iout.n622 VGND 0.23929f
C21211 Iout.n623 VGND 0.04775f
C21212 Iout.t143 VGND 0.02304f
C21213 Iout.n624 VGND 0.05124f
C21214 Iout.n625 VGND 0.02606f
C21215 Iout.n626 VGND 0.04775f
C21216 Iout.n627 VGND 0.23929f
C21217 Iout.n628 VGND 0.23929f
C21218 Iout.n629 VGND 0.04775f
C21219 Iout.t180 VGND 0.02304f
C21220 Iout.n630 VGND 0.05124f
C21221 Iout.n631 VGND 0.02606f
C21222 Iout.n632 VGND 0.04775f
C21223 Iout.n633 VGND 0.23929f
C21224 Iout.n634 VGND 0.23929f
C21225 Iout.n635 VGND 0.04775f
C21226 Iout.t12 VGND 0.02304f
C21227 Iout.n636 VGND 0.05124f
C21228 Iout.n637 VGND 0.02606f
C21229 Iout.n638 VGND 0.04775f
C21230 Iout.n639 VGND 0.23929f
C21231 Iout.n640 VGND 0.23929f
C21232 Iout.n641 VGND 0.04775f
C21233 Iout.t234 VGND 0.02304f
C21234 Iout.n642 VGND 0.05124f
C21235 Iout.n643 VGND 0.02606f
C21236 Iout.n644 VGND 0.04775f
C21237 Iout.n645 VGND 0.23929f
C21238 Iout.n646 VGND 0.23929f
C21239 Iout.n647 VGND 0.04775f
C21240 Iout.t63 VGND 0.02304f
C21241 Iout.n648 VGND 0.05124f
C21242 Iout.n649 VGND 0.02606f
C21243 Iout.n650 VGND 0.04775f
C21244 Iout.n651 VGND 0.23929f
C21245 Iout.n652 VGND 0.23929f
C21246 Iout.n653 VGND 0.04775f
C21247 Iout.t138 VGND 0.02304f
C21248 Iout.n654 VGND 0.05124f
C21249 Iout.n655 VGND 0.02606f
C21250 Iout.n656 VGND 0.04775f
C21251 Iout.t175 VGND 0.02304f
C21252 Iout.n657 VGND 0.05124f
C21253 Iout.n658 VGND 0.02606f
C21254 Iout.n659 VGND 0.04775f
C21255 Iout.t223 VGND 0.02304f
C21256 Iout.n660 VGND 0.05124f
C21257 Iout.n661 VGND 0.02606f
C21258 Iout.n662 VGND 0.04775f
C21259 Iout.t17 VGND 0.02304f
C21260 Iout.n663 VGND 0.05124f
C21261 Iout.n664 VGND 0.02606f
C21262 Iout.n665 VGND 0.04775f
C21263 Iout.t161 VGND 0.02304f
C21264 Iout.n666 VGND 0.05124f
C21265 Iout.n667 VGND 0.02606f
C21266 Iout.n668 VGND 0.04775f
C21267 Iout.t23 VGND 0.02304f
C21268 Iout.n669 VGND 0.05124f
C21269 Iout.n670 VGND 0.02606f
C21270 Iout.n671 VGND 0.04775f
C21271 Iout.t84 VGND 0.02304f
C21272 Iout.n672 VGND 0.05124f
C21273 Iout.n673 VGND 0.02606f
C21274 Iout.n674 VGND 0.04775f
C21275 Iout.t215 VGND 0.02304f
C21276 Iout.n675 VGND 0.05124f
C21277 Iout.n676 VGND 0.02606f
C21278 Iout.n677 VGND 0.04775f
C21279 Iout.t249 VGND 0.02304f
C21280 Iout.n678 VGND 0.05124f
C21281 Iout.n679 VGND 0.02606f
C21282 Iout.n680 VGND 0.04775f
C21283 Iout.t100 VGND 0.02304f
C21284 Iout.n681 VGND 0.05124f
C21285 Iout.n682 VGND 0.02606f
C21286 Iout.n683 VGND 0.04775f
C21287 Iout.t193 VGND 0.02304f
C21288 Iout.n684 VGND 0.05124f
C21289 Iout.n685 VGND 0.02606f
C21290 Iout.n686 VGND 0.04775f
C21291 Iout.t156 VGND 0.02304f
C21292 Iout.n687 VGND 0.05124f
C21293 Iout.n688 VGND 0.02606f
C21294 Iout.n689 VGND 0.04775f
C21295 Iout.t202 VGND 0.02304f
C21296 Iout.n690 VGND 0.05124f
C21297 Iout.n691 VGND 0.02606f
C21298 Iout.t36 VGND 0.02304f
C21299 Iout.n692 VGND 0.05124f
C21300 Iout.n693 VGND 0.02606f
C21301 Iout.n694 VGND 0.04775f
C21302 Iout.t109 VGND 0.02304f
C21303 Iout.n695 VGND 0.05124f
C21304 Iout.n696 VGND 0.02606f
C21305 Iout.n697 VGND 0.04775f
C21306 Iout.n698 VGND 0.23929f
C21307 Iout.t127 VGND 0.02304f
C21308 Iout.n699 VGND 0.05124f
C21309 Iout.n700 VGND 0.02606f
C21310 Iout.n701 VGND 0.04775f
C21311 Iout.n702 VGND 0.23929f
C21312 Iout.n703 VGND 0.23929f
C21313 Iout.n704 VGND 0.04775f
C21314 Iout.t181 VGND 0.02304f
C21315 Iout.n705 VGND 0.05124f
C21316 Iout.n706 VGND 0.02606f
C21317 Iout.n707 VGND 0.04775f
C21318 Iout.n708 VGND 0.23929f
C21319 Iout.n709 VGND 0.23929f
C21320 Iout.n710 VGND 0.04775f
C21321 Iout.t71 VGND 0.02304f
C21322 Iout.n711 VGND 0.05124f
C21323 Iout.n712 VGND 0.02606f
C21324 Iout.n713 VGND 0.04775f
C21325 Iout.n714 VGND 0.23929f
C21326 Iout.n715 VGND 0.23929f
C21327 Iout.n716 VGND 0.04775f
C21328 Iout.t152 VGND 0.02304f
C21329 Iout.n717 VGND 0.05124f
C21330 Iout.n718 VGND 0.02606f
C21331 Iout.n719 VGND 0.04775f
C21332 Iout.n720 VGND 0.23929f
C21333 Iout.n721 VGND 0.23929f
C21334 Iout.n722 VGND 0.04775f
C21335 Iout.t217 VGND 0.02304f
C21336 Iout.n723 VGND 0.05124f
C21337 Iout.n724 VGND 0.02606f
C21338 Iout.n725 VGND 0.04775f
C21339 Iout.n726 VGND 0.23929f
C21340 Iout.n727 VGND 0.23929f
C21341 Iout.n728 VGND 0.04775f
C21342 Iout.t3 VGND 0.02304f
C21343 Iout.n729 VGND 0.05124f
C21344 Iout.n730 VGND 0.02606f
C21345 Iout.n731 VGND 0.04775f
C21346 Iout.n732 VGND 0.23929f
C21347 Iout.n733 VGND 0.23929f
C21348 Iout.n734 VGND 0.04775f
C21349 Iout.t77 VGND 0.02304f
C21350 Iout.n735 VGND 0.05124f
C21351 Iout.n736 VGND 0.02606f
C21352 Iout.n737 VGND 0.04775f
C21353 Iout.n738 VGND 0.23929f
C21354 Iout.n739 VGND 0.23929f
C21355 Iout.n740 VGND 0.04775f
C21356 Iout.t35 VGND 0.02304f
C21357 Iout.n741 VGND 0.05124f
C21358 Iout.n742 VGND 0.02606f
C21359 Iout.n743 VGND 0.04775f
C21360 Iout.n744 VGND 0.23929f
C21361 Iout.n745 VGND 0.23929f
C21362 Iout.n746 VGND 0.04775f
C21363 Iout.t250 VGND 0.02304f
C21364 Iout.n747 VGND 0.05124f
C21365 Iout.n748 VGND 0.02606f
C21366 Iout.n749 VGND 0.04775f
C21367 Iout.n750 VGND 0.23929f
C21368 Iout.n751 VGND 0.23929f
C21369 Iout.n752 VGND 0.04775f
C21370 Iout.t122 VGND 0.02304f
C21371 Iout.n753 VGND 0.05124f
C21372 Iout.n754 VGND 0.02606f
C21373 Iout.n755 VGND 0.04775f
C21374 Iout.n756 VGND 0.23929f
C21375 Iout.n757 VGND 0.23929f
C21376 Iout.n758 VGND 0.04775f
C21377 Iout.t95 VGND 0.02304f
C21378 Iout.n759 VGND 0.05124f
C21379 Iout.n760 VGND 0.02606f
C21380 Iout.n761 VGND 0.04775f
C21381 Iout.n762 VGND 0.23929f
C21382 Iout.n763 VGND 0.23929f
C21383 Iout.n764 VGND 0.04775f
C21384 Iout.t101 VGND 0.02304f
C21385 Iout.n765 VGND 0.05124f
C21386 Iout.n766 VGND 0.02606f
C21387 Iout.n767 VGND 0.04775f
C21388 Iout.n768 VGND 0.23929f
C21389 Iout.n769 VGND 0.23929f
C21390 Iout.n770 VGND 0.04775f
C21391 Iout.t220 VGND 0.02304f
C21392 Iout.n771 VGND 0.05124f
C21393 Iout.n772 VGND 0.02606f
C21394 Iout.n773 VGND 0.04775f
C21395 Iout.n774 VGND 0.23929f
C21396 Iout.n775 VGND 0.23929f
C21397 Iout.n776 VGND 0.04775f
C21398 Iout.t44 VGND 0.02304f
C21399 Iout.n777 VGND 0.05124f
C21400 Iout.n778 VGND 0.02606f
C21401 Iout.n779 VGND 0.04775f
C21402 Iout.n780 VGND 0.23929f
C21403 Iout.t241 VGND 0.02304f
C21404 Iout.n781 VGND 0.05124f
C21405 Iout.n782 VGND 0.02606f
C21406 Iout.n783 VGND 0.04775f
C21407 Iout.t140 VGND 0.02304f
C21408 Iout.n784 VGND 0.05124f
C21409 Iout.n785 VGND 0.02606f
C21410 Iout.n786 VGND 0.04775f
C21411 Iout.t252 VGND 0.02304f
C21412 Iout.n787 VGND 0.05124f
C21413 Iout.n788 VGND 0.02606f
C21414 Iout.n789 VGND 0.04775f
C21415 Iout.t38 VGND 0.02304f
C21416 Iout.n790 VGND 0.05124f
C21417 Iout.n791 VGND 0.02606f
C21418 Iout.n792 VGND 0.04775f
C21419 Iout.t166 VGND 0.02304f
C21420 Iout.n793 VGND 0.05124f
C21421 Iout.n794 VGND 0.02606f
C21422 Iout.n795 VGND 0.04775f
C21423 Iout.t43 VGND 0.02304f
C21424 Iout.n796 VGND 0.05124f
C21425 Iout.n797 VGND 0.02606f
C21426 Iout.n798 VGND 0.04775f
C21427 Iout.t185 VGND 0.02304f
C21428 Iout.n799 VGND 0.05124f
C21429 Iout.n800 VGND 0.02606f
C21430 Iout.n801 VGND 0.04775f
C21431 Iout.t210 VGND 0.02304f
C21432 Iout.n802 VGND 0.05124f
C21433 Iout.n803 VGND 0.02606f
C21434 Iout.n804 VGND 0.04775f
C21435 Iout.t96 VGND 0.02304f
C21436 Iout.n805 VGND 0.05124f
C21437 Iout.n806 VGND 0.02606f
C21438 Iout.n807 VGND 0.04775f
C21439 Iout.t162 VGND 0.02304f
C21440 Iout.n808 VGND 0.05124f
C21441 Iout.n809 VGND 0.02606f
C21442 Iout.n810 VGND 0.04775f
C21443 Iout.t62 VGND 0.02304f
C21444 Iout.n811 VGND 0.05124f
C21445 Iout.n812 VGND 0.02606f
C21446 Iout.n813 VGND 0.04775f
C21447 Iout.t87 VGND 0.02304f
C21448 Iout.n814 VGND 0.05124f
C21449 Iout.n815 VGND 0.02606f
C21450 Iout.n816 VGND 0.04775f
C21451 Iout.t2 VGND 0.02304f
C21452 Iout.n817 VGND 0.05124f
C21453 Iout.n818 VGND 0.02606f
C21454 Iout.n819 VGND 0.04775f
C21455 Iout.t64 VGND 0.02304f
C21456 Iout.n820 VGND 0.05124f
C21457 Iout.n821 VGND 0.02606f
C21458 Iout.n822 VGND 0.04775f
C21459 Iout.t52 VGND 0.02304f
C21460 Iout.n823 VGND 0.05124f
C21461 Iout.n824 VGND 0.02606f
C21462 Iout.n825 VGND 0.04775f
C21463 Iout.n826 VGND 0.23929f
C21464 Iout.t5 VGND 0.02304f
C21465 Iout.n827 VGND 0.05124f
C21466 Iout.n828 VGND 0.02606f
C21467 Iout.n829 VGND 0.08168f
C21468 Iout.n830 VGND 0.49611f
C21469 Iout.n831 VGND 0.04775f
C21470 Iout.t51 VGND 0.02304f
C21471 Iout.n832 VGND 0.05124f
C21472 Iout.n833 VGND 0.02606f
C21473 Iout.t224 VGND 0.02304f
C21474 Iout.n834 VGND 0.05124f
C21475 Iout.n835 VGND 0.02606f
C21476 Iout.n836 VGND 0.04775f
C21477 Iout.n837 VGND 0.49611f
C21478 Iout.n838 VGND 0.08168f
C21479 Iout.t68 VGND 0.02304f
C21480 Iout.n839 VGND 0.05124f
C21481 Iout.n840 VGND 0.02606f
C21482 Iout.t230 VGND 0.02304f
C21483 Iout.n841 VGND 0.05124f
C21484 Iout.n842 VGND 0.02606f
C21485 Iout.n843 VGND 0.08168f
C21486 Iout.n844 VGND 0.49611f
C21487 Iout.n845 VGND 0.04775f
C21488 Iout.t97 VGND 0.02304f
C21489 Iout.n846 VGND 0.05124f
C21490 Iout.n847 VGND 0.02606f
C21491 Iout.t136 VGND 0.02304f
C21492 Iout.n848 VGND 0.05124f
C21493 Iout.n849 VGND 0.02606f
C21494 Iout.n850 VGND 0.04775f
C21495 Iout.n851 VGND 0.49611f
C21496 Iout.n852 VGND 0.08168f
C21497 Iout.t148 VGND 0.02304f
C21498 Iout.n853 VGND 0.05124f
C21499 Iout.n854 VGND 0.02606f
C21500 Iout.t16 VGND 0.02304f
C21501 Iout.n855 VGND 0.05124f
C21502 Iout.n856 VGND 0.02606f
C21503 Iout.n857 VGND 0.08168f
C21504 Iout.n858 VGND 0.49611f
C21505 Iout.n859 VGND 0.04775f
C21506 Iout.t167 VGND 0.02304f
C21507 Iout.n860 VGND 0.05124f
C21508 Iout.n861 VGND 0.02606f
C21509 Iout.t11 VGND 0.02304f
C21510 Iout.n862 VGND 0.05124f
C21511 Iout.n863 VGND 0.02606f
C21512 Iout.n864 VGND 0.04775f
C21513 Iout.n865 VGND 0.49611f
C21514 Iout.n866 VGND 0.08168f
C21515 Iout.t130 VGND 0.02304f
C21516 Iout.n867 VGND 0.05124f
C21517 Iout.n868 VGND 0.02606f
C21518 Iout.t110 VGND 0.02304f
C21519 Iout.n869 VGND 0.05124f
C21520 Iout.n870 VGND 0.02606f
C21521 Iout.n871 VGND 0.08168f
C21522 Iout.n872 VGND 0.49611f
C21523 Iout.n873 VGND 0.04775f
C21524 Iout.t232 VGND 0.02304f
C21525 Iout.n874 VGND 0.05124f
C21526 Iout.n875 VGND 0.02606f
C21527 Iout.t102 VGND 0.02304f
C21528 Iout.n876 VGND 0.05124f
C21529 Iout.n877 VGND 0.02606f
C21530 Iout.n878 VGND 0.04775f
C21531 Iout.n879 VGND 0.49611f
C21532 Iout.n880 VGND 0.08168f
C21533 Iout.t42 VGND 0.02304f
C21534 Iout.n881 VGND 0.05124f
C21535 Iout.n882 VGND 0.02606f
C21536 Iout.t57 VGND 0.02304f
C21537 Iout.n883 VGND 0.05124f
C21538 Iout.n884 VGND 0.02606f
C21539 Iout.n885 VGND 0.08168f
C21540 Iout.n886 VGND 0.49611f
C21541 Iout.n887 VGND 0.04775f
C21542 Iout.t245 VGND 0.02304f
C21543 Iout.n888 VGND 0.05124f
C21544 Iout.n889 VGND 0.02606f
C21545 Iout.t107 VGND 0.02304f
C21546 Iout.n890 VGND 0.05124f
C21547 Iout.n891 VGND 0.02606f
C21548 Iout.n892 VGND 0.04775f
C21549 Iout.n893 VGND 0.49611f
C21550 Iout.n894 VGND 0.08168f
C21551 Iout.t54 VGND 0.02304f
C21552 Iout.n895 VGND 0.05124f
C21553 Iout.n896 VGND 0.02606f
C21554 Iout.t218 VGND 0.02304f
C21555 Iout.n897 VGND 0.05124f
C21556 Iout.n898 VGND 0.02606f
C21557 Iout.n899 VGND 0.08168f
C21558 Iout.n900 VGND 0.49611f
C21559 Iout.n901 VGND 0.04775f
C21560 Iout.t30 VGND 0.02304f
C21561 Iout.n902 VGND 0.05124f
C21562 Iout.n903 VGND 0.02606f
C21563 Iout.t236 VGND 0.02304f
C21564 Iout.n904 VGND 0.05124f
C21565 Iout.n905 VGND 0.02606f
C21566 Iout.n906 VGND 0.04775f
C21567 Iout.n907 VGND 0.49611f
C21568 Iout.n908 VGND 0.08168f
C21569 Iout.t108 VGND 0.02304f
C21570 Iout.n909 VGND 0.05124f
C21571 Iout.n910 VGND 0.02606f
C21572 Iout.t121 VGND 0.02304f
C21573 Iout.n911 VGND 0.05124f
C21574 Iout.n912 VGND 0.02606f
C21575 Iout.n913 VGND 0.08168f
C21576 Iout.n914 VGND 0.49611f
C21577 Iout.n915 VGND 0.04775f
C21578 Iout.t227 VGND 0.02304f
C21579 Iout.n916 VGND 0.05124f
C21580 Iout.n917 VGND 0.02606f
C21581 Iout.t27 VGND 0.02304f
C21582 Iout.n918 VGND 0.05124f
C21583 Iout.n919 VGND 0.02606f
C21584 Iout.n920 VGND 0.04775f
C21585 Iout.n921 VGND 0.49611f
C21586 Iout.n922 VGND 0.08168f
C21587 Iout.t47 VGND 0.02304f
C21588 Iout.n923 VGND 0.05124f
C21589 Iout.n924 VGND 0.02606f
C21590 Iout.n925 VGND 0.08168f
C21591 Iout.t163 VGND 0.02304f
C21592 Iout.n926 VGND 0.05124f
C21593 Iout.n927 VGND 0.02606f
C21594 Iout.n928 VGND 0.08168f
C21595 Iout.n929 VGND 0.49611f
C21596 Iout.n930 VGND 0.04775f
C21597 Iout.t19 VGND 0.02304f
C21598 Iout.n931 VGND 0.05124f
C21599 Iout.n932 VGND 0.02606f
C21600 Iout.n933 VGND 0.04775f
C21601 Iout.t1 VGND 0.02304f
C21602 Iout.n934 VGND 0.05124f
C21603 Iout.n935 VGND 0.20242f
C21604 Iout.n936 VGND 2.65139f
C21605 Iout.n937 VGND 1.25122f
C21606 Iout.t159 VGND 0.02304f
C21607 Iout.n938 VGND 0.05124f
C21608 Iout.n939 VGND 0.20242f
C21609 Iout.n940 VGND 0.04775f
C21610 Iout.n941 VGND 0.23929f
C21611 Iout.n942 VGND 0.23929f
C21612 Iout.n943 VGND 0.04775f
C21613 Iout.t137 VGND 0.02304f
C21614 Iout.n944 VGND 0.05124f
C21615 Iout.n945 VGND 0.02606f
C21616 Iout.n946 VGND 0.04775f
C21617 Iout.n947 VGND 0.23929f
C21618 Iout.n948 VGND 0.23929f
C21619 Iout.n949 VGND 0.04775f
C21620 Iout.t141 VGND 0.02304f
C21621 Iout.n950 VGND 0.05124f
C21622 Iout.n951 VGND 0.02606f
C21623 Iout.n952 VGND 0.04775f
C21624 Iout.t239 VGND 0.02304f
C21625 Iout.n953 VGND 0.05124f
C21626 Iout.n954 VGND 0.20242f
C21627 Iout.n955 VGND 1.25122f
C21628 Iout.n956 VGND 1.25122f
C21629 Iout.t200 VGND 0.02304f
C21630 Iout.n957 VGND 0.05124f
C21631 Iout.n958 VGND 0.20242f
C21632 Iout.n959 VGND 0.04775f
C21633 Iout.n960 VGND 0.23929f
C21634 Iout.n961 VGND 0.23929f
C21635 Iout.n962 VGND 0.04775f
C21636 Iout.t238 VGND 0.02304f
C21637 Iout.n963 VGND 0.05124f
C21638 Iout.n964 VGND 0.02606f
C21639 Iout.n965 VGND 0.04775f
C21640 Iout.n966 VGND 0.23929f
C21641 Iout.n967 VGND 0.23929f
C21642 Iout.n968 VGND 0.04775f
C21643 Iout.t135 VGND 0.02304f
C21644 Iout.n969 VGND 0.05124f
C21645 Iout.n970 VGND 0.02606f
C21646 Iout.n971 VGND 0.04775f
C21647 Iout.t93 VGND 0.02304f
C21648 Iout.n972 VGND 0.05124f
C21649 Iout.n973 VGND 0.20242f
C21650 Iout.n974 VGND 1.25122f
C21651 Iout.n975 VGND 1.25122f
C21652 Iout.t208 VGND 0.02304f
C21653 Iout.n976 VGND 0.05124f
C21654 Iout.n977 VGND 0.20242f
C21655 Iout.n978 VGND 0.04775f
C21656 Iout.n979 VGND 0.23929f
C21657 Iout.n980 VGND 0.23929f
C21658 Iout.n981 VGND 0.04775f
C21659 Iout.t120 VGND 0.02304f
C21660 Iout.n982 VGND 0.05124f
C21661 Iout.n983 VGND 0.02606f
C21662 Iout.n984 VGND 0.04775f
C21663 Iout.n985 VGND 0.23929f
C21664 Iout.n986 VGND 0.23929f
C21665 Iout.n987 VGND 0.04775f
C21666 Iout.t74 VGND 0.02304f
C21667 Iout.n988 VGND 0.05124f
C21668 Iout.n989 VGND 0.02606f
C21669 Iout.n990 VGND 0.04775f
C21670 Iout.t144 VGND 0.02304f
C21671 Iout.n991 VGND 0.05124f
C21672 Iout.n992 VGND 0.20242f
C21673 Iout.n993 VGND 1.25122f
C21674 Iout.n994 VGND 1.25122f
C21675 Iout.t86 VGND 0.02304f
C21676 Iout.n995 VGND 0.05124f
C21677 Iout.n996 VGND 0.20242f
C21678 Iout.n997 VGND 0.04775f
C21679 Iout.n998 VGND 0.23929f
C21680 Iout.n999 VGND 0.23929f
C21681 Iout.n1000 VGND 0.04775f
C21682 Iout.t153 VGND 0.02304f
C21683 Iout.n1001 VGND 0.05124f
C21684 Iout.n1002 VGND 0.02606f
C21685 Iout.n1003 VGND 0.04775f
C21686 Iout.n1004 VGND 0.23929f
C21687 Iout.n1005 VGND 0.23929f
C21688 Iout.n1006 VGND 0.04775f
C21689 Iout.t247 VGND 0.02304f
C21690 Iout.n1007 VGND 0.05124f
C21691 Iout.n1008 VGND 0.02606f
C21692 Iout.n1009 VGND 0.04775f
C21693 Iout.t147 VGND 0.02304f
C21694 Iout.n1010 VGND 0.05124f
C21695 Iout.n1011 VGND 0.20242f
C21696 Iout.n1012 VGND 1.25122f
C21697 Iout.n1013 VGND 1.1235f
C21698 Iout.t88 VGND 0.02304f
C21699 Iout.n1014 VGND 0.05124f
C21700 Iout.n1015 VGND 0.20242f
C21701 Iout.n1016 VGND 0.04775f
C21702 Iout.n1017 VGND 0.23929f
C21703 Iout.n1018 VGND 0.14126f
C21704 Iout.n1019 VGND 0.04775f
C21705 Iout.t116 VGND 0.02304f
C21706 Iout.n1020 VGND 0.05124f
C21707 Iout.n1021 VGND 0.20242f
C21708 Iout.n1022 VGND 0.23244f
.ends

